MPQ    }0    h�  h                                                                                 M�Q=b ʅ��������Mo~�A��']h�ӋH�@�ZW�@�!n<w)��v=��}s�s��'QI�<K�m��C&n6��<��I
Op�5�P>��a��."�KZ6�
U��BHdgU��J\Q5�Z|���譳�c@�ش<�G ��T�so�#�va
��W_,�im�Ti#�R-<P�[���HO��i�61�kc?�K �%��Q�z([��V������w�x���T�wx��c���/���݅)�=�K?���\_�)=��S�UH����B�� ݇���o�a�R�śG�ۦ�����`}k�2�馭{ьGY�����ZWC
A��&��b�ʣ|�d-{&��0�h-*�d�\D(���J�l��5�����SI�,B{�k��՗�߇t��SQ
�A}֩�H��Ҵ?����wTM[��ؙ��+�3]�8ٕ��
��Q�������=W12~ '�~���3�.�� �C��wFYY�O{��>����V:B?�ʤ�n��ӝh�R�$�+81�KF=�d�oO���1�`K�ͅ�@�b/ҿ���e��iX��m7����$l�i�|p:U����5�S�����]��^�-.�t!.���o<7�<85�G�wU"����c�I&�Yv�a�W�˛׍�۾-����d���w}5fv�If'�J8�^@����!��x�+�݇
�V"�p��
�}ϟn�j���U��FL:/�J�bk_פ��<���s}����D��7X�cZ�V����U����6�]��n�������_���.�Tdl�x�6�F�%y���%�$��u"�:f�2|�ho��$K������CXffF0֌M2V�x�Gh��Jh��V@5���6�hu���	��7b��p0D
�]���U��Q0�NmW��j��$Wni�sTE�_G׿2#�݁rH��0����
�M�^ YS��h�o����~��@Wh"�&|D$��"�`4t����� �)�!E��;Ԁ���4�m�s�X,� ��>��A�J�ll����g"5�S����1��@�M�_yxV���A�{�K����g���kf�-��L�R��tPn�gӉ����ǪLK{��q� �y�\K�"��3�c5�< ���m,N)	�6Jv���./`�2��cxl���1���9�K$jޠ�hW6�dM������_�l�⚡�q܎� �Q����{��2Ӹ�.Ð`c�IE��?�/6�-�n�y�2��,��;����q��fk��q�V�J�b~d�;��b��n�I\kZ��Wr�ъ��^���
���Q�S]m�g��h�y3j�e~�z%9Ș�BFK<(�Xj�.�'��oIE[>>��|��Q�38�Vh�݉Z@p��no4�PB2�J������'C[XD��*�lh��@��Bo��YڑX��1ė�����x8�n�.<G)�7�Tալ$6�.t��a�}.}*]�A�
��""X/d �W�3��#�	;�@�G���x���'@�i>h�x�x$��>=��oPJ��{�>X��b�,n����y�9p��U�D����;���\�O<���/e�s(�Z�������Ӧ�4����j/A,�P{�u�~��f��!(d�֛��{� 6����Y�g\̒ޣ�ey�-�@��f=���sҟ�*TN��!��|82�-�^�Y��E��ԭR}Uq}"�"(,�_�J��>D�� ��
s-.2��o���6ܦ��4'������f��^I�G7Z���*�ꟾ��H�qj���
�Ë�0ꍠ�|s�U���� �Z�~ct� ;د�K��	���8v��/�� �8z��l��L_��8l�5j+�|�=�QħH
��f(��Z,�Զ��
=�x8�z,��-�r��%��إ7�V��i��0߰��>#�>� BRN׊�Z���P�f'���*��|dD��B���Z�fs�]�Y���kk'�պۉzx�pUP �=R�tV�ܡ3kg�n�9.����H��~�sJ'W�&�F�d����q >c��q�Q�)j�U��2���t��gq�C�4��ԇP�(E2�*�&���yI��?�u��!S`]1��w&/(�����d<.Q���Ы���Iq�fe�^/�j> �b��
f�L�U�?�<W��j0o(��� r��l(��>^Qg<`ҩ޽�mv2`8�!�u_�Hq���O���l�����!8+E=Y���Gi���=4��R�$�Y:{�Z��ʤB 3# �Bئ���;5�)���8�VZ���.N�rE�pm����o���2s;�!�3D���F�(�����,n��Z�˺S$���Z@�� ˦X.Gv����6��N��eq������T���]&{U�R�~[��$��r��]�ħfjE�����&0�%,|�z�3ܒ�	��b�Ǥ��Z���u�#��k�(?G��Ϩ=Lח�����j�f�p����*��34b���˹^�O؜5�k��#vK���Y�no�TfZRr�0ja���H���E%�{�ʬ���]�`uspbۍ�/R߱.����)�>���)D��u*�!Ng�	6ˋt˰y��#�NrK����0:V,�*
V�B�p6;�wS�+s�믽`�X�8���:˶���b�t߬���-�[r��4�p�xxㅓ\?_'��LiI�7� &悔Y���u�.���S=�""\, �O�.�+�%�z2�8�'����V�Da��p�	���_M�H
���:O��Y��X�+$O(|��l�a�w1��=M̲��h�Qd��1H�4*��'XH2zvrR�N�E���lm�©����9o�H�Z&�Hc{^&" �������������7��Y�T�y���0	��$%����1��� ���y�0a���v�U�?*؉�vp����ʣsu
&�v
Y �a_�|M�6�V���]k���f����B�r#,r���qc������O��NIk��^��O\�=�_��2�9}}7-���m�K��h?M���R*��Yv�Flw�Ч�C�.]��"�ni�#�0����g��P��q�pds~fby��zJa��S6���	[�%c�ڝ���(p��tr�%(���I� �H�!N����* a�A��^�w>qeFԡ������k�^��W����c�<��0:AE�RG��qԼ��k,c ���p<9Ho�bJ�3�B?��J^�y�&H�+���ހ�5�:�O�B�G�(\Ėƴ���6E��i�n�]�%����*ؘ�l�_
_l[+;썊�w0H�� ��%":j[�e��q=*L��z���|��i9X�M���'6/���b4��/��O^��A�r�]_�9��]�藜��iD�o!7Uq$��b�� �%����iKn���I��X�����n�:�0?9��j����D��xC�d>�;y)�u5i$�V7����9څ����FE,�$�:�>�I��-~�ҡ�����!Q�G0<�!�[��Fv�v��{օ�M�7����]<����`$�_o|{~��V���j�h �8z�>o��8z���г����(M���k]�Ӿ��v��\��Ǚ�],�cfS�����~blQ�K�h�W�$ �ɞ-��8t��r�J[�S���~�W�?�"�T�j�塨%Gh����)�5A'ф ��s�^;���K}θ��+,燅��V��"�A��v�n�亡�콶+uLU��J��~bFN����4�H%�sx���M)����/X4,jZy^)�6*�*+h�F�R6�m/�B~W�V��F�_-+4.���l?y�����F� �y4"S����$�e"�Ӑ:A��|"ToY�RK�/���,QX!w 0�I2��������@␯d;���A�th0[��$�G7�18Kv#DE�������Q���m�!�&h>���D�rT��<GrS�#���r��0�H/��R
1Z#�9�cY���h n���ݪ~H�@@�سAP��{���WS��t[&+���	)�VELWTԛI�ү(��N��,�MC�����JZ�=Z�����	��$�1L��@�M�Z�VW��gj�fp��T����*�h�
L,���oNQ%���Mw�Ǜ��anxT�������W "����Vf�W�k��Vm��	���k���h.nB���;:c��V�8&�{D�̆�$�n�c��ٿ����&v��
 ��	��|�F��[����������ߛd�xÁ�4������Ez���ߩV��n�n��� �縍;�����LfFAͤ����$~_m�6"=�)��\*�Z<r����GFj�%���?�ҮG��"�!hg�j �?�������3�FF�E޳42��v�]o� �>B�|�0��ΥtVc���������4��2?7	J�xj��=3f p[S0g��C2h�_@��B����w�ˑ�lB��u������x�>�I��G��f��Ti����.o(�a<?�}�I|\��
w&�"�N�d[��W�.�3�'��d'�@��.�
A���3iyE�xm�t��V����P�Ö�%����֯�,NV���y��\j9���UO��� %��pn�7�v<��/ ;8#�6ZK��P������.���Ag�
PYL�y'afXp�('H��"�{�[��L���*\���ޞ?b<�-�닼�l���E�z�5�bhY�I㖋x2:o�����6G�O§}0u]�(ǲϦE�O>��� A�sH
*�svb��M����4�Z��i� �v;.C�b���Nvתř �4~�߹M�(S
13���D͠	<���h1UӐ3�ZΜ ��~��j��K�Z�sӨv�J��7L;�,ߎ�r>����ݼ1lrj�a�����U�"�ޓ�+��/�P��8�x�z���-~l�`K��@��V�s��DL����"#�G{c2N��c���h��	�f"�V`1�F�TD�_�B�Zsb��\"���Bk".��6��x��P;�R_O&1Dšn�d�	��.��eƣEZ�֥��i�W��J&���d�[�5�>^��qׯ��ۡ�_�n�2ֈ�tVO�gCC�Ǜ�E��P�[�(`'�*�@��-y�Lڈ���L��
?�`̴�X#/�|���<i��5F���I���er���	����'
A�^L�?���R�ej\��(�� �d�硲����Q� P`�5޸bvy��8b� �� ��5����i�2lfռ��-�!���=�A�b�[�UMd�Q($�3�����B{'� }���k ڶ���y�N)ȡ8����N��{]��������\uPD�z��AzB�a�f�Z7�G���ψ�.$���U��;ˡ����~#��Ծ�� eL;L���}���j�&ot�5q[��l����8%���w���{��5o�8�*�o\�|4�pz]��
tԝo�?�%�U���Ї���-0�C8p�n��='���+K�my�f�RJ����oO)3OF(�R3(^k��p�(g�v����)G"T)5PR��j<�+�����	{i�������R`�-�bV�
�j�i��fy�>�Q`ք椘�b����g�Ȍ6��
t��y�KNmYA���A��j,&�*���B�s��q�Rw��zS�̢F�1`�\�8�L6:F�y��F���H��gg���%�X pK���?�Pq�t�L�����j&��=Y�6�u�7�+7�%ȫj&_\g��O:�F+�_z�\8֙�B.�>�����a�r�pp�������H�ԫ�Uv�*da�3�r$J�Z|3���\Y�1�M�m��7' �̹��M�4e�C'��uR�H ��i7�=J���<9S�H�m��C�^aK Gcݓ�^0���(���T�h-��'T	�,�%a�j�L���|V�ʷk"��x��P��*31�1W�����E%u�ֆ��X ��X�w�6�U��J�k׭M�����1ԭ��,H��l�t����BL��i݃�46��jV��xϮ�|�]�4��)��k���NؚU�[M�>��@���K�v�nIǞ��b#_C���I�"nD�a�k�'��\� Zv����,%�d��b��z%iH��9ϯMt�� !���M�����p(�rm�%k����Q���tN�o��ȿ���2y-Xw��TF��ل1���!R^�����/<���:�?R�O]�����&uc�g
�p�cH���J��.��ޙ�y���(&C�ʾL[��7�U�O1��" \�Љ��J�6@HAi.Y?��!��:�W"*���lҤ_H�;l���QHI~ ��"�o��@o�qxzz�MҮ�����XHC��:��'����~�4��[� �RAUHg]vG�,B�c3���D �&7����b]�� ���p��1�kwoI��UX�����M�n�e0���'� �8 �X���d��柲���5$#v�q��CJ��`�>6$��/�S:俬�h��H��������!�:?0ה�V�Fџ=�Ek{�������M�䘮2<Z�¾[��Fk6A˜�p�+4��C��s'����3�s�
�n��-�\��]ًp�!*y(w���|�Y7�u<�S���`z
~=�>��b�)�Y����$�Oh�t{r�w�.�̹w}��w�O�'�	i���5v��Kw��j�5��ѿ����^6k���+;�?L+�8� �KV�,��|s��<�n�~��@ec�q0�LpG�J�db!];�� ��VssVm¨-��Z�,XO��Z�Ȉg�v�e L��5�6���Ν�Ӑ�+��_��'.{�lzy��l<F��5y�|ʕ�1$�m"�3:��|]_xo�SYK��z�O��Xܧ0�-2LJg幜%�WАJB�67R��w�h���?�7XȊ&��D�n�-�i�g"Q�cDm���A������!T�&�Gh#�`r��F0f���
����e�Y�*{h������ ~�!U@�s�\D����]��Āt����~Z�)E�E?qԶ(~�*���)��,!��.��1tJ�[��}T����k�w�1�3�@4���U�`V�C��e���%������?��9�L��m�jl���I{ڬ3��B?v�<�x�T�V�!�R�V"t���j�rú���m�f	M	3�;y��]*.�u���8c�8)��qG�V����$��t�^5�����P��k(�b���W�����χT.����:%ָ3x$�O����"EUVI�Dk�=иn��\�O'Ȣ��;���g��f!���纻��qm~ZM�����V�\E<�Z�p�rz۔������Ͻ���n�	R1��>�h4t�j{�/�~���{ ��FA?�jZ��W! U!o?C>���|���i3$V^L$�Ⴅ>&�4��2�}J��R���[N<K��Ηh�V@!��BrJ�R�m��H�gk���a�=\�x����d��G~��J�TKPI�Z��.j��a� l}�V�w3�
�M'"�eKd��1WJh@3��D��3�@IW�����>�ݣ�i�Bpx�]�����t�GP�8�ñY��W�3,�^ �S�f~_�9&X�U
����i�1y$���<,�&/����bZ���E�T;�*��p��A�vP�>�t�f�(�(��=�O���R�Ɯ��Ϲ�\TM�ޙ����-|:{�ȒǺy�C�U��ʖ��x.㑺�2�q��s�H���H}�<��(bٗ�@�>�2� �=sc�����������&4]�@��.��[H�A�}�I��@���R�o�"�TJR���
���Ȧ�0�$��r~^U�U�.e 
�~�zIu�%�K����3�v��p�r�n����\����w�Sl:�j!^��
Z�������⊷���T�x9>�z"�K-Yޖɛ�i��h�V�/?�W'�#5���>N�L��Љ��7fz�������D��B��HZN~����.wrk������xb��PVp<R�&D����V���.��H������:���mW�&�
;d6	&���!>Yj�qh�.����̉��n32���t��g��C�zג�٫PL��({<*�w���sy��ut���e|�`Ӵ��&X/�
���?<�ͺ���N��I'>�e-&����X4�
KLW�'?(��M�0j�6*(>�� �:�b;����	Q��6`N��޳^�vԎ98嫫�\>���jTokl����!��2=Ͼ��}�"��| �pJ$%.��,���B�; 8b����1
��TY#)��8/���A�NK�=o�q�8}{�eG��<업�D:��<���5�y��b(#�P��	D���p
�A�-˜������9Ls�-�	|ve'1�r�����&���� �[�"����X��Q��{&���\ѓ���*�x|O!tz�����+���H���l��P+��+���C�^Q��(�=O��fR����f�TN�PFS�*�53jJͺ^F?��q��� uv�Ď�rm<��>�TD$�RhXj�ᬾM��{�{�b+P�UC�`�bѨ���&��k����>Ӵ��ߨᘔp��sg1�6�[GtAw����Nh���Y}\��K�,A�1* ��B����w$GS�� ���%`o�g8 �:��H��0���)�I����v��p�u�?U�(�� L�QȤm�&܀#YH�hupqtF���\fEJl\�>oO�,+���z��b8�^K]��������a81p�9�����H�$��p����s�l�$���|�#�WIm1?}�MBHR�RY��G/��q�4�Z'���p�KR7c��u������
t��j�9��H���>On^��r T>�-�������an��2�aT7���xs	>��%h��gtԲ���ʒ�����N� �K�*�����]D�.u
����u�� �� 5)��r�X6kò��܄k�v��\x��������j,�&��g�]�D����hҌ����m �E}h�����/W�EJ�&������MM�c�QM��U +v��"���VC�"|�ĝ�n_Ь��e!^��l��S����d�Hybo	,z ���\S������
�S�O�h�p ��r�7�%�=�����~��N�A������X��x
w4�PF�}K�l�Dܡ�^�a�j�E��m�<�1�:7�R�xp��<�����c^���(�p��H���Jv����5�ި���&>�ž�[��Y|�p�O�A���\:+A�*�6;8i���ӡ!�:2!*�́l
5_�T�;�9��H	� 2��"0���D=q��܀�I_��2Җv�RXY(�U�',��w��4y܌����7�A�=z]���G�����ia$�D;\�7����b��. ^���
�_8ƭFMbI9�X)I����nM��0��ˣBf��Q5�����[�dT3&�If߅5�d�Č	�¾�H�;�q�|B����:?a&��4|�c&=җ�[�yz�!��*0r�m�Q�F,lo�{7TT�C�զ��z��k^<�?f�V��>z�#��٪����@�����t�&�.����\�)t��SM��_q]�cr�\��ñZ���:���056S4�ѯۍ~R���@�������T���
�t.v'r�矊	4���`7�u���J� �d���D(��1k�K5��������Ko^1Z���g����+9�҇{�V�����rw�N#�n�8��^��,U�L��J� �b��դB� �~��sn�x�Ry�>-XjZZoStB�ө�5D�|�6��7���o��G�FJ�_#��.V��l����*�F�jy����V��$��"���:��;|��1o��7K��+��W�X���0'e�2ǵ��w��N�2��?i1���G�h��t�ZP�7�~�b�D�MT��^��QA_/m�j�\�D���f�ǀT�rG��V#�R)rY�80!���4
'�K��@�Y��hV�/��~�rI@�~�wX����޳��&t�Y��y7�)�/�E�F���'�ҥ�N��b,\8��	��J��s฀�Cy�R�v1«E@�,�ProV�r����y�Jq��n���޼�Lb��e� N$�N����������x��Dj�M�"����L�T���"����m��]	��P����1.$�H�c��c��#�˔�16���$;��YԌ�uh��M�����x��2 �2�`�?���"뿫�r����'��L��jDO�v}�E05��U�s����n��|C$N�]X�;�l��/qf�4|�"����V~UM��� ͟Ab\`~�Z�rUb����[�����d|󐘴�hO��j�v��^/�+W�iEBF<��i��_X�;mo�7�>�7�|P�����VY���kḁ��O4��*25�J��ʌC ��[IhK�;z�hJm�@<p�B~#&�-���	E�����z_��2�xi1)�g$G�z��֜T�W����&.e�ta�!�}[�6���
m��"���d��nW��3�!�`�@n1Ij-͸��i�_Mx�f����4��P{{��������,Ćx���y��9��U�ML�6�⬡���0�<g��/6PIzjZƞ�1�-�a���K�gA�?UPLD��oy�f~(�η�!���qS�wH�
m\�Gޔ'�#�-7����Ⱥ��m�0\�X�TK�	�2�C3��m%�2y�EK6}���|c(���;�E>U�9 ���s~"R�i���jK%�WdX4�H���鶓�-C��썒D+ժ{��H���f*�hn
�q �aZ��? ���7U�:�Юa ��|~t��O����K����i��veJ���B<	�����V�]��2s�lU��j�ذ��E�X�H�X3��-����8�;��xT�z��-4�Q��m��v1�V�����_���#P�hqwNh�<�6b�!Q�f!ǙM����DR�B�@Z)�ޜ�/���k�3��=�x�Pq�WRU���f��Q<�?��.�*��Y��LU]���W�#u&s��dq�[�B�>Tr�q��͍N�}��d�z2��t��*gB�[C�Mϒ��P7�(�qJ*Pݡ[1y��S�[��h,����`����Ax�/��{���<߻�k���j�I�Ƃe������Ӣx
�V�L��+?�}H�j��(��~ �0�����d��Q��`��ޮ] v/mF8ؾ��Ƣ�f֠�U~xl����㡐!I�y=��̘mQ�K��i�\$`HlL]���)B1p� �!���-ڬ�^�/C)>�8�\涪�;N�0�*�S���,X���B�ҵ&D��7�7�����4愤}���g�䃃�5�m��;�˗��X6����'�4�W����e�Yl4���Z���=&%�1���[��f���0O�X���؞�-f��� ��)|jo�zS�gl2����uP�K�d��ٰ���y���d�e=�:�١�I��ef�v�������H&3�nďHbI^!�Z���:�^��v�������şVdT_3�R�J�j� ����!�30{�-ʽ�Ɉ�`��bL� �����`��xd>�7}�:�^�O��*q�g���6\��t|
�̯��Nc����םa�,\��*{p�B��j��?w�{S�r����`*�b8��:<�#�o�%{F��������Pp�����%?���qL,�#�&�/EY�3�u+˽a9\m �I\���Op�i+�3�zC��8LC�x�4��ŝ��as�p���_[�p�H;����$V ���2$�n�|i���RY�1���M�B;�m�����'�¶Z4�:+')�gk�RR���v�����#�3���Z�9�ЪH����9��^�* �d�HE�w�ܾ<	\�m�fT��|���	�-A%�^����r#��m�����i�F
�*�[<规Q�Is��;��u��*'�t м�m�6Ʃ��F�>k`��ׄ���(~�#��,C%��by�៮�������e�*�#� �����(ײz�*��H����v@�����K�8M�,�z�����v�|}M:�ب�C�̇�?�xn��n��&��\���|����բ��d�ݮb�Az��ּ�+���t�� ڮ��#jDp;rc�%�0���j��N����;y��rL&���w�|XFeM��3z�<�^��ԑŰH���U<��:�1�R��3�"�%�\ήc
��g\pm�rH�J��	�Ӻ�p8ݨJOi&9������<}O'��\u��ŭ�66�i�aⅎ�%&���,�*illH�h_=�O;�6��U�H��) M��"��d��8�q�zs�������M���?X����po�'����R��4K��V��FAS�]�׎�b�N�Yʲ<oFDv�7&Z#
b# :�����^��!C�ItʄX�!���n�L0p]I�]J�.Ã��1�)�d�v�� 7:�5��fħ�$�9�B�d���w�>�7:�"��z!�~����Tqe!�
0�G�LU�F�X�*�{RÇ׾Pw�`qF�I�<�ġ�QT�pU��&˜��!O?���c���N����)��)1���_�#�y�RH&]�[����F^
��C�n���M4SO��V��~��i��>29x��+�ɯ�7�ŏ!tI�8rfԊ䁛�/j����E���Ϛ�Vs~��7�����5ҙ��5����^,im�\�T���k+T�����?V�T�����)�n�ڡ�w��L���J	�ub��_�}�ԗFsi� �^����2X�!�Z����@��jP��B6�]&�Sl,���3a�|_��.1(nl�ټĢq�F�QZyE�y�ݢ$��"	5�:�/�|��>o*��K�Ḛ�XRi�0B�2BA�or������]
,�ߦR8ha��u��7NUT��D��Μc���5Q�z�mC� �w"���T1�GC�}#ɹ.r���0��3�
�?R��<oY?�Mh�)���~Y�@CT����B5ގ����t,#��t4�)���E}n���F�� �\��-1,���dQ����Jk��nõ�ӊ��	�3�-�z1�C�@j�־K:Vh�-�ϋ����	2�IKX�`�L����`Cby�쓬i���8�Q����c�����H/�"*!�������y�Um���	�[l��ܖ�%.<��x"c�F��D�߻�7l�$�L)�T����4�����X�̚<��zi�Ͻ��������Y��A�����E4��p�s�pn��u�ؑ;䡗]��f��k�]eq��j�~Pm_�G "�ZL]\{��Z���r0e_���ŧ��Q��|ҿ���SJ8hj�{jqgs�^��fRX��GF7T���4ˠy�V��o5s�>��.|��ԟ�kVT.[�����]M4�2�j+J[ӌ~�7J�[D�g��ECh�5@W~$B��-����Da젝�]둙��(x$�D�`�G����T�~����.`ngaMC*}�i�ۈ
��-"��'d�W�;w3��U�u��@��L��͓ͧ�vi*�>x>K���^j�*��P6�{�����Y�gVp,�����t�s9�|�U�;��Q���'���Ȉ�<�M�/�
��NZ\��� �HTp� ���&�ZA��P�i��jRXfi��(Pҵ�<%E�����R��El�\�N�ޏ˷sF�-�7F��>�o���rw@_�*P��x�2K���J���M�\���o}��<��(��0�6�>�f rg�s�^���TŞE�Tܒ�}4�v����8�l]I��Z��5&�VG'��݉ߊ���8�
BA��d�Z!�h	�Ud?3�O� Q9�~
r�I�؛51K��,��T�v@�����S��D-�����C�lp��j��"ēa��ѓ�^��@8m���xoĕz��-ʜ�/-��V�E�U^ ��ԥ#kw5��NC�1�F�伤�f�5�g�ǵw��D5�RBw<Z��I�t�d��k��GaxأP�x�R�5����4����.ʇ�ƴ�.�݃�߆�W��\&NN�d�å�ݒ�>O�$q팍	�!>=ߩn2g?~tؿg��C�@��V^�P��e(��Z*�H-�|c�y5������&��W�`I��\��/���`��<ʾ�g���I�n�e�m��*$�N13
Ҵ�L���?^]C,jm�e(�� �F�X�Ƶ?�uQS!`��'ީ|�v�k8����� 4C,�{����Yl7���ދz!��=EH�̳Y���;}�D_$����������B�� ����'_��
M�)y�8eIE��!xN���[�n��[2z������Dp!�2���rj��ۑ��b��Fa������p%�w��˒���د-@�O=����e����N������&����>�a[	v��L.����ēk�7���ً�I���U|���z�9ؒB��N!��TF�F���*찹2���㛊��=�F���@��>eTf��j�)�����3��.��)�^�jf�!v�����v��(��Z�TzbbR^]8j�b~�4hğ�w&{����c�˨d`�4b�C1��.����7(�>��%֕��
�Ev�gb�67��t��O�J΁N^C5����� ,w�*�c�B`<��"tdwZ�S�O��WQ�`�'�86~a:��
�>�`D��8����,�Yp|s���F?K�z?rLU�C��~�&���Y���u�D�|������\�NO��+���z���8H!�������x��a��*pAj��5�˞(H�#����O�C<�Ŀ�$�ck|=�M��1��M�]H܈9�=z���4;m'Ħ�f�R���1��� F�냝sj�9ܚHRe��4��^r{C x�,�cM����ĝ����Tm���z�	��J%������:���HQ�&������Af@*D72�b��d��¶i�uv�b�� kp��h)�6!���`�k(i�R���r���^,�C��]kC��߅�s9��Y>��<���*5�)6T�M��%���ނ��^h�ً��Ʋ�M���Ǟ���\v���ԮГC��;����nո=�~W������	Z-�]��dߒ�be��z�@�?X�t-���	����pV�r�^]%�C��5ٝд>N�ʈ斁ܨ-`��n�w*klF@�ބ�C�ע�^��� ��O�_<�5:-kRy*��]%��ٟc<��xžp( !H�~J�����ޙ�ǯ��ō&4.о]N��œ��O��	��&\�?��`�N61'�i?��I.A3��F�*D�fl�4�_�͋;����4wHz~� h�"&@���M�q)+>�����h��,�lXy�ˋ|r'"1��-^�4��ٌ�N��Af��]K���}�������D���7��rbnl� ԥ����U�N��X�I���X_3�� n�\0+Tk�x���T�ΰ�d��d�����C�ғ5UH��[�´������y���J�ٙ:���5.�ЙNDҍ�G�/�!=��0�᙮G�_F�d��X{mRC�9ä�;3"�IF�<+iu�L:��ˌ�gI���������$�����$�c���П�}�>�m��P�]jsf��,�����Lɡআ�Sjd<���~η��7](�]n�ĳ�
O�S"td�Qr������j�g��	/�@b��ب�x��]˂ǰ5����p+l�Q��^'�4����py�+o�އq�Vi�-�9�P�n��Q����L�ۺJ���b�Iڤ�+����sdE¹�q���:X��Ze���ݽ��p���m6��ή��B�|κ_�.�hl+:�=�QF��y�K�����$&E�"���:���|A�o�k}K�"�`HX��0]�K2��7�J�
��YS���'����H�h
sېV�7�K���D10ݜ����;�Q���m���������^���OTlk�G���#�@prb]0�O�"�7
̤��XYz�uh���e+~�u�@�ך������iR�?Kt���oQ�)V��E8�����қ��꺟,�B}������FJƱ�)��������خ18��@���F��V��ϋ���@��$]�T#�L����[�^�ZzՆ���F�����y@_��'P��CxD"�����eS��w����ms��	�4g��2��9.��Y��vc�Z��޳���rP3$q�צOrH�+�+�Í��	O���Ś读ܵX��Xx뫏�Q�K�k�dVe��|J�l�E�R`���a�5�n��1�,���w�;4{ߗ��f��k��jj�Q�~K����_Y�w|\�b�Z�`�rڌ�3ǡ�����㫝�18� �h�[j�w�a~���m�ȟ*%F2*T���չq��o��	>��(|�	��:�VO���!�ߥo)�4+`�2+OJ6�k��BWҢ[? ���0�h��8@r��Bt�a��s���8V���N?Cx��$�y�G��`NZT��-�+� .[p�a��Y}�<��ߍ
c��"ij~dGc�W�F3����@z޽g����n�Wie�Cx�O����;��$�P�`��Tx���B#W,:7ń$x�o(�97?�U;I��ly��R�� 4<��-/l��Z���<C��cg�<��ٽASpP��X�eK�f�<(�7�W��g�z�-Ľ���\%�8ފ��Ή�-��!��C��F���B{��k-��2� �����h;��;T�}��tI�(3�1_�>�r -,@s���_4i� �t�͘�4.Ŷ�=��l��'�S��Z��:`�1��� �[�% ���'�
�0$���3�uD��~�U?d��F� � �~�Zd;�V�!K*�_cvʪ�#��?7�����/�ݨ4kl�Ҷj�������7��:h���f⛨!��g�x��'z�T�-��w�Lmج"�V�#������#�U*g)lN_֌��+�W�f���¹ϵ2�DP�eB���Zߑᜄy����k6?�� x���P�,�RKm&�ɡZ6�u
P.����u����%TWw�&) �d���xG�>J�:qy4l�����Zw2B�tB��gx|C�S��BP}�&(�;3*a�W�uyp�FP���v��`/��w(/�J"�;�P<U�\���I87e^A���uA����
�2pL4�?���>�:jȰs(ous �|��%�˳Q�Q$`��ޤ��v剠8Nr+���n��>�V����l��(�ٕ�!�Y�= ����e��A�]��Q$�����m��B�8� i!�-�{ڢ9f��v)�vH8 V<���PN\O��憃��8��WH�y[8�Hv�D���-f��4E��⤳/&���u��cj���0��ˍ&���jμ�j���zN)e�&(� $�E�����&�����#e[�޷S���������L𕞉��Ѥ_W�[w:|�knzI�ŒN�ԉ�Tǫw��A���<���tt��\�Z�
=�r3�����f���a� �[³3��>^�Ab�\(4����v��ީ�r���T��xRُj��d�o%{�Lܴ{��G�s����]`�UIbB��v�z�Ud�����>ĝ�����Y�`��g~*�6��t���DNY�>�j��ե,��E*qw�B;��]R�w��|S�����`���8Qy�:2O��`>���-<�������%p7���ҥ?�6WU#L���>�C&��<YY��u�ޜ���^�ut\S�|O�o�+���z���8�lb�^�*��S�a�ەp�a6�I��&�OH�����R���柙1$6y�|����H�p1PaMs�yܣ��ڸOQ�x��4Q[�'_�#a��RHr�f���0�)��N�T9?�H����/��^� � 3湓~���m�9��O��(�T����+�	O��%M�a��z�hpE�#�-Wgb�[��<�*�2��2X�Ϙ�1k,uQڎ�Ga Do�cp�6|�I��Q�kC�����F�M�ԙu,y���X}@�U1%�.�m�� �n�ֱ��d�s�譻� �(�Z�Wf���[�A�FM\F��5��&�Yv�N3|C�N�,C���5�~n��<�W�X�;���es�d,���Qd�grb�Iz�ȥ�z�د�^��Y��d�����Kpqh�rY"�%ovy�pg��O^qN��&��;��*�Rw�y�F� �F��rc^�}
�{7/�
J<'��:�ėRT�ʔ�ɚ���c ���C�p�i�H��:Jy�����vV��\
&/�߾�����%����O�c���\�����Y6,\i�ꅅa:\�kx�f*
ql��_s:`;��^�J4H5i� ��0"���լ��qd�<��p���3y����X4Z�˦��'�@�>%4��V��\fؙ�A���]�f��"�O��d_D��7\�P dZb�� �1���3��%�׎�I�X�2{��=kn^S0�j1���3�$�΋�*��d%^'�Ό��5�g��4J�/|��[�"��M����{:P���Z�д����
��!xæ0C;d�BOuF=�Y�d{��״U^��cZ<�-�G���&�g"�[�*���~�����_��E������Z}�Y�*�Hy�]E�X�7e�!���$O��a�\S��ͯL�~��U�r��oc �}��e'K�;7�t'sr�a��}�̥�ݿFzn�;�4�u����0��7��Х5��4ѫ���}�^"�7�%o�+s�+��P��5dVD�ϔh0Y���n�&f��
 �]��L���J��6b��D��Y�O]as_*���FHX��Z��K�Q5��M�06����	����4���_���.�ѓlf����`�F�'oy�%)��E$A"�"��:�/|I�Uo`^�K�Mg��6XȪ�0x]�28�U�%�������4"�]�yOh�E�۫	�7DbN���Dl���X���QR�m�^���>������T�Gyt#���rj�0R�=%%
�xC����Y�Gqh'G���~'g@��ų�TQ�s�D9�z�tb'�j��)�d�E��"��5�1�,>�����oJ!�F䈧�	��������1s�l@�k�A�VM�����9;绚������{L32�V$V��5�ݬ��~�.�¨�{M����>�"���}��ނr�o�<mN�	9.�!����mJ.5��𔕜cQ�����̭TY$D��Jq ن���~7O�$0�N�
��C���gC��n���p*���]�����H���E�����F�	n��Ta�Ȏ7�;O2��S�Bf��{�ӏw���~F���������\��ZvF�r�n�n���,�Ń��z�u����՛h��Pjg��<���ܨ��:��F- ��z�����u^o+J$>`��|Po�թ�VJ���|���*�4F�\2��~J&�����m�[:���L<oh{q�@��(B������Ց�����9�¶�u@x����в�G0�;:qT7-"��-�.V�aa�h}��|��
�+�"D�d���W���3��W�+�-@5�k�%�A�I�Hi�w]xtt��������P��������n,u����,j�&9�!�U�v��^`����~��<T�/�
�Z������~�E�z���A���P�`d�fJ[(�9>�r{���!��'���\���ޅs	)�-h���4k��e}�������`���}�>2�����ȃ��ʶ�}w(}�Z(γ)�,��>fX_ ��s�6��3y�����c�4�����������b�������l�[<�[hA��|C��7�
�?�Ȓ�'���_�^�U�#�� ��r~ �Y����!VK4L����v����^��ډ���pn�n��cE;l���j�1�_���	.��)���} ���8V�l�x���z�t-�5�ɇA�GKHV�_�����C2#�SG��(N�O+�����8f	�Ǚ����ƂDk��Bm`Z�-����z����k	Ϻ��xN��P� R���xfb��X��tV.����j3��}L���[W��&�d"�u�p>EJ�qԛk�9�8r��dZ2Y�t}(�gA C���c�P8p+(���*����2ӏy�\������[�ѱ�`��%Ӓ��/
�W��6<�F��<r6�e~I� e5��f�D��
�МLC��?�>�94vj#�!(*�� ӜNᰵ��Qɵ�`�w7ޟ�v@��8	| �*��1zl�lmF��Կb!ZÏ=�Q��Nʼz���+4$W3Bs�ܨ�BB� $!0�H�n�4����)��8��˶���N��[�+���r�Q�®TP���D�0
�(���(�e'x��b�<b/�uV�����hˈ||i��%����͉��)=e�q�ǜ������&6��o�[9oO��y4����	�H�Ș���+���r�N�|�z��ޒ�����y��F�t�<G�7Q�/����v��Z�=n���R�~�t�9f������%��P3֚;���^�8N�����/��v�8G��^��]fT� RT�j��[��F��`�{��>�����A�z`�b�^VQ?���L��m�>����K�U���{�g�6�zZt-�3̀c�NT$��r����,��q*�4Bb��P
w�l)S�!N�b�`[Om8l�Q:����;����6�n��N���Jp�!�'�,?A �0�L�⏤ٕ�&��Y��Gu\�2��j��I��\��~OAv3+�a�zT��8}���:��?9�.=6a$�pw�z���^��wHl�ѻ���x5�z��$q��|:�u�CI�1�z�M.��ܾa��3Eh�SE�4���'�\��R���L��-;��Lĝ)�"9zRwH��F�*��^(� �V���=���J�͙q�.T��8����	���%���Ӏ���F{��|��g���5�7~�*�M��ظQ��-�¬��u,+�س� �7��^�16���wck^�e�Hj�(�
����,ᣮS��ᰢ���0��������X���׃w?��%Y����Ę�����M7���=�����v�[�C��	azC+����n��k���g�ۓ������}��d] b[��zlp���)��Ti'��ڿ�g�Td�p�H�r��%JɄ����ӜN����L����� �$w ��F����X���D-^�qO�֪��(_<BJ):#>�R/\��Ӎ�-Q*c��k�.��p���H�>J�n��dV�!FѨ�&*"K���E���܀�O��)i�F\&ԧ����6'��i��W���Jw��ە*���l��{_��;��\��S�H�s� �K�"k{Շ׽q��o�ThR�})��G�X�������'���=�4��'�'�V�O�AS�]��h�i���D'�7�b���>b$�  Jݛ�2�Q�K�����I%��X�k��ى�n�^0����������w�f�W��d����K�#5˫���-Iª��ڧF]���j�}�:�&��������҃|��I!��b0޴��=�F�� [<�{��R�/���
俠�<a�B
�[���ٜE����� ��3x��P���l��,�:�&�k��t'����] ��H��/�(�����X�S�dG��+~��s���p
�ʖV�����:�t���r����u+I��E��
ƛ6�~���4���Y�!
̂��5cD{������y^Vw�ms��挤+�2�g�hV c���L��n�`6��׽(�L�3�Jz^9bh���. 
��.#sZ/��o#k�=YX�6�Z[���q詌���$�6�m��dz"��r���._L .���l�ZS�s�F�yV �BN�$\k"z�X:cߩ|�w_o�p#K����-�X�{�0�E=2��_� #)�:�D�Qv���c�.h�����܊7���m�uD����4A���Q��mtE����2��Af��T��1GiC#���rŎ�0^X�Z
E.�[��Y�Ah�J�i~j��@t�Գ��?w(4�@����t�?(�e�)a�E��?�=dґ���p��,H�5�G���4J|���V�$id�z9k��q�1�̌@;k�<~Vy��^:�����6���W��	�LΜ�Q�)s5;����힪�P�
�[��]�<�9j�";���8�b������m)?�	tG�>'����.�V��O��c5g���p�������x3$��ܦE����[�9Ǆ?1�������V�+��ώ�w��Z_��/��߯��4�b{&E����A' �D
n|������I�;j	��YKfh���՘����~A�!�X>(͋,'\���Z�K�r�#x��G���E���!��e}��˳h��gj���(�#�ՏhF(6��TŠK����o��*>;�l|<���p�VEq�ע�� _4aF(2!��J��L�/b�w[5Xe��g�h6,@�h�Bj)N��_��u�n=?ܖ����xU�0��%G���FXTr��a�{.Q�ha^gX}Gv\�G�
Y�b"��d�g�WQhN3����QJ@�-�E��`�$MJi��x�������;�^PgƮ�8�\nF����,�g�Z�ieN9�#9U��T�c�☃��YP�<S�/���r#Zm�v��������~�A�x[P����[�,fz��(��ț�V��]K���!�g�\[��ހw\�p�-#�żO1_���Ҝ<��{����x��2\=��{��Ȟ}��1��}R�U�9�(iz��'s�>�1, �,s�҃�US���Ƅ�CM�4dO˶���"�`��t�I�0b����];�[|��g�
So��M@��{���UU����\ "��~��g������KO�|�U�v�����/u�_��6�����vol�BCj�F5�:q�DD����}�x�/�Q�
�'��x��cz�a]-�����2��⓴V׻��f�"��H�#�q�]�N�`0��&��_�f��x����D��cB�2dZ��$���;�5Љk���XC�x	ZqP���RA</S��К\����.�^��ŏ�84�0��Wmm[&�#�d]K����>@�;q/#��:��S<�PrR2��t���g��|C���g�P�mt(�<*�F�;�y�8�|�5� x�,��`z ӭ8/�qy��<˴��ק\�NkI�'�e�H��'l�򿜫
c�YL~?/�z4��j~�o(�� /IE�h��|@Q:G`U�ޚ�v�&�8ĥ٫2g��pG��A��l����	a!�LW=v8���7Jc���$L�]�#��׽B��� �`C�c��ژN���*=)*��86��a�N��\��T���/e�쾶DDA��#�L��)� }Q��)f����PÑ�!�C�H�˃��Ko��oⰠ�j�p%=enܶX��A���2&�}��o��[TRȷ��ɆZ���DI�������ZV.��D�|���z?�$�ӯ���U���`�7[����W���P�P7�=I*�ٍ�8�q0f�>��m
�ѻ�3�>ޏ4@�^�O*��������v�+�9kuŋ�T˯=R�T}j^Hb���$���{����) ����`2*lb8k,����T���>���֦TӘ;���Egt_6Ȓ'th����PNOM�  ��M',��*g��B�$m��n�w+R�S����hl`y8���:(l	���`��	k��w��=�3p��&�B��?��R*�LĤtQ�&�+%Y��ur�ͽ�#����\�:UOܜ�+�[�z��l88��6� �.�	��a_PHpe7������k�H'��� mC�U�q$�1|�ҋ�>�1
PM�mH��3;ڮZ+�.
�4��k'�}�WS�R�ƖbR��H�]����ZA9��cH#}��%�Y^��� �� �����c�F����Y�T>������	�h%òu���^=���B��I�U���2:�*U���_�����'�Du��@ <K˞Y^�62���2��kyDv���5������,�_��NO�4��؁����cj����ڼ��a;�����X�����*�M�7��M
��xo	�\gv��2�*���3�CF�G�+�5nf�ʬ�G�(�-��Z�1�Վw"d0rVb�c�zG8����կ�h�5r�ޝ�M�p�H�rO	�%%< ����Ѕi�N�EW�Zz�^[?��w���F����ܨDn^~���1>���'U<] �:��LR
%"�r��ȼ�c�x2���fpY]�H,b�JoSP�?�/�\5 ���&%��n��� ����,O�[Dھ\a�#�1��6"&PiP�)�z�_��4nVQ*�}�l4��_�s�;��� ��H��� ��g"�0��bLq��ր���x)��=�tX�����c�'����]�47�L��A�%�Aw�z]|���r��Ex��8Db��7�P^��bM� �(�M#x��8���Z�I`��X0�S���Un
O0\�������v�A�4I]d[�@����5��y�G��%�"ڂӷ��+��~�S:h��f?���[��U����!�G0yNa�8�F�I�4k{���ת�u��8���f<���=�����q|�`��o�e ��ոC�{܏����z���xr�����>*�]�z-����ʶ8��;��	;���S���B��~_���w���l�O��8_�^=t�=�r���P�M�φ�|�5�1N��+S�Bn@�<����C5>�q�!���"��^����ቸ��?+����>�V�#Ɣ�N�U��nͺb�b����iL��J�=�bCV�iʮ�� ]sUT����瀼�nX�}zZ��C�땩�J���6�]�οi_�sM��e_���.��yl�C���F�}ty�:ٕ���$w<�"�v�:>��|�B�o��:K�9��qr2X>l
0�M�2.�U�۝��u|��@=̦�9�hM���χ7:�xH�{D�s���I�}/�Q((m/L$��ڒ���wA��T��G��J#���r U50Ȥis��
�1e�6l�Y+�h]�l��~��0@/�ǳ����_a��fr��Ht����`hL)g}�EiMu�X��K�,�
��cR�� �J�';Z�)�?���֕��k1���@֊�7��V���e�#�籫1��*L�-[Li'��L������O���M��$��^������]�4"�����0��z�e�Sm��	���W�Ŗ�5.�I��
3�cP�b�yj��x�?�#��$B�3�@�$�<������ZRE�DIy�y���f���)����d��\�ḕT���@P��
�Ewo��|���߹�nw�c
*��;� ɗI4�fC�ˤI:��"��~<-E��ݿ�F��\��ZlqMr��5��n�b��Ԍi�+0��?�h�bFj]i���R��pr�F#l&�0J.�<q��mo!�>ζ|w<�%�V@r��2ý��Lm4|��2��JǱ��j���lM[0$��h�@���B�z�tઑ0��	a��-۶_B{x:]���GI�qT�[���*�.L6�a�(}C �
��L"��"d��W�a�3��I��g@������u����[i��x�L��~Y����P"���S����n��I,,�/?���_`�9HF�Ul2佈�L'�4(K<��)/=5:  xZ�]m͇�Ի�����AWPS@O�V��f�(<!כ�Q��ة�ƾ�1Q�\��W�{���-޲��j)�[���w�,p�~%�st�2�@�6.�ȹNkʬ�N}-��8�(a��"-y>+� ^:xs�T�Вݞ��t�~W�4�����lP�}	3X\���ے�������rI���L���
����@|�ƚ>�T��UВ���^ �~��1ks�؇��Kj&ҧ�v���������� �$�����lܪ�j�$�L��z�_���sb�⬹?���x�PzR-{!j��s��}�8V�7����c���N#ׯ���&N���2s!�(3�f�CJ���g�c�XD��NBc�Zp�~�5я��k����Ix��P��R���.Te���F��.�;�� L��;G�K�W�Os&�U�d����I%�>;z&q��ʍ�>n&h˟�2��t��gI �C�L����P��([m*|j���´y!CD����^q����`5�B���p/ 5����R<C8�r�zWTIIP�e�|5�B��:��
>l�L���?ʟv/�Aj�J^(�Q� J�DtK���Q?�f`�'ޕ8�v���8�V�M�	 >����|�'l�SW��s�!��=1���JUʲ9����$��|S%�����B�U ��Z�~-����v�r)ef�8�;���a�Nm�)�F��)��G���
�����Dܿ��g���S���n�W2�2��+��\�K��H��~�w�M؛p����3��@)eIg&�s�����qe&��M�*g�[oUI�w&k�5���p���z�;ѵ��[�|���z�?������:R$�|���2��MĶ���� �r��3==$���ȝ��_f� ��rn����63鏯� ^h����P�e:�v�2������F��T�^�RJ�j9*y� ���{�0ʄW��� `M�yb��+9��}~��&3>��!�א��b%�ʦg�Cw6��Dt��g̶x�NJ;��{�����,㉂*�q]B�F���w�WkS�s͢��``��8�*b:�*!���L��������"��ϼphn��]D�?7��bVLAk��-t&�zsYj۷u�k�����wg��\��Ow��+~u�z
.8�~�R��^���:qa���p�l���x�7��H�����-_�0�)$�x�|p�9�9��1a��M����%��)���	�&4|~'0#R�zRY��xw�cՠ�-5���9�H�H�o� �^��f d���ϭ��ފ/������MT�W9ֽ��	`�r%~�Ŵ	�h��Sʴ(��.��T��-*��J�N&1��I�¢/u�,NN�
 �~M�T�6�	����\k����>����y�J;%,J��Is`�f�C�_���&j���Z��g��׹j�������=1�EH����uM�
�<U����v��D2��&�Ca����nA�Y� !�z��~�uc��I�pdK�tbQ<�z" 5�+�R��ށ��Ҵ�u;4��UEp�h*r�,�% ���!�\� �NԮ���Y��6��we5F�Ǆ��2�Ce�^y�-���;F�<x�:��R�V�Iv��cH�c�w5��~�p�HGCJ�W`�^@��DC�Q��& �6�ɳC���3���O�>�'\�蓴�UK6�/i�'��5@x�Oe��*�g�lo	�_D@n;�k-�[�Hf�G �o"��=�q,r�����sT���<�Xe{c���'3����(4r�Ō]��6Aҝ�]7{�����������D�! 7-^��F�b�-j ��9�h���A��h��I� �X�<��ρ�no�0o\��Z���ڡ�6�P��d��!�|s��5A�(�.� 1��]���V�:����I:a�b�!�E�4�y�1��#<!)��0��3��FN֯�K${�΂�%�Ӧ�z2�5{<�;��8Z��7�vSC�{����Bi�@���A��l ��\�Ћ���������]����	e� ����5���S��򯽢F~: �#�@4��gg�vp)�l�Nt��rx���+���Vx�����,2fꆀ��<ˀW6m���5V�\<��F^���#p7�\ �+�4X�]�UV�g�����*�n�4롽�&����L-�Jp=�bE%���G� 2sP���%�d�w��X��ZQ2xd�S�U���
6�m��y��.H��VC_W�.x@5l�fĩ��F�Xyu��97$�y"pW�:��|�-oo1�)K|�_���@X�|�0�u�2��7�8��r��ѹ�}��mh�����7�e #%Du��jr)xk�Qc��m�rG����w���.TX�yGJp�#���r{;�0�V9���
	>��Yf-]h�����m~ �e@�
��qUm���խ6+�t3��[k)¹�E$��s�v҇���&�*,�7�k8���h�J2��!!�Z��p��t�`1$i@q�q�2�4V/���u�>��,䯶�r��@pILұ�G�e)��f�;��͗��7�9��,�����v�/�J"�j��t��/d����m�Z�	���|��ɉ.F]��ű"ck�M���SY�^!$ݦ¦;.�ٗ������u�F�����T�2ܡU��d�{����ft�P銐m"�X��ER�����z{snr�le�9ȿ6�;�'��.f�����	J~7���w�bb\��Z綒rw�#�H��TY��{҆Ð��h�O�j���=����uF�$ދ_����\ݝ�o�|�>�q|��Ԧ�V;� ���[��4���2�VJ��n��G�>E;[+��]�h���@ޤ�B`���O��k�Ġ��C��A��ظx˛M�!�G|�̽�T�"����6.G��a��}�/�40�
O�"Յ9d3��W�{63���<
�@f�����)C��p}iQ�"xE�]�������HPݫ��n0da��,&Є�v[�59���U'������4r� �<���/؏����Z#v�(���S�J-�m��A?UP���QoQf0��(��i��lw�S(\ƙ;�lZ\�=�v�V:�-�������y�RRg�1��n��2�����k��?#�'�}�v5XD(�g���>wDf �s k��K�1��DUܹ��4����n��M,��:�P�&J��T��kߑ����'c
	.��Úܠ�L��ϔmU�7��2P� X_�~������Br�K���KW�v�I��&"�A���"C��|ݔ7l�2pj~= ��FBĺ����s�n3�������x���z�R-Vǅ�8�5���V����D�t6S#��S�gN��J�m�0��&�f���.p��iD�(�B��PZK���p�:�kmbk�=��txs~P=�R7��	�ΡF���p:.�8�{����c��f�WcR&���d�EE��Y(>6B�q�*���s�0�F�F2��^t.��g�]C���ڍPi��(8Pf*����j�y\棈����F��X`����خ/{���0�<A�8�s�z�9I��>eJ��]��ٍ
j�L�Xj?e��*��j4��([0 e���Z����Qz�:`��sސ�|vQCV8:Y��h�x�ـ����y-l>
���q!k��=��U�:���-I��|$��FU��G�BSJ� U@vؙ�xڎ��Q^�)�K�8l�	����N���Q�����-:���d�4w�Dw�U�R��9�%��Ф�Ƣ��$��������~�r�y>�z��V�����f|e$�y�U�����&G�m���[�xҷ��Tĺ��2�u��ͅ�G�6|��z54�����un|�Fߣ-,�򨺉�`�J��܊FP�=�a���(�En&f��}�͏t�G5�3'�[�*��^Cݲ�H1�� ��v��h���Y���T.#Rřj,��[Z����{�����F�rV�`h~/b.���匱A� �>v>��v�\y���P��o�gj�[6~"�t���Q3�NEI���z����",�g*]�B�
��I�wa} S�L���`��8���:	E��5����?l ̟�����p#��x��?�����L|�H��(�&���Y�)�u���@���Bŋ\?~OJ+y��ze��8�?P��^ſ��a�D�pH������H���-/)8F�A�$"�|,��4Y�1���M_ç�8�ڤ����4=�'ˬ=Mi�R��ؽ9�~ҫ�Ο���n9+�8HY�<�yV^9�_ iؓꕺ�Yv�^Jx��ATtխָ/�	�/�%9J��$�ȲT�eʏ.QC����=��(:*`a�	��3��u�ݘ��� r��Ő6�?��X�k�voǹoU��o�ԅ�,弼�D����c��ьA��r�B�Paz�T���Bj���C�m�`�`�-_�M�M4��)���p?v�.��Y��:9<C|i��!��nI�C�^z���q2�еU��df�Zb�4Dz�'�f�#�%Is�����и*��~pݨ�rEp�%ہG�\�.л��N�7x�]���ԢdQ�w��F�n)�	���ޥ8^tǑ��}���-<�,�:�j�R�:�������c�t�?}�p��HbD�Je|���!��s:���m&���$���v-V�-��O	��w\�"��g�66p�i|΅���&d�l*�q<l�ND_�,�;�����q�H!T� �1?"����WqP|A�%V�n�����X q���)'��T�t��4�W����8�1�A-s�]�������;��^��D؇�7ȋL�'�b5._ {����	������C��I֑�XfՌ��-�n�@0�������������!|d��:�w�	\B5����I����[�8���������:�J���M0� ct��rz�vڝ!dLP0��>�.äF��w���{���נ߽���^�p�<2���32+�f�-���͚���=�K�v�)��CK_��F�����4["]��B��C� �������D=�M�_S��$�8��~fn�^��۹����J���s�'�t��Ir����̑A���|]�'6��p��+��r�y�|635�oїH�X,/^c��~����+�����>V����T���Wn��ϡ���I�kLH��J�\�b�SP��~ԗ�c9sK�\��2��X'l�Z̜8??!�=J@���.6����u�9��b���_��.S� lR���D��F�Sjygω�sߺ$���"�W :��E|59uo�h�Kw��']�X��$0��2$&��눕�"�+?+�tz�h�t���70����8DX�Ӝ��s�Q��m���������^T��G�##��=r�A�0>(����
�j����yY�d�h���ߤ~{,{@�gZ�4e|�. ް�fV�t�|��V�)�E���Ԏ�q�/��Y,��
-0���,J��Г<�ug	����OH�1_u%@*��-hV�V���ɋYN��<��k�&�{ӋL��@�B���m^!A#�np����=gFj�.��*ł"Ls��i�X�J[��m��	%S���J��},.�����PBc�ia�o���.t"̙��$x���6�9��\D�jǄ��:2�/�X�����_�^�v�&����N�'�\�ӉmE-����d�]�nm���ra�zv	;�N�?I�f�y\��du�XV\~2�`�i|Oͼ,6\��Zb�rRB�Z����P���H��$F��l�h]\jS�a��k����Ȧ�"F8��� �|ݬ��ox�>̃�|��A �V6Ԣ��cҥ4���2�1�J}�׌�I�=A[&`���Hhg��@�rB�}��*B@���?�?ͻ���x��<�G��l�)�T#
=�2�.BZ�ao�g}x<TO��
�	e"��@dn��W"�^3�|,���@!�M�:k�͵2�i���x�F���y�L��P��&É������,a ��+�sV�]9���U�m&��2��	=���7�<��/s
�{�Z~J���T�����Hg?Azs#P��v�L�f�k�(����ާf���2�t�p��\,R:�qC����-T0
��C5�Qcg�-'������8�i�J2m������P#ʢ}�w�p��(:�=�y>�}� ��s;g.��q�g�%���e45�Y����3���ŔU�M����x(�G���,���巃
d���~a����J��U��E�m�� ��w~�P�!�~��w�K��էƷ|vb���J��F��HB��i`�O�dl��j��ǂ�a���Fe��.�i$@�b�)�X��xW{z��_-1�1�sVZس-�VȏY�w�Ű/��#�L�0�NeS`��k��^:�f�1���y8���>Dב�BYx9Z&ݢ��-x��Rk����i�~x:0�P.�{R�bg��(��!8�|Z!.�U���dۈi����!�W�tG&pd�30�y(�2��so���N����@��c�{��~-��I�)��mQivސ�#�f=\�$G�Ѣ���Y���}atlf�&��;]���{��R��k�*G�<�g���@e�fp��K�ox允��(��a�
-���8"p,Ś����	���S4>��50��O/RZn߱
C��z��Z=NR�E_�!�^5�g.�s�����1�:�,� �Ĉt�lw�7ZmgCDl�}��|Zu�y~�A�s<_O�tX�hjZw	�(�c�����/��AC}�������f����Q�(W0F�S�7��Y&�B����$(�ݕ���Y�FĠ Em���,���Ķ�6F�)(&�M�������T�O�c"N��<��]��5H�����v0P��G�O�h�B�|����3ԣ�ܕD��34~��1p�i�n! �`jPC��j	_��O���N�"nz�HM.��63�D�|!�(ȼ�@*N{����o����8��ݪ�6�}��AH�9g~䐧tJ1|f������'�˅㔬�]z�➨�@��狵�?"=W�GP�r�(˲ME]%{"�<b/��o.���7��l��{�Zp�O��������DB�e���7ƌ�<������n��-�_ �#*D�Q����[���<���5����~� VC�8�	8b��s���t6�j�0���9�M�5�i�i�ހu���-�̤pm�%=w/�����şq/{&����DC���q��'RU�3�R��2 X���T�����g��b�� ���R֓��kdvG����)�|R�/ɽ�&Lo�V�0��sy<��:�߬�!�Qg��>���-�Z�g}�yC���_sK�|��X��S�[�T:.��lC�a]��/�7�w`��-5P�S��_ػ�Q��&UdM�o-5�?n��;`�/ۅ}9��E/QD֍�	��#��-��#�я�2/P����TO������o��d��?�k�d-\5�6�	�\-��Y*�d�ۊl�Ԣ��]��H���Y�n�_����nVFϥu�x�s&�-���2u���V/мw�nA��Sr5�
��!�ȝyIi9
����@z5,�EC#�:�a�ov�ȃ�^���.ZY�Ź��"}�}?8���kZS��g�ufͯ�o��R�E#�"����4�b��=��|3[F��oRf�t����mhF �J�IG
h�|��!@p6����G��@N�7>seIR?���!�v&�k#p�$W�M�TQ7����ɦ�0%�_ѭ�\#�4!��!@u}
4�������>�#C0��U\-�B:�!W��`]�kTf������]��q���Y�׆��XD/���n���8��;0�r.^�Y,��܉E<)!�h��d�tq�r����/�T�	vAvU�	>ܓ�Fl<�3l���O���k������z[�7�>؏e#��P�
�os3����9�(����GM�݄�����e��֦$H����.�(��*�&����S�ţ��$e�r�*�(R79j]6ƅ�?�dg��Z\�#(W��p��G��N�L"G�mN�+?5	�D����DO��<Y�P�7YpLL����=~�R����Ɨ� ����^��n�&�jj���2��3���+*�Ch�q.׍gr �����M���2xUX�E`�8ω����'�l "�(%e�0�e4�}��Zwk�;E7�������˟p�����y��(�EEZ�n���?lу�e���AE��ZJ��W��1�מ8=N��<�B���S2 Y���F�9�%�Hc��o��5��\ƁOSf/�F��[\̧\ʴ�/���| ���?��h[l�	�T�[%a.����cl��75��v�w|h��6�{��AY�K�ª� }5��L�����f�?�ߏj���'F���f��s���șs	R�KF�Ǌ�pxC?�ކ�m�$�������D�29쩑�G]��f����qm�O�2ڡ�?|�>jGG�ZB�x���;�_�K��@T�V(uz�;G�7�L.���S���,\b!��IeT�������懎'��3��~�K7$�!2"�fyŻ���r���������������C
�P߯&��"k��������;i�M�'Wl��s��(��-�XD�2�����b�3VCU%�'��f��k����D��z�0�1
b��{�Ug�tjx�Zg�<�(ݶ�I��6��$i���-z�w��'�?!~�0��+��O�Yc�*	��-Zڡ���ܐQ��l�(�|�u��uX������ܞ��:}�fbb�j�����{��:Z*�����:���f���K��sx�o���B��WƖa2�w��+�8����d���l��p��B����>��pr�R��R�y�%�ͮ�0萍ie�R�o�_ĉ�^��Yg��b�Lh��ifK,�Y~� m�tU3�����g��\l"���X��\�$��s�gc�8���G����&�=����_x�$ѯ�R�RѲ��Ȃ�����W���pR-�_3�^V�g�<��[7��g85S,��ˏ+�t�Ñ�5��g7Ql1tp�� E�w_A���T�t�gh�������>� �/�}�A���,&)��)�g�b`Α4���#�� �A���(O��ŏ������O�m�i�,xD����Hh�9��+�����pK&�G�/�k�UB��$�G��}��� �-.�<K]e��/*~�4s��5���KP�	�,����<5�����7�������M��	�+�NZ������Za���SC�)���զ{2�y���|����L����|�?Fh��5!����%꽧������z�<3���и�J(�+{���T��H��po��Gӗd�DgJpV{�|��\n�t�����������c�ڜ��+�h�k(�[q��2(��ܢCIt[�6Y����5����_F��q+�M����C��3��nK�p>L����Z���[�h/#F�X�02�1��K����ֱ՝R\I
%�)f��cX:8}�����SIצF����T/% ;�#��`�����)��M9��fk�+���rģ�c�\�
�-.Ѹ�n����QI��>��DY��:����xJ���F}���fo���>ע�06)OYH���*ʯĳJ�0��Sf=�K�<xH�0C��na�u��8U8e��hFQE�VZ̛<{��U6����2��P&V�"A��F°�1��'m%}�m��9���sU"��b�� �d��]Dy�~���Z���	6��"V�>q�5_bn���uO	��;��tڃ�o!�O�ϫ$<�`���bI{���p��=����Sš�����v�SY6���'*�O��R�Z3uU��4{9��>a�=?O�V���d�" �u|RX�6�edxCL�J���q�>8��1�=�h����mR0]�y>ϫ:�.�	Q)��>������g?��yE�����fKK���dS�NT|  �G�#�4��7G`N��k�S�a:���~��$d�2-7bhn�}`=I��:i��VQ��������|-�E:��X{������I�V�U����CE��J��Ȍk������5�8�co?�Y�S"�����w��ţX�G�]�?�p���v�n�z��g*��z��&�ֳz�_27 ɻX-��R5�n�VS4�b�9z��07�q�i��i����@�A��)�<ޕ<�{ֱ� �A��\Z[���,��"���ٸ����Z��g���f�ۚo�s���Gc"����� �4�7l�i|�x_�G�VoT�_t��U��v� N)IIyV
U�-|a!�=���I�6�¾�7 �BI �̎,�bX~��/�#rN{$�y���#Ȼ���觘*��0��9�o{#�`�����u��~4p�����>� 0u�qU^��DHr!C%1���+kͲ���7#-����P׈��X�@�j�o��X��/9;r����Kt�������W�)�w5hn@Z�vtxr/`��6ݦ��zvC*�UG�>^P�����5Q����n�)���x��a�O��>Z�(#��6P���o��G��W9T�L��)�Ū��ɜHse����f$�T�ѽ� *��މ�h$�5�����e��Q*�7���6�I`?ʠ?��<�l�Wg^0�Q��[�L���m�k?7'D"k���������	!�y�JL���E��T��V�	�i������^!5���j,�?���u��M�g��R��p���� [�����դjx���E�Uq�����$i� ��%'��g����8Z��.;6
�n|����2��e֧{Ay(�ͩZQ��F�l�<���Ӵ�F�|��vK�譲�Y��8���!׾B4��ՕY��FօW%���Voi�:��ټ��lPS�+$�s[^��\�k�{��Ns �O�?Z"�hݓ�	mlx['q���׭-|�lI֡5�Ųv��hck���4 ����Y&~��,i��M����t��l�>�τu��D��~A�ms�`2�Sv?��>��[G�H�Ȃ�w��Ú_���߸%�&�RT7�}u�DG�OL8�m���ض�_!��0�S�WT�̀�ǒ�Qб���a�ȳm��,!�8�f���K��r0��yV������4M/��P�ې߹��1���4���~׀E��MQ�|᥏�=�Z��W�\-;G���TdW��u�;����jQ	1dv6��a����L�W?j�Q�ݣ�(��|`����<ȫ}F�]u�by
��R;�X�UQ�CH�~D3H[�����V���*�'�P}P����!��Cy��;Y�IPW�}w�*�@S�a�L����KS���0 syA��:S&I��g�QL��>2�\��l��g��YyH྾ZF�K8��=S2�6T_�cB&���� ��7i�Q`��_�bSs#���W��d��s-:-�nb1�`��ǅ�ʺ�dP�Qi1��΄���{�-�c��]7��wI���L��ۈ�FE���a'E��9�k`J-���5��L��R��Y�:E�@mb�;��M
V�B������!��4�n���
���}S&=��=��2Z\����5&�nd�S�A[����3�3��g�i�:�\�@�9�㓏̪���?���'��3��T�Z�@��"B�iu6���0Z�*<g_��f���o:�;�jѽ"�u��)�
4��"����|x�:�j�o��tȐ��2�y �)IL/5
�u�|ң}!%{*%@�,����`7�h~I#�v���MݭΚ�=#� 8$|�D���Wcp��Bn^0jR�ђ�#���#�u��Z4)���!>7�a08.�UAR!���!&���%��k�����f�϶L����=���Xi�.���5�a���n;����9*��yא��ܮF�)�BEhtc�y�r�����`�9.kv��U�h�>��ӟ��Q�8L��Q0ۃ�`�Ri�~�i�2�>��t#H� P��o���a2�9w� �w�GlM8�I!���e�"����(��n�c;*!�m��#��x���ye���*}��7~��6�b�?M�F��+���W
Q�����7�kLg�m3z�?�7�D���	3.Сhj����bJL�5��D���92f���$�^��h^��v�k9jO;2�w�O�X�Q����������^�2� ɧ&����X.�xzV�E%L�4�=��q��� g�%J'h��63��Z<#�;��O�
Tx�g2{����5ʾ��W�"��/X��R��v�3[UT�7>���D9ޱ����*T���4��J��{��J�>�#��5PaU�o����Z��9�b���+�����������eS����Ș�&�*Z~d�j���� e�y�*V�7w�6���?����0H��a��W�Ζj�6�˅L`SmL�?��D^ӑ�J��:o��|?ڵs7L�aQ���u������% ����w0�^]���dN�jh�H�=����	�ǋA�������j ¥��亵󑎘xӽ�E����FJͨFi�x� `%c�#�1����Z�ި;C���њ�@gퟮu`����7#[(��Z@𿻞�l���������X�C��T�$C��R8;e"��2EBp��МY�?/F�_�%A&���o��l1�����STb��D��[Е\H0Xm���� ���?��+h��	���[�B��Q�+��ql�5n�v �h��;�\ÊYbY��O��J5q#����HV�,}�?Y��]���({'Dj��$�'s%Ҙ=�=�;��-[=�a�����Z�ު�j�	5��/3׮����_�qv�6x��d���{�.S����7:�&�����NZ0v@g[R�B��e��}���qݵsä�H@Z����ԭ���X��b�Nu��+|�b(��8�*����x���be=uom�n��w�h����*����<�<<*���ض�h���swH|��Ɍ���3^QH��5�\��.)jX��+�����%j?�?�Q��ʖ�#�Z��M`+=�F,�� ރ�f��7�����`8�(Kف��+����w�}Б<F��I�zFL�8�5�]�P
��)&⒟�st�3�ʟ����� ���e�`J�0�� l��s䤟9C����}���}��C^� 1pI�p�Kh���Gz?�M�G^9�H�]~�3�]�~�F�����5���l���gǋ�~z
z+@�����<�F7IO+#�0X�w�h�����A�>:�w��m�V�k���N��m^����U��{5ŴX�2��N�5��",Q�dm1�2J�
?� '>��|G]t���\(�q__}�E�Gʫ��T]ĀuꬡGR�L�HS�Â�؜�H!s�4�T�Tc���!Q���;�Z["���C���!�S2f�$u�q��r�R�T��5ծZL���4����u���WྩH����7��p(Mw�����.�Ah�}��-!4�����[��b��C��Ն�˚d9�S	"�.ٯ>4�0��b������t�i��yB���g�&dj�`ⴔ�&���@��ى���J�1��F�)a!�]N�m�-9�c��w����Lλ��[�7&�"�bc��d�\��l���g[(���G���p^lHU^c
nT�Y�ڵ�=�t�Я=��~��pl�����	�a���yի��}=d9c���+G�� ��EV�uT'�AZ=/~��ܟ�{�$l��E�n"U���'i�MW�mٶ�]-h��5v$�lhɵgn�ʄ���~�i|�G��\}6�%� B�d���>��S
~�J�c$�������ys���*�Px�����mX�>4<����ˮY�I�j�J��%2M�������j�V�wrZ�v'}�QHB d��2�5����D������|<��l������6�]�~�9Y{�K�ӌ�^1�O-\m��E���@��G@�TYb@����+ 𪋞f3<�4��+�d��������S��D@��MK�y��Lu������v;ݟ�q xd�2�jǗ��Diw��8[�/~�����8������ʪ��yY֏�����1�W��wG�YJ��ԻGT��Y�t)��pP+��$��z03��4�����٥�vY��_N�%�@Qk�[��3�Kt�'���0�D��!�N���@/�%e���1�u.�$L�{�-EX�g��߽����t�7�h�v��K�R=��+KJ���S-�*����+�'9��x�2���a� �� �S�B;����le��{NГͯ�j��k9�����#g��"��E<��Y�N�
�3i�`�V�����FI�x���� �x�"Z�Ju�s�~��n�o�F�b:|��iӜ�f㺞�u0�A:B�wG�<F��5O���Ф�XtUg[\�$N���\ޮ}��.O5P7T���V��V)����R�\"�'���b-�&�ն;�a��)QGlny����ez�؋�Vw��/�)\ȸ��7�p`ϱT���h���vU�!�0�ݢo(��>TB5�4��������j��TKK;���Т��˯|j�x���Ƀ�8�YTjc��e|��?��]/���w�.��8	|X Hc<���~R�,e�?6i{��VDB�55_�l.�K��>��{p�cR���E�k��lL����Z�0��O"%x���yAYk���e;B��O|�r�E�􃆳�
x=����
?�,i��>Ҏ��K�Eۃ/
G\��mP�K����j���3S7���ʹ���h,Mu]M�{�m�$�}�q�W+�3(��Tg�fNZ,W���?:����ǝ��2�b�Z畕��k��>�	��nnJ�����Բ@�&�<k��Θ�s�|�K�N���{P��S�X�+�%��y�e�(�]������̡l8grHlѼ�:�'��vԭXŎrq�_��~ѵ��<����q:ʇԟ�]L����{N�� ��!���qn�����ٲ��t_a2t4"aW˔��a9tk�&W ��ߚ���O��ta�i3����3A{~�ͷ�;��<�,4��4��
+� ���G�;Hf��T;h��rM�&��L^�c�)V��mH̰MmX'���8G9c%����_0);E�v+�}{!�%���hi���m@�W�4�$u.�4�X̎A�+ު~�y�6ڻ!�b�G���H3�1��w.x>��&����<�<S�[:�����%đ��aA���ʖIE6���t��)��q#|թ�]}��4�u�K^Zȕ��0Wѹ�h�,x�5�C"P8����g�^v�CE\SpI���H��ʊ�YAu���H0�J\�Bɫ�ƚ�[��Ʈ����)ݺ�^Jr1��!4S�ޏ6ͱ�?Td�w/����m��b��X�������X���Ҍ�;����N��Za�����̲)���hd��P�rI�f䐒l��A�v��U26�>�"�����"_��;��zZ�0�վ$�i��>�:�#?�nP�o�@���B9�����&����`㻜�#�eq�H���i���ӽ�?*x����0��pe�|�*4nS7[�6"��?��������&BWd�
2��/�L�S�m�0�?��D<��� j�И�Z���ړ֨L( ��4���.��p�����@i��^;�����j�������U䦧~����������R `�k�BI���$x�[�E<��+�������� ��O%��G�AX��4.ZS��;�2��H���L,�F�|�U��(�kZ��(�l�Q��[���ն�v��hu����a<8�l>��%�BNB/�/CY)ƛF���%��?fTo�遊bF��S�R3Ң�[8`Z\&Į���o �-?t@Eh7u�	y:[��/�O��zl�l5���v�p�h�эm;��z��Y@�g!0�A�<5���x=����E�w']�;s
��Q�'���B�s`�%:=38����9��a���	� �x)�x���۾���������=�v*�l�[��� �.�X�Q@2:���#��,�vޞ[�����nK �~��q;,���*�H�2C
U�'l��.���c���U�,��P�QS���ӎ�C�l���f��:K��xE Z�Z����a���h|H8�fP%]#�+����uγZ6�F(-�!��R�x�jd��j�at���w�R�v_Ut^g�Zg�f��=� �>��,F-��q��t�͕�Xyg���l�Ĺ�<�٬:ATnf��<t���ʸKi������'>�/`�A�׶�)�;q��m��3��lγT�0H�tJ�d�(@���'�:1���m���,d�O�$�!6�Rd(�MNLV�s��Q_��o]c���牷4�9�)I�-o�ş>�[�_���q��v��IC��/ ��K�,�L`(|���,��x����/&=X';����dK�0�Y�*��I\II�%��f�MX��}KQ��7IZ����^����%���
����x��G��c��E �����`�FGc��m6-�`�/��3�Q�e�?�`�l&V��P#W帱;�͞�Q}'��fR<�ǁ##��
�R���2k*�eG�m=
�HZf���K��x�H������ia�i���8踻K���Z����/�p0�l�i���R`\X�м�"}��G~ߍ`��Ru�J_{�m^M`�g4����:���#�,칈���tm��}k[gIR�ly�v�.���A�@�%��t�ع�Q��]�UD��M��/���AI�tV�aK���@W/(w6���0�jC�H�v���(fP��q�rԠ�+[mφ,J����u}6�4(���M4w��/�ە��x'ch���t(�Oc/Ǣ���a<����3Pr&���k*�Cp��>3���)h�y�u��OV�/�!���`��ߩ�4�j�0d�����Y�n��WM���6���¯��.��b6{@�����W���&��U6-����H��gES�-ˌ1.�!�+U���Q�ٔ�m�]�R	�n�;�[d��L�"C�����Z����]+�"���/:��.�{t7�ڸ�X&���O������̊.D�
�e溟7̎�<V��y�k�:Te����K�D=@���C�ah~�I������
���7bV	���L�b��y7�왃s��m����S�l�/�|�d����ҘDp3�=�<��
�ť��Aj��z)Bݵ�ܗ<��gER���3����8ML�TQΗA�^�ھ��h�� _*wR\퇷��}d|�o�Ӭ��%��?�5�������v
0�&�yB)�:t�׬��Q��>�o��:Tఱg�)�yI� �{_4KOu�ʞ��S���T ��$8Y맙x�Q7�i`��R�>�|@�|���1�}5T��Pz�>[����P��Kd��𳾢٧�54yH��z��߅���?g+��ԕ$<�2�Ǫ���<K�X%���2bb0��ǳ^yŉ-f��EC׷.�刏�����l��a�s��q�^�{xE�|jQ�.��/<'@��_� ���)�0{aĤ ��5�o����(XU�h3�i娈�	�i�
�p$y�d(�#�M�wU��t�'�&�q�/�b�����i�G�:���@��7�<�T�]oN/t�44�^���dq�U�	I*e�L�<�P���͚΁���!�����3���	��N�؅��Zki`��C�0�Öf�f{<C6�'��ǂ���AD������R�hB�5����쏽�c�E��]5Foقd~��Z�J�0-+�۽��|���	��|����h�%^��J:����\���)o��*)��V���]�c	�2\�(��yq���2��f��eI~��6��~p������_P�qu�j�&��CY���RK־Lg���i:�����/��X����;�K����`����!\��%W4�f1X�}�T{�=�Ia������^�N%JTP�:S�*������)���L3���������c^��EI-8]z�V{�:CQ����w��E�q&�k���@�4w�}.2Tf9���H���z���.��X0�*����0����f��K���x��ڗG��uBak��5D�8�'h2L3�ئ�,�=Π
���Շ�N�zR���c�w��U�{�ш(�)�<�V|2���/��&S:����7([�1��	�8�H�%���R���H�id�VMu�5^�`�F�s�/��$�"c<G�퓤k�7lu��<7z�{�0�O�>xp>�bi�k�������Yo|Fg�EQv��\�*x�����
H��i�����x糴��Ed~�
��M��V*�T����b��'1J7%���'>e��ׂ,�M�.:�}�$Ȏq(�K��'3�mAn��>, �C�(ƴ����ܹ�������x��$�>� ���Y�J�iJ��m�ۃ.�ov*kc�q�,�k�%N`�9@���O��NrX݇�%��κ���:���3����UO�rQ`&��>h:�AF%���r��ĸ�~����E���HU:�)�}�]L����.�u��
\j�zT��@���R�ta�6�"
k��gCe9]&`ߍ˟��f��O'	�a*�6�y�3
�>��2�;ȯ�<��3�s�q Jgv�$�H/���k9;qb���׍o�~Lǩ���VQ��H�d�mAT���x9�0�Nh�����&ڴ]��:��d���pg@�nRm�wo���$�M�f�(]`��Z���%SR>�_4&~^&��g-���s=��H,e�)�p��t�?��V�LgB�
l��Y�;�_�1�Asz(�%@t�Tp�Ds���nQWΆ�/C�AֆH�p���GPfs6����%�oj�����c�X(@��>Lْ���J�mO��,�ϩ�C�6���(e�MŴ������1c��n�Rj����[�:S����P�W�����u�z!�33%9���3�R����*7�H�!�0w`	өp�jhϱ܎3�m�nyv|M�6�z�ө�7b�{����7+��Oh���z6fP�0�<H�&�g��T���1��^�Scn�Պ�N�Km�]�<��9M����P"<�"�&���1��Q֧]��"3i�/�|.�H�7����ɿ��0OZ�����ۛe��DT��e�P<7���<o5&��	��i��Ǣ҂ D�����!�Z���q��+��c���yV���H]�b����rZ����)3`�`�^����ȕ��u��u��ˤpL��=6+��cfn�Y��D�3��ou�Ռ�����Rş�3R�bű��I����W��Aßa� x�=R�-"�B=`d�._e�Cf�͛�ܟ.v�������0:�Ky�Ę:����QQ��>�B���COg@y��k���K|��wѩS�&�TY]�� ��zb27#��`�p[T��S�':ؚ�w�Q�-d�Zc-�ޤnI`�̖�2�h��.GQ#ߢ���ԛ�z-/���2��q���ށSǓ����X���%�Z��k_��hP5��e�L��Y�Sr�z�2�{]�9�繺Pڦm�ꅈ0�n�g��D����G&�Z#�7�T2��f�UT��;�n 1�S�����ԟ�=���![iX�ǻ~|�@Yi2ݺE���r��m��΁|��28��6ZXڹ�1�"<�����A�Z���gYvf콯o��}�$5:"�P��c�.40�Ӝv|rp̝��boQ��t��,CٖUWt����44^h[���}0�L�Oؾ5x��� Dk�����a���_|��E���i�)x����%Ҝ
5=�i<���G��ME��
��.����_Av1�G�h�T{�7�B���=���l,Ç�M�m��T$U�qU�2�i4���绺@A,ͺ��uq$���x�il�����w7�a�Q>�Q�ˇ�7J���u��hsR��W�k0�O���
�2<�����C^>�̝5Xj��%h��>!�S8�B���r>L��r��:���ں�N�Ar'pq"9~EӇ2f�[:@S�J�L�Gq��"��W�(�gzs�[$��(��o6a(��"M4�g�9��&M��X�S��O��a�$��F�3�=N�ɋ;��<?cE�?B�@� ��@���H��[�G��;^_��(�����L�xY�QV^��HB��m��ڷ��9H�{1�ҽ<����3�Xҳ����S�p�"����i�ϱS,�1���?�E� *�ѓfAl4��Z�[�凤���=�ˈ%�N�Ύ~um�ӌV�p�����<\�2֛V�b�/�Ϋ礅��VSJ�;���hDP�7-g�c�"Q����_�
(W;U���´�3�}�ٮ��p������J�B�β�/w�
_���"L�}�G�B̗vO��N �|We�����H
g�oK�h�I��d1�M�@�Wj�\�� �p��zH	1~�[� d�_	cP��ՄFžZ=D�E�1Ro�v���f�+���X��<q�����g��A������[#Ź��q��ڐ�.]��'��H&�����=������	��-r�r�S�%��fY]�F� �wr�ԕǿ�v�@a��r�+�!��0F�U��)��E������/l��0��)y��?:7@�7�mQ0�>�`�F��E�g�R6y�",�>ըKr���!�3S�ІTC@iǿ��Md�7M��`/b���S�_���:���_d���-���nFU`-�!���P��h:�t�/!��f�fF}2ӦCHR���Pn܊�@����s�3���إ����k��˼P�U͓`�-�����1е ����G�q�e�;zO��٤�B{��#�=B��m�z[�(�����8��� �B;����"T�mG�'���a��w1���s��%���� ��Gi�!*���*�AR�B.�se"ǉ��јW`b�i�%S�3�;�|�3�C�]�D�w������4X,�v'��P�3��Z�C2S�ұ��8�T$oV�)^��kP��u�[�����A{O�e"��ew������z�?����\Gxޏc�������[�"ka��%d�b����C.�IZ�n��zi\�����#\�&�ؖWD�u���^�?g�(�W�Y�v� B��9H"�Hū/�D���^�C�gUp�ȏ}�O�jrY�ԫH(�0a���‸��q>�����N�D�@j	�Z/J!ש�126*�VYy�N��J"��W�,�V��_^���3���w��$R!���Al�E;��\�_�kcdZFɱ8��59�ʬ���NlRJk��(f�ݮ�����'a�59��~��
]!����}��k��
�D����W�Q ��[�����Ob�/��e~ $��x�7f.v5 P�EW�����x�Uz���[G�"�K8��̞D������J�����H�G�z-�>�ߖ�7��+���ԯL���?��D����V��X�ơ��vb<�[��Uyo�fjy�E{�.�	�T�\��a�s��>�R�{�|D/�.���+@�"k_�ME�)(�)=�r{�H� n��͉���)�U���CZ`����ðr��y���⨰ç"U����"�'&��&Q?I/�OG���9�q�G(������ y<�Xs]���/�4�$�����}�	�Y��&�<���C������:���g�!nc	z��N�5����Z�d��#��
����.	{�['�����\am�0��1v��|��h��5����ؽ�������I��ޗ���Y�4�
J�:+x8������q��|��� H8}TJT�;W27^0�B-^���Q]3�~Ӹ��;��wGSUM/u�¦1��;O�W\��u��G��Dv��e!��7g��<Q~��n�����6�d
D�+�#����!���Ҟ���M]�}2V��z�j��b-Y�P��Z�K����nCϪ�?��!��m߳p.*(=X����5���9�	d�U�  �wI���L�R��3���ST_��;B��O�4��ݽ ZځR��跤��d��L�\�e�����O��6s��m��7Q�0�L&y]�:�.��Q�^�>Nb�|�};�g~ڂyd�	��*6K*���ىmSN��T���h�bա��7�m`����pS�n��|���ssXdN��-V�In�͆`�������jQ�?��b�$�-�81���P���,�y\=���x�����
��]��j�k��[Ť�5J�b�Z��Y�l���|����:m7@�S:��J�jSn��|Ϧ""��&�ȳY �2��K��$��� �n"��SsS̀9�=���p��c_i�@T� �@;��=�Fҿ�[A�ְɠ��v�퀰�Z��蹫�{"^�?p����Z��g{d�fN��oV���`�"�����4�4����~B3|��q�(�o�td�-�N�� �,�Ih��
Tλ|�a!�j{A�����!�7?ƵI?��+
��u���	�#`v$�J�5λ���a�
oe0�v��.� #"�`�i"mu���4�)@�Ѕ>Ӝ�0T�SU������!��A�VkU8�e.���(�Β��'0X���I����L��;q���q�3	�׬�r�Jٿ))�h����ur.�=�&��EWv�&U��@>��1�Gex�T���팹�Q�FQ��<P��,`>�=�#�Q�PĴ�o�!N�}~�9� ���Atj�e��\�e���e��3Kͽ�o*=
�H&n�	�%4e�>�*yd7�¹6G�g?iY;�s��ɶW�F��AW��O�L�p5m���?��D�F�%A\�=:Z3�w�xuL��A�Y�x��5O��ȫ��	���d�$^ G��Q-j�VM�Z���	�����D߸1����{� �s�g���t�x�EAn_�
����hIT ��%���~��>�ZX��;F)?�&�O�KA���0�k����(R�Z�����l�F���䴢TZ��E��ox��g���v�8>"p�@�JB3����oYN�IFu�H%�Y�D�Vo�5��A���cSw���ڽ[�YO\��B?��~m g�?Y�h��_	,#f[��U��U��.�l���5ы+v�b�hB5}��:�?�iY��
����5�L��]DXy�& �{< Ő�dm��oE'G��ԇ�*s�:�2��=X�Ty��O�a�i��u8�Q�]��,)������fHq��)v/��� gd�4�.�ᬻ�B:rm����đ�5v�[[U5w�\$�S���Eq`� Ç�FH�%H�$԰Y:��[޼���q�`��mqb�Ie�{[�*/���s���ifb(,o��rn�Bwͽo�^�o*Wו�?I<�-3ۚ��1M��DP-w��|D+U�/����MQ����~����)��fȋ�0�nފ% ?�3-Q
$��W�#�s"�м�+ }�,~,�&�������w���8��z���+�@:��z}sw�<I:���YF<�85�];4����)���B��sw���.�b-�� ��x׀���q`�㷒R�����ѤO�C�젡��2A�����Z�1p��
��<z_��j�8���G~� 
]/�FV4���O��I���IU
�Zt���Ք�X�F��+&'XG��w�����AAۓZ�n��B�@]�Q{m����;=� -�7.2���xaS�Ŷ��g�Tm|�2]�?%&>]�`G@-J�+2�����_�# �ʫO˗T�[gum([G5��L�Y�f�U؟4�!���|&�T2m]�p�ڦ7ŝV���P���5!,f�	7�e�r�� ���Dñ�����_���|�����z����2�6���J�^�.Zk�d4��2�[ i*�R��1�s hdFU2y���G#�L�����S��\��&"0k;Xy�5:~��^4%Q7�>}��A*9gM(by�Ҿ�( K�_��('�S}2HT
�Vn7^�1���7���`VUQ]�S�t;؋i��b��d��-,2n�	�`T����Y;�lQ'z��/���C-����
����f� �Rt�Q��*w��Q�a1u���0ևan�X"my�ڇ�90�&�^^s��YOzca�3��3}Ė��(�;�_`<E�t��7�ƙ' ����uH��	�̈́H;����.��b��L����KVd��H��m������9�$�Aw��X����������>�aÅ��Up�m��a����ʹgES2h��
B�����/�ׄA2F߀��=�+#Њ��������?����m�jzV�蝷Vcɂ����#��eW��`P���dV((;G�%h����=}��)K�QB���,�(]��]����-}'¾�f�w�'�p�B�N��5 �
%-��.[}�z�B�3tOv��N�7QW�RN��!
-mo��[��$^�d�H�����W�ԏ\�ǂ���� wT1Y}��a��d��M	���e�$Պ�6� ���1�T�v�D�,����V�B����QJ�7�ЇO���O!��&9՝���P]ɚ1[�����	&�QWЯ==8��@f�	�rx�(Si�@����Lc��=�Z/g��@#@g��rh�6�y��?&#��c̸̦�b�ڿ�^��	�P�8&��p�Z��9�P��qm��^w�=��&,7��y�#����k���~�s��th�^&��d�G�8�`�WT)���)!{�qs�.��	kŤ�ㄣ�MO��������7�yI/
��q�T(�;	���3M��7u�J�'���E1R���?�P6�5�ƋY�4�5�UoK#'s0�,ۛ�y�=P�����\�f��4X�;�a����j�w@����{���FvZ&ӚϷR[�'� ����%��\�shX ҋӿ�ں�_R�?�~�Iډ`���-�3�[� ������e�6&�zC�����Bo#:�͵���z����1A�)ݏ�qX�oB/P{���T�<Z��U$��P�| }�m�5� �%i���*��0��:nA��-.�P��Br����WԊ�ix\��	�d�\B�8��a��U8qMlK�m�H�lj)~� ��J��i�$о������bvR��*��QdW����cb�w�oݘn�wZ͘��պ*$�@��Y<�;C�G� �~�1��wU|q	���]���YQ�Wn��A�`��)t��Up�]���WF�?6nQ�{���#�2ᢽe}+�C ,5��S_�r/B�&DNk��8q�����+FD��*W}@�<������F��8^�](�ʏ")�Hi��hs䋂������d���eW�[ju`�+���bͤ�?Cj���Te�O�h�M�"�1��gpL�й�z��G�fj����~&i]\�F#C�n�\	����L�2��
걹�fƔ�F�y�+��XT��wE�/�0A5K��L��F��H.��8mm�v�~�A�mԢ�$��2�s���b��<���+Em�2�+�?\��>J�G�|�X����$_��������T���uZ�G��bL뵙3s9���!�i�)��Tf�l��g���mx�^M\V�!��fY�n�� r�����H��q������#���ߏ0?�h����p��&��c�M��'7^��SK����ߜ-�:1�����jb�I�C5�o��4���0U��q���~e��x�0g�bbf���5^tJf��J��`ݖJ~��s����T@=�[� k�J,[��%�a�9iN�V-���
Jw/��7��+D�[�!ڒ��c)}dd8�^ݷ�#�(���GJ�>pΔ���czr�����b�t�=I��~SO�pܰ��m)C|}nab���S
�.]=�e._}��O)c� *��ʱ4/�ͯ��o{q��$��*EC���k
�i*~�����9^�n�-$^U�%^v�:I��D�~%
F߷��̙06n0<Ðd�B�
�2S:�n�~a[[c�$��|�i�ta�E�]y���k��P�VN}��w�D�����e�;����+�jUɁ�h�02��F�'�!PMjY��w��v�3��̾ ���2ms�>kDE'��S�3����_�anv��A�����@��Y�B9<��u:�1*����������vG��^Y�\h� Tl+�������3�j�4���6B�tn��icu��@-mb�o�3���v�%����D@�u�AN��R@#�ev��Ҟ671�ޓ� ��{�]�ߓ!��lLߙ+��;s�� `h2|h��y���	��e2K�����j�Ĵ��x�g�9�~�xn/E�xC��s���t_��qF����e��N�|ïo;�G��COf��]�X�7��c�+3�N��3�cM`��06��Y�I��%��= uN��tC^�x��u�{��Q{�J͢�):Xe-���O��"�wuљ:�O�G�iFPvO�f�� �y4��g��� ʳh��\��}�)O�'T>��d�a�^)v���(\��q����>�8͂�ɶ*���)-Dn�����"+z$S�݅��I������=Ȕ[�瓢9LD�����������U���!t�~��=,q�*�5?������z�j��\K��ݩ�d����X]����X���J8?��j?��/3�|�������9>c�Tbӷ
$k�d�	Xu�H��ґ�R8l�[j�i��V �M5��u�	9�F��F��Kc.��`g�k�yHl�`�9���,0��O~��x�R���k�q,�� ��[?�|9�vE�-���x7�Kw!
�i�>]�jA۳��KE���
� `���F2'FQ��g�Һ��7�N�z�=>H,),&M1�tK�$��q�찏�����l��5,3e�ћhľq��Ł�>�����GG(>J�)��\!J�������V��C泌�8t-s �2�]�`>_��#����ߦ��H��TY
l�����y&�f��uX�B��k�,b�C��'3�y%�~f0�#E��.G����t�q�s
�L�~S{�|�|�t�.3�+���@z��_(�وo��)C\�{�[� �0j��uv�/�U\���0��^��(,[hwy$H���r�í-0UZam�'l�&W]�/w.g�?ZU�N,G.���R�a�+<E�]ϙ�/�JJ4]��_t���Ԗ	��Gʬ#B<_��Iy����A�������'k�	@G�ND��);Z�t��q4��+�ƈ�{�����I�����v���7,��B*"h��_5K����Q1��k��=[�:��ĵ��BuJR��+~'t�\�$�����C�K�9��b2��J������B\h��R����{g#�λ���-钫�(V�\qVc�2+��I���6��7��X!_��Tq�����C�r��G�UK{��LǙ���I8��9</�2X�d���K4
a���z�6��\p��%��pf~ϘXd6�}�_�ꝄI��u�%�	��lG%�{`��Mh��28�OX�������βUC���M�clѩ4%�-�(�������?8�-�#ݼg��}��:�d˸_��O\㫖��T�32ut�G+�L��j����&=�!=S��l�TY|u��d����dh	�8�1_�!l��f��󻫊r��U�����U���6�=��K�<�)�B�Mu��^'�R�>��QM��\Q[hխ�IK�����-�4�l�7�eҫb`E�CON��P�b�n֬������<�p�0��b@�O
�t�z-��R��<}ݰ8-�����������@W��z9J��n���ra���Ns��-C��䮿wI轉�h����k[���ڬ��c���d�Oi8���=E�(Y>G�Rvp�����c�Qb�c餵<<t9��=��~���p�+�����a����ë��?=.[���u]}gsZ}����ʋ��/���i"�{Dl$���E]�0"t��iJϨ�^.�'dвF�$8~��?�ᶔܕ���~�)��lS�&~�6�t�j��B)�ˌԤ��G~;�kc�_א�{���.�S�y����
�P���(��ܑ���W��f]��5����j��g�i�2��X`�v�{b�j��w�ov�_�|� n\�2Ga�0�D����;���Q�y9��߈��5�ѧ
��YE(�Ӎ��O�1D&���On+�^oGʌcY,� ���+j�f�?�3H4��c��ˎ�v��]��.@f��у73'uS�w����DZD5���N�;@�U�e�o�����1y[f���{i9�]���s���U{c�L�h��Қr�\�Ȏ�D�eK@+��G(��\�!��9��x�.���%\�=���U<��m��'Kse~�RN�:y�2���e��v��x�rh���s�ŗ�N�3�V�`!Yx�Q��^��I�7��0^ ��Nux����u#�q�tm��$�DͼT�:���_=����0^�uf��:8e�G�2�FjZ2O��SК��s�g�1�Z����\��}�qOk��T�I��>��x�@)��3�pq(�(,˓�b�Z�չS��"�^��8�fWuZ<�g#��f���o��q�ɳ"�vX�m�_4z��&@�|<kJ��/�o���t����Tu 5ȕI�$
���|��u!i�+�e�p�|�ɳ�7��I�=���W��x�*a�#���$����/X���V�n����0.�n��#K#�ۨ,6u���4W=r�x�>{:�0� U�}�T!j����-Ik�Gw�þ��F���z�@�:������X��Ċq؍�CA���/;���{�� ��T���Zj)��{hU�m�=��r֞ ��_�}eVv�;�U?��>e�,��ϱ�����ʋ��C�'���By��v��>aD4#�-�Pl!o\���%�~9�Z�;���m��Jr�/`1e^�3�u��ۍ��Q�q*�l��Gu�<l�ӽP�e���*�.�7B-@6嗢?�-��GBWN��u
��{-�L+0mw�8?~�|DI����/�嵢ۘ�� �LU�X��fޛ:��}b\�pؾhC��'^�t��/4j����;����˅�T�j��ݹ�����vѩ �&��U�nx���E��x��ͳ��? + d%���������$Z �f;�DL��Y ����y,H��ç¸(�-�ZXd�fL�l���N�&�J��Ճ��E�E��`�8�O��pB���\��Y���F�e%,��n�oP���wJZ�j��S���ot[�v�\3�!�%��9� ��l?cuhd��	�r�[nD��</��4=�l0��5y�v��sh�W�:�<����w�!�>���/f�T�>JJ����J̞��sN�O%���kVH����z_�*�$�i��Ӳ"�X�%w����a��9�a�Q$��%�7Or$W���:n9u�$�4��r����A�~-Q������:��ԟp�cL�ۢ�O,t���ϵ}�ӇM�x��َ>���a��"��Y�z��9�>�&3?2�����_�O�ya}�ܦ,�k3o��)'�;�2<��c�f�� ���c/HB���m#:;D���m�NL��v?`)V�]H��Am��uڝ��9�%�ᱝ��J\"!�g�-���� �yp�tt�.9����i�S�t��W5\:=��[~�w+BA��M���{���Ǌ'���1��t;�d�0m\��V%����U�"�9sl��	��X���0�+�WV��w;�lh*�Ňݳ��U�Q�k�E_(�����j&�"�i}��s�&=�YD���B�!���&#
�'^�H}+}��Br��O�NF��WKŸؘ��
͵>oq������t�d�3��fWP�\^.h�� 4�.1����<idY3�	��:��`�*��������18W�vA�F�)���7[>T��8��<�=�װ��'�����w��Wt��*��|]i���6��<&�,��:=������	\��r;�S	���L�w��j�������y��s�@B�r����c����#'̪�Fw���1�yԔĴ�'���P1����bZLc���C�q6^'�=i�:&��l�3h���'�s�kKo��-Fs7��t;)&0|8��8�×W�
�(��!�Vs��R��q��D�[�CJKM︊��3�F"\�����qR�+�ۋ��9d�M�bS��R�i '>���wbڳ��?2�r��ː�� 4f��U
6'�",{�sy<���1�^����4��1�F_Ƙ,��I�G=R�C��F1��:z�R��#۠{lX4ު�@�ܡ}c�3֬"͌���Lڬ$?,^Ӛ�CBR�p�����鸧�Y�����+0~
�����i3���v��U�} "�7mZJ�:n��`����]��K�!J�QKW�{V��g_�I.�)���'wd�$O^SÙ�4l�����	_h�odw)d��~��+9մ��^��lW��H������˯zƂϦ'��9�+�~&��R�[��eFfK�Ɔ-��b;���t��d� �)�����gJ��L��e;��$ ��(�.��� �ӈE4������zr��[�
=�H�	�i�<�������
�:�2��/�Y�g�a�]Π�����⪦�G��j�;y��Ǖ�k}�vQ*�	�|�]iB.�?\L:��M���0P���{��;��+i�"0�x�yR��:��T�$�Q��*>ËF�؍�gӋ	yY}f���.K_]�ʮ��Sù�TO�4������7���`��9S�)ؑ^�(��d�q�-Ḱn���`|e�i\��Q�ֺ�l��y]�-ƃ��Y��ȱP�N��j�J����W�{Rj����?k����5�����Y���1R�]j�~n�l���񿦦��D�IWn������Ꭸ|&n
��+2�q�lђ��[�n�O�SȧN�.��d���3�~i��a�� �@P�@��̛���PER�EL��L8�U,:Zo�E��_w"~9Z�q����Z)�g���f#Iso˓��j"�$��4�A��O�|�W�ۭ=oh�tyJ���" ��I]W�
�|#�!��F�����y���� 7��DI4�����.��W��#��$-������H����0�D��9	#��[�~@�u�v\4!a��g[>h��0��U�o��X�\!��c����k�����3�����g�_ל�,X:ʊ~�<�R�Ӝ2;HR�oq���!���_��)���h�e��J�r���J�l����vW�yU�	->re���p9�I������=	T������㣓>n�3#9�P�OAoIᘲ��9�]8��o0Z�Zf��q�e��k����h��~��*���]'��I9J�j��e�#�*���7ϸ�6�?ްw��)v��fW�e9�K,�h�+L��tm��?KD��ϑ�.�В�(�]�!L�o�.K^�h����}�����bp^�u�v�j�"#��]�	�aw������&���c� �<�<����>x+��E�
�%>�� )��_ ��%��s�{��S��Z#�;����̒�lV�&�@����I(g�cZe\
�FNl�.�;�����հ%U��R%�|��m8����5��BȠ���0lY#��F�5%��B��qo�\���s��WITS���ҜČ[r~�\��s�T�iJ� �F?�R�h���	�[;���Mw�A)'l�%�5��vo]Fhw�=�g.���!rY�,,�@ꇣ;��5��j������Ւ�;���4�'�!M�|{�s}�gՊ=-���;��uaqޠV�<���/�a�����ŮۥA��5�v�I�U�s�)�.j�*�$O:�y��KݮĦ�v��[�m�Q;ק�y4�8ݙq5����~�H��m�T���˝��Ql�Цm^��$b^�z��6C*�.�Lh����b�b\o��n�� wB���s�*����0<��	�/ֹ�f�ʥl+wgf�|Y�I���A���Q�U��fӄH�k)\��=���E�-�?�?�>Q�A��[#۲����+�]V,m*�ۇ��Z��oS(�8�X�����+.ƻ���,}(.�<����ZF�r�8F>�]d��w�)�o���'s�"t���(k�Ln��M��C��`��1�M���J�����CRĲ��t�vl�PrQ�ox1�mAp4����Zz����[���~:�]DP�F٧V��D�t��$	���
Ҟ�N����F�u+{,X<��w-����A�j��>��u���T|���|m��fW�U�d�|�2$���x��z��ۼ#mq+�2���?D�>2��G�ڼ�@�`�r͝_��O���)�T���uB�G���L�Q��#��n!�s��J�Tg �T��O��Ų<��F���~�!���fA���`�rnN\�wB��Y�L��0�����K/�w���08�r�F���F�M�h�W�;a��n�w-ygQ��|D���Ibn-^C8,�޲ޚ�k���	!�������0OZ�bN���@t2L#���-�~G�s����m�=�@%�L���J�6\���ay��N��-��z� �w�z�����$[鿁�z�/c��d &�Fa�lj4	:2~��ֻ5q�>���0<�U��x���W!��ʊ)P�k=�e�qG�-Ϻ��zqd���X�ꊱ:V�����Й;Y�I他X�sה��2�%)ꁢh��h�},Qr������o<vʍ�U>���/C0�< d�Մ���E�g������ؐ>�f�#̗�P��o��B�e�h9����{�L����M�3�o
e�~֦M������p�*%���0�	�|��:�e��*��7���6/�:?Q`g�[�[��) W����||���Lk�m�>?�}+D����
��% �K��|i�\�v������lg*�+Ծ���ģ`BW�д�P#2��L�υ�ඇ���v]��A��B�1&��l�$8=�5�	�	���r��iS�~����몵#]���Ƕ�5����@P��rq	�ע�҄YO�#���/��m��T��?�f\P��^�?�Z_��ٸkq1�^@z=��l&5�Շ�V��f���<��k4���'8=s`c�tQ,&�- �=8>�Wkx���*!$��s�f���jŭ@���*�M�����Z[�/"�"�.ӏ�q�^��DXw�½jM3�����*�(_c'gj��.[��?���~�;�³/4OR�U��'<��,�W�y�v��:M=T��C�4�4��
.���C�`���f�1\s}F�;$�#�qRw#��}h�瓀����s�䇠�J�����l��s�hJ`qǏ-��N�/��]F|��n����Ͽ�z�u���Bx�t#c���Mz��懥�����4��q�}�[B8f�C��T�C��8��-��O؏E���>��D+ +�	iʙ*�/ќX�"Ao�o.��/����1W��ri����?�;�d�PɊC��D������֮i�O'��P0ݩ���C�Z��_y���aT����^��eP�Lu��ⵑ�A؜>�^�s~��÷�Ġ��߂���T�J�x;�Ѫè:<��R[�c	� %�y��� O���+Ipd�HhѷoG���=@�!S�䷚W��F��;�m�����'���T�������8>�)��Wd�M�'	�lԉ��s*���
�=��{�\�d�a>'G�p��w����K����t*�h�O��`�v�����v8�6�r.�ûXS:֒g��0���:ve��[�7�^������Ѕ	q"�hÉ�HŠ}����r�i��u��.���p��b�F����G*�6�i̝��bjs o�nƽwϜY����*�~s���<����C����D���w��T|��ɱÆQ�Q��L:1�����)I��.��r�^��A��p��l׍�������ds�%���7�ۑ�`���-8��죪��\%��-��_#n��z�&D�`�>B�~�#��Ƶ�y�z�Їd���[� ����Bw�bc>T����e��O�3������Y3����� J66i�%�*�;@�.sAN�.26���]���W˸i����к�;B;Ⱥ�wEC"��DM}&��!��Mh��'ς�P����CS�Ⱦ�y��qzT̄>�D�^�3�P�!�u����42�A7M��Z>���	��m�h�{���_����x���4,[��c�[����?% �)�=ߑ��#�I[�P�*��ѶU��si&���K�����ul�|^6i���ѕ $Sp����"��z�k����}"^R��C��Kp%o��9(��UgY`gZ����0x$��y�d�#�7-q�
1��|ɰ�V�JN?ө}��nӦ�������J�%�WGV�ܝ_��/�ȭ+���w��`$�yFø�l�э|�_'��d$u�>���zIO9��}��lV%r'-��d�Z�j�/�-'*/9��?~E�4Q����
�%���m3��̫�7X�RV%��E ν��t�:&����{�e�*$m���L7.��/ ��SE%˲���4})z�I/[� ��h��ꀿ�ad��uf�SHg~zi�kߛ�ڌs��+K܉�닛�Hfǀ��̜Ӛ�m�X;����Sb�:��yۑ]f���E�<
.=�'��"0���_槡Vs ���tq�{N�*| �.)5R��@��P_^��e��)��{7�� *\�Ŋ���yU�چ���j�I������yZlz����c7jU����Vh'bQ9&R�/�ٰuT�DZoG��R��"y�MP<;�S]���/J�s4���UK��k��	�����<Ur(��/�W�ح�_^��| ��v	��RNz]��3�Z�k2��V�ƛ���{R`Ǩ��y��!�lN(��x:��h�!O5A���Ϳ����m��52��`�\�(�:�
��j�JH�y+45���R�-
5�9v�����>r���J�l���[�\����{J��p�1�{��������3(�	q�S2=*Ȥ���I�e6y>��>�I�_f�"qK
�����C��\���pK��Y�j�^4��	&�;��ra�шn=Ɍ��M.�~#&���� ��2�f7�~`��8�Nni�SS��ɀ@�Ɵ�K���ia^s���
@�3WF��mk�b�6֗Hȫ�3�'��Z�P=�5]"���,"��k�Z{AugB��f�S�o��,�mq�"E���;I4��6�e��|[�t��joz7�t˃���#$ �jIo��
;2|��!hd/���/��h��7f;�IF?�e�-N�)��#�%�$5��|\6�I��͒	���0M����#�����uA0V4����ͩ>���0�U���j��!)힊��Rk|&��"m"nhϙe<�9�>׮��XlmR����$16�|�;Xԇ䚅Xڕq�3��ܱ+�)IȬhԥ����r�����|�<viߓU���>��n$�[)��Ա����&A��!���5mo> ��#H�P�o�o�=E�D�9�\.�k%o+�ݬ�����De�嫦L�0���{�Pw�*ć ��T���h�<�re�'�* ��7a	#6�	�?�m�ڈG�KdW����A���P`LJ�@mv�Z?]��Dcl�l��d:�)�_jLt��� ��zx��<\��
z���<d^6��N1j����4��[����kR,�8�|׵a� ��͡����wx}&aE�L��E���O&Q Jg�%��ƒ��b�)Z�� ;m�=�-<$�����"�J(���(�cZ�Q�����l�Ф�Ĵ�i|#Ղf����3��ɡ��)�8e><�G1�B��{+Y���F���%�e���o�hR����Ʃ�"S>�:�ni[���\���W�V�;# 6J?@�h���	�h�[M�
���b���|l���5�qXv�	oh	�{�97���DY����C���5�I��D�@Q��M��(����� 'n�Ԏ�Xs�����=�K� C� a'Z�����|��Dr^�1X�Y�V����	Q@vv� �'<�; �.�dໝ"�:�J��]���0�v*ǟ[|	��c_x�: ���Mqd��\�H�:b��o��dݝ&`ޣDm�8PA�U�cbpe����"*v
V����AbmxoW5Ln��HwTp5����*�G��f��<��ہ���t��wy�|��5�v����6Q�A��ԍ���s).@�Ol����:��Cj?��Q�I�>O�#m]P�w��+���,o�j�m+��,�P� �5��g8�u=٫��+@O��H��}�C�<p�����F�v�8���]���ʉ�))M����s�����G�I_:��nL�P�U)*`��w��F���v��	w�C�,4�g�H1��b�f��Z91Z�*p��� Mz�~��1�T�r��~ ��]��'F�\��(MʹVi?�0�$��=�
��&�`�ՔU��F!m+Mn�XN^qw����HA�dg��sMf�U��x�.mȊۮ�@U���(��;2Kb�߁!��'ێ�,m���2�X�?֝>-�G��pȒɗ�s�_�0C�ko�6��TG� uqG�
LH������x!ݷD�c�T����&p��a��ܙ�؂��:$!�f���[c�r@����1A���o�D,������s����}A��D����i
�UPMa��vg�M{,�A�g�w-K o�P�&�b �C�	>��*��z�=b��X~"��oH0��^b�lb��e�tDJ{9gZ��t}�Pd4��e�>sqqf@�����JN)P�0ʀaKm�N=�-���V0w�C�1x��e��[{nh�L�c#�Ddr#����݀F(���G���pH�9�%ct��]��#t�s=C�~�pV��'��v6�a�ٹ�c3˫��9=����>\����<��9��+Ա/����	�A{���$V�|E��!�����i������ǓE��i $�9��-T�4��1�~�w��q�b��M�6�c��
��Bɴ��,t�̨V�~ۢkcN[ؐv멯�.]ؿ*�y���eJP"��Ȟ��1L����=�jص5��sI�jO��ng�P5����V~-��)X2��������w�<�Y��m�!�2�c?�j�>O�#Gr�lȝ�	�o�s_r���"��t�T23�u_��Gg96LS���Ttؑ�t!D���!�T��@�qT�E�����CC���!7�%fW��Fa�r�^C�4V���y8��'s��z�����T��,^���V��	R�`��M���z��x�Avd�Rj�-���j���bk~;C����7T��wӧ(������Sx0��bK�Ǻ��to���?q��^oݛ�c�0v �I����@��S�E�J�\P�o�a��mN���-�x�w��<�\���i�[f�ڗo^cΈd}�[Cf����($'DG�>p3��kcS����G�~t��=nt%~_�pA���r>!31a�k���Q��=z=�e�$�� �ha<����*�}ʖ�]/s��4+{6�$A/EHtjt�^i[Ѩb�r��㚲3��$�#�*��}'�<�~
��<ڬ��s63�����B����\�̳T�~Fb�cQ��18�9:�ت�y��N��YP-͇3�G������9��*��ؠm��~�j�|*ɭ��2�,��R�FN�jt�wGv���fU� _�2R�	��@9Djz'����pE��dP��܄��oѲJ,su+YJp�职��1/�2qT��fJ�lmG5\#Y�Y�����+�؂� �S3Qr�4Z湻��������p�;�@��z���3r�㸻eS��C�Dŉ���+N�Z�@p'e{r�C�y1$�,�叛{{���҈����Ĭ�@9�症�hw��}=x�3Jx��GKkm��A�(�,5l��7�9�Wx�$���铂8z�a8t����r�-e)_cN�j���[�l����d�6]W��:iĜp�YN��3J�`�R�ބ���FI�t�C0 �}+�Y[a���u� ,��������ͧ��:���
���Н�@`u1˓:c�G&�}FUz�O9���E�g<O
%]�-��\�,}�b�O�7�T��D�I"��ܶZ�B�7`Q,���t?���Qd�;ad4��U��'zm,�y�w~��C����HZG4z^���ƚ��YM���g��TS�g�FX�ӼL�R���ۢ����' ��Ps�Z\�tڭ�n���є��^7��N`jD-�j��?����o��Eu�Sz�����B��#�P��9�Izs�}�>���ud�aE�vNMBQ�"�|{mTm��}��w��M5q�VÔ�v&��{� dȠi#��*s������A(].�(=xX��0W6�8i5�j5^;	�	�C|H�D�����K�
C���+'i�P�
P���YC�R��X`���&T�w�G>^R�P�c/u�7�RaA�x�4���<�WI��=���U�y�����fx4�I���u�r�k[0�\w��%:U4��s���C1I5��DX������������6���<Uu�r^���   -  5  �     �+  7  �?  bJ  �U  .\  �b  �h  *o  nu  �{  �  7�  w�  ��  ��  `�  ��  �  '�  i�  ��  ��  N�  ��  �  ��  ��  6�  x�  ��  � >
 �  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�?����~��璹W�䑰L|�� *�S�<�g�Q9 \��!+F!F����SřL�<!���d hxc�ϖ(��h�K��<Y&�7f�O���R'&�����X�{s<e��650B�	�S�QA���1 �\ ���-E�O��>YM>�&��8�P�S#%W�{x�Yz�<��N܀�1�j��r�Q��bN`�G{��Ox�I%������U��$@M�0�OH�����n�@>]�t��"�08pa��1 ����9D��pH��d}�t�C�&>��k@"�Ą^�'�1O��;�f�}�ZC�"n�h���B؟��	�z����h[.�h�6Z�]����O��(��|Bd�	�ܕs�m�0.xx��� \"��O�#~�`ʻh�&�öO�={�N9VnEv�<��H�-�ʉ��^b�8#d��u�<��L�0~6�k%��sT��%�y��d2��[4�Q�s� 8\Ȣ,�fo�(`���T ��> N,:4'�ц4��}����A"7�T5F���]��^�N���
�m�>i�c��|�n���Ϧ��Y�<���!z'`H�bj$h�`%}R�'���2���H��``��]�z{$���� ��i���{���%�5x���"O�T)u޳Q�ʝs�O>p������'[�'�^�I&�0*&�ӗ˹C�"	;	�'Ih}q�&ԃ�D��✽CU����d���O���q���RE�ȉ��	T!U H0r��';��Kѫ�|ˬ���3S<� ���V<��'�����O��:cΑ�f�yB�j�\�*��x�
�O�c�b?��Q�16R�ː	�/ZA��Sa�v�����|&�&
��8S��1�n�d(���'��zQm�*-��c� ~�lp�ի�y��'��X�`��- �:W��$2���'�E��'x>�w�&���p`@�kv$sK:�O�7'?q��5k����  B���s�Q1w�jY��H�)#ɧ����CB����
��~�̵Zc!F��hO������E#��
 cۊ;��q:��['x��	�U��	�q��E)eeE���cP�ɗ?�@�'�Q��'��H����dŨa����lO�0?q+O���į@$���cJ[�K�́ʡ"OXYQ�*�"1 RqU	��p� x����Z>Ғ��2k�yyR,�$ �q�
7D��C��G}1.\�lz��ђ�E�O:�=E��ܤ�A�y���a�܂S��B�ɞ-��X��z�(2f��7nn���Ķ<�Ot�"��K��Y�$�L����"O�@���S�F�� ��E=!���"O����	>�������)HK*$� "O���]�@� �
P��
p����I'���'e^�S�`�ƮC�C�Ɍ�4��G�2�Ĭ��G�_>�C�	�@��IҍB���d����-C���=�
ç_���8���=1.9��L�7p�-�ȓ�����L��I�Q���A�U�ȓ<��JQ�ϝK�4������*�ȓdشP���Q-�A#��>'��E��_�(���E���`��7z.����I����*r=ĬkW�@f�6�$[ PC䉑/�H��p�� X9)GNp�Ң=	W�S���|;�l_	B�XրL�.�B�ɲ�� 	��̞`�D���4X)�C䉅<�(�y5��P2��g�G�xィ?��4po��?�Y�gʥ���@��KB�0��4D�L �+��Y�aO��K|��8�I�<�'=Q?� +�<X�ܨ�SY�	̸Ǧ4D��8���p�xhv�9O� ����.LO:�(6'z�>E	p�]+��
�"V=�y��E�\FP�j� �!ehA;����y��%��<N�>vDR���1��x�jW'N�j�@$lӌV�x�-Q4
�!��X~��0r��*(�Q��Q�!�d��%�,�Q�H�0H<�I1I��}N�]�ȓc�T��'��4��ai�-��0
Շȓk�sA
@8	3�gb_��Y�� ������5�����8L�	��	x�N�pG��a� ���'��Đ�����V>��]� ��u9d��GL/���d?ц�	>��/t��YӨA$Iň!�f7*�˓�hOQ>e���#:�HV�b���Ta�X�<�{߾���^4�^�A7d�'<�	��Iy��|b8OTb��xR�4Jԑ@'�Y�zE
pF]@?�瓡y�C��,4�f�m�()d���IrX����̭3] 3c�w�q
��"D�H�P��_Bx�k���82���4�A,�������N&1���rB�Wk�	*t_�pF{��W�@�	�� �/�2��Ee\.>�I\��� zd#D��.?NV����K�ri�1�|�iT��>ap�
JG(UIӑ?����&D��y""�-r>�tH����_��A�/�<���4�Lc��ȤN��H�X�IO�2.�iAD�5<OL#<)���79)����/ˠb��PQg�'I��Fyʟ<|�/H��1ȳ)��0�G�'����7� !����%U��1��\0!w�D �IX8��Yua*e5�T�����fHZ��+?����~�>%>q�)�F1I m�}an	S�^�9@�P������;����S	9
��!�g/3#B��%�S�O�6]��KN�'*IA���k7��	�[j�	�=����b���b�aBؑ�ȓyY��hƂ-4�d��iG�RNT�>��yR�I{�p {�i�fg�P��I +�(H	��ITX�t�� ��O�*(k�됑(�L��� <�<A�O,7�;�ɛ�}gk̇^.��e$�
qa���Ɠj�hyH�ȋ(i������%WK���>���8�Æ,�NU�ԫv��yEV���M�j.��:�.�<h�@�2AΥ|�L=��hO�>�X�_4h]c��.?T�ݪ��!�I���=��"��E�%
��2X���'�"�'��y����[�ٿ5|��kF���y���/N$u00�Xd��y��'���,�O,=B��P8`ݨ(�ˆ�5�E�g�'���� ��O�!6 ͈�F�I^��"D�4A� 9���j�剮7�e�eh D���bd�E���g	�B�ͻq)>D���Y�b�(�r�ɾ�uy��;D�`�d�\�0Θ�
b
�4r!IAC4D�(z'�LV��pӄ��*6�R�0Ҩ,D�t9blޑ`����Q��n�R�G*D�3�mӯ$��ea"c�&n���$)D�r�K�W�v	���Z��� �&D�X��P��y�AN�	4?��$�/D� ɦ`�;�p���bŊ<QԤ���/D��H�<$���P,à	�hc��-D�$�VJ<e_�%���"�R؊��!D�[�iަC����	z$�j��>D�\�E+h@�<���8.��ѫC=D� 2g��E��m��o�F����-D�X�Ц܆
�����9>���66D�4�G��JHɳ(�%k|�t0�!D��ɛ��&A0���Z6� �#j*D��s"�/p.�KO� ߺ��%c-D�P��"��<G(����M�g���EE-D�T���u*�%R���>���P�f=D��ڂF�"8������>+_Θ�(D�tU��&/�-���/8x�ܹD&D��p���;.=�RF�{�L�u�$D���M�~I�����*�`'� D�� �O]4��]YpJ�W�h]ȧ=D�����ߖ(��AP!��H�z�l6D� $@�	=��=�P���n/mkw�4D���!��)L���CJ��T��\ @l4D�P8E�?h��Zw��#� ��Tg2D�PP�B�t$2��!�Ο�����(<D��2�o��f��;i	�O��� �,8D�h0�
��t1q�)?%t��X �:D�hqGG�.M�cǋd~9x5B;D��Y�a/_�#�L�����awB:D������U#p���E=x�4�B�G:D� �W�˝*	Z���C�*��|�C�"D�X�Ǔ�`��%O�L�p��6D��C�X9@@�tҨ��5D�� (��E��=x=�� Q�ЫRL@�3�"O0���%�G8p+ �W=Vذ�"O�Y��匝A��H
�JԼ����"OT˷ U�X���:i�5X�%�"O h���#�x���bM���r�'�Z� �	؟�I�4��ԟ��I"7S�=cGj��W�0c��7"4��	�������h�	ڟ��I���	��P�I4��a�ң7� \X�R�����؟��Iɟ8��՟���ן�IҟL�	�W8-XPo@Jk��q��'jBI�����I����I���	៬�Iݟx�	�K%�-J̖�6'��h@ǂ+Qߴ��	����Iߟ�������˟��I����I;B����&�e \u(���9"��������	ԟ�����d�I�H�I۟��!L�mq�_.L��b��9Ѿ��ş��џ@��ȟ8�I��H����4��=.LdE��L�g:�!�B/��8-l����l�	�@�Iޟ �Iݟt�I�P�	f�:��c�Y7:��oF�C�q�Iş<�	柬�I����ڟ��	⟜�ɛ��LZy7�_�Z0����<�IџT���������L�	���p�b�2G(m�4�jw��
Z��	ן���ԟ|�I�4���4��˟p�	�!��X�n� /x��/X�|��L�������П,��Ɵ��	������\�	9>�I� L�2m�2������[L�@�I�����՟h��՟��	ݟH�ߴ�?������B,vBě6-�?H2H��&Q����ty���OR�nZI��E� dFK�>�[���D���A??�d�i�R�|��yRhr���D�#;� �G��\�e���H��=�	�O��$??)��
@�[#=��v�|@Ѓ���sEB�qF�Ƙ'DR_��F���J)Th赍�"��\���@R06-�
L�1O��?�
���s��O�^걈���'Rv*g�#����c��	T}��$B�&7Ohȳ"�[�f��A(λg��0
��j���af����K�.Lc���T�'�Q1&)�Y�5��睍Tn:��'��I^�I��Ms��|̓P-�\# �Gk�X+̈�����D�>!6�i
7r�@�'~����Eo�8d��Ͼ�$�8�O&q���A	~Q����\Dqr�]��?�Ń��[	�0�r$6"���6�����<��S��y�͌3T�@���(�4��ԃ�7�y2�|�:��䕟�Z�4�����J��f��Q�͏t�RU�����yLv��mZ�� !� ]���'�RՊRł�j��9��ZO��R�AKq���AA�)==ў��vyR����Xt�=*$I[)c�>�y��	����M�� ��d�'���@�bD�`*�4���v����S�Xٴ?���?Ot�>�)�O��Iu!G��j0���(U҂Lr��')vl�S����f�!)�ҳ�bФOM�'��	3Ⓔp��]yvN�)�r}�q�'"�Iyb�|��gӘ���3O�M�oG�b|��h&���RN �-��d
��Ik�i>�I��M��i���5;���R���W� A�E�!1�Z���it�dX�kC��0Ѧ�od�i�O��DG��8͊֘
_�fu�SK�@e��Q�HS|�	П �'��)�'p��y����b�A*q�!P�L�<�i��B�OZl�G��* �cR�;t��xy̌=�f����ēۦi��4�?��KΘ�M�'6j��7Gti�Ef��Bm��J�#�.�t bb����x☟�kyb�'����L
���RIZG���'��'��7-�<Y1Op�'I�b-�נ%�j� �M�t�B��'#��ʛ&����U�S�?B��ǛY �	� _*.��ؚ�(,t�d��b��X����,�uw 5��_9)�:@�->b^� Â�Oh�D�O �$�O���<9��i�44�(S�L$�񒇄@_.lk�G����C�U�?�CR��ڴhh 0���9d+�сĖ<A���i�6І�6s����0�t�Xs�'�� �'ո`"J��.:��+�.�ڋy��'/�Ih�O(L���#֙F�~���I�|�Ь�$m��*'�$%�S��M�;/;�(����t\)����D�i�7Mg��ק��Oj��O�\��6O"����ۻu�܈�G���P*�б>O�[��
|<ԁ��B ��|���"��E��5	�<2r)�N����(���YH�0�I��>|�T�ߩ~U��F)Ӟ_���?� S�|�ܴ3��f?O`�de���RN(8�:�9��ſ7��͓�?y��y.�s�Ub~R�O�H����!�ɞ#h�J� X5C���$֪�*�����|�I��IO�Oz��=�)��c�-�i�* �Y�	��M���^~"cs���.�4�F���Ĳ����B�$��L[�8O�nځ�M#"�i�`{$�iv��OjJ*դ@�J�3�(ɋ"�^eH��` E�Z��u�S&�d�<����?Y���?Q���?A�Ό�j�������,�"1�
��$ܦ9Bw��I��T'?)�IΕ�"0��}��AJRgbI�������ߦ�iߴu��$�OA��舌gUIS򩏵T�\��&V)z�A��� Z��I�X�R�3� NǺ���	�'N�R�;4�A�2�ڴ�	py�S��'�x�4e��9��
�=XQ2�B��Z�� ��&��4���ߦ��ܴ�?��������ǋ�8}H��qI�%'���rش�y��'".���q)�]I�O�	��� >X %�W;f!�UQ�j2"H���7O|��<))O?�2�(���"|�d���D 4*�	�MA(�W~rOb��$�<�A���&4����q!���t�Δ�yr]�� ٴ;����'� �2'�i����O,�#�cID1qh�)��	Q��/f<�p���8���=ͧ��D�O��Kn7@�JQ( w����7O��O��lZ>?nc�$�O���SQ��(X�	�V'O����O`D�'��7�����̓�ħ�"t�K�vtͫ���nh@�J7N�F��y� �Q0nHY�'�����\���w�	�5���0#X=�� )d�R2y���'�T�b>�%�n� U��H6㓶V%ց��ޤ�v (�O��mߟ@'��s�@�ٴM#�	A&�!oO��Z��V�J1��#�i�R+P�]���8O����L�­]�rq��>:/��J���w����oK"��c���	by��!r�]�cN_�8��a���aw��aشSt���<��'��'SN��w�>=���X�|~;�Y�C��R�s�XoZ�<Q�O�i�����M$O�6�t�����*!��ڢ�[�K*b���Mt� �KȰ( J-��'y�����'�x��T���V�NE����ә'��	x�?�Mc�bf���dy�Q [��W�̂wvRU*�rh�>y��iv6-|���'���u	�::�l SCd�z��C�'� ����2SH!(u�A-������ݚ�t_wv��\�D�
����ߡ![�%�Pg�]����D�O?牋Xetd�㈖�h�n�xc�83�N�8�M{�n~b�g����5�4��ɘ�'�:`�8a��=NO�8Z�;O�-l���M���U�:mC�4�yR�'��� r�Pc�h��C]�-qN (a�Z�f��<��N`E�'��i>��	�������0�	;f��#�ܙq�	��IN8���']�6M�}�D�OH��-�9Oh��A�Ӑ1Ύ��gI�#24`q��KJ}r�n�ToZ��?YI|*���2�Ǟ0+��m�5#ޤ5F�� iÃf�)���W)��D�-Rz�
'�bݕ���D��i�8*B��Um0��AAܑ�v���<�,Ot�OF�m��#���	�5D$I���8k�4p�,�r	T��M���y��i�4�oZ����� #�(:1��p1��t���*[>�nZ�<!��q��%��!B@��'��T�b�QӲj��B��H�3�	~ �� �a�|��Ɵ��	ޟp��ey��Ta�)(��I�%��4�����H��yR�'��h`�Ja�G���j�4��FA�I��
��0�*�9_Q��$�i������������,�	�M��'~+ȣ]ࢩX�ٚ�2�z�)=U)��JT��i6��됞|B[�����������L�dG��C���:��Ų~�*����PƟ@�	}y�	k�rY�W6O����ON�	㟪��bd�,D��P�a�5+Ą
����`�OD�oZ��M��'��Oh����p[.�� l�#{��J��&���E/ʌ��yC _�6��L��fq�!HL>!�_%��zK;n=���fV�����O��S�g~��m�ҝ�Uj˃��5M�t�!�-ۙ����M����y��lӚd�+�+�p*�+Qk�����	�ɴ0��nZ�<i�c<"��@�I�X���'EP�  �S��9��.*��h2�'#�ן��Iß��	џP�I���C&St�k�
�6|%��	�
4G��6��9B�d�O�d5�9O�`oz�q�b����E��'`"|tX���M�Ѵi�t�D�>�'����U��Y�ڴ�yR��E��S2"p�	��IX�y��Y�e���a眴��' ���|��.g��x�o�0<qn^<����	՟p��ԕ'n6�U�P�ʓ�?i���_(��)�l��I$�5��'A��q;���~Ӷe�	r}2B��J-�6�	0������y�'$pMkO�~�2�;�T�`���E��"�瞐q(i���QN��Ǆ�u{�	cy������Zc$������v�p�q�^���Ď�=b�>?�E�iw�O�	�))�Z��E���	Y�̓�S��ͦu��4�?)È8�Mә'��OȲ`�D��f)� b�j5a����Q˶�@�d^��1b�|�Z��ӟL�	��t�I�t�EKZ�a���$%߮�����jwy�y�6ĸ��3*ܼ���O^�S�?���Ovq���N�z�nI�"�y�ڐ����<���ip"6����x'>9���?��s��ZV�����h����7艰h�|���Jqyb)�0	2r�y����g?9"`f�0��m��xc>�7əf�L�r��$D� �枷X��U�#lJ�G�E��(?�� ��k��̿k�X��V��Z��#�.S�(��� ���J�	����ы��.��I�!V�^��������8Â���:c�5H��(pX1J �4"�rX�t%�@=@�0bZ�<�!r���\{
Ы��.?�u��A���I�`
 p_� +S�V0V�Y�	 ۦ��@9w����M�+�*=�ƅ7����O���+���O���ˀ:�����#�� D�-y|�j�#R3p�lnZ՟���П��IПP��,z�K�4�?�+l2�@�s`����W�G�X8[b�iGr�|��'Fra�=^���'ZB�%N� d��k/<� "0D�^��6m�O����O���N<���~���P ލ"�" 
s��-�Ee�?de�M>����?�C-�?���?AO?-)Ǝ��W�T�V�\�e-�8	'�}�����OڝId��֦�`��\�$�>`�'�|dk�f1#�>���F�,�0iP�4�?)�&G����?����O�	PAU�IƌL�(c�\���&�O���"��7}��m�U-ȂT�xr�
�%�2 �m�9�S�HP��y
� xaފ/ϰ�X��z$p"sG��M��2���/�б�6�*(C��9�cۀ;��)�s��f'T�b�E��Y,��J#�@�H��I^E�6��u&��>� t1�r�̵1�FS*(
��E	�h�HJY�_�D0�����*���ǧ��}}����L�?z�>��D�	�M�u3��Oh���O��d�躋���?)�OO��@"͒�!Wle����0@���)f+�����bÒ�r�z�J�n4,O�e"�MK�vz.x����vIrl�Ƃ�4*�l�hV!��� JK]X��P��տ�8Y+5o������QlM�j[^�DE��Mj�4��'�b?a�!�ηL����Z! +�� �3D��7,�#D�HCe�}�]�dd/�	4��$�<	A�7g�V�'�r�ʹR���%V�%��;�b�'�����',�8���!��2pcV%����+���2�_�^W�䑳/�F����`e��f�2]�6���(O��ɣ�Íf�0��3㌽v���Je��M�^y q�ڷ3<���G�G���٧�X�(O��q��'��6ͦ��	0XG���Tn�sե�3_P.y�'
R���=P�Q	��_�1p>���)5�#<��4��oڽx�@my7�O�KDF`�W�W����Ivy"B�
y�\7=���d�|*�?���֊�Z�iI�3�z��2���?���-�P�A�,���ň�N���R8�*��ʧ?����H"s�Ή@���:Oz��O��r���e��t8a!��c킠(gnZ�%F��\ꠧ�%P���@ۛ%nZD��>�c������4r��>���2	����_"(���[�t�:)a�94�P�R˄)I�(�i����u�j1��h*O��Ez"��8Y���d�[&	��Abaى2lZ6�OH���O��`�>d|���O����O䰬;��9��d��s0�a k	9��a
ՊO#&I�U�Q:�8�QcL���O�����<�p*��'  ��C��+�>mɢb���HqHQdާ���R%&,��}B珇�'�<�	�#z�����n	4�FX�f��I���I�_k�y�)�<y�{e��B���A�����2�'F�b�E��?-HI)P��7R��'Z"m+��|���򄍡,(�%#��5!�4��d���9�,�c�G]�|���d�O����O�!�;�?q���?� +�oij�8���B�%���_�b
�,�F痎+���jP
@<.��ƄV�QEy�T�'���㑂�YP S�ς�d��-�?-	�l	榉��id�Z�ߜAFy��$3ݬ����	А�B�ϖ'�F=X�kI��e�\�d�<����'r��d♊F��0�o�� �򔉘'4�y�|rBN�&���]` �������|�iw���m�lyR�.k�t7�O��D�{"�� ����q"Q����$�O�M9���O�ds>3���X�d~�%���J+-U���k�R�^ĉVB�)7fl��CG&ֺ�<A3�Wd��ę��֡5Q&ܲ�EJ%r��$X�'e��r�I.i�&����ږ'L۱�Ū��%LI�Iퟜ�'$ ��K'[>"�(D�tA�0��'���'P�O>��Q�9L )
s�
��Q��h=��hO�i��i���V�%B��u���F�� QB�֟�'�H�beuӲ���O �'vϺܻ�~�2Ѣ��2<$ڄ)�M�y�P���?A�F�q�^H�y*�|�$���BL���=��d�|�h4�O�e
Q�M�
�1O�Υ�ǧ���3���r�RY���>1w���L�Iǟ��	u��=Ā�R�@�r~ ��$�.J��<Y����<�)P�͸�r��-�!G�����d�yE��U����\�+D��=E�hdhW��On���O�H�ώHH����O����OT`�;H��$�A� ��p�$�V�r���w�Pjk��~a6���ڷ����T�>�:Q��9����&��3*\�;f�Ǹ+�J��N%=�@`D�r�g�\�I���N?`(�9JVoT�w��(��4A��3{���4����<�I�[d@�3��xCP�t�B��=]Ŏ����0^DT�B o�����C�� K�O��\��-q���;��e��/�%f��
�iT	U �s��?����?����D�d�O��ӷh@����m����6V o�.�-�a��D�Z3đ�%*\�)�(%���ɂ#����,Ɩ�Pe*C�Z(���sf��4����r�Y&��U32)�P�L80��I�BՑE�*��!��ȏ�][B c�O(�lZ���?	����'X�%"VF� %�pP ���&��r�'����!H�Gܘ����UR�4��y�dtӦ���<�q���<��F�'��	�R'�	��o��<A��A�,8�r�'d<���'���'&����'L�'B�Q���I@�i����p�%�
Ǔ'���� �G}�T�'*F�P�Ȇ�"iX�A"�[=Yv�J
Ǔ@���IҟL�O|���a�N��d"�%�����'4O*��O2�O��}�A#�+P����gͺ����y��C����M�3��) �>��e� Hq��,6pq�&S��2 ���d�O��'��Uk�p � e�Q�2�uy��!]\�h��?���0������A�@���]->]��n�d�׎B�Pe ��֯!�Ɉ`��2��	9n1���#G�u(�tC��1<�
`���n�7Q�A�ND(
R��i���I	Q*���֦UP������}�J7,�͠�+J%X^��.?4�� � a�'T�)��0±k�FL�lK��'^\#=17/�:!�y���*$wn�|�6�'k��'��u���sN��'(��'���ݦ'6�M��o�;g��DN��6�v�Ka��-�|�[U�^=S鲔@���f̧a�pD	pmc��{�)߆0�Az�l�#d�T#2��d�|ѩS�$������ ���>m"cB�g.�>:O�uc�(f�$$p"]�r�o�	���A��O|����R�)W���n͚|�D�K���*]!�d�>GlųV�m}�)�S��*Q��O^$Gz�`ӄ���<��A�<����ՊY��UspC�(;��=�����?i���?1��3��n�O���i>����<]���fF�+�5#���-�|�0�M�(��1S_�v����	
}Q������EC>��7O�!H�;�ʏ=��1� N k� ��(�,Ƞ@*�scQ� (7F]�s1� ���A;~��jL�V���dʦ1	ٴ��'ZBb?Mcg���H�)R( I�ã(D� ��g�F�f�R�GN&n����%��M3���򤓵���O�r�)�~q��2"@�����'���C��'��6���c��T"$@�-��,XS?s�٣H�*-� ��U&I�P��F8�����0x�9�I� �~"�X�6�0�TZ�*��0!e�Q �p<9�Lџ�
�4��I�yL5{r��2^
vA��2	;Xc�@��vx�ԢF��V�6ՑW�ċ9y��ɑ2�(Yٴw�x���D���H!A��P��ϓ��D]+rO~�l��t�I@�T���u���h��[Pk׎SmD��V&ߟ`uR�'��QI�@@�Y1O�Yy��Fƅ��a�R9�]�Ȉ���ɧ<ʼ�4�>�)��&��kY���ڑ��48�^�#@�>��#�ȟT�����	V��%ԨM��b֘i�,���d�
��<�<1����<����61R�"�F��Dr���Z]�Hr��d��)��L���P�#a�@�f�@;Fp-i���Oh���O6���ņ������O0�d�O4)��sY�x��타H���Ge1�43���>I�>�X��Y��T��'H1��*��PP���<i�&���d+\�b�>�����M9���ٴ$Ѧ-B0+X�a�2�#��DꜨKp)̓;�<zQ��#� �ȃ\G���Űi}�7��O:	���Oq���ޟ�K�K4t�4�q*8���qy2�)§`�2P ')T42*p�Ā�<Brq��?�4�i�86�/�D�:�ɠ<g�k��<�$	��Uv&DG��XML�C-� �?9���?�d��.�O���t>)X�'��G�l�0 �5���8��N�$:�C�Ip������A(1���� �7\�vMHB3���Ћ�#3p�����tE��`u�
F���Zh؟�9��G�k*ِ�~X��5�1D�D�@ ��n��M��hē7�1��	;�	,Ȱ=y��c��� ��ۅ"7�䊦�\M�<Ig�6\���숸|!��*e�c�<��a�#�v@q#� �tv���'��x�<Q�(�4"�9E�ƒW7�d�Tj�z�<i��_k���ĊIK"=��v�<9!艀w�D0�ʪTBޠ�B�|�<�Q��=g��t�pO�R>d�XsB�v�<ɓ)�E��̙6�'-y��h��[M�<ѣ��V����،|��EÐ�I�<���uԸ��w�������F�<�V.
�@�8%M���@�A(�I�<I.ٟu� �2Aϔ�ePT�("(�[�<�c�HԖ�bNS�6e�q�Z�<A�Mՙ}�b�c����bN�V�<ys�
��8�u��C��8TC�F�<ac��1U�]P�H5R�Qc���A�<���R�$�2��Bnֽ�d ��E|�<�U5$���+P�<!ی�"��_�<Q��L8�B�J=��LZ���G�<�c�F������E-}��P�aBB�<	�mV�1vn͚���'.R��Y�dS�<!w2Ѽ@��ռe������D�<��A� _>�a� g���F�NB�<!�MM*O5H��b��&<x�#�e�<�AT����e  ��KP�\�<�p�Q�Dv٣��Нp\���"EY�<qwN��E�F�c��[0�n�xW�L\�<��[�Ex�'�eА��Ub�<� D@���-8]t�e)^�'�Y*�"O�ԋ3�@�	�`iJ ��p~�h0d"O6��cI
	�A��1_`j�"O���E�"���($	�n��$��"O���.إJ0�}���
x�Z��G"O𭠱ƛ"`�)j��Lk�� f"OP����1?�1IB"��k���"O�`�`�xnz�Jb�,p���I�"O��r��SѸ<`1��9It(a�"OХ��Ð�zI�u����\b�"OY+�ٿ8���ٶl@1MJH[���;V��{�'=��,T�U�RR������\{"�L"x�R�Atd�ɕgB�%�c�>�5h�v�\V��y�+�$�y�O��t�`3�Q��]Q�
���M��M3A�f4(���k�Z��s��T�?�:�ȩcěi!���B��#HU"���X��M	�E�4z�@��O=-d�F{�)��d	C�J� 
�6����L�
K�(0��\��u�*�T��V�ȱ���-@N䱀A�:�`$st�,O T:����#��("��,�e--�x���b%?�\� ����Q����#�n�Uc�!@I`e%S4���x�s�),�Ԉ��ė�P $���!�>Ic
Lq��J��VȠ�H7!�Z?��D*����Y���X ��*ͤ|����GD�J<��`�!�Ta"#��#wᛆ�J�G��2,�
�d�y�&���S�'ݼC�i�!E��-���)l<����TqO�]��Y��gk^t�]��+��K;�!�� �	166��I>��w�˓H=q�8@����+f�"�1��I�ĩf�m��` "OJ%s��ռ[$%�c��в�o�֡�E�R(2�U�����:5��O���k��C�W�By8S̄�kR~�#����%t�4���*!<�+bJ�i��	�3�z�1L�*U���8#�Cʂ�<9��sjz�5D�
4��:+�CJ���	����p����o���JB�H�.�n���`؊t�4XsU��ZQ���Q+4���֮grZ!䇋\5����5 ���D^+!���r]wi��=�S�
��l��kФ:�J��ӄ�{��:��	N�t��I����%8:�Q⡄ �d_" J3 �~OL]��B�|�0��ܓ�Clä�jŏÖ?�~4���d����wG.L���&R>5��'P���a)��0��3i7}����� 4h|h첐L٦HZț0��W�Iv�`��/K ,����r�P'kS��F|y��O����ɦؓ-6F�v�@kӞd�ɫL�" S�� S�&�Y�@�06-M$$J�!db�p����H���$+�f��xB��p4b_< i۱CM��?�#�,����.ئ�KR&��hO����#	B7-��9D���bͬA�^1Dr�O��@x�������� ��v�Fp
�g[
HI��3�ol�����ML�l�8��VI��Q����H5��h?QI�p�O�� l��>FRQF�W� [��CE&��h}<�Gz�M?c��)!��W�m�� �OQ����݀g�>�pTϋhe�����;O��'��������H�ɠ'<>��>��ai��]��{��'Ц,��J.#����h�	xZ��Y޴\��al�!VS�3G[2sK�L�=�#-���y���ct�\��L͊�te(3h�	�� oZ�v��[5˃�L��9�+e�����Ԛw����x$jii��O;o�J�{��p�o-Ɲ��'��$���)H6��`��O7��ѵ��'m�du@�.6��xRO�"K�`
^c��Y��(��k7 �l%�p��5�����'��֐:����R�����(�ŁM4R� �!J7^��<Br�2ғ+�	��ȒZ)R����?� �'�y`�V�>�eh���US�(OZ�X�L��?���F�ٰѮ��5��%��I�4{�-��� ؖ��R�D�Qؼ�&�#bh�6�x���1�}@��b@�=W�������E�d���0��׻k�y�$阺�?I2�,Y|��2��H�����U\�'Q&���Ō^llP���ן/��mҊ.�X�?��}r
)\����IN
k­PF�ǫ['P��q�1I�x�J	!^/n�BYcN:\h����El�M8�	
OJp�{���d�T��+g�.5�O�	���U܀�X��S��g�'d<�#��$��f�#?,H���O�DHn�=tF`ڧ&��x�q�$��x�ݴHIR���({�7�uw
�O�i���Q$g���q-�^<�|2��iu�=���Ɵ]��D�҃W���ш�d�6��A�JMA�(��lQ��9�Q>��VX*��
��TC��_1���e��"Ia��ܱB@4qB��o��M��"�6��) L4��x2�G�H����aj�U�a�G&C��X��G$W�~���ŏ����Bc	3�FL�'hԱb,bQk��΄�HO&U��������0�HV1�4�P_�<�fQ1
A���c�̕
�r��eA1�o����{��]�t'�<�	�lQ��Px�"��D(o6�j������
�R#J~���&�����sF���,ջ�칟�ړ$��d��b��-%O�QÀ/�U`��c�E_�Y�=��͠!T^lP������� ��#ݞL�H����b�x��YB���˰�'�|ɡPc�/�i:�" �^߶�
�Ƈ<J������>�>�o��s:=3�AJ�lyr��3��r�<!'o�< �*I�5FO+1�܉dC��-��Ji1��k!�'�Pq0�-oEv���ꑠ/����R�\<�퐾?8H�d?��H�-��s&̶Ƙ��!�DS�:e���s���px�r��)�O�݁"`���K��	W?qS���uf�s
��c ���!�_!���q�R�K����!/����^�.�'�^#}�'��S%,Ĩ*)�l��)� R��hc����:mT	5�Z*k� u�3�D�Z�4=�-�4.͖%RH�1ubͨp#�����јƤ۶L�t&N�ft����J�9��"�D���DQgcw�XX�6��� ��)1�j�hjl�'�I�!\������&U�VH"V垆��I5MV6�X�J�jw4�����0n�Ȣ=I0�L��q��� ��K�N�Dì0#��'b�������eR��7jF�B#щ[	:k��'�ܩ1}��re�]� ��a��4�)`�+7�O���aLڵQE�B�GX(\���X�D_6�����䌤b�J��'$~h�B��;DI�I�2�r�;1�0H$9!��ڔ {�>)� �SC: �L�3B��L�O@ǟ���a89���vaT�\�x�#�k�>�/WVP.��s��4O��q[E�	�pE�U�Z�$ DH��ͮ4�|�ɸ8T
�")R�v�#�W�b@��=��BֆE�0Ų��m��I�eO�h�dlZP�'E(|�4T�Y��ģ�S��|��U���@4��'���ʃ3�i���=,���+[;nf$������	�T��'_?"m�T���@�� ��D.������k�$#=�"A\ 1�B��F*������U}r��<�p+qeާp�Dl"g����ɜa���2z7A��)�R�2@�2f�t�'`�ehԔnN	"��T`�A	�4|5��V�ݩa��@���h��F~�(�6�: �4�
}$`gn�:)�R�b��À���'ff����Oў��*� +P�`w ^�%Ը����0+Pߓ{{���9�`�hrD�
�Z��e+�"R*��֮f�t�񤇍d��I�;]�hjT��z����X\��F|��m�nJd�D �`��(9���J�U
��ҞF""=)	[䔝I��"eG*�HTa_C}� ^9 ���J��1�"�?��P>Y��̠����	�'2 ؛E%�`�^�S���O(9;E�J��@�N�3m�E9B�i'��"R�N<1��٫s�'��Pp�{ҪF�C$�8l��+�tȚ�� 4�Q2e�9���ɴ_��鞲i�Θ��õ7�d�=��d�f��8��	6]P��g������D3�$�>����@����C�nh9�;4��p��ѿ ���eb�8_��C�%�/�	Ǔ]b|hZ�6��	�6kB��V�QU��^U0 ��C��Is���hMu���=�̘��L��̪G'�5<s� q�8")��P�	Q�'Ȉա�
�yÐ�B�
�T�F)�O���A`�k����C7o�>�hQ5Of���L*N{Dp�4�k���EhvӖ@�a�(&|3ժ��H�lΰv�j$�4�Ij!�MZ��xӒ��fM�$F=�E%T�	����>yԏB�S�* ,I�Y�p������O�T(�d��6��=�O
���A�
jpj7�30Q𕳱�	?[� Z��|��8E��C<��1�����?��X�agD%$�4�c��$lBc$��S�^'bG�Y���pB&�3B*�~��xb�G�s����;i�V��)kӔ	���E�轒4o�0`�j��4I�0,o 7�m��.����7Rf�X5�W/$�Xt"4`׊3
L(�~�'����ң� �:�cU�Y�&��O��T�'[�4��-Ⱥ7ʢ�9��iՊ]�f���]7:X�BQ}�29hQ��%/vzh�I��D��㟼2d�S%��a�C��8�l�Lxh�,�,[�aj�	@'"�{a����ֈ��D#�ƈ/�RU;����c"�zS�0�.E�S���U�v�2M0i���#>>
h9$GL�j��r�oI�#�x<�竐���$גt��y��W1MGd�Ȍ��m�b���k�l/���C�/>[���%/.0�x��F,)?��ݣ}�]�q�׵^4����0iH�=�#���[W�]�GG�����dj�iײ.���Ԗkɚ�ȷ�Li���J�cI/WY�ipbە$�d��p.�>�外.&��p؄j Yʥ�q�Ky?!��p�cR*��<qVCs�K�)���Vf�O�!�01!Ij達`(Aѷi�&�!"��	- <�����AH>�'P�@ �6M��m<l�cg
�h�x��Ҙ4���ɶ��щB�ȪWk*�K�E��Y�<�=�W�Ƴ)D�-wJ\�Z9����?%l=�F�|��o�$B�"|����$]H�����)no
0��̉?�hHЁlM?�p<)Ġg~���<`2��@�>�q�O�!q��YċƦY"K>E�t�O��j�,��b�t,��l�9tC�PrF�LQ�'�5K�F_�	�@z���a�(8��Op}qw��/F"8p2fe��U폴�~⃁(��'����O�ƭ.1�����OX������uyg�_8S|�C��i���%� �noL�	cⓏ2�T�K>�g}B
M-S>�� ь�D�>�H�`�;�~��&<�$��aT�DC��!���	�hO�����H�|5�aJGaD)^�5�\���K�xi"��qO�Sz x�A�.܏nƭS�n�z>`ģ�G>dk���� *%�e�}f���QF^(m�C"OV񣗬M�2�H�{� [��)"O)�d⟢E��d@�@D)�R$"O��pW���n|�p�	q�1 7"O���a��H�JA��)V�A��"O��If�J�jM>tScח2K�0"O��3VF�Y=\�i�F�<yKF"O2	۲�_�d^<��p,	lj d��"O�����������2��v80�t"Ohe�&��-��)A�S�2H6�&"ON�c	d�z5o�=jBn�q"O2 �D� !����� &4*ΐ�"O�q%MT��m*l�@��"O�S�9R��<h7,��;rF ��*O�3œ	}@��(Ѝ)�
U��'y^�
����="�E�GL ~�H�!�'89��d\	��E*�Cs=�"ONH��� �iﰕh�"g�8`@"O� �"D��d�B��;���*�"O�!(f�� H��(Y.F�H�;�"O�YAeB�#	�`J�m�|��d#U"O�\�e�6,��E�^=2�L�0�"O����=8(R*ӎ�D|Q�"O�"VN�-#���P��d����"O�I&��Ym.��� 3L\]�"O굨Э
=�$ЫS�M�LY.�$"O aH�/S�Zڂ,G��DF��"O��qA�*8��b��)s)�d�"O~���I�JA#�Ӿ��"O<�1��i���ͦ*օP"Ol�ɁC*���҇��RB,YQ"O���O�T�"  r� \"G"O�d��d�%|z-�6N�3����B"Op�x`���^}P�0p��!Kb"O)�Մ	*1��qVnF��>W0�y�o�"|�
}&r9����-�y"�.�uC-Ki4���F�zw!�όd�c�c�;P��,�)Da!��*C &UR�`�42j�� ��R
�'��Ze�	����@��3F���'��ё�'E�=X��g"@�mr4���'������K=7���+�L\�.�,��'b��j��Wd^��
!�O�;�����'k��2c�e�X��CՍf����'K���P7H��u���,V�T(!	�'�؈H-|���$� �SH�ժ�'�<����:K�����,��^D��'���⎣G�t!�A�����'G��3(Ky�8�sh��.���'��sQ�_�)���G8 ����'�B�:�BY)UB�0�8�tC
�'(��dQ/BxP�˱h�%`��<�	�'�  Z5�N�?`�zQ	�Y�܀�'����FM:Q��)�u��J�
�'r��&
E�#��E�	�;|�T��'y ��S��]��Qt��2�xM�
�'���I����t�Z6mX�S��X
�'�$1����>rf j���8�r
�'��\(��T�`��U�Q���.�z���'�\��c-�n���N�8&�9�'�����G-~"t0y�����0ġ�'R�8#+T+!��L��摠	d,�	�'$p�Q@䌽l#�!�����L#
�'�~���ș+M�88�W����1�	��� �ڇ��e�]��,V�&�����"O&�k�'�=~�{@MD�|0�}��"O��3tʇ-#�]0�ᓈN7H���"O�����8��T��Es#�H s"O6�����HH�S K�N��"O�`̀3$����=z����e"OܭZ�B��Բ=�5ٺY`ȴ��"O݋1It� �� I0[ ��"ON=�ff�a�\Ui@�)���0W"O�R¬��NP���ܵV����"O�`O:IQ�E�6?�Z!5"O�]�H� V�h3$ϵ+�L�"O��s�,ȃ]�r�@�H۳3�f��$"O��@��H9Ko"��J�
�0 r"O"@;Ŗ�K������Ye�<��"O2Yrf(%�ʐ0��V$�p�+�"Op���)֒&�P��aD8����5"O\�cZXūR$�3xvX��&$�qp!�$�	Zb~q)��ń/du�a����!��4p`��^�P�A	u�M1p!�$�/I<�0xfJʫ�2�ǩW�4}!��͹���"^L�x�f)�'��1O���:��{5��2����"O�<�o�h��gI$��͛"O+�A�*�(�H�,`�s(�"�!�Qٮź0�ѝ"�ĥb�9�!�DD�z���	cF�Fi���$l�!�DR"ĺ��+�F�ҡn�sx!�ĂE�Rm�a�Ȧb�&�*��K2b!�c�ꔱ�@�-�"U�v�8l�
�'���Rc�KX����v�D�]����O��=E�$��>Q�� ī >R%*G7�yR��*�|L���
�,��F�-�y�-�6Ш3gS m�"���iU-�y�B�����L!e,*���б�y���F����B�_��jU��3�yr�_�l��88#`Q�=b� R�����0>ё��F|�\� ,�:A�X|b *[k�<9�l�!(x4jg]�i���q��q�<�W��`n���7Z5N�m�ȉo?����S%/��<q���nÌ�*qǧ<�hC�	�5�(y�ES�8_<�*�J��BC�ɅJ'Bpy%�V�_�x��@­V�
C��,�`Y˵�^:E$b�̠y��B��2H	��NۮiM
�CʬlB�I�Q�PyP�	�o%$E�=t|�C��6��r���h�b@aVB�5JR�B�	�
$S���0
�r`K��\B�hB�I�XU,�VB�9W�~iZ䙖����y�I�i�YaF�NC��� N���VB�	�b��t���p0�Y�g"�PB䉖	Fl�(3+�`���ɝ�	��B�I�U���!U"�����ݭE�B�	N����(M z	�<Õ�H�d�dC�I�F�Ss��%/�QR2)ѭ�BC�I� ���S&�m�j��'\I�jB�IM/�����)})��Z�,@B�	�K&PhA��B�LA�hλ:h~B��']<��3�Uf�
EOM�~� C�I�
�0j��<qf���b C��<u�d)͋nq<R��M3�B䉚v$��C�J)��Y1s���QBPC�I�.����#c�
��0�V�
�rʌC�I+#ٌ(��	@>r�~�[��'C�)� n���-U�wz`"0�H,T��'�!���Qw��U7!��"��\?EV!�D�i���+n������0}6!�$�;i�Xm���I�v�a�L��:?!��ңm�T(��aIvVƉ�����l9!�䘰g��قc�B���3��=�!��١�B�R�蟀K��'A�:!�ĒD��A@��4���WED�"�!�D7O,%1"蔉�: ö���!�G�\����pH�5�Pa�a팶!�!�D\�vX��K�I.�1i"��9�!���6,��"�k�E�e
0#�!��PJ�Ju�7@�>I���
�<&!��8M��4E�<-����UI�/a!�ۡrҮ�I'j�'��j�HE"Od��� R&q��Qp���
�j�SC"OhT
�*�����(HTbܑ��"O��+�fȞ@���$E'0Fڔ��On���%�NX���o�#?Hq�A�L�<���HSW�B P"=,�8���G�<���N M�
��3fҲDW���W���<���!?�U�s��2(A`9��B���0=��ܠS�F���Ń�KJ�P �X�<YsGH�3�Ȑ3j�6L;�P� Q�<�A$C������
H��-:5˕N�<��*'A����hE���DM�<���^t&p��I�8 ^vy�5�	K�<�,	�b��x��I;6��x7
�G�<�u� *����֎48����j�<yB�ʉ1��]���1j�Ps��Jh<��!
P�b�%��'^����4�HOL���Dª�K��SGB-�F�!�Py�g�23��x�t�M�xT�ŌȰ�ybn]�7 �x"�L��m�@�E�Q���	_X�8��M6p�!��·I�dKp�<D����Q�F��r�Q�@��q��6D�л��M'�a� �ϐ���@+6?y���SUEf�`nǖH?�LS��^�L��p?!Bk�^z�����<>ިs�c�a�<��C��q���)�� ����y�FBYn��qaH�漥vD��y�/J�5���� r��8�,���y��42�L��6lT�c�fU��)�yb D�D������X�(R��%�y҈��tš`Rw��9�y�&WW0��v"�o˄� Ѩ܊�y���nd��s�W+b�F�i�a)�yB�'��ݘ��f�~���BǏb	���'�Ha�I_*9!>5�#m��P��'���UI�XI�"�fW���	�'gX$8�cAN�6A����"JB�`C	�'�`�)o,�Y��<|�"�����[�>tL�����57.���D>D�$�&M�K�f�tL�Pml%��C'D���Gɏ*�<��#� Y�8��&�#D����͛P�Je�Uj��"�Z��,D�dC�	�d���Gሹ=vP��)D���D� -t@ʱ���h��$��i(�Z���ON@dI	�<!`|��©�q�<T�	�'�Q��&�dxh�
W�
�Y�jy�	�'�beHdO�[yJ8
�ˬb��K	�'�hu���9��lH@�O�Ul��9	�'��5�F+]�x2�җ\(��0	�'�Ȑ�uI�(f�Xe�g��+�(�{�O2�=E�� �����ݙ"��h)T$[7^h�B"O�`[ n̓ng�9b��ҴZ�MKU"OZ|4ɟ�h.s��:fB��j�"O�@Zw�4�z�I��25�΁��"OL0�q/��%i�c�{�,�IW"OD����.�QF�K�>�zU��"O��؂E�.������ǪP����s"OB��G�/������; �y�s"Of�wg
0�����Ş+��ʧ"OLy�Tɐ�`|Z����`r
�CW"O�5�h�22i�y���)gg��"Od ��%�B�J��_�R3�l��"O�T�g�Yc�n����I�V&M�'"O��!l	$-�����J�"jFI�"Oq��%[3Ek�ѕ�D�7��x�f"Oʕ��+s��@8�G�#G�Q�V"O�-H�ҿ��\�0酕7(D��E"OP�zp�Е?��K�j:M'P`x"O$��E�7!�n�Ӗ��>10C"O�9Yt���T�|	;�C�&7�8��U"O�QZ�ݓ<<�8���"H���8R"Obt�P�x(xPaT6?�4�X"O@��U Y9P��pb�.=��3 "O�TP���r�b��D�Y�'BX��"OZiñ��\�V���E^ ;&���"OZ@Y�L�1
�4)Y��"'\͑�"O��CV.ƾ{��`Ս��](�44"O*���%ԃ�zq��k��,Du��"Ol�rEc���-{����c�P��T"O��!Va�hKt�_�[Ǩ��p"O���r�P7/qj�`s
�k�Ƞ��"O�i�QA݅#dF��B ��e�ꝙ�"O�$òo���Ƞ@��t���"O�i��$J,=Pj=�D�	s��ٺ�"OЛ&IϺSQ|��'C�D�̄2d"O�5pA�� @h��d����x)%"OtY�cn�*-2��6��m�U"O����%A�9 �L����e"O����S�	�6�DK^7"�0sB"O��9W�۞l�`@�I؍}vz�p�"O<�h�U+^x��i`j)\4���"O�Xȁ�T�5Ϝ���/�+����0"O��W�L�}Tԑ��E2��8�"O�-��Bó:���IsN�a~2��"OP���J7����'�)g>�r"Ol�!
@/��Va��`�a�"O�p�6�׊r�6��"����"O�Q�$̜��2dp��=h���J�"Ob�C2�'6�B@�UM3�ruR�"Oj��K��V�Bl�#h���"O���4#�/�Je�2���A��t� "Oj�J�!�9r���_�|�p9��"O�L�A�'QK^II�+��fORtRP"Oz���� �4��DԱ'J���"O�d�F�_
�n�a�$��?\�0*B"O�5�T�ڈ�2q#ՂǷB���"O��	�&2Eh���>^$$�0q"O�ű'�N�==�<�f�/{2�J"O$`A���:�PX���,V綴��"O�Y#1e�3M�][�%�R�|j�"O���#9 �~���܅�����"O� ��O�'��i�A�ڌ��EK"O��֪��L|<�v�ҵA�J��7"OJ]�4$�Bh1�r��&{vѰ�"O� *YRF�N�Si2M�3��2w�j$"O�l���QzX�+��@</]	�"O*9���N! ���"�L��ٳ6"O0T�'
�a L�Ն˖f�Zx��"O`��c#�:U��
��U�m;"Om:���)%SDh����+B����"O~�0�[�&��iJ���)&-�W"O��4D\6O7\H��Z����"O�%��69�mã�� ��؀�"O�U猐G��Z���)�n1��"O6�ȔjE�P;� ���2}r�I�U"O��h�B�.7��T�UJLvm��K6"O���
�x�R���_4��|s""Op��㍓;Ayb�g�.�渘"O��֨���A�%Hj�
Q"O<0Г%�$��hj��7$�N!6"O�Q�1ICG��)ᑠ?s��A�"O�r��x�H z6���
R�h�"O��W�M��4ͻW�ğ@6L�A%"O6�r�<+��sG�I)^H�2"OД��BC��@����A�M�����"OƱ�aJ>Ze+�BSA���"O^�[�gKYF�����3{�0E��"O���f�/���P����"Om���O��NL�d)�?���e"O�h�!e�#���1��
^�r�"O�8��l_���]�/�q��"O�����: ��h��,���e"O�(����~�n�lP�Z*h#G"OZL'g��4�H�!��<
�y""OHT�AÀ�F�T #fK��߸<Rp"OZ]��gK�6�%�C;HAV"O�@�WE��옡�Z�.8
���"O��`S�ѹ5����fA�CP��Bb"O�)!5�)~�8�h��Q�2.��3%"OQ5h�������i)��z�"O2Db4�%#a� ���L�9�"O9X7�{���s��O&q\��`�"ON؊�ɥ�8%��J5q���sQ"O@��uFS0��a�U�:�$��"O��1��.�V �#È�W-�P��"Ov���7k�^�y$�� ^7�U�"O2��G٠g�NRp�� 5�|�"OX}� �ݙw�	��䁲f� ґ"On9zB��4@�� ���1#���U"OR�Z���Ƀ�j	[�\M��"O)0��I�\T�4���;3(�q�"O�k1@.Wg$�#K�3�`��"Ot�k�L�F�>�����8sP�%"O�}��ɀ�^��#�W�#V�e��"O�h��.E�Om�$���;�}�G"O	�E�$7=40�w��͐8�"OD��fX�gbPpE	�?
� y��"O��#���F�@QpGT�:�Y�3"Oh�$(gH���&����I�"O�@����`tŏ�Yl.M�U"O�8�sÆ�{C�xh3��<��"OV����&m�	��E�]]�`��"OXhٖF�QBi�2%ΰA�	�6"OXX�IH�V/��9�JE��(1b"O��+T'G�b9t��2�j�;"O�xdd��5�e�K�I�(d��"O�XA�n�H��+��� /aD]��"O��D  >��A�$�,�F��"O� v��r�_�d��ĩ�r�ʸ��"O�� 2c�f .A1�@z���"O΄[�딕L	��P+o�ұ��"O�}�"+��r|�m�Pm�,G�b$��"Oh�x�	*R���xuk��T��"O6��-ӫNAx�H�
.n�6�i�"O�a�FE��~͔Hs���?yu:�!V"O�Pɂ�6R�q%NԝW`<Q�"O��J'��:+��SíI�Cp*ݣ�"O�X��L�����ZP���"O�lp�&ڎ&����Μ7x���i�"O�X�b� _����τ	�F��"OZp�p&�1iƲAXS�2e�}j�"ObU��� �MM����4sO��b"O�t:sJ�Vɸ����O0����"O�q��o�`���HM6CY`�"O�KE�8i�U�įj9:��"O|kP,�%g��Y'�5�� r5"O@+W��&,Ch��g��j9�t"O̼RgܡH4���$��c��}2�"Oj�*6[�!a9Q�jI�ފ�R�"O��`�,l|�
 �O�+���@"O�pÄB�y�*��C�ܝ@�4(8�"O�9�l8F���i�AC�?�Hö"O�)C0�¬C�@����Ѓ�"OJ�	a�J��D 	���s"O�)q�ϽV��T��Ë�Vd$ej�"O����i��8E�j)G�j�^P;""O$��ˆ!����ԆV�[�yD"O�9��W����Ӆ���e�"O�����R�akt9�Fʙ�x���"OX$����2]䲂o暈��"O�QAV#	YT0Ͱ�n�+�P*P"O��S���q����qC��k�։sT"O��S���k�A(�bV, ���3"O��PìW�Ul���R#��}��P"O~,zlZ�, 4cP�MX&$;"O ��T%	S,LcA�XRp��"O���'���y�@�I����4� �"Or�+r��+�6$�N��_3�� 2"O�1�ӣ��S���S,�3s �)
""O�9*w�'w��y�+
+CzA"O|I9�!G8\�
 )�� $�pC�"O�,�g�2TP� �H�C��:U"O�ap��!ـ�l�>�����"Oi@#�ݢ�)T�JL>���"O~l��i�5���a�A�c�4 "Of��,�Q��\&'�5n�.�9�"O�hQ�� ��Tza,	=_�U�"OD<�D�0ߴ��U��'���b�"O����c��k�E"�yz#"O���L�2j��{�D�%x�v��"O
ظ�!�-09n0�É�W�(TbR"O^X��M>;�D�ŉF!T��cQ"O�}��K�AB(ꧩ��2"O"�1�m���6�C%(-貘3""O6)[�Ѝ(��uj�� ~�~��$"O�0�Gˈ���CtF��R����"O�Ղa��)T�d�� 썥/��x��"OE;wg��Bbٰs��h�A��!����"�s2nS�,ѸȲ�J�\�!��D~T"�h@�X���*�l�0�!�$���ɓ�W�ה�k� 6H�!��U,�����i�b�R�h�Dσj�!�� �	r��y�i��}950"Ou�ҧ�<(��!�/4�D��P"O�9�K�%x�\ Rh��ks"O޴ ��(�qJW�Z
�E�4"O��!��9eZ���Ş�2,҆"O`lA��71f���A��T;3M5D��C ǏL����.wo"h"%�0D����ϓ=lt9��W���Vn;D����A�Ε�#G.&<�w��%�yB��Et�ɤ`��B��8�c�%�y�▄#s�}ӔN8��d��5�y���l�������=�DS����y�JK�p�0�e�j���jW䉢�y�EI�8�.a�I�K����ah�y2�3�l�U�GH�V��PiD��yr�1n����=E�B�S��?�y�܅ r����G�+wX�q�m���yr�ͦ$t�!�ݘl����EZ��y��l>�����Y�)���Q��y�:�}hr�ݞ~��Yt`7�y�m�R<0��r'6o���f܍�y���-[j,Y�I�yt$x���;�yҡ_��6�: Gs(���U��*�y���m���U9g�@��H�y��WRhqHF�Z�-1�BGn��yKuO��C��?5Z[ak�,�y�χe��a���
�͊�P��y�i������C�� n�e�B���y�C�$r"C�!jA��p"����y"#P5'��@�7�6�<�
�yb'J9 :8A���?��c�Iؼ�y�f�B( Y�&�
��y�EW��9�c�H�m䮉v����yr��*T��H v��]��J��yҬ�>Đ����Yɾx��D#�yRgD�Y����ԁ�!I�����<�yr�� D�Ȅp�� �>��3D �yb�#��(#Ug��f���Z�._�yR.B�S46�P�@5�u���ڞ�y�Ú'M��H�B�ː(�Ę	�!���y2@�s��y���9X�z�Ѣj�y�������⓱Nd9q�����y�=Hb۷`A�\j5bBL�y"���=��;�d�)P

��K��y��ɏ>�XA"4�2^r>����/�yr,E]�d�@�"��S���J3䆰�yB�M����"���?;@���>�y�a�;Z�`�%�$`��nK��y�@Dq�ְ�6��ʰ�p���y�l�r"�8�$��m�é�9�y��&1�X�K�yTp�;4�P�y�W�bœv�U#tR�pH�U!�y�*���Z`�B
^$l|���B*^��y2�H6e��0Ư@�]o�&��}C�'�N}Y�����m\�Y>�\��"O&�C2NߴtJ���r��:(�.@��"O�����g|��(�C�`�`�"O�4�Ȓ�@�Ju;�D�2�Ձe"O��&	��0�z�!V�Y�2,���U"O�=Is�.V��q�tHB����e"O���'\��&�����YH<��"O��9�ď"Y���!�ה�X9�"OZ��a�:!K歑�4�b�"O���R�АX@ cPdA!�D���"O� FMX7/�� �THat�\��vQ`"OPt)F� � �XaMr׺�s"O��ƮN!3�^�c�n�UӀ�yd"O�L:��q-�1�R}��"Old�f��e
��D�ϣ%�h��&"O0��2CˊZB��a@�U*�1a"O�!����<d&x
 cF6sO>\�U"OX���E�H�B�Ѧ�H+Q��"O��M�u�h\�Q"�.-�R5�"O�)1C��G� �34�8 �j�b�"Ob�cF�
��p,���Ҙ�$Y��"O�8��aQ 5,�[SO̰�� X!"O�!�i��y����4�@�s�~���"O4m���
_�|4
�nO=9q����"Ob��ԅh@t��'������"O��b��&I���høH�x���"O�PK�/�P,���U��EP"Ov�vȚ�(����Ҳji�8 �"ON8QЌH���ع�&�rgѹ�"O8!�#M�X�����t��"O$=��%!֬L'ɝܸp3"O��n���H8i�JvJYk""OV� %��+o��q �(�bq��д"O��p�4yH5{E�4�
=�"O!�*V$����G�C�>�Ą�3"O�H��OR�Nτ���@�'#��@{�"O q)d�ڨZ��r��N�V\0"OԄa$���\NX`%�:\�p"O�� �
NN� +��"ʰ��"O�ѻ��%ŢL�D��xJ�@`"OH�P��J�2����%��Du���"O��u�}���H�e�:�:�"O��;�EE����/^>I�z�9r"O���ǁV!J:"9�Dώ_>��B"O��Tn�<:��V�Đ^$6��"OX�¡5	d~�k�b]`��c"O�<Y�FE�b�~qpu/�>4�q"O�TY'�E�K��A���!��i*D"OH�D��<#<�[rH��{�h��"Oڙ@��N�+vtm��g�H ��"O��2i�*��1Q�E"3�I�"Opx����9g����i׈ h��S"O.]cG�,z��=)׉�b	��S`"O L�r�܆�R-*$��-��,�"Ol�֤V~8˖!�7�N9r�"O�*%j�9�l�����*J�"O"T�ΟD�"�+��W�Z�^��"O�8�e-V/ ThɈ �[-'�. j�"O���c	9�Di�4��-,~�՛5"O��$$A�WF�tbգ7vh<�*�"O� X�j�ZR� 5��4 ���`"O�}���A�]Od�3�#�.O~�}�"O�YIPt0!2C@�XL�b"O�]rN>N��=X��/.84,�v"O5#}�Y��-'��"O&݂���4Z�L�0I�n}�)*�"O^�H��ܭF��:cj�p""OĜ��OH�[V��g,�{�����"O*Q`O1;��1!��TՎ��""O��bŅ����΅:���A"Oz�D��>,X$z�GCS��9�"O�[ �&�P��F��N5��"O)i��G�4
IIL�5��� "O~��qn�/[1H�æM
�[lH�"O� nh���~LdQ�w�@�]��{�"OP�`Ҋ	$z�r��D��Vd�(�"Or3���7�,�Z�jAm���J"O@PI�j��"Y��#\�9�4�a�"O������)^���QA�ظ8�"O��F��|��hu	Tnɪ91"O�07(�-0E1EMt����"O@ �uf�N��BQ��/�|X��"O�xgeė@}��CF���?Q�1"O�x3��M����g��Ldp(0B"O8@�/L�d�E:�畗G�`2u"O��D��:��ER�g�)�u[a"Ox9�©0i8�4RÆ�:p�:�c "OX����q��$¶G����@"O��KF)��3�l��2gd��sW"Obɡ��J�br�%��E��|�q"O*q��G@#W�~�u�%O��:E"O.Q�!��!T�Q��5g�(ʷ"OR��3�
�~J���r�OBT�X9a"OB�S��]MD!��F+_@x���"O*x0�Z (*�B�	�7F�!�"OtU�AF8 �a�5-���	x!"O���f��`�����X~$vP
g"O�QZ�KF6GU �Kb��,&"�7K4D��(`�"�����U�'�Ni��3D��H�ъ->�����y~�R2j0D�ܚ�D�*T����d
��i-D����,� ='�!�Nϗ
dH��q�5D�X(t.O�<ԍ)�Κ%�lT��4D��W'�:�2h�Ҫ&3d�E�A*O�l�d$M�U`I�B,pe�ق"Oz\q��9_�J��@�=s�~�
'"OZ�0��C@ډ���\P�� k"O�=r��-g傡1$�T9J�X�"Ovm3�(��	w���/�'8��5 "Ob�G'IuX�a� =
s��j2"Ov��Kҽ����ԙTpNx��"O����\*$B~�isnO( � Y$"O�\�� ��:�(	�5Yޚ92�"O�X��i�M��i��Һ"� J`"O�����Q"*��0҇��!���{$"O���m�.V=�Y�G�X
&n�y�"O�A�/\0o~����W<gj���"O:�S�b�0q�|8y���k�$�ї"Of4*R�_�l�(hi�LB, @�h7"O�k6�J�s-
t���D&Q&"<�`"O��`A;!����
G0f�쁗"O���mOHI*�qF:L���"O1
4Ȝ3k0Aa��ӝxS([�"O��9F�ũ�M࢐0__�Em*D�$`���#}�t}��fC�]F��*��+D���&�>ݢ&@��-X��`1I,D�X��0����D�t@��n%D�,�Q�B�~1�=���@�5�*e�,$D��Xâ��<� h�OI�/�5C�*O�Gi\�J���ʄM�T���A�"OrȂ��� 5yȸ�j�$R�&"O"�Ju(]( �3���1�q��"O*�WꊭwĜ0!Pɛ�2�n�"�"O��e �%z�D(��W�b���"O��5b�/?���Gm_�;��4�e"O�Q���^5(,��BB�O����"Od-	��Q(QȜ�#�fՀ
�	��"O�X�A�{���򤕨q�z� "O� ��a��߫�Y�d��A*$"O^�ʑo �&T�M��,��Ñ"O�]��/#i2&����3و��"O�IÌ�f���*Ow½�d"O�� g�.�Sri	s���"Ob�
7��#����!˓{B5�"O����*$�Ƥ�A�*�ͫD"O��#Pf��X�)F�1 �(�"O,�④ �-jrH��;2���"ON�8T��D��e��-���+�"O��cvj�B_(�@�K��鱣"OPY+%!�E|�<�ďT'u~�0H�"O�4��)G#5�C�M�wf�yjT"O��
���<6�Fc�8'uV�	�"O�8G)C�Z�H��.@6�ik%"O��2f� Q�z��&��X
����"O��c�Wj��0NA'=�D���"O�	E]�X���u��$��pҔ"O\I���X�kc$%�!^*'t��"O���i�-?VR��g�	a �q#�"O�,��E��!���&��00�nqzc"O~4;�"�>
�D�̇�(�"O���LF�ar�Q�x��0�"O��J�gЁ"!�}3E�2z�5B�"O|!����1"��-@<q�L]h�"OE��oƣ%X�tZA���ȹc"O|�5č�Nt���6�){( )�"O��SeЦe��dq���}0 �H�"O��G�'\�t�!� _w��Kf"O�y�g�<�D!z�kX�Y�����"Oƽ`N�8{d�C땁#�z���"O�A���8I��R#����j�"ON1I��\'HP�� `�8Ugn�)�"O�R+B{�$1[ɜU��h7"O��8���kR "fB�g9z���"O@=BO>`�"�0W�*[#\�"O��a �،�Z)
Dʝ(bu�P"Ox���(��To��c���D���!"O�k���i������^�@���"O� ôD�9]�M���%}a�\h"O�r��ϘWXH���-;l��c"OVdy%�R�0E0D��֭]���hW"O@x�ph�_��GC>]� ��"O8AjSN-b�B9i�Ή}�
�ۤ"Op4�Ղ��$����,�:�`g"O�])u�Ӵ~�Є`��*$���0�"OX��F�!Ԑ}_�bU(���y�lʯ?ƀX�d������#�y��� ��*D�ւ�ņ��yϟ<O䀰TK�8
*<�灷�y�ʑ>U{�,.��! ��y�GQCN��J���D���)��y���	xB�3&��Z�ˈ�yN�T�U�%$!<�j�w���y�V�9?��gÄ�:�!�5F�y�kǼK}hpʶ���Z��`3�`߱�yr��̦��3��3�zI����"�y��$�z��5h�*r��(�@`¸�y��H.rl��$
0�"�H�lɶ�y�#G'Y�0�T������S�W.�yB$��1I���/�n,��a��y2�!��`����y'M��y� B4����N���*W���yR�ğr�<��ឡq ���)W��y
� ��6�I���@����Ҕ�"O��P��X����3Y`�l5r"Op\�"gD�%Q����ًTz�H G"O�����I='���׀U�NE�UY�"O��ړ`�������@�^4>�@g"O�ݓ��Q?��}�+ݻ4
�Q"OT��',�E4�q�Kϐ*��w}�ȓ.Gv�St(U=GWd�g^>Jb��2�Cp�Ƚ(Uv�J0O��H#D��ȓa�fܲ%��&-:e3c��?+�P݅ȓn���Ee��Po<��RH�r�ͅ�;m����	�dLp��ޏ/��p��Y�(�A���
��	��I�'vr���rٮ��S�J\��R9r��������L��	� �<���ȓg�, 0Ä67��0�ẽ�B��L�ȓh|�P�#��U���`%
�0�Z��ȓ����͗#O��ru	Ǆ>Ť�ȓU@̂2��`ڨ��(E=vg���9��㕦Z�r�ؙU���t��iƼUå�ͱHt����gG�H���ȓhid��w��ml����ԏjPpĆȓ�fQy���_�F8;�aیF��a�ȓto̙����*x�~�r�E-pZ�8�ȓ)����MƦve:�Jӈ�/ͨ	��{����WN��dU(�0KR.sF��.4z�gA5~N�i��L��D�ȓTҊ̠�ǘ�;-x)3�
)G��|�ȓo��@8ak��-����Mo�A�ȓw�ZL;��Z\����u��"�p��o&���g���t��;�&ɝj�40�ȓ0ְ��k:h�@�Kқk�h��{G�� H^4D�,����6E�y�ȓg��q��	�e�4� �N݆ȓL��s�Ƹ���������ń�16��W��1Ň�]�.�ȓ��4#3�Vt��ش�>��ȓc ����b_^��x�ł�TD���o���P0�ڇyit)�Sd���ȓaPa)�D^��q��zuX���)��nŢ�
4��i'd| ���I^<)'̘ �y��'Ɯe�ޔ��[%�p��ƾ(2(���^ê��8�(p
��ڄSt�L�����E�ȓ:�<=��M?U������ȓN,0��A��Th�	� �<ą����2�.� �z�U��>aІՄ�S%�:�NX�Ae�� (_�!���7  �D�#��xt��!�9�ȓ
�(-����e"�@�|�ʝ�ȓT�4�fE�#�Va`j#G"x�ȓ��!򯐢i�L f�GB�d��,4�xӖ@��? l���W&t��,�4�I51�bQ�Џ�� ���-��!S���`G�$�0��<9�G�!>B*�b�zD��"]`�<!ê� \hK�� ���(�j�W�<�2mة�Jiy��a��d�	R�<	�#ݔ�2�����I�4�PW�<t ��:�v���bQy0��d�T�<�r��6K���F�c8��e.QQ�<�%(Y�f��5S�D�V`�r�D�<Q(^� �Ȩ����V��)Ys�j�<���d�xvNX*5���8V�f�<� ]�3-��XHɁ`kFx,.�pC"O�kf�������]<Xbى�"O\غ�o�<m?�`ȷNNZ�Vt�`"O����0 ��R��1���"�"O*]a	Rj��(aW耖X�,�"O&m��o��K��;��14LT�3�|��'���bC<�F�H�jG�L��	�'^&���g�cJ>t:��Bl��K	�'+�e�!��<%C�+g�])4ώm	�'	�u��t�tV�,|��)%�.D�p��bȨ��<�1����|�G�!D�ı���h���1� 	��*,D�x��n�~.(�;卜�Pa��)�e�<I����9S�e��E 5���gbޔ9TB��T>���EA��I�$皔�C�I/Y�%qdd��/ـu�#L՟Qg�C�I�l�h��P,ŝ#�tZ֋�06N�B�	  �b�B��-����Fb[�V!�B�	�D���o� �U�#i�Z�B�ɉ%#F<��읚)It8ը
��B䉨\�J@@4[����r�ɷt|B�	�kT�l*��V�)�!�4n�tCXB�I�yz����5o	���b��e�TB�	�*R�K�	Ì'��&�S4@��B�I�~
d����5p�0���`��B�	
Fa�Ay�b�?Q_�|��צ>�B�ɏR��D�ƆQ8B��Ȱ%�`���䓦h���U	c\�؃҈�G�T��鋁*�!�5yZ4�æϋ7�}�F�J�w{!�$��al�d��{����?k!��]�t�t/����s���]Q!��N���!P	�4ՙ�ꀡmM!�d����%~�ؐ�*E�W�h�	
�'8֤�G�i/�0�Q�/R������hO?�ՅI�/{��2T�k�U��}�<�2�N��0�f��U�Z12�m�~�<�1�[9?�ԛah��}͜E����y�<A�F
�Y}t��3
0yb-iTiy�<�DFH�!vx92 �M�9����QLJ^�<9T�۩pzl)��L]3X�l,�fg�t�<�ǃ��o<�Ҁ)�/H	���	Xxy�|B�����ɠ<!|��U`J!ڨ���%D�tq,��p%
�x�iH�c�̘��7D�(��ڞߞy��`S�N�^Đv�1D���unҏ~���Q��cTJ�� 3D�@�A��]�bE��]>D@�B�+D�(�%h�
Q+:����	�
 ��o>D��x�ڳnjR,�cLZ@�i�Q�=D�� !Ǔ�|h�l:s�?>�d U'?D�0� GJ�o���GNS�r̠sN D���"F��"����VF��+��y���tR�ISVB��j@i��^�y"гuF�p� l��$��j�9D�|r
�
\Quj݄Y�UH�1D�  ��Ń�������4�Efϣ<�M>����OLE[�� J19@O�
��D�`"O�����@ae�j�(��\�5�t"O���#@�Wq�2�O�m���rV"O�BrD�rGHI����5�`�e"O���#IAhc���b�ZȨ�"O�tß��	`�ҾM���"O�u�@�Zm8��6H�8��=��"O��v�^��q���8/����D"OՑvE�j� =q�S(KJ�K1"O� |Ԁ4i+/���Gj@�I�!{�"OA)�`�/)��]�i\ d��pQ"Ob�"�� T�0i�ꟽh�J��"Oڸ&���}nl��) a��u!C"Oj��1X=�h�%�= �̈�"O�p�u
��)odA{��L����Q"O0��ġ�p}!d)�o����"O,�w��
5x�J&.F3j��d�D"Oy�3�.l�aQ��Bb���ѧ"Obe����&󶵙��5^:��Z�"Op�:��P��Y`+CD͠i�"O�x#� ��`8��Duά�#"O��;��<.vH+Wn�2X�"�"O�J��p�ʽ�Vm��C�XR"Ot(B�۵75~I�Չc[TA��"O��Bu�̿���c����)R��@#"O�xk�#�8	 }�r�֞t����"Od�g[1)�n�`@/��	��"OMJ7�\�e�8a��#�#�RU�"Or=5�F�E���spA�+�4$ct"O��P,ә ��� [�jܪl�"Ob�k#��{f��i�h��."�`��"O�M��B��]��%R�D�#8��"O&���Z�~�D��Ӆ��p@��"O�Փj_7��P�6#9� �j�"O6!x�AB�)��`��_�6z�y�"On%
�C��c5lD�R`!���J�"O��(B�JD�2qN޲9�z���"O����,q�	񍇺$	QQ�"O|�(��?`$�݂�VI�>t�""O��s&ڕ*�|+4�D1O�h�r"O�I��̱E~�Y"P�[���"O"����E�)�0�㗣N'��"ONa���в@ <,�C��z>x�A"OJ�#0A�TY��U�]$uճ�"O0@#�� {�N��b�K<�YA�"O���������˶1 z� S"O�Cc���1�����w��q�"O����,y>E���.� ��"O����j�%���D��"�p���"O�p�G�׻ZJ�dA��%GV��y�%�,��0/D*�1�⥆�y�X�bp����ز@͒�S!E��y"�]$g��P�
�-���D6�y�nL��� F�J{����N>�y�kV�%5�`PQiT#x�� �dN��y�gߠ9�L��B�T��  ��kW�yZJv�s1	g���,EYr�{��=D���2��g���҉(y���BD�:T�,؆&Tm�r�J�`Z�Z���"O(���G� 6k�AS�ȉ�#��!T"O�頦�1o�u0�팄����"O���`hƞx\6����(p��q�"O�$SV�M,�a�KZ�>&�,��"O�jPb��ȼ@Ŋ�����"O�@2�Q�+:0� �6 ���0"O
L��Û�0V�RS��{�zE"O�!�!]$i�,��dg���  "O��@�F�<�֡1t��t�~�ѳ"OАH&T�E�FԙucR� �J�"O2��"�HtѸ!(@�� 8�P"O���Ŏ�'肴���W޸b�"O4B��8V�0V�Ow�JQQ�"O�xBvO�%C�r�8�L8���!�"O� ����Ş�x$�(��K�B���b�"O��PW�F�k��ԭQ!� (�"OFP��JX) �1͝*
�����"O��`��o�0�B�� �b�� "Ov��F�sVf\�r͆�hb��h "O�8Rc���r�ڱ?`ȸ�"O��Z2
H?Xw>�A,I1x�X �"O\�a�Ǐq��aQ-`� ���"O�\a����l+���b���=�쬲#"O"�(d��C��@t��!)��Uʃ"O��/��"h���E@��L��"O�*Qi�6[Ѭ�P��e�\D%"O.�n�e؜Ѩ�@V���j'�>D�� �q�����3SР���8D��A��T�X��l̴n
���4�5D��a��O�H�<!�e_�-o4@�� 6D��9֧��!���+�d�#Jc�3L8D�������l:���8i�Ȼa�4D��Y�E��l$8�:U�
9Iȴ��+0D����ʝ�v^��h�.��{��,��n"D��Z%�ȻT��C��8m�J���c!D�t�6�ǂvL���?:	�e=D��hP��$|�@���A,�� .D����� )`���!`j,�
�3�+D��"E��V�Д ̮w
���"d(D���6�6zH&i��ʓ5:���&D�p(�	׀F0�aĢۏt�.r�&D��k l�.,3|T���VH��K�	&D����'��-�ֽC�-ײD��A	��'D�̰�)��p��lT�$���h��1D��A6C�"�������!��O1D� �'�:D�p��ӯJ30�P��<D������v�F�{�
�5fts�F9D��X�Pz\ ���j�6
�*4҅�3D�y&��V;|�xCbI) 3xbp>D��K1H���Jj����7D����ގC�H��OG'}�R�B5D���2$�%��"#H��;o���t"!D�0i!lœl"D,����9knxd�>D���4��
:��ep�C���>D�� cO�{+�lg�L-w���J��;D���iՀ<p�1�i�,]?d`w�>D�X�pl��o��Q2e��	�b}��E>D���Gm��,T5��P �X���;D�H���֛<���C��@�.=�7�;D����醍r ��#�Òc)�䉅E9D���K�8R�a�9'_���G9D� a�ŝ�@,�#1L[=:)���4D��'_���
C]:>s���P�/D��Y�'�21��!�z�
1��,D� d%��}J  �7"]-����b'*D������	�ʼ�V��P�l�4D���F#���&�ڗ�M�}�ެ��1D����A�1`�Hc��	O�����-D�:V`�fHވ`�@�2<� ��#�+D�|�g��'|��qvB�5:vRIc��-D��cʁW�����
�S�$�[D�?D��y���vk� �L�S#عc �0D�3&��,>:$��4E	,(q��R�.D�����]��Z��ꆉt �Eñ�-D��
P�E����SÄ# d�����%D�db�my)H�O��C%��#j#T+!򄗥�1����5< TPy&B�!E!��׹{!f]i�K��G����!�d3!�� ��x��͙[=�PȢfˀ߸�"�"OH0k��#��9B��31���3"O�:�`�>�@��h�_�=KT"O°�&)�Nk����h�ve�h�s"O�L�s��d���F�Zc �i�"O2��T$�4R�F��P ϝ�@=�A"O�a��	!��0�'�@��d"O�bt�B)4�(�2��$V U��"O�`8����4w`|�rʁq!�w"OPy� �<- y�H�g3xMa�"O\��˄($�(Њ�'ƈ�V\�T"O\�ag�vP���K�A�h���"OP!FXX,��ԭ%����"OP�Z�n�"7~���S���@����f"O���l԰"���3օT���5r"O�����EXC`����j�$�Q"O�����+����gF�h�4�C$"Oƥc[�9yؼJ5�Bۈ�{�"Od��ǯXte��sd�&ʆ�a�"O8�N
6���s�
��h��"O�H1��<�D��H�HϾY��"O6UH�����
���0�,�3�"O���j��MqC���\�`r�"O�m�3�;�F�뗆�?+q��"O�	W�
1V$�ȀE1b�"O��4K" �N�k��zjfa�3"O0�e��Y����4�J:T4���"O�1���ŕK��Xǆ��F;����"O8(�B/X-���W\.:��b"O��D W�cM��ήC 4(A"O L����i��R#�m�ƕ�T"O�0G� oP���fY%L��,ѡ"O^EhT�˒Ij���$ڲ<�"O���5���)N�"0�P/�Z�(�"O Pk�зf��hZCh��{��Ȁ!"O��U,?y}d�
��C M�� �"Oj`��͗<��t�`B��ﲨ�p"O���#LҽX����AbDk�zL�"O�]�� �d\E��`�	8��AP"O&`�Q��$I
�R7)^A��:�"O��G^��N���˳��@�"O�I�Sj<F��I�&g�v�Dݑ�"O����H�$,�|0#���'~���s�"O��Q�n^ m�5�I_�fUҳ"O�����3v�Ģ��Ľyzt�C�"Oh����'T�+#�O)1��"Ojq W!����U���96���"O���׌����h6GE4D��2E"O�Ey�9`�)"�d�ICʖ!�!�$��y!6	sw�*U�T�A���:i!�B(4$jiq��-p$�\J�-���!��ŁZ�.@��S��Q�O@�!򄌁nĘ!b�$/ T��׀4!�).:p�P�B8<��(�( K!��J�y*p]�s*�5�T� gI�7�!�? �U�ܢV�<��ƅԍv|!���G~(H!��q�ƀ*0�"Ud!��['+���bC	�f�3���)W!�dX51b��Z�◅�hq���Rq=!�dޙ7#����g�E����3"OhD��l
�#�� bś=uE���"OLi�EIФ;
\y�  X ��"O��y���Q�<��Ud��L�Y"O���'ŝUL����13D"�a3"O� ԰{�
��\�]����>ST	W"O�i�$�����ڢ�����g"OH��Ā/>� d��"�;^.P�e"OB���Ɏ{h�
�A��P�es"OvP��hW-$ٲ%��:X�c�"O�(�̊N6Q��7bTT���"O*(�Rm�M~i�B.�#=�|U('"OP����4$�As,�_� �"O�h���3q+�4�'��I0�"O���!�	;*����[�k*u:�"O��GlS1X�8�au�9A �ٷ"OH]�CM	1Q�h	�!�/<���"O���ҊJ6�TqT�լ	_���v"O�[�ĝ�Is�J��ĺ^IL<R"O�Y� ��D��i������lR"O4�:D
U���	Ȓ�θ/~B\p�"O*\aЩ�7��L ��=[�aS�"O�%(t�֑)9NH��Րb�xE��"O��	`@��$��,�p8S"O�t���۩7�����5u"�(�"O� Q�J/L�`�*�D0��"O��XT���q�Z�0 �l3�9��"O�xW嘶��P�3� � ̙�C"O*�i���BO�t:���xp�x:C"O$�Sd�Ӯ/ʔ��KO� RD$#6"OD��2,�0�FJ�J�A�!�>9��pw쟛o��A��`O�D�!��b����d避]�a��ϟ�!�$U�kT.(@դ#X�*Ĳe�']�!��Ń~��V��?��@
�.̌4m!�&�и7D,{w�y��l�^=!��	1:ԪhPB ct����K3*!�I�}�ԕ#��Ks�a��͚�F?!�d�aЂ%8��ݵ`8BIqNP�A�!��T���ᡊ~RM����	4�!򤇗��!x��V���𦔦b�!�ą��D$�S@B4Nb*eZ�K؁L!��L�v��m&��s�Z�P!��U�U�K\�[T�]���d!��2#6 {P�J�dh��	�(ɤa!�$�%~��k+۞j[�{	B�E�!��$.x)p
F���h����+�!���q}���r,F�"W���نȓ��a���-D�����R "�"O�<s"��CS6����:�麔"OJ`I^L��yk@h��F~��"O`���=Ԁ9��H_��h�"Odh12
O�?��X�VA =>�����"O���@[� J=�F`[?�ţ�"O��`��l��ؙ�HԴpݩ"Oz)�$�t3ĐI�Fǂ�t��"O��ʇ"mV-R�E����ɶ"O�}"��J��E���7]�� s"O��x�K��.x$s�L��ĵ�"OH�î�9M�jE[����]��5ʒ"O�A�W?(�1!&�
6�ҁ�P"O�tzW�!;�l,�Ċ��x580"O���Ó�;�(`!��P�_�9 �"O�b߼A�`I2��*�r)�w"O~d��V�9��.�r����"OT9���C�/TvԘ$��$�p�"OY0®�&�B�`�MM0pp�"O�j�Ӑ��]����7���"O��)$�[O��:`Z����Ѡ"O� �}�'��G��/�@P "O¤�F��!;*��֮��\6�x�"O�8�"F���}�M��	S��P"OH���E�H{eꙃ'~ɊS"O8e�MͺF�K� K������y� ڢ8�T�P��B'HC 䛰%N:�yaƳQ������X�8��M��e���y�տ�:��kC*��bjH%�y҈��+{0Xs)�P>@HzŃE��y���`{���S��#BEp\�s#���y���
r�����b�\��S�Ў�y��۰h��%�f�S!^^Z#g��y2
�
bt}���M	edJ��"���y.L-M[:X*#h�,_�\�ڡ�F��y�`�"V;B)���c�1��oԘ�y�B�,(d��K��[��*v�S��y2�Z#4_�]�hϲD�lQ�@@2�y�x�|U�󭎉;�2ԲG熥�y����& ��D(��0�@ܐ�E&�y��VP)9u`�7'D:�Y' ��y��^5�~�qvgι��������yz���Ƥ�L��2d��y���r�4D�=������yR Ti�8Kr)ƀk�.4�`f��y"�U��@I0 �i�d��- ��y�@Ǖk>`p�$�\a�*�9�A��yV94�LL ��U�[�2I����y�gB&tkla�qb؀W{6\8�Z�y��|ε�%g��N�|)ӣ�E�yR!�!T8]�%��Fe�9 ��y��+b���,�Bjp���y�.G;J޾HQSꋱ=����S+�y"�J�:$��*�+.R ���+��y򯝀(�F`��.��qE��ѯ���y�ʏKY,T��kǮ8���۵��*D��
��ڀ���j1�xaV1:E#D��ѡe^%���3O����s�� D���D/ �:�,Q��!���L=p!�dΐ)9��B�kGS��7�]/a!!�dP.u��{�IL�yC"��X�?o!�[#�tAW�
$�4�Q�-��QU!�5Y�r��	Q����1�9:M!�$�����
� �/cZ��0�J˅#�!�$5u8�0�k�fNt��#B�go!򄎯|�Α�IܥWD�lA�_�n�!���5�>�`�*Ԅk4�JR�2�!��U�Sm�rP�Ť{,Lٰv�V�Q�!��(I~�9�B(���r�
�[B!�$�	ȴ@�;I�h��� �Py"�9c�l̙�OC.i�jfI�y\[D�R@º�d٨��V��yR�'���C!Ⴂ
�b1@U�F��yrC���ɐ��Ҍ��T������y2JC#`����dMy�0 �1�:�y��|n�!��H��2)s�<�y�i�Q���b�)U�bY*#Л�yrk��) ayrK�>wF,�%�F�y�D�0��X��5=.X�%+�
�yR#߮�$��8X�5�t]�yR�O,��=���*��l�!C�<��?y�'4��	��
Q�X����S5H�����')�!�)�gڮ$��a�G���`�'aRf�*��-ػ9�L��G��yRbu��P(k�����1�y
� ,!�,Y���˔#A�%�#�"O���� S��� X�%A�,��"O��7�Ҵd1�A w��3"��Xg"O���G�CU�-�2��7��y3"O�m�J�F�@"����s��U"O@��#�S7) ��Q��^�9+ "O\
R�)�"�8��26�����"O�<��h��z *�,��3tV�yҀV�NFt}�P��WHN�����yB�O�{P�m`B���O$�s�Ҍ�y������H뒎��θ��n��y"nO0'���чf
�1��1�y�Hƒ0�$,dC+x]d�c`jT��y"�@Gd��	D����Z0@��A��y2g�Ȁ���0,���K#�yb�Ǒ0�ʴ*�BΊy��L	g�[�y�"E1���*�
�`$���!��y���w�bU�S�n0h=0CBǥ�y�/^�4`��J�g�(���gޘ�y���:@����!��/�r5��KV��y�a��l�₝n~�٤	��yҌ�+�[D��.u���梙��yR.��^�֜S���Id� fᓠ�y�b��v���"U�Gqb�P���yr*��v��0ru V�p�D�4+I�yB�ΛaX�%����Ri��24��y�L^� A���b]9K��P���y��V2m��Y��E��(��yRg,o�)�VfR�:yvY��ƕ��y2���y�"�Kf+�0�����M��y�d�Ep4�Д�'R�0Q����y���*F��#�عQ��ۆ���y"�B�b�\-�� רw�@��m?�y2	�&G��:�����+ۇ�y��=+�y�_{98QiR�
�yRd�{	�ie�W�b�x�!!�L'�ymX�g?��;�n��` ��!q ��yR�A(1_��c�۷_��g���yBiϋX�, �&�8$�$��fL��yr�R�j̼��Q��ܑIn��y�',�1��
	ǆX�� �yB�
���)CO��:�(��L��y��߾sN��Q��S �f�qC���y����sJfš��T
�)�pmB��y�g�-T����ǈC�R�6l��O�8�HO:���|P��#u-H�C�����)-m!�^��"P6� ������!��^���,��EM���Dj��*Y!��P� �`���7d�p��>7�!򤔜q��i�s$�V�i*d�*}�!�$K�,�(������g&������l�!��.]���d؝��H1/ !� .�zc�f-*cFp��!��+m��5ڕ�U*NL9#6F��$!�ĉ*[��#s����Q!��? �!�Ѕ1ִ ��",��z�`�v�!���Fdpk�	�b$ږ~�!�$Ċ�% "%ҵc֘;�K�C�!��#-hU��͕9J:\Ѓ��(�!�X98P�D�rPj�nʃ
��C�0P��iEH�!��𺣌�B�C�	�,oNq!��@�,M^PA�C�a7~C�I<#��%jV&�>����;T�C�	�!D:Ab��w��4ʰ����C�)� ^��1GF�Ě����u���B"OV`{��x�X�@1����Aq���T8��2E�ʱ*y�)x���"(�"�7D��I��ǎSʄ�f�^B/�$�f�3D�D��Jy���'ő�I�d��0D�PS�ͦ={8��)\�P8R�-D��q�a�jU��C5eǔjR|(��f,D��A2��[-f)��!�&o��a@�(D�@��d�(�>��3��!B��#�j4D��Q�X�M�@aq�kU�F�ht�4D�<���Ν��{6CS�F_*��i3D��s���\�؀��/�����2D��P��P�F��P�a��驥g/D�<��0g�t|���H[����W*D�kR��
g���J�� �	��A'D�x�i��^�"pcD�I��qqR�&D�p�Aj�� 6����aVU�z�x��#D��bC�΢ ޡ)�e��r�B��!D�\�UCÊD�`@�tjڬP��:&g!D�4AkH�^ F�h �׉IpB%�a�!D��[���a��囵��.
)�2D�L�q��+gL�Ӡ��{_��ȅ�%D��h�ρ���c��P�g��<H5$ D�L���� _����JҷC�T���9D����,U����df#z�����6D��	4MT�QKGhA�!x��20�!D���"#Ԏ���@�F��YE2ep��>D�D��O�l9(4['ʑ�T"��z�0D���"k�"~�բ%T�%��k$9D� #��ʓ����B�3�CI1D�ذ�j��3k��M,8�>(��/D�ܚĮ�,P\=�CC�#(6BDꆄ-D��)�)�Q>0U��*�쉓�.D��I��L�4p�AR7���,D���U��~੣�7��*�-D���¥�J��`���OO�H��@0D�[R�-��0�%�x3��.D����R 8$<��jF4W�y
�)!D��	E�[�0��C����QB D�\��-C�&�ɡ#o�����D�<D���t��B��!��mf���"9D�(ad&~Z�yC.B�"b�p&5D��S�b<��J�'X�200�7D� ӑa=KlܤYu�4���qc�4D�\A�‸���G#�%���a1D��1aN�eؽ�U���]Ժ���+D���S��?�Е���7r�l4��)D��6nR ��q�AO�-5�  +;D����!�t��"�.�Խ�$�8D�|� 
]E����Eڢ�`�b8D������h�E&�'@�6�YF3D�XSm�"dbI6k��[�2�ڤ/2D����cW$�Z9��/>y��LB��0D�\8鍳`:���!�B�R�8�M-D���A'�l�A�� x�-D�Л4�S��mSVm�+�4��6�,D�0��
OT�m��Vi+D� )�(�+��1Ӡ�U�]�6UaB�3D���v̅i��Ip�U��H��@�0D��ٴ�Y�huxeǎ�?/�9k�)D���t��_�(]�Ŋ��<|���e+D�,� g�'\i��ʱ�60@$�RB>D��� Z�6�~t�!HB�(�2�jw<D���-A��Cu}<`�<LO��pfL99�0H�.�'of� ^y"&)_!�<C@7��	�T"O@"PeǏf��ڳ&C9ME��"O��@!b��9,��ů��}$���"O�� m�p�`QiS��s3M�"O���q��:+O�M�u�	:Բ��Q"OP!��O9n�ĉ1%m0i)K��y"B��-�AB�!�
f+ 8@�M��y�.�p$:���Z8is�E��y���/v�y�Qe��U�䱋�E� �y�Ƈ�.�T�#�@R�TRa,���yү��5�-j��K'(3��Q�-�y�ں�1� -]qK��g���yb��1�u��(q� �ǯ�yR	A:W�Bu�O�`�J��5B��yb�J�,��F�5[��pY�/�yRm���"6�V�E� ��Q����y�%����%��<��1�Ľ�y�TJ+�� u�Ҥ="�AY��� �y��ݛMu�8��?$"=+��C&�y2'�)j���g�'Gqj��1�ч�y�)����o�1q���@ņ��yrԙXu����c�6+1�� @4�y��Ƴ2��,� B�+$e�5Pcԅ�y�+�-��9��.ޟ �<=��*�y
�����ٳɴ`9(-G���y�"A�4�jِS�ՠ�\]CC J�yFJ�*D-0�d�zg��I#)��yr�I��eꥯB�@[�ˑGצ�y"H���=���;>�dl�����y�dW�w8(;��14ĈlЃM�4�y�ԕ~J���D'K3S�h�I�٩�yҦ�:/���bp�^"A�d�'��yo��B����2�ڄW�2�#r�yB�_�c�Z!��F}<TP�b@��y��ކ1ڔ��&/�m�PmX�Ƥ�y���"OGR�Ҡ�\9X��Q��-B�y�LCk{��8�o�&d?�$t���y"c_�8�.`�D�n!�>>@��3
�'o@MRӠq!1E\�:p��1�
���y�B@0)L��o<5�d��r��9�y���1q�yS�KP��@��i�+�y�ŝ�)h�pk��DO/, ����y��-T<�G�]�I7�#W�X��yr��
ll����M�Hd���O#�y"�4�	R�&]6b���v! �y�h0\�B/_8)[��N��y(F\��D��#xɡq���y��%��)�Q�4�89p�@ض�yRDB �� �0d #;z��!�ڦ�y�@<�-��B��b 윪�E�y��)�r�I��X �(� [�!�^�&B���!�
[�"pp�� E!�$�]���P� %��%(��1!���?V�\�r���*��D�F�ҷ>�!�DV%"O���p��%�n0���$a�!�d�-�*�e��e��5�r�\�D�!�$�>(`�X�hӫY��]Zu�N�`�!�$�9ojU`�M�(�hPZ��˳>�!��L9&� �1f��Q'K	E�T��'��Q�0��3z�sfo7,�u!�'�f,�F)8�� +%�Y)/	v���'���E�;���D`	 	���'h�d�Q�=v�,�Ȧ�IL�~�J�'>.��c�}o��HF:\d� 
��� �P�P���_����U�`j4̲T"Oz9��B��v��@"��/�ֽ!#"Ǫ��i�g QCǗ+�⑹F"O|�ue�ϲa��h�-K{,��"O��o�5 ��9P�PK�l+�L;D�\����P\V�
�ʈ� ,��Rb
6D�,+U��t����a�*��M��5D�l�	N.6, �Cp+��0� �"a2��<)�A	g҅���L8^xbL�1,�d�<)�ǰkh�'�W��`2���x���"[�<�$��h+Z!����0=�"C�N��j��V�g<��͍��y"S(@�:��b��^�&9��GA���'�ўb>%�w��5E@@��e����Y��&D��0�@<*`mia$�ٰU�p�%���<a�L1G�<� �6p"��Z'm�D�<�3��2u��0�o��j�����y�<y��Z�>�tx���®;�Yca�p�<��̐j\����X��Uv�<Q�#Q�D�pP[� ��P�Չ�H�<��3B{��	�-�^v�Tb��J�<9�,+� J�)ޭ8L�	�'�~�<af
��&��(بZ�,�����t�<A���f���S0�@/A�,@:�Y_�<�D����Uۣ	@?~Y"�K3��g�<�A�͌c�n�9�lJ�!�bቑ$Ma�<aC��$REd�B@ġ@�܃�
]^�<q��ǲX����CR5���T�<Y�?bά���MD�p�ɒ�_�<Q�.�_01+��A�{<��kg�A�<��h��(�8\s�B�I&H5j'NCG�<9�C�=gp��ܐ>��	[��h?)���-ް>�q�H�x:��I7�ݗQ�>�Y$ Ig���I�K��fZ�a@��8`(uE��!�ɣ���s�`�=ۀԅ!�������DQ?��ɞz,��z5����8 7D�l�u/	�}"���_�x J��'\z�3���I�S��y�KG5!�
� �gْ$���e� �y��:p]d�������'.��y�E��k$"���I\��4���\)ՀəK|����
(K�H��'U����W5G�r��d�
����'XH��ϚE>��C��W�stx%!��ė0[L"�V�{�R8c�+�c^��,�W�<�S�`\��eA��>1��
XD�<a2jE�>]0(��쏐c3��5 �D�<���eKRe ��� g�M���@�<���$B���7	C`|C�f�<�B�F�Lڗ*
1~���hO�<Y�
��dsTD��`�CO�' �}�����&�� ���@�{���r�H�(ߞ�"��Q+!�d�@�ɪ(�6����܀:�Y�0�^,�t��u���?�S�>Q�'Ҙ�z�U����j�{J}�<�Bw�l1;ǆ�)��-��@�1o$|aG��QtdX���2	3P���*.A6���n�>._�1z�a�`k���d��.�-��17r\a)��;0xH�eI�O�����FƑOnh<,���=+cʍIS-Ӓ_~�Q$����_z���5Z��ȃR��D네W ��'	�dM&.<EM�(#�D�h�|�ȓd�4�G�T�N������Ї_�&�bv��!x�B��D�޹i? y��̒h�'Bz5��'P�aqc	�.n����߯u��+
�'u��pP�K�y��p��8�:(���S�4�W@0ֽ��K3N�ihes�'ju���
���b�D
Y����)~l�KY�*7tfK�CZ��a0�L2&�`���@IVʺ�C�6�4{2*6�Op�i�h�A'Tm�V��7��I�����v�
�m3b��L�>�0��E�nӠ��v��~��M./��c���l�q�_�y
� <�8c&?M�.a9�n���`�G��
7l�؃D��7�d}`��L�xA>��taP� L'yC�.ς$�d�V�C���#N$U>!�O%��(:�Y9�T�I�MX�2���P�
�A��q��/�aҒ-x#��s�0�8ړ=�6`���_���q�C·�����F�v��EL��E D$�b���A �$�2Q"4,����!�%�S4hrN�ex�`&��DW�(k��˳�}��(?A��Y�d? ��IWj��a8C�K�a��iI�C����i<	�ĢԢޔID@�G�5G!��ܑ"G  �cГ.[nHsG�ܾB�5q��Q57��G�v���s��<��F4u���S�4�}��f]+a�0D��c��ؠ"O�q���ƾ,C,�f'2F��g�an�ӂ�A kzH�i��E�;qT�)V ?/K�=5%ހE㾬���<)%��GM}�$��ŵ$�my��	�;d����/A� �;b�NS�<k�-�#l��q���<1%`I��ɮ8Ѻ�����9����SHľ6���,q�I�G�
yg��Ň�Px@���g^�y��/��0ҷ�Ց9�!y�*��KG"OF5@G�Y�E���s�M��~:\�@�q/��:4Z?�D�C\
B�� d��C^	��.UV}�S��9��Z�ў�!�ă�/Q�U +żA�
,��l+�B�*�ڵ�@�K�������a/�(!�M3p+$�^z�@���>�
Њ �S /����I��-�7`Vt�()1���
�^�� /CZ-�㋸扬�I~,(�KP�AJ�}��U�}!|��B%�R,�h�w������ʔ�P8�6!�Θ�%�VV�\)
l�l�'+8��	�8c��HR� �cM&=��pӌ�j �E"5z���Hc�83G-��*J#��;�ʝ1fj@rܧ@��+ y�P�a�	e�p�2O�/۸\�5b7�p��dA�z+��%胸b���"cͬs�̚�X�^�0���O!/4���A�x.�@9�c1#�F-eR5t�<��",,O0�J6J%h��a��˄+atX��EWd��"��%��<��
��|V�`e�.�O<�3�/_�����(Oh���|�GL�N`��U>��	��{yĈ&>���d��_���F%Ʈ��x�*D�)a�� -�*	*0��oa���H�r�b�! G8%�6�p��A�SLy2��B�"4J!J0 B�sV�R��y¥�)B	rU� �~H
��"+�6e\X �DQ U���$@-.��e[�Dۈ��e"\#I���N���퉠\�R�9�I"v��Q���N�j��E6f˞HiA�?.b��r����6��;~�X�U�U�i�^�Gx"-�x�0E[-%w񟺵�f�0:m�X�c�Ǭ�HUQ�"OEqЧ��6lSl�P��y�q"O���F(+4L�rƜ�}���B0"O ���9<x���Zd��j"O$`�U�7O:��P�1�
Ei4"O"�J�CY4_4@���?�6-	�"O
1#fAΝvS�u�򎂳l?.L�Q�P�b��a'��X�@�"�g~"�Ħ��Ѯ�?����#F��!���4��ycw�̈r��m����!�!�$�K{��aF��4��p!�+s!�Ċr|�ɳG!|�d��dG�t_!��"g��C��J?���`�F;F�!��'8�V�٥�fOT4"���**�!��6�nak��̌D6�Ѓ�&�6!�d	ja� 3�I�$a)B�)A���!�4y_@����N`��I��,j!��^<�<�K��E�zt[���MB!�J78�p3��&`q��H�!�D�S@��"ѯ�t�����k�!�d�F�\%�%oڮKe�����!�$�?�T(���4M_h8��̌�Y�!�
 NQI�)�!3X�k�8!�$�Z�a�4%P6K^r,Z7��U!�dG=w�DM�p	ћ�0\�W��N^!��ģ~�
�J����FqB0��G�OB!�$� '^��9�n\�#|�pIf�YO4!�ē�+FmR���308,��a��;!�$�7Qa�@*��Ӏ"���҄)v!�dA���$kɡa �r�)i!��:�6�ɂ]��"�!'6W!�� �9�$���P����Y.YR"O:0��J�p�rpAHU�x��"O
l��5Y�b�9%�,�F�A�"O�@=1�zl1jI�r�2�X"O*m���B-G���!�Mr�~Lb@"OP	)RJ�0, �X"���nł�	7"O�P ݻ/����G#I{nx��"O��2�)&/xd%���l�� "OʽH�O�04j��@A�0�
r"O�� �B�{�Qz�J*��a�4"O��Ja�b�k��[������"O,2@!�>r�(K��u$�\�G"O
���c�4nD�i6b����"O��螣��8 @�!��hq"O�\IƬI)�|�y�	u��Z�"Oy:����1#�+Sv��6"Ol����_%%�<9�jG����I�"O4-� �u�����r��<AQ"O&8����>
�`kC�U<�U*�"O��2�Fф L���'(��*��Q�t"O��� $DY�l�WꞑŔ(�C"O�(fj��$*a���M4e����"O�0��Ը4�.�X����&�b�zB"O��BS-�%n�"��P
߾!�\Ȫr"OȌ闂�,P�5O��$|�a0"O����3
t cr е	$"O��"@���Q�GME�	��8�B"O���C�Y��-q�Ļa�F��b"O��rp#3jZ�c�/���@Y��"O&�8U�P�t�B�M�w�8�"O��A�,�Y���*� ʋoJe�"O���,��"i؈�B8S�|�B"OZK2ǜ�O��0�D)H�x1y"OP	@��&,��9Uj��	���d"OTasH��Q���^8��t p"OV +T�1��	�Ț+w&��e"O4t���^_�tS�m�/lH��"O��xp�M�4�
��t,��[��0�"OI�A J/^��e��fY��ڨ
�"O�D
��[�q�z�CqO�	�j@"Ox}���3�҉ ���/�Nlہ"O��pӎ_�>���O6��h�"OV�ro��7�H����<x��"OV$rU�_>K?�IPU��n��9�"OBE`�E˖`�Ƒ��/D��H�f"O(uI�/'ߐ4�Ó�g�$E��"O\���1��[�CF�Xɢb"O�QA�؋#2�a��+pn�g"O�ɖ�A�ʤB��@)xp(�V"Ov0�[y�dxCe�Pڰ"O©BB�4��X�$KW-.=���0"O4Qɤ R�*�l�U@ K"��h�"OaL�/��+5H�fv��0�"O�5�c�_�9L��X�I�"O�ň��J25��!�0�H1�R"O<
֥�i-\Y� ��l��I�"O�\����P� K����.�Ct"O�����|^$E �mDCО%�s"OQ�b.W�=c`�i1k��l� }Be"O�����H�/���5�Lc���6"Ofu�E��#�J�[b���F=��d-D�d�f�C�lj8�AD��x�,�H�
)D�yB���q/N��"�]n�}p�#D��S��>�(@��攡m�1˧� D�� bd���-9R����9o��"Ox}#$��?=�Љ���/Ff��"O�l��`J�c������P�*�"O�!����6e�)AG�J%@����"O����"_@ H�lI;���P"O�5V�]�ꌹU���6���U"O�E�A#�>�Zy�c��<��hz�"O"D�d�ϣY�R)��H>���c�"O��¥޲mT�d�	<S��"O&\���U�S��+6������B�"O.�) ,OAל�V/�/?�*"Or�
�-N.k>�T�>�	H�"O �:r�]�LiX�Ц.�4	�5"O�!��>P}@�!̽ �"O*aqע	�R�2h��b�>)j]0�"O�1�'H��9�`L�L�|�Qd"O&]�1E�iW���eY;Z׀t:R"OL8�R/�5����`$R�(�jg"O��c�${���qT�дD���+�"O(�a���#o[�G�ۺiB\l��"O,(B����yKه�ܸ��"O�!@5I�lw��C�$a��EBa"O.�	;�>����
�"O>��lF7U�t��1J�l��C�"O����;< 81���P�J�c�"Ov=���p(B�9xt�%"v"O.�j��5I֌�臍�ftU��'@�9:R(�j2�l���Т�\��'[V���2b$��o�j:����'�a�C�V�T�2�A��ʮm�jA��'�\�ҧѼ"ٸ]Pg$ءrf� �'~�3�A1ת�A(�}�H���'r��Rg�={�NТ��@����'�Jr��#�乐'aӑ?�Q��'��bF�L4�b��Њ1��P��'��ȇL��]9��L/5$Y��'�^���ŏ3p9rw#��F@�
�'�Μ��L�2y�"9��bF~����'[1e��6�>�&L	4�B�'�"�'��8E-	�d�H�'�lU!`��v~"�EDL�L�Y�'�pyr���,
����u)
���#�'���G A!]��t�� F�R���'P 0��4&)��� �E�a�NĂ�'K�;�$Рr,h�\!,���'
�]�Q��lB�L�5��5!2�}��'-D��B�@�j(���V("; �
�'�,#�J��u�~�`E��"@i�h �'w�0[�E��h�zR ������'�v�v+��(�Aj�:�=��'u�T���G�zQ\XXf�B<[q�_j�<I�-��%�x�Fm�;>6Ux��}�<9��jb�Є�ʶ��p���~�<ّK���RD �(�0<���t�Z�<��.��j����Q�H~��VGu�<�2oE�yo����C+��`�I�O�<Q6��K����Ά�(6����]�<1S)f:�;dF;�&�fKX�<�p��!;r\c7��5(�D �E��U�<�mo�2a��DӮo]�D'�W�<鐥��P�"�X�f�,rA@ɡ�S�<�w�Ѡp�씉��I�m{,�1".�O�<Ⴀ��GH�2�L)rv�I�E�<��k�*�:�:�U([5����*�{�<� �!a�ϝ��.Ya���^���"Oh���#Mr��0�H=Nx�� "O��*�%�cx�p�έ`e���"O�3s�ĝe&�����{g���C"Ot()���x �un
�p%"O��d�L2��u)���R�"O�E+��
6w��`�A�Tބ��"O�4 T	^0�6ݳf��"��(q�"O�Q0BH��S�<�E���S!f�W"O�d)�*abT��ϫ{,!p�"O\���'�>uc��BVh���͢&"OE:�Ή�}׀��6�_�F���'#D�����b�H�e�[�4Fdq���4D�`�n^$0D��I�����i�N5D��Ӆ��1$Ad���������Yv`3D���3.a~a8��
�cWd�Qe�?D�Tpe�ئ(�JysV��a� �14"?D��ps�_�q-�4J�- �	���.D��q�f��m�n؁���1tͶA�h,D�أ��O3p��	� �	;nr�IY��>D��Վ�2��`B��fq���*?D�$�0G�¢����["�O�C�I:h��9�E��d����B-�Nv�B�ɤi�4#SK�%-��X:�d�m��B��#d�A���O.�uhV@C��B䉌o<D1�*�!W�Դ�2�=P�C��s�b�H�*l�fu ��8C�I⎩�fk��G�H��b�P�;��B�	%eKT$�aIN�s��z�&DKC�I<�AQ��>%�� ,�(g�B�IO�ڄ�&]7%Ŷ���lV/xxB䉆Q�䅑�mU�\V\l�WeFBB�I�_�F����A4�F��%���>B�I
5xf񰁦�Z0%h�O�7��B�	�_a9�g�JU�w���HB��/`�DC�i��?a�\����9z~nB��,j|4��fN*�l��� T��C�IR��5�K�d�|��T�^�xC䉸1V�ʓ ��s 4���>e�LC�I5��!�h��N�YRiL�vv(C��-p
 �0������/t���T�1D�����:���Zy�`�B&�/D�\�P�ñR��9�7#�d/r`;��-D���\����_�~ņI�łP�ҎB�:�Z�X6W�9ژy�'�"�^C�	'xu�uYu��-,rE����?9��B�I65`eI�gI�qV�	9��S5I��B�I/2�@�&�`���%�J�W�C�I=((Z\��́S+
�§�p��C�ɵ"z�ZC�	� ��3V "
i�C�B��e�š1낍�DR	I�C�I��2�Q��Y
}��ʴ���nC�	�inP���N�&;~�H2�ѵ'�ZC��:e���X��Y�&��i�7�ȯFB�ɗqq�bT���5��0k?�C䉊-A�hB�B��s�D�PK$B�IM�T���n\=A8��7(��C�I�-Q�@ �K{��@�ŢA+�C�iV\+$�Z�Y-<�a���$XV�C�72��l�c��.�R@h����B�	>/Y@�1e�LM/�j��8_�B�ɘa�䌀��P?]u���@�H*��C�	�)r���$&ژ�Ɇ@�����4D�x�椓�@hH !Bq��bCJ4D�� L-3pF)d9*�"� �5UH(��"O~ԒƉ��"���ACNZG��!�"OJ�ziu�0M����y����"O>�:&&S�`rx{QA��e�ŋb"O�Yq�C�ZR�dbT�ә\�P�"O@m;��V�)C���V����C"OBH	v`�6%�V�{�����1"O�I�F���}c���5,�2<S��'ʠ��*�J���÷}��AjrHF�?2��Q��==�؃	�'�����i.ࡠ�[�;���?�I"�MG�ןb-��.�-�|���ϝ!l�� ���P�A]⟒��#�]�3�t"�Y2y���>�T�G2���u���5i�e�D��c-�9���QK�K�B�
⟢}�c��	�Pe��$ �w���C��?N�P��:�p��V:�d��1ϛ�k�4���b��F>���k� K���p΄�Bp� � �.�	�8il�?%?m�acK�
��;ci�8T��u�8}b撐@p�O��d
�m�|�h�9�$�;t>c��O�T�.�)�'q��� �!�Zi�1X"%�|Tj��
Y� �O�?1�7|@
�S�$�Z�,��F�}R�O��?eh�/�sK�`�R��U��!I
"]�p��D0P��9�NG��(�EM?�J ;�3�vP�>�|�U�cY�س�ݍp^q�D�D;���?�p��b�Ęk�"ŇV�b)`���4�k�S�Oy��S��4\�n]���W�z�����E�"��'��O|RE�_Ib���j?T� A!��#�a�T��-x��a�.H���1�ۆ�y��(бC�w}��)��?��E��
D}�ac�6��.��������L"���	�RjDP�S)��~A<O��O�>�c���*L����ǥ|�i[�&Y�fN�ډZw'?�zS3q�]��J�ut�Qئ��+��'��|��( e��24!��=�Н�ϛ+A���ĈߴA��O��QA�$�D��,�� A�b��'DW�<�)4FDXҋO�Zr���]�<�f�
�l����74�$=��a�<)�,�*F���"����>C8#�� Z�<��.J/�T�2�
&3�0�#�R�<��B�oČp�3�UN��m"��R�<q߽:�p��*��S�r�!�DN�<�s9H��J@.ڡj����PA�<���22�j��ghj%k���w�<Y�,���L7�/��Q���Ј�y�MH4.,lI��� �Oᨉ` ���y®�EZ�dSe��tNB`�w.�*�y��p�{��M.o�Z�b̎,�y2�U4D:< ���F�<��@��y���� �W�4�t�� ���ybn�f͌��U�Q�~`�;�*Ӂ�yB�H��,��k��?�PyKB�y2G�3�ȡ#�M�5�KW�3�y��e��԰ �N�c�Z�kg�yR�(!4�%ҵ啙be��#��	��y҈^o,+���V�T�)���y⨁�ir��b��{Τp�R�@�y�C�\�J���w�ޔг�V��yB�ʎqeB�A�Κ!�h�[��G:�y�~�xt�� �m�D�G�y��!8�8��^�1���8��K��yE_�`Б�[#9��|����7�y"�٩:|�K���5/@���F��y2�L�0l��yU��,%h(l	�y"�қ2 �!Y"l<*��Z��F��y�k�+
�+��%$����?�yr���C�qyr/L�rkڅr���
�y�e_&BXc�J�k�@q@�o�y
� �A�Ċۻ#pƥ��F��N�x��T"O�(�T<5f���b� C�ʍ��"O�a�V���O�����C�9�&ٸ�"O����,َ3Qf�93�P��T� "O�m��/�&(1��NK3�ŰF"ON}�V��{4���ț%���BC"O<�ƣ�Dn:�[6H�9^��h��"Oz�h*٦QԘ)B�D V���"OX̹�BE@|����fсvR��g"O.��#,Q �P&�<q��"Ox9y�.j�q�-��*=b���S�y� �+{F�i�-ʴϞ��C��%�y��&^E����k�-�ȣQG��y�6b���Z�E�7iv�qj��y/�P�չ�e��Nt�X#0.��y��P�*(]�G��#MB�Pؗ/�=�yO��e�n�Z=�v������yҮ�.Y���pJ��@����Μ�y*I�>�TaQ�Q�1e�p0!���y��D�`�)q�ғ)I,9���y�D
�xxb�+2��E'��y�Ɔ�β���܈�֩H���y��o��5E�"�
a����%�y������Ю̽��,ئ���yh��찁e� s
 ����ʟ�y�ܜ26΍�$bFq¥㗕�y2/�6�<*uHtL8P�)�y��к,��J�A'{��l8�*��y�ͳ܆�8$�K^΅���Q9�y2'� ,'�|���B1z��a��y2,>r��N((�!q	��y�m�xil����?7U�ߛ�yN�U���A�6�tb�f��y⋑y���:`�:��L��#A3�y��"�DYvmC0T~�GD��yb_,$�����!N�)&�5�'���y$J�r2�\��䒢icj�KB�Y2�ya�'~#�\9a`E�[�����̵�y�� �l���NB́���%�y�/H�&L�8��2L&����F���yr�ݬnzR�"���3Z~TR7���y"�X�y�t,Zb)�z��e�֬S�y��I3p�В/_�)����N/�y�+\��"$��J0!]��5�O
�yB�����Ɗ÷f@�bա]��ybAY7��ۓ��(����n�t�<Y6� ��W�]	� �1�A^N�<��aR}�q!�)ۈ	�d�����H�<��GH5SD��;�J�J���t�}�<Yւ�	�ƴcv��1
��FUz�<1��ҿTU�0���a!��2bf�u�<��Ipɚ(�k�;TXb���K�<��O��
U�|�P*�]�5��
D�<���>������З!�����Xh�<��a>P����mZ�ΔY���e�<f�	�l���GS��лr[Z�<��H�w]��S�`�S���4JZ�<�D��y�6E��,�/�d��@VR�<!�+i�h(���-+~iZ���d�<	����Eh1��lHH�f=��,^L�<�3�I�'8�c�h� ������]b�<Qiö$u�4�1��2L����g�H�<�F�hGrI�q�Y0^j| �g�O�<���Z��� �rz�4��`�<� @\���SE�Ft;C�X�sF�ݫ�"Ox�8�j_�ɣ5���
?��c"O��C��N�0��G�>.�M�p"O��K'C"�\�@F�9B��Y�"O��ۖg�H<�#GcV6�X0c"O��Y���ir@&���H1"O���Ȉ�@Lb9 ��^Wx���0"O���2�3�仡��JH��i"O�ؓS��s�1�ҫǷQ(���3"Ojٛ�JV0���T��2X2���"O��7"R�Y���P�9A��h"Od��.|"�P���j��y"O��7..WL���rnO�j<$���"O��+�,�+	��	��"F~4~m��"On�2� �a�B�ӣ.'f���"O�Pz��S�C)�ţ�v���W"O�Ђ�'�V�H�[�.��pS"O����o�( �5h��ǈ=�N��"Oh�xS�2lf�:A+��y��"O8�yED:h�8���P�g�A �"O����/u���Ic��e����"O���vo��$�xh��j�:�a�W"O�R�-1o�X�%'65���"O��K�D���٥ޣ<��)J "O����dTFG,�S@��^�p�0"O� cX�[�`j���I��\��'[�A�ɖ����`� \r�	�'�<�z�$�'W��q#����r��'��,�#�N	�R�*T�Q�'�ft����Hv�$�1�ěyC>1�
�'(p��g�M�V3fQ�@OI�<�!)
�'$�xaK˲Eob���ś���	�'�^�Ѕaϕa�޽��n[~~�PP
�'J>�)��S�VXI��ȥr��l��'˜|h��3\��(�E��k�%)�'UK��ܙ��3Eր��Td�<aww��(cCH	��c�!Y��X�
�'�x3VÐ*�����bś\��	�'\�X��=Mk�$�@���Pބ�`�'6�� #�w�����̓uD�#
�'7@q!ϗi�|rg�6q.�EQ�'/>	r��� )�5�6�.l��J�'ݾ�PCi�b�P��/-)&�CK<�	�L贉��&Hp
� cU�B�@4�ȓnުu���ԉ9��� ��4�@����z��֙"0 X��ʒ��Ȅ�̢T�D��(S��4�_�`)0��ȓ?}$L�4N���P��*綰�ȓ=�x��
V%�0�i�A�)$|>Ԅ�`�JD��#Ĳv$���aƤa�T�ȓP��8�%��4)/U3�@�6J�h!�ȓI�8ppӂ��B���b�f5O\��m&�E(V"����Ҁ(0J�=��K�TɄ'�GdDӧ`�=����ȓw��i@C#R��0{a�AK"D�P(N:o���hA�׭YoV���@ D��!�5�؂sc�#��Ai;D���2F_�TB�tR"mբ!i����8D���6�J�	�$Ԑ� ��-���6D����J�S��$��c����p�5D�� �!�rא{v(�V�@�4D�,���;�����C)M�4�1D�T8��KB�~B���G��`���+D�؂Q��9��r�n�p9��(D��  u�vK&*:Z4K�75��)JC"O�1J���p ~]�����""O1��}�`��@�@D�	�"O�)D�!X'��R)W,�$Y�"O�����;L�ܑh^ W��0"O��"�Z&/��)�aD�
x.�ʡ"O��i��� �Z��M]tLd�p"O4hd��/<�F�k�� e\≘�"O�M����4X|	Pb�9*���z&"O�٘���R������U�ء'"O�Ar�A	5^�y:�[x�"-��"O�0�d4Jo4�P�b d1�Lu"Of�c�u��QӋ�,
"��[�"O�Q�EW3����)
,5n�pz�"O���GŖ�w��9�EW�P"O�y�O�M�^�q�eS��dQ�"O��#%�mcDA�㣐��ؼ"T"O>���F?��Y�פ�5L��D1a"O:-	��0��h���+G��lG"O��e�S�a��(�d�f�����"O�a�F�Y�n�;c��.��hy�"Od�cB���h���	��',�lRv"O��2�@#݆�c֬�W3��"O"�y� �kE���<�b�"O�=��қE=��B�n?�Q�"O֥Q�\�n�(�CXf��d��"Op�w�'k��iz_�v;a�,�y�'P�}���y�
ֻzz�-[q���y�/�./B��9��P�?��X� �.�y�i�.Dƪ�3i�=B�LS��^��yBa�;[f1��K�G�hH��V�y��5 �ȩ�1`T568
�YUa�<�y��U&����,1���!畈�y�G��)�αj��:wY^Lb����y�dI7ց��F�iL� �D*�y�"�1�$T�"�>g����[��yB'�x��'h�Sp��c�����y�(O�K `  ��p�(0Ě�[��)�A��p���Q�'�4�z��L�4�n�3��_�u\�	�'��M  ���'܅#��ۉ'qzu����8h3p���'��C��ךk���A3G�j�6����� �͛�ɤ��}��cT���E�"ONШ�4m04Za������u"OPm9w��ld��RC�6m�r��S�'�O�0U ���iA��Y*���R"O���+�%z^��	�X�Ø�y" '68Z��,x����f���y2��LQvlE��e`��*ܥ�y��kEԔ{2!_1sR��E��y\*u�
TY���%�H�7&&�yb��>�욥g^0��6��yB�ތ�8(�p	Z�+3X)�(���y��2^5���#.��X#5	�%�y�m�y|�x��/����I
W�yRɱXHܙ(�)[���L�
E��y�A=2����+T����0�J��yC�0�Q���0(�Q`����y��\�h��p�v�D�R��\��yBO�y���jVj/h��t�F%��y
��gʤ����+^ξu�3���y"�C%F���#��UZ�t�Ђ
���0?�.O8Y�+8s����2�$cI�IS�"O>�2g L�hcU��r^�aQ�"O$L�%#µj�m V���TQt�yT"O��Z��-lc%Qײ �#%T�!�$�(j��@)p�[�ـ�Zpd�p�!�9�S��V?j�Ҽ��Bܤl�!�ě�w��d����n_`y�� !
����?.�T�$	/6��|��F�9L��@T���&�!�Ć�V4�i"�*)be�a�-w�!�D��� q��C���(
�S;+�!�dJ�Z滋
����Z��a�qÁ!kax��'4�O�4�f�^7�dɤ��88����(ړ��|8��,�C�zq�p�Z�ex|�r"O.숦�	>��q��ڲdƹ�s"O<�M��'�~��2c�<|GJtb�	Tx��M��5�@��e��"�X\H�*D�4���4���t�%n�JD��.>D�$��A�#*dY�a�8<����/LOR��ѷ�] �5�g�^�vPct ,D������GP���N�-n�(�S�>D����>�P*� G�v���H��;D�4��5J�jD���S�=Qҥ,D���Ri7 �J���h]�B����=D�8��`N�#��נŒ/�ʹ��9D���(S!z�qHV�Q��TE8D��ɀ"Q�$ ��� f�0��1f�z����	�)XH�	�E�/0����ƥ�	gˈC�ɸq-0��di�}4x��%TLC�I=H�@AvE���,�9�T vRvB��.4V�L�*nQ�P��0Hz6B�	�t,��Rt	W+c: ��!]"T*B�I4C�`�g}�,� �YB�	1.v�����5+�,�L�8C�4��Ig�S��y��J�11��?t�h��*�y�'ր;^VAP�ǟ����"��E��y�b #D� ���[�r����L�"��d7�O�PrB�*5^:��r`��r&x��"O��� _vʼ�/S�
���"O��G�k]����#�\PT
�'��Ol����Mw u����X��<!���?��'o�I(N
��k�H�T�C�\B��#<����hO�)�~tPD��	��$1x�-ۯ\!�d�;U�.l�1�y��������	���OH��.��"ړNY�`c։��y�YZ�gϋVw ���S�? ��Æ�@�#d9A���;!�x��"O��7�c����T'�� �b)�B"O)�Qʬ<q�iz"�������6Ohʓ��=�2��;UZ���A�..40jQb�l�<��kO�y�FA{Ʃ�����#�@���'@�O���K��'����o�(?�Pzp�N66��M��OL��䅇VЈۀ� ��h�$���!��)PT��#��;x�LaA'jݝl!�D�#B�*�x���~���;�b�/3!�ٷI:�4C�h�	04�b�&|��'�)��R
4Ѱ�ɑ���
!�_[wV���&�ɎGW&93vF۴o�&QU��D6B�-�A"�h�:�zb��>&�8B�	�_��m!1&��I�JTrQ镣B�tC�	�t�(q�5��V�Ӂ)A�eS,B�)M�$�����!x"YJ&��!�C��+yR� �F�3F����!x�F{��S�IBt�P��H�J��J�K�'���*��Yª\��'F�:�L� Y��'��O-��ă��"9h�-~�@���喭�!�
*�Z�b�'s��؃��*�!��cКpB)����{�D�2�!�npkî;a��v$�7U�!��5GX,�"jN�HC���V��8N�!�@��T� A��A.��@��� �1O����E��B�ŝ�'

![��T7��(E�� E��	�x�hTF[��yC1��s�n,�!�㤃��y��3�p�q�Ӹ�uSvd��y�BҹT�uB��Ͽ�����䅐��'�ўb>�3��T�����F
�[r��!�!D��:%�	=���$@E�T��Q�.!��<���ڦ��y�I_�c��y�C�U��d�<���|�+� �d�<a3A��C�Aj�W�j�^�C�Zv�<�� &�`L�0�݁~��c�Y�<	f��kK�=ȵ�<�b����Q�<Yd"�>Аsbeو`X훧m�V�<GG��U��^ \{zy�TcR�<�Q W��Ǌd�Gu�tb� ��	�l.����K�9����b��1aTB�	O�Y��΋b��j䈀�n/PB�I(2�ɱRP�pa�f���RH4B�I�X�F��@@�0Tȓ��Q�}�.B䉻yS�(��	P��뛅j& B�Jel�I��c�a�bO�<G�D{R��'H��� �Ø��<`(Ɋ�����.�	+jV���t��F��ɀF.LBO�����<a+����s���@�l4c�Ҫ]F���"O�9���c�L�q��r2��"O�uzf�R��$(ӪY3/��D
�"O��٢C_� �L�{C�
|Bp)P�"O�(�jɥq��th�g��mK"��(��r���O�"AP�d$\�T&dK�r���'�ȩ��ա!�咦$�s�0��'�H$;wL.a1�ur%�eZj�h�O2�=E���	z��[�0N��1�?�y�閁-������qgVАu*�#�y��&I� %YîD�mdr�BeJ��y�����M���`�иX��,j�!�G�t�)�I�Q��`r!�$�	Uv��KR�$2f�A�.>Z�ʓ����O1�~��<Q&���G��j���X-3�P~��)�'8���Qb%C��B`(�1Z���ȓ@�T���AV..n4�GdJ.W����S�? $h��B�/!�:���Ķ
��mY6�'��O�����r1�!�ϟH����A����S���<���`�<��U$�p�"1Bv�<�B�������+L��r#Jk�<�i_�F���V M�m��|�pȕ|~"�'O�O>aBI�7&����*W�i{,�3��9D�|�/�(H���B����{�*��r�2D����m��u�X8 ���;"�!��4D�H#�� ]�� I���%F��X�"�4D��)$�)w��P�$.@5m��Uq]�C��!b��
��G9a������=��C�ɿ5����e�?h�2�[��C�	w��<xw�S)Fc���)H�C䉀Dޜ!�t�Ԕ~p�p1��Q�7��C�ɤ(��=	�g��[��}���)C�,B�I�s��)ӰbK�LZI�Dk$B�	Y�\����S�#
J�`$�M�a(�B�ɀ-Ah�H�ձ{�I�&��3]��B��`�X-8���#Y20Av�� :�BB䉼1���!s�&PW߻$B�`���aU���/���P��� ��B�� 1ɚ�(�<q�a��.7Y�B�I���̻QdY�@=x-��W�'HdC��e�����g4�(a�`g�2��B�4n����`��"	߸�q h��m�B䉢�*y��,(�FMӥ"@fvC�I�&<����-Y%:W�ԱA �C�XC�	5Vth	Vk��2�v�㞔X�B�ɡHӪ)1C&�**�\l*s䟈@��B����C@ ~������*t�D{���f-j\�p,T�B�Ԉ7am lB��6CvQg��x��+�JB�ɖ&�bCo=c>�ЎѰf�BB�I����`��x~��ŅT(W4�C�5nnQF�� ��(���&E�^B�	��޴96�̎0����)(��B�Ac��:��߼'�|�Q��� ��B�Ie��X
b��{9>�rG����B�	&�	��A�'u?F��u�U!F�C�	 d�z�2Q�ٙS~���&!��P�C�I��G��;}�1�Nå9��C�	�߶ ���	�6�@h)��>f�pB�	��<�e�3:��� �K�B�I��*�:IԒ��+�@B䉺t�p�����a#��P�B��B�9��IC�:�C�	 L�y�u��������H����>q�K�'n�yh�l�-�� �l�<���W�0�n�����D�0�S7�`�<y�m� �Nc���E�j|�&Ze�<��-�Apf���j4T���Yh�<��S+Q|%2��@ F�R��v�@g�<��̥����Q�ڿq&���	�f�<��1��8X	J�]?�}8"ȑ�<Y
�)����EE��{ Yq6h�<X��ȓ�B��eÛ/+4��ӧO ZM���6�ց��mǊ"�Pp`cL:b̤��2�����mXOIH�����0��m��D�"'B�뱨Z��(��������i��&�q�!f�d5x��ȓN��c%.1`*8�S�\?ʴ"K>�����/�b���	Q�n%{C���N�!��o"�ࡳ�7j�<���ט�!�V�H��l�S�٪Z�U{��	�Ze!�� 2�sǩS�2�|�H�ʲ
� �K"O0��Ǉ�c��p���)[��k""O��q�擿� E�զ_�^Uʩ �O&�D�=c�UJ����j:R8��B�>�!�䃭Lw�l�� -�E�ڥN�!�
�0��Dҥ��
VFܺU��b�!�;*�\��U���e��r���4!�$?L���4IE��X��ր9!��I�W�h��*r����L<�!���Z��{�P3���0ak�)#�!��ǃrKnQ9����6xk���u�!�dC�f�Q��ٗ^�ʱ�����!򄁮M�����v�|A�*		 �!�d	W�ƙ�D�Ҟ{�l�%@c!�Ą0dZ,�� ���ԇ���!�d3*AJL  L�	&�s5�U�!�!���+`��|SE��.W�h7J�?�!��X2!�se�B26����*}�!�D� ��<�Se��;�$ �c��6�!�V����k�Bַh�$)X�!�$C�'\XJ$
�b��̓S�ˏ7�!��nza2�o�,��T�����!�$�8[�v�{a�1qC���^%{!�lU�2�jnO2?J,2��]�$K!���/OUp�����76BU"D��S�!��׀?�*Ix'
J0�iV��� :!���)kN����d>�qF�y/!�Č&�(�y5'2o��`3�E!�$ k������; �����,�!�dEQ>l����:_�A�I
]!��#*D֕��a���� ��U�i�!���1�H]q1B��6m�Qc���!�Č�~��I�V�n��}V�[�'�!�DS-9x� T`ŲX�:t���L\�!��$hv��c#��Ҭ�p� 2�!� �y�ۣ��!X@)��BE4�!�ށR���c��<:f�bw� e�!�5(����	S@쌀|�!��$� 1{т�~���
�t�!�$E�̝q��A�)���@?!�D�+�!P�*�)[�x�C�R�C$!��C�p�~%ǩ�4,�ĕ�'K�Py��
$|�񪠢ʓvJV��#�Τ�y�V�/H {��x�vS#�9�y���1�0��R��
x�+�&��y��Z ��\Je �	�����ڼ�y���w�>DaCԣr`r�2�S�y���{֌]Q���f#x�S�+��y�MT�
Ly�$�G��1�D��y�k�&��)�c�V�I�����'�x�%�]d~]����pe��'�ʱQ$��pY0����3��DH
�'�*��p��8s7
��ᯂ5A*\� �'hR��'��=sBC�'/����'6�Aq#�Z���EU�''\��	�'�t���ȁ8�ܠ!�S4,ஸ9	�'�0*�#2]�Z�[7�X���'����8y�4�J4Ɣ'�:�'�2݈��ܚT��5Q�B�� 5��#�'#�pё(Ե�%�
����'H�)��&�����C�EW�fd�'	0�+�(Li�mE�?	�]j�'>�{�GTL-9#ǂ ����'�VT� ֤`�^P���ҷtT��C��� ��KC >}�|A����$H"�"OEѷ3lpn%Gc^
R����"O"�0�L�:@q����0`���"O~L�3��=7CLy)��PYGN8su"O�����2�IAv�V!8�('"Ox��@%�0H.��0��2"O� ����'id�[�P������"O�b��'o�����CȚ ��"O�a�9����2,�r�dը$"O�UjFΤE͚��_ki+�"O���	F
D�8 !�2Mh��3"O!�'$��t�Ae@Ȏ%�8B�"O�ԙ��L!q�y�rHN1a�����"O,��bA��0�ʨ����$4�dJw"O�1���A�a�V�xB��<.��$3A"O�DS���m�C�f�:q钬�"O�q3�@��E�*\�Cg��H�2�1�"O"���̠PWpR��;O,���#"O��I0f  $�Y1��P�"O@@!s5C08�Dĉ"��r"O���E��DLH9S�K\:���"O �h
���R7������'�,P�&�C�B2���:�Ɉ�'�Z9K�B�}�u#2)ż,�� �'�E2�ax��E�'�DѰ	�'�����U�y8��l���'d���'	D9s�3�����c�'ը�֤ԝr������;38���'�X$�3��o����`���3�'�xPd.�c�~�@�L$4z@�'�v�C!+X!q$(�@��'аI��'�sd.߁����u��5ajh��'Pp�NB�%L@�r&��07�z�'ƾ��g�=~�0��	ʜ5���S�'4ܵ)�T�@*�A�u%��,��d��'k�}��f(����a�B *����'����*O/gv���͘�M�����'�~�#D�%e���ãΙ�E9&�"�'��Dq�!��5�޵4�W	6\��b	�'��� Cht�����S�4Rt���'8rp�A'	u��<jщ�33�D4��'�TP(S쟄N:�S��:'?8L��'�T�e΁*ӄ�ɦA܊&��ձ�'o�p{���QPୈ�Ȳ#� ��'���G�Ӄ?��@�%d�_�4�a�'?��Rk6����ݸV�&���'��y %�^h��2�+S�̔i�'��h�B/؛^�c!��/])����'k8�D��m@!3��Z��i�'S�q��D�t�z�A7� 7�`�'r�Ȃ,i�<��֪��|dt�	�'�Q��E�Q�N s�Ƿ>�r���^��]#��/C74K��72�M��[�r�����"ڰ�b��ɼh! ̈́ȓ3��qE�O�+��ce��Q!nt����l�7M¡P����6N�H�ȓ tք��a�(yDh�Ҋ�(������=a�"Y*+��A���I)TC���I�x*m�4���c�("�Շ�%Ȇ�j �6}R����J���`�ȓ}����#D�;f�9�CZ%d6��+��xX"KCr���e������#;�	���L��o��X�ȓHv!.u�5��m�R�1Y i D�� H zE���J�p��(�u���aD"OŲ�L̊H�&��FN'_���ٖ"Ox���%D&"2��f�N�W���"O�pI rs�$�Q*@�bQ��á"Oz��v�8V�J�
ߦ<Er�q"Od0��h�/AnP�H+5/lb"ODi������2�Fлm"��q"O����T<ib�z�NܨY*���"O��#E;�jQ`��֎M�Bu��"OD�p��L�I��h�\<�"O��ۄ-�&Y��(E��*N̄��"O�� @ȭ$8 �g�с5`�$��"O>���@��Hѯ�V��9z"O�1� .�"%R>�P6/ث��=)�"OPuyR��**UB�p.D#j��t��"O$���7gJI"�L�1w�h)"O~���;��l���T�s��,�W"O!�0�f\=����EQ��r�"O���Wb�%��RC�G0EQ�"O8�"��1�DQ��fÐ4���"O�8�cC�u �@��cgR���"O� ��Z�#b~����4[}Zlt"O%�S(�$^+�`��Ğ}^�=p@"O��
Pa��Ό_j�a"O� �����YhY�9#A�]�"O��	���{p�U��B]6yS�qc�"O�Ԡ-�Œ�Ag{��J�2�!򤐰2]N�*�&���1�A�3�!�DL5eT:V#»4�PA�d�ĵ1�!��]�}�(�ؠ���S>�$[��J�7�!���q���Z �R�{��l�&DD�}�!�E�0�t� 1��',�x�6C���!��2�D�,@�<�#�!�^�t����A�K�A�v�E���!�����ԉFF|�`m��!�?1�,u���FX��8�˷�!�$��}�
 �3e�,?fA##Ч�!�dт
��0Qp�ؓn<X���+�4v!��E���4�B�UI�ը�!!sj!��S�[����"*l+>E�0A��X�!�dY�������$b�s�,M�!�$�s$Lzp�D��Y!�Z!A�!�\�8&��r�����r�M�o�!�d�.s�B4��C.(���C���]!�\�s��cf�o�\���Ɉ;!�Ę6���1%hќU�̔�cg^c!�S���%G�.�8 0�!oG!�䏧���)�tY�t	hc!�Dc^�tB���,���"���IK!�d����R���N��n@:!�_H|�ԩ�!� ِ��"���!�D@�>�����"��v������f�!�?*��R䊺m��H�',�!�ߚ7�P;d��TE�ĘU�!�$�/
9\���ۘ	���kb˷+�!��K�.�g,�:*oP�Yh�d�!�DK� \��N�1{@���$2�!�d�'JtZD�%�K!Hц�1f�C0*!�6o`I�5�/�"����!� Y2���1�%?�x[ e�/�!��^�<��1�Y��̐�c�$,�!�DC�8�Z��д(�(P6L~�!��)|��Bp&�7\�"��D�Yw!��Ƿ6p�
���Y��iy0J�]X!�� �5��ūk^��rsN�/M�pU��"O	t�Q�E,`��MK7�싗"O��xQMǦY@%i֬:���C�"O�-���$R�H��K��+��"Oi��Y�ẑŐ�*�7QꞱ��"O"x[�O�6 �pUHH�*���2�"O.��B/�$lr.}�WD]�f��cC"O��S�$Ȝ|�1#���X�"O�UۦARK��� �GL�ޭ{�"OxIa��X�C��"�28���A�"O��P��8{�yc���*X����"O�`���ߵY	̐4@�2��Q�P"O���)^� �r��ΫV"t�"O�%���8>��"s.�v6<�'"Ox�uj�+�\����d�t	c"OPQaT�]'(hJ9�U�m��p�"O�e2��b��Ѩ� C�J�6X��"O���}�̀�`�7�vu�V"O�d����64`�.X;�� ��"Oƥ/��~�و���9����"O�eq�kN�J,��ӌ�>4����"O������0erLͱ��y$%��"O��� ��0.�����ȝHb �9�"O0�c�B)?k�̩/X�b�)�"Oؠ��;f:D'm+U�YQ�"O��Ig�r��ܢ��۶1���{�"Of$��l��"�8V�_�*����"OĐ�fV�Rs�,��]B���R"O١'E�'�z$�
Ch&����"O�Q�N}{�Dx���7Ab-�A��d����a��[�OBs%|M�#��6-�!�d@l��XP���E���V���N9!�*'�TUZ�!X�T% � ʽ
6��R*�I�>�g�G�r����F9Y�4k��>b^�h�'��6orb�@���H��(�H>���� ���#�8��=I<4tITJ�0p���q�x`���V�As�]���C4�HE�_�O�
Pڂ�	s�� f&����+O�D���m�P�O��M�wD>kh��2��!s�B���'Or�+�/,��<@�>�P%��y"�/���3f��ʊ��0��
�Hw^,nT؟\oZ0�l�acB�t �
��󓑨O.A�%�x2���S��E�X:1RF�%�0<9����-Z"��! 8Ev�9����\R!�ā51��1��/ޟOb��M�!�$����6A�
 p�����=����'l��x:W��h0p��� �(@����?D��P4�
������J���e9D����AQ�fL���Ih�8����*D��b�,��z����F�.h �m=�O>6M��~B�O
Bj��� Ӑ%Y��SB������p>yA�Sg$��dN'a�<��c(Bw�<�a%V�͖3&��<_��g�M�<i�C�Yk8���'�#�:P����OX���O�}�B�;��I�����0��"O\l��E�$@�p�G�W�X\
L����<�M�(%>1�&��$����ٹy�xt�Q�)LOX�4Q.���NŐ�M
xD�2e�eӌb����sӂt����*���e�P�^�G�|�-�OZc��>1j�
�$^A��V�T��Y��H���'��)�3�@�(a��'Ɔ�	�����Ӑ|��O���d[8l"��72�D��ל-�7�O�H�c	*,BD��Yl,BZ�`�O��$���zr��Dx9��gJ'�<���OZ8�0mLy
� ��0������e.
Ue�K3�i�B���AW�B�ɧ����L��L�ܑP�I��k���c7#���O\�:�̘3���{RG�)o�R�8pĊo~Ҽi�a|�.�B,���M^�\���֩V��ēӨO@�M��dʒh������|�fY[r�Ut��T�'f��Gc���*Q쀡,^�9��'����Y�q�1Q=0<�4q��D/��@f��Q1@V�88��ė�(чȓrMF	A���'�"�uiF���hO?Y�`W�i��4�ggлJ��5�4�:D�L[CO��L�v�Z@�M��~�ؔ7lO�ʓ�~"��w'@}�4Iܷ-ֈ�
LU��y��K�.�ѣ��"D ,1#��y¡^�eIi� �By��EY���O�����D���a�΄(l^<��O��d�0�L�2�a�m�E��N� 7!���.7�֍11�C7h�4���D�.0!�;Ȩ�e��6�:m��"���F�tLa�\6������2�$V&|!�� � �0���g�0�cZ�!��ۍ<�P���دu���b�-K�"!��8.��!pq�O;R�ʘR�fM�3�!�ɆM��IC%��_.h���)fa}bO0?�)׊H.xktdŘo���[�	�A�<ɥ�V)��갩��cb� !��y�'1�#���5�P14%-�E�$H[�<��^�H�ٲ#�N�Z� &G�S�<��K�=�X [ch�\�^��5��P�<i��ٛd��hbiN�����v�<��
wEF=�֥N>X�D��v'Js�<��G#�\�Y��#6M���k�<y�
W�2[ޕ��VY1�'�g�<�͍�	�P��K���@�Wb�<��';;���C藘I���"�_�<��A\��\���[�kZ��X�<Q��D|*A��B�\�,��jFz�<�VMA�Y�X�c`	�%�� �_^�<Q�Խ ��d��`A�+� �3Q%�\�<�%D4Tr�Q��[�S8n�1���[�<��*E(Ha���aF�03��X�<������:d���~J<��բT�<�t&̆����օ>��kF��y�<�'b�_
�;K�8�2��[`�<	e�S�24]�&$ҲK�:楒e�<1�jN�-w&Ś��²s���)��\e�<�&'ӗDX���'Y؉���^�<٠��/x�h�d�r xt	c�[\�<�LόV�V�S�hY��Z a1�\c�<1p놐A~���O@�B�ؖ�v�<)� ��D^�18�C�"�
Ő�ʚV�<!� -��$+�h7�����BS�<�箔8 e
�&��A�B�HL�<y��H�B���o�p�(HWj�`�<�`�1�҈Z���B�&)R��H�<��	����hR�D^\�l*�_L�<Y���`.qzr�80��mYA�<A��էa�=!Qc���p�
��<��ޯ |��,�@�(h�̓A�<��#Q�Z �x6/��pOd�[q.�<�"�_�$-� ��D�>|^��Eo�<�Ef��&�*�HoH���EZl�<����</&�mJ�BZ�}Ti���l�<i��J%A^�)�&͗f��jcd�<A��Z�cق�{�_
=ʬ�a�\Z�<� �x:u"<]���������p�S"O�ZqHHg#�L���D� yz��$"O8�5fK��ԎZ~���"O84:A�9=6p�V 	G*��*�"O"a0Ď��]���b#�0�B�` "O΍���3D:()[��D�C��I�"O�4�G���4��Uk�6	c�e�s"O�)B��R>%��yy�	V�a.��"Od3-��2�h(��B�礌��"O�]���@�	�dp����;p|M�"O"9�g�GnZ58r�  o� "O�4��M�yΜy	�*غ3VP���"O ���34��I�h�LB(�B�"O����=Y� ���F=`#f�Ss"O�I�5��;t�f���f��7�1�"O�����j����wD�()P��f"OX@4���ܙ��^�[�XU"O0-�2�k�lE{3e�G����"O�(��C�xeِ֘DՀo�y��"OV��ޢSS|�9pIر[���"O� N��]���^��@Y�"O������L���A��/�f��6"O�+VNM�-���"@>ɨ"OX��V
��4�d����3� �"O�%X �R�e��(�,@�<��"Oi÷bY��Q�R[�Q���0#"O~�;�	r!p�b�DD�F�����"O�x���9��	���U�%�؜��"O�Hq��
;�ĤK c[����"O�u@u,܅�D�Ӣ�֓=����"O�q�c	�g\���׃H�l��"O �`���B�R!	"���(7fb�"O�$�v���D��b�P�B�89�$"O�� ��:g4q�� ;�"O �[��]>|ĭ��
qp80�"O�!ʇ	I�QyԨ�O�#'~�=:�"O�|�碀� O��#&o�+���"O��g(L�\M<��O� 2(�Hȣ"O��:��E�
�0�����^�Q��"ONx�1h����#X���� "O��`��8>�B��J�6�0�Z0"Oz�2CI=gr���N&9ӠQ�"O�a���^3<���a�� �Nyzq"OFpk$��*���L$��X��"O�pi$P
�����T"�-˒"O�\H6n��'�P�H�j�#9�T1(#"OF$*T��<@Ǟ؃bJМM����"Ou
�gēRߪ�
U�G�3}�" "OZ�	�B���9��U| ,@ "O☫���F �bf�X�P]F�+�"OBܠ�E�L=<������13"O`E��(Ĕ��fL����R�"O2a��/f���3�ќ��i�"OB���/@	��`qËM��LQ"O�1�SD�<�����ޗ~��C"O�ܒe�Z�46 W�L&5N��
"O<L{G���,!&� �L֏,� �'"O.���nG;WUƍi"4��2"Oy���G:7�f}Z&�]2��@"O�!�wM�%J^�$y�B�P��H�"O�a�V��h��l�� PHlʦ"O ��5n@O�0	�̮!h���y"�r�P��KԶe���bݝ�yBZ%X�Bd�qC�
VH�n��y
� *$R��^�>�;b[%0;�""O��x��Ӹ%(�)�oI�pX�zd"O�̩�-�nP�ŌJ�v�B5�"OF%�2���@�Δ�jvt�se"O�*2
�Ϥ�!f.�nGlt�"OF���	pY��e/�557�h��"O:�aF тA���@O[�v�t-A�"O�P�U-1"�r��M�]p:]�"O\@2!D^7a\hL�F�Z�Ag��1�"OjU���V������Y�_ȵ[�"O~Hӫ����Q !��nL��!"O�i*`I�7K�|S/�>zF�!�$"O`���B�4��7��l4��r"O�D�MC�\D�p�S���|�&���"Om`��Ԯym�){R*��ЙQ�"Ozl���9{� ڷ�U69�\JQ"O���'��q�U��͘ $ Z��c"O�%B�۱17�a�r��0R���"O�H����Vp2pA2���C�$�P"ORQ�q��A��pb!�FوXe"On�� q}����L��%�`"O�9��7�49��A,��\�"OR�QVa�av������Mj�"O�� E) _��ˡ
�S�D@)"O�a��E�+y��������"Oй�!�$AM���wiK�.h����"Ov������ ��@�=��<H�"Or��G�&)�HY�E�m��yjG"O����΅	D�
Y)3Ί.,&0��"O�K��Q~Il�p���=Q,$��B"O`PP�];��ieNW,*"I��"Oz�p�l\�u�@y�CS��lP0"O����1�t�S��	��8�3"On5���?4Xh��(�p�="O�}�J�
'u��@�aK�HX$"R"O Tx֯�"���[��O�@lX�"Or�w�ݳn>����`L3<.��"O
HjS�I�2�vQ���� ��`"O▜{H4��X"
!��p`����y 	24���a�%�EK�O9�y��\q�ҕ�B� 6pY����@,�y��[���2�o�t۲����L��y��UV�L ��4@����3�\��y"�_6}x�[aJյ&N�� RJז�yE	�a��AcI��bHzQ*W��y�bP�x�ڴP�˰L�X�C-��Py�M�?|���(�[�����M�<	���	;�H��@�#[�f��Q��L�<�7��$8��m+�Ǝ�9��0u�1T�����3��}�!'R�oa4ؙ��!D�(AE��<)#����*P�1@�]!Ŧ D���aՓ�:�(�;!�%hwj D��	��&��s ���f�*��!D�X�R�ڗfz:���� �/���R�=D�H[��[��l*�B�Od�۲�%D���V��>S`H��A_�1���J�#D���7��4h���`�GA�Z|�,!�@��<2�A/t����,:]6`��Hy��=E��4K=���G�e�0��Ӄlj
���n.�j2f͸�(���aֹT�чȓ9�������a�ٱ�̀�1I��ȓm���1��\�x����(�qC�i��VD$D����+���uI�,��k�Jh���S����b�-d�&��S�? �� ��;J&� ��L�2��Y�"O^�(�䇈^r�)������d@�"OZ�+@�R�`r`��*�<�"O>͋g�>1%Ed�x�2 h�"O��`�,..��=�Sb݄
�x �"O��q��3>ﶤؐ��sjL�i�"O�Ӑi1+䞐�� :T��G"O���W��@�H�"#6@L�̑#"O	�n�F�� p��X6֔��C"O�d 5�[s�z�IB������"O����!G*X_�\�"部�*��"Op@��;�°���N�k���#B"O(�R�垔΂�R�߀,���Y�"O��-a�	�O
$���T�!��C8}���`L�2��]�Q`A3G�!���&��6# ԼĹEj�1N�!�/o^���Y6�0�2��;}}!��&S��l
�L�P�6%����*�!�d��c"���	A�om���&�+\u!��P�V1lL��$�.S|J���e!��Th�<<�MjY����	�PG!�$@Q�5�͍�NP�ǉS��!��H�E��ʆ��
Z�8iź�L��7z�z��O�lg<$�$ql�E�ȓqB�<x�qR!)�#jJ���e��,�j�`�@�[�#C�c�@�ȓ�,t�5τh~�(��	17�X�ȓ�tkԅţ$�(���/H7dɆ�s�hę�@��1G&�)fG�L����ȓT�Ɯ��;<�|̱cޥV��\�ȓ!M��(�ȂM8A��P�L��ȓy��ux���,F�R9����- �9��+��+�ȸ��l`"l��%]���>��SL�	Blve� ���ȓut�ˠ![+�D����!����ȓz��%��a�O4�mՃ;����T�.] b��4*:��AeM)	<��ȓv�6��T[.�aC������ȓ[J�l���}��V�& p!�ȓC�6M���ڪnN8���H�P��ȓ6�[!��3](܂e�<Wq�?q���~�ӌs��kB"�%~�L��@�]�<i'�S	���!�_+zm��`PA�<�B���z�1Ï����|�6lQz�<q�E�{8��#I�V�h�歀�<��(�_@԰�a�:l��-��g@�<!�	p��z3o�4
��mۡ��{�<a'�ѣ��!��(BJ~�As.^�<Y�N4"Ƥ�d�ܧ�� �E��Z�<��+'�13�kB�<�bik" �T�<���U(\kU��"�(I���Sv�<A��.�٘�� ���*�'Lt�<15��K�Y�ՠ[�M��z���q�<�*����dx7B��It�L�kT�<�����
�p�u	֯{tr�� g[�<�%,�B�×�Iu^ؐAV�<��S>w�vX�D�]�h������}�<2�J�x��L�C�ѵ%
�Df"�w�<	�\m[Xxq��	�5r`G���yrj�l�^��&*F>��Pҧ��y�aC�~�
 J,�1zV���y�"�)��ɺ��]�&+\ӕ���'�ў�OCh$;2a�\e.�K�[�\x���
�'��dؤ�'<N]�a 	Mp<��� (�贩G?K��S��$$�DbB"O�<wO�_(�3'�G�/}�	��"O�Pз牚
z��a^�;@11�"O�܃�����qqEk�o�t�"O`�h�i�9���p�5�%��"O�ĩ�΍u2@Y���9�R8w"Oʅ ֡�FCH<�؂,x�"O�(8/D�_y4��U�/�@&"OxQ��Ȱy(�x�Q�]:X2"O9�c�M�-�\�9�ë�
�h3"O&�z�L�D_`ؐW��u��9y�"O�x��Ժl�| H�ӶV�*Q�w"Oޕ��N�W� �("�2����"O6�{��,���5ᛱ4�� +�"O��y�jE�UB>,�C�ָ�(�:t"OR���A� (�y�A僖LV�%��"O�����L9n��EBW_��	"O&!y���p��T`I�%D�u��"O�z'� ɖ��� �8>$��v"O��4�Nk�PJ�m�)5=4|q0"O�H���H�z}`��c#B=��=PF"O�5KE�88�Pst�ԟ'r��{ "O�5��$�afZ�+g �b	6��S"OR�����Y����e�0>��*"OF�&C_=�PsEX_�$4�"OVL:�L���ꡤ� &��E�f"Ov��,7�~�+ ��pNA &"O&)!�#�:*@����ެ!&"O�t�2˘���D�4DӘ8�,
"O(�I��(NpR� 3��-zx�y�5"O^y��ώb���Y���'>th�p"O�|��HφI���9�
�5H���"OBlh6� ��Ze�T-9��=*�"O�̊3e9m�ؤ2v�A�,f2t+$"O4l� ��Ew��RS�D?mZ&�v"OT�K�7�^����I	 �$�'"O.�PhC�X:�x�+{�$��"O�yӂlO�b�j�µ��$aDe��"On�HF�#��t�]�o7F!s"O�@���4h6��r���<?y�飗"O�8��/�t���s�$ �M@~	("O�a���@3�^���ő&*��B"O
���_�bg��ʧ%��R����"O:p�-��'�F�x�n�&�jp�&"O�I���^1X9��s��OC����"O���U��3{xX��k��@0J���"O�$IT�<0�1d+ґ3f��"O���	,}�t���p��p�"Oz� Eˑ��%���j%�@9�"O��j㥍(Fv����(�v��"O�45���0�`���c՟"t���1"O>���KfjP�r�W}ц�*�"O�,P��P|��M�B�ޑ����"O2����)K����(W�(����A"Oҭ(&�O�8\��8�fX�HO�\;"Ov����l�6U��*�
�E"O��#ߨ;���Q���U���@"O������= �X�׆`�P}��"O��7�O,�V�z��X.�d� 2"Ory��埠V1v�K�D�q#��$"O�;�E�h����U��dpPڷ;4����&�lP�t�^\WPA�BD D�@�#��"y\J�
�-Z|�(�sT�3D�3�nN�)�\�AT͜�e"�`/D�� x� D\�h(*�/V,Eq`` "O�X�q��V��y�qǅ*�1�"O�4;VΓz��)�ҭ;█��"O����I$Y&�u��E�{��,�y"e)e� ���"I4y����yr� Ж�xc`L8	D��@�9�y��пolD��3O�:BԄ�dh ��y��L75�Xp���0gؽ�$�W*�y��	"N��צ�3e�,
d�\7�yR�%*�"�"��ʪq/V�yᨙ�y"O�pf�[��j��la�� ��y2kM�-��hq�H�I�`����Z�yr睿Ϥ�Á@,AJ��ef��y��[��,P�ti�o@�i�T�X��yB��
Bi `��m�	b]�!��&ӷ�y�HN�F����t�P-[;�2���y��ٚl�� #�@�B_< 1�J&�yR���&�jP���9��E�U��yRk�#��(�� � E��p���!�yZxd$W�����V�D�^���+�'�8H3e��٬��Z�v�Y�'�D�Z�)��A<$�b��<[f�a��'?b5��ݫ	s����9�0�B	�')��$�T�� �8@�V���c^:�y��
�h�����F)~�2�e͛�y� A�)��u�q����pb2���yR��-p��hc!JF#����-]!�yB�y�����Q70h:w���y2�[�<L �TW�ؐ� F-�y�ŝ)N&��j5>q�ԒSJ�y��Қ55�yx�M�0��(6�E��yk�My�(��@@�G���+F�y�(��-��0�dɉ|5Y��J-�y2�#.�%y�ŀ(Y�9���D��y�*�'Un�K�D%��8�c�#�y�
=j8TD�����B����.�7�yB
t�r����
����NN��y�#V�K2\�)��L��v�Yf�y�ϙy�8Y1e]�
�$`Af����y���yzm�<��yzv�Q.�y�o�s��a�[�@ūfM7�y����T.T�q)�I�,8�d[ �yR�ڧ_�±�'��;�px`��B��yb�M�w�Va	�C�6� ��4�W.�yR�ݾi����O9!H�Y�����y2�ѳM�<����$!2.�ۓ���yB\(9�`���1%�LY���y�`�/n�(%�'��yaSˏ��y�ɖ�lEB�!r��a%����г�ym�<*�T�@����%>�Ӕ@�(�y"`���j}��.ӗQ^����)���y"�F[�p����8M�밂���y�^$�a�B�F1�-2@L�(�y���#'J�a2��N�5yس�B���y2���9�^�;Rtc5oW6�y���a�q���8)	�С�b@�y�M��1��`���,+�����y��� ZL��s��)5�[ ��y��O��YHB$�.$��`IDˊ	�y¢U�N*����l&K����lϚ�y�KR�W#��UA�5	U���+J2�y"�[9	Z��v�?kR`�#��y2Ozpݪ �?�z)c剋�y��=3���J����y
� 4=3s�<3�U��BD:��""Oa(�f�QKD��ū2�y"O����Џz�֡b��v��|1�'�ԥ
B�Sw��x93O��s#�.O�����:�����d=�S�S(<Ϡ�"�Oًq�T��%f'!���'��H!+�OA�����^ő>acɾBVr ��ޔf��AA�:ʓİ<Y�(��kV=��h�-�e�r�ǲG�J8�f U;��p�b�Ѷ/�v<�|�<1�Œ./n6��UD���q��.[�~��D�J��M�v&BԤ�JG)��Xd�M�K�%ib(�8��v���U�$5��G~D!9�ҏJF���lM�4&�#?�J	�>�t@���em��LG#>��VK�&E��
���O��|�C����'�ў�� �����* -@H�cH3����OT	x��dՀ"�b�����FQ6�V��,�l�(B!1���<q� �98��Cpn͙|�&H0�g�F֙����ڜ�J�OT���MKCV?�fN�}ڠFG,rW��
�h�x@ԍa��'�;�'�� ��]����Ԉ�N��K�ȏ!���`I�ɟ��&����]3>Pn�z6�z`��`�4O�ў�R��՟�7��Z�4��S��CE;9<����޹R��{�M6�"i��ORL�S��0 �TХkM�[�9�v�'��P�i�p�	%]�dЂ����aJ4��k7���'b������{r�%��CV�C�ɳ,�h1����W%(�+w!��>x�2��9��hu�B>sf	����|���U��uWA6?1D��Ky˄�ښpd�e� ��Vx�l�@%�C5���X�޸9Ʃ��^:;��9,�e�5�̙g��9��eðaȝ�b��ݸ'�������ہO���R�(�2o	Ȏ�dۅ0�1�F@ӡl�@��ƍ�D�] �� �<	��mN������˳2��4) �3����G�h��pb�[%6+�M+�
�Ot��Vi &ղI"7T���򫇈i��PR�;�	�!&�(i	f�bUI�"F�3��C�/j&�$�qE�=T�	&F13U�ڶB� p^�j�C՘Sals��|R!�VfF���O�-rwʿ)����R��0�|9�'�zfl]�vRT��"���Y�@�cm<��Z��-�b}��OE�;��i���*d�axR�;Q$4�[��R`>hl;g
S3�hO�����M�-�GY�ڵ��l��j�Hڱ�D�w�ԬX��9T5����^��NB�I�2�� �agΆE�J-��'aݦ�� r�lP�+��;��XBv�7����·G�N���$�7��f���6�!�\p1�9D��U��ײ1;s@D=tW�X��L(T��P@m32D�[wŊ4OF��'l��8YwU���ȜZEl�{���j�OA"��p��	#��dmZ�R(j1q��P�9��D��\���"Vd�0E8EؒHI��)�E	�0<�$oT=F�Ҭ"Uf�'+��B�c]�'u"��'�L�y�i
$���Q��L�ۖK�D���!CB�p���'.Z2l� ���S���z��+V�\I�GN;l5(��w���4z��f�R�R���	�W��>M0��̂;
����]� ���2FA.D�T1&
H#t�>L��l��)޾@pW��b��0��j̖�����5ϟ���~�'��̱����-�pLC�M+#3*���
�2U�sg�pI
�0Q�F f(b#���	O4��9�d �RbPւ�0躔�˓a�ة{�d�A(��p�M��XIE~�]�&ofj��n�,�����1F��-Yw���(�`�=&p �D��3}��B㉍b��*G��<y��!��J��˓��5�7L\� aR'#�98���i��I���PS�
1�z� s�N,?.!�לD:��CAH�Mɦ�� �p�i4 S;��ҔL/	&�Xa���
$����ޟy���qn�ݐx���*8n�a�O�'����X;/�d�$��<��� �d���Y3#�R�g�2�p���{����	g�6�`����z���a��%X$$Ƚ�P[���>Z�Ą�
�bxD@�0�'H�y�$1�ȓh`p �)�:�ly����>;�9���Z%2��K�`=0�͓#2,��My:D����>W�`!��G��d���Y��x��pU^$�a�[���d�ȓZ�a�_}*�(��9��ńȓ^����1ȏ<);"Ԑ���?0�^m��Zx6���l��`-�$��2Y���ȓ ^����l��Z$�Ћ	�ll���v��$��ћ=a�5����1�RP��f��x@7ʌ2`�`�IW�'� ���S�? �,���Q�$����	��L��"O�Q� j�z�×a��0�H��G"O���r�FK�$����u�&�ZR"O��R�)J�3tڈ��n�.Z���"O<�2EYv��TH��� c�H���"O&D3���mX��)�6�Fm�G"O������+rJ�s&�ߙ
��<"O�%�^�@���0�JS=Kܾ�%"OP��񋁹��%�$��1
����"O&��c�����1,���0��"O�a{bPv ���N�t
���"O��Ӯ���L�3��LW2�a"O�a�`#�������:d��ӣ"O
�˖�ڙ:7�����l�<$*�"Od%�tA1Ѻ����Q��t�!"O�0c�Y/`�މc��$��d��"O:�p�Cq�ݠ�dײ""�S�"O�!G�V{�`��O#' ��"O¡�ь2U^�̃��&��4c�"O������P��W
0hNī5d�T�<��Ò�D�� �φ8�V(d��[�<�aIG\8�f
�;P\՛�IBM�<��� dˊ%�#�6v���KíJD�<ѵ)��^R��"�,W���c��B�<�&��^|����ƖI�"9�R��<���»���5�_E|%i���<�5f�'>��9`�-r��8pm�P�<1 � U<���f�.�$<����R�<����%G0Ep ���'�n�c�Fg�<��J�<� �
cNX1G&��Poy�<A�ڵJ����e@.	�Z�[o�<y�p�����*�����d�<BM�{�"0�2W����4�\�<���k��q��	�y��yW��^�<��jS�rz.���J��*Ѐ`��n�<��UM��6����qR��h�<�#�D��2�0*�1zXp,
��H�<��hJ�{�
(0�C��71���e�A�<�Sˮ9���1��2F�����[�<F)
�4�2����D$���I��YO�<���F�o�l�t�����G�\@�<a��\7z���*5HjM:���A�<	a�W�'���@K�$yX�FC�<��M:b�Lt�+� P0.}
�k�x�<)b)�,�H�j��a5����r�<Y�A[3D��tD����p����n�<i�b�{�H``�¯S��x��Ln�<��J׷9a� ���_����g`_b�<�ƌ�~-��s1��&=�][� �\�<��AO6}��M�L�>X�4,|�<���_[sx�+w��p��RP�W�<Qs�	T�0��oF˒ ��DY@�<���<R��W��"B���0.}�<�T���C�A�B������i�<t�-�,�'��r_�bt��W�<�A��:sk\���B�=�\,"�kX�<Ac��6  XÁ�Ky���Z�<U�0#GJ�8�/.���QfC�<y7�׉o�<�1��ƯE�bF��y"��*� ��D��;N~��9S�yb$ݳF9�ta�"̦��(肤�6�y��H���@�P|�MX�� +�y��-V(�,��F)$HJ�9�yb���m�H�s�����`��ҭ��y
� �MB���v�9dB�(�"O\ȋ�Ċ@k2����2�0!H�"O�D�M���y�����&Qp�"O����Ua��/!.?���"O*|h7h��b��q+TM�Wp��G"O`�����I��+ �]�tH��"O��`D��;sx%��� ��xe"O�����d�X)�Ŝ1�0�W"OȄæ��	��%� #Z��<s"O���Gꁒ5��mk"�2ͨ��"O\t��ʞ4�����~�Ld"O���W�L�!���'����4"O8�RA^�($$4����"O��9�AD�hϔ�8�U�#ku" "OY��Lc�T��� ��KB��"O��9Gf�	�P ���ĶDO����"Ot4�m(lv���oǦ;?�4�P"O�x���Ӣ+�N5b�o7��9��"O&�*,0)" ��قl��ɒv"O��q�Y�n�:`���U*
�T|I�"Oe���KB���W�ˎ���"O^�#��G�����E�a�"ORł"�	i�t�Ӷ�ʡI3�8�5"O�����7�ޘP�b�v#u	�"OH<��.N����p@�/	��܉"O~T�G���R��tAI�9�U8�"O��AB�^����Qʈ��"O(I
��Ed�6�B�I��F;���t"O����� \�v�����:kR �a"O:���dT~�i��\"XR �P"Ob�C��@�&�x�[�(�VK@�"O��gS�&DTTk�gILJ���"Oᘤk�?�>��@'��Wnة��"O� ���'l���@E>,i��"O����#�:f����>x��`"O���"ۯ
��G�K1\&���"Oع�����-P�,\���9B"O��S�HV(,N hG�X�gpܱ��"O��C$�q�̳�h�i,9�"O`���D^ =E�B�V�-j
��"O����7<P�
ejˑ]]���"O
�
3�A�!"vk��p�<�"O����N�#T��u���gjH�2�"O: ȃ�ۻ]������ԛ=q�m��"O0Q &�>�"Aj��߆
ކ�"O��MʼL%འԊږe$B5��"O"��/J�r�I���d"O��h�M�#Rp���.t� �"O0e{��P`�QE�[7':��A"O����R��"ht��% �h!�䆰!:]rDd��4m��p�n� jX!��"|ԌQV(�48mD��q�ȁ5\!���rU@�%��;I4y
L[R�!���:5w�,��Xך��ULB�P�!򤆤MOp�t��#�y@G�!X!�S�������/|�z�j���P3!��#�X���=���\��a��E�P2ffˏ, ���e:/c�I�ȓgi��[�+o��ȱ��ޏZ��ȓ4,=rf��Oq�m` 		��T�ȓ,�9�%���D	�d�R�LSܬt��*.�2�Y�Wʔ�;kFH��}��kh4d�`�4��H�H�zD�ȓZf��Wn=c� ��S�U6h�~���S�? V�`�i�.�B`ĩez$��"Oj!ɣ��{����b�9D��2"O\P��ہ	|d�C��-r�y�#"O�5��e�,A� K�#Hh!y&"O���u���)�n��U�Y�X�ʄ"Ox�Ra�>@��Hf(�>`�n�"O��r��,� ����"0a��"OD3� ۚ:��#a,¾Y�M��"Op�2H��E|"���Ώ�hŮI(W"OVܓ����`@�Cۚ^�*���"O�A�3�N�68`�K!�^o��"O\`��N�/NT��/(2��#�"ONp�4KF#>�4ؓ��7��@�"O�9kb"F� 3��J�׳ vy�"O�H���iI��T&Fk��!"O��JP%�%-��q�tJE��䠚"O���vf�0o�!h�!U�n<�5"O��z!�:��-"�G�V�[*�"O�-�#;c��Da�ƅ_�p��"OX�j�Ï�g������'4I�� �"O���e�͜,tH:����� G"O���ө
�\�P����WRz<���"O��Xd��E���H@O�m3\P�%"O*����=)�����-�5<u:�"O�x��#��,��T�	���"O"ܩ7�E(^R�R���U��A�"O)J��B�I~Z]��#ΡY�T c"O$餁8QȸA"�E�&	��;e"O�}�o�g�`�S�
'(��i�@"O��Y��$MP��
��νaf"O�ي��2�(p��v���!�"O��X�����Q�m�:��,z"O�m �� ap�"��3mA�"O�1Ȱ>j��J������P"O�QI]*2���6
��f��=!v"O��Y$�K�q��qGɎl��h2�"O4 [��W��T�qH��݊�"O>,�/�\��iV���8�\07"O(��݅�NM@6��Y�h�7"O�=)�K�RUp둣�X�j�d"OVl�#M�T�����,�5`"i�1"OT=1w��9r�z��AT!f�5�#"Ot�Q���xj	�F��+!(�B�"O��Y�lA)Z�P-��-T_{`8��"O慛P�P�PW�M	}���!"Oj����ќ3���cϩP��1��"O�U3�8qӺ�Bu��d��ဢ"O��isJ.|KZTB�BšB�\�s
�'W�(�T��"�,�'���
���'8N��3!� ����yyt�:�'�`��⊎;��͂�n}�|�+�'�X\�!H:&*��Ha��3i�@��'
|1&�1�<���݇��
�'JAJ�T# *���D%��
�'�J��Rcٌ)c|�aP# ��I
�'��
2�5d-ܳ�%ۺ{&���	�'���5F���~@��'ص9>&�		�' �P�ߎ1t����ES9 �Hq�'XZE���[�@��4 �Y���'�.�vdI�U��-���Σ*[��'�0(qgC�w��̃��	?	�0`h�'nT}H張C�U ��D�P����'��]���E4n������z���'��� bQ�hp�9��Aix�y��� �AV��=q"�3l��y/(Cq"O���m, 	��#�mW�1x�5(�"O����z貐�0%ԓǂHxd"Of��@B&�`hw�כ�6�2"O��bg&+I�ı�4��Y��+C"O����B�\��1İ{�X{t"OЁ�3��T��x�C�{c|HS "Olp�@�X�T�`�蚪4>ܓQ"O���A�)�DA�S ֻ>�h��$"Oh��]?�!˃^�U��"O��9�b_d����T��1F"mc�"OP�R��8<H��$�"I"Ei�"O8��f��;'%ꠃ4LJ.mJ�+�"O��$��S�D)P�יU&�Bw"O��H�e��}�����0mH1'"O^�Ӏl�p��Ƞ���8��2"OB	[������-��.�&�j��"O|�H���b²��!���T��Ҷ"O� Y�`�do���m
�c^�a"O*�æO@�9�l�t��!1d�1""O��c��|$E9�왻0��SC*Ozhs�BX\ �����!C	�'�9Z�E��n���9�J��O$���'���[ ,�>)4��$�(k/ر��'p ;r�Zi,"TR���`��\��'��hբ� 6�i�I�b�����'�J4���_6R��1f!Qw��
�'�xS'`�&]�����Y�^��'��c�gЪD5*��w�	�PH�@��'e� a+��n��8b�QI��!J
�';x�-	.���2��.2n�lh
�'�fx�N���d;�傴!@�1��'�`����3(5�ćJ.2*���'�>�9��	e�,��'�� H2I�
�'�z�S6��&b��P��L� ,��'��ZF�T%��myA�
}A`li�'��1�!K�@�ڃ�F; �ٛ�'����E�%r�畤}}H�#�'Q@n��1��O=�f�3�CY�yR�
 t��B��W937�<bC'�6�y� �0.�%�G�&4f��R腤�y2��+WP���͒�$����y2$[�Rf�y[bHX��P�ːgص�y��O]��ÕoD�4"lRpIZ��y� -k��ڷΠq��-�D����y�K>g��9�ub�<ɺD;�j��y�%�*��g#�b
�KSN�6�yr�X�TjVe�0M�t���B��N��yb��q���
�1Ή�� ׹�y�	��5��A;�&�r�\�藤�yR�Tq ��ٵ��w�p)B ,Օ�yB�.o�IEJנo]D��w�4�yRk����u �6-v���%�6�yB���5s&=�soP��0����?�y����&�0P1wBʕ�(��� ���yr%W�'�Z��a�����F��y��[���Ea1؜]�4��y�ƍ,~Z٧��� ]<U�d!ܟ�y"�ùs��F�X�I��b�l��y��S!��� ��ŸU]�e�I+�y�jR /C�xp�9@�^8*�/^��yBɚ�6y����ߘA����-��y"�;�)S���61jn�C2둭�y�O�LH"y8�
6��Z��F��y
� P�1C��)p߼%��D	Pw���e"O�P, �<J���p��jFd`+�"O�S�lO����AC/+O�䨆"O�$���-u=��`��. ��"O�OS6&kB�zWU�Ipa�s`04��Ag�h���I�P4��u{�ڝDq�L���IDA
�H��i� b���Ze��cG�J��i�m��0��x�#۬#�O��|����-pΙ8v'��)�J� �[�h�s�q�S�O�x�1Ɂ�Ҧ��B���QRݴ6$=�����Y V�L�B�C}_ ��U��1��j6��*��AؑkvĀK}2����Lg���t���,̛uB\	�Rw<
�
��x�E$��O���k�!F��D	vxv�2
�>�p����H��1���2��I��O�wW�t�w%Vئ�HЃP\�S�Oj峄@�2 ��}����2���b�~�YYa����g�s��0Z�;aO���'�Lܛ��%��~8ې.^�O`�ݓ������u�E�{�d���y2U>۪O�p� �Z!u.��7j�> b�YQ3O�*A�R�~���'�"~��*P-O�� ��(8�b�0!��{� ��DkЈR��0|ʤ�J�W�.�s���&A�p���M�L�0s�y�m�B�O���r̆�҄e"H5��A��gK�����)�,�K}:d��H�em�1!���y��P XN���=[V�ljf�њ�y��,w� ���V�Qm�i��F:�y�`��SB^D�C��A�ɀ��y�"�&�0�S%�̗ �NA�c�@��y�jV''{��z��]�}�6D�BN�.�yRNWH*�	�eÌp��%�%�yңgY�=��/��j�T�A��@��yr�64�N��S.�i嬹����y���5���C��N؂	h�	��yR�GVp�Ts���F�+��C��B�	�*x���`��jO���a�|�tC�	�H�mZ����t� q׆C�ɵ*�T�,
�$��P��f��w��B�I�N�P����[�#QP�H�G	���B�ɜX�lAh�Q�X���7��'��C�i�<�SBӚ|i.]キ�F�L�	�'+� [`�T�d��+�/9Q�Y��'mL�1��V�5⨜�1�*i��'��u���_Uś'J	����
�'���#۲rD���k�����'':Y8B�ۺ,_A��	Qg�H�ʓH�٩��$���CF�;�P���x�d[���wA�Ykef��$���ȓ6�^-����i���v�i\-����Xˁ�F�rbԍ���̊(^�H�ȓEY\�i�ł�xt��0�
K��H��j�:��-�\��C�mH���ȓ6g�  �9',(����<.vd��1���H�8�,��޼idx��ȓcE�3�M�0���;CA:\ \-��Td��+��Bx ��3
�*\<�ȓ^��*�BΥ���F��#1�8�ȓQ ,���k--���z��Q�tv �ȓE[�<(b�k����G/A_��U��K���E�lQ��bm��S�d�ȓq��qE��C>0|r�O_�Et��B�8� c�c�F���X _���ȓ73�HT!�� \p��,$C�نȓMz,��&�A!
�J���yoX<��!b���#i�L~D	'��a�y��8��1�Ro��vQp�lB�$ߐ1��'�ޱR�Bίcھ���EE� ��,���� \܀�i'@�Y3�dL�0L\��"O�(BA��n��Z����B�"O�����9v����Ś!Ba �I�"O�<H#�N(:4"t��DP0\QR�[C"O^ݺ&��!/���H��23l!��"O2	QqN�?2�\Y���=C���"O�$�B��3��DO��k����"O��2E铆R,��Hׯ�" ���"O
�a�N���r%�ь�  	!"O��ďW�,y�RБY�&��"O a�f�֨P��E�&�HiJ�af"O|�4%�.���b�55��"O�a��o����;8Dt]���:�Pyb+B�*��$Y�oE�*�{Ќ���yb�׀:D4h�u�9������V2�y��T�g����D���=�eLĺ�y�ƛ-w�0�Bߧ����A��y��۳V�t���?����\�y$�!Z� e3%Ei�`P&�=�y�ܠ-������^E
���yb��j�Nh�l��{bʉp ���yrg)T�X*"�`�U�6�7�yDT�c�=k�`�̑Z֮�y&6<��T�'"V�,�2K�y�dۘyy$�飫��0敁ADM2�y���V
|���D%W�}�w#���yr+U� 	J(��3~X��J�nڗ�yBꝶ4�dXa��h�ڔ����y�PB�hh�A�8g}B�{rM֜�yR�\!Ѱ����$cM�����E��yҥ̗[�0-���Y��`�K��y�	7R��R&o՗��� �
R%�y" 	[��#*p#���@!-�y�&�1�h��F鉼d��x #X�y��S�"1j1�F��]ڦ�0&�G�y�-Ђce�����,g�Z�"� V �y��Z�/�&(��Ñe��,XEڿ�y¯�`)v ��fT�
n��1 
 �y�N�5>q6#{���@����ybj��?�T
p
�q�ܸ�U�^�y�IM�*9��gʒo4�|C&�ϐ�y�l۬+���аE�7fHH!z�HҢ�y�Բ=41�a�0\N�H`p����yrB��F5F���&��@r�d��y�?�Pi2(�3SB]��H��yb)RV��rf�C�=\�3F� �yb,� b���4:䝋QoO�yF��R�&� (;�0��S
��y�m-\Ą����"���e^��y2���O븭�+�qd|	k����y2,��~�)���۠bqT`��3�y��@>v���R�LLC5��:�yB/��t�6�w-�7c����ĵ�y�-�(*$����G�:���,܎�y��
y�д� �l4�D�;�y�F,|H~E�D�|�	�Ɏ��y!��h/�K�B��X�jSɇ�y�1��H�Gφ{y��
b�S"�yb�ތ|�:�3�Z�
� P�6̙��y���^԰l�ՊL.e覅��yi�4Y$ �Z������I�6h���y��_�,�
��!�U�_ԍ���2�y��)RL4p�D�$	��M��y���8�'dY�|��"sfK�y
� �8���� I���Em�}ja"On)��AC��|9B�e���p"OH͸�K�g���"��PAJ��U"O���7&�n� hP3⃦97���"Oȝ�	'O�Z�%!91u ""O��8�n	j\S�OP/}@H�q"O���'�E�	�>��b�A�1��"Oj0��%�'lJ6%C h�8Z/��i�"O
��'���B�l0��ı�ȵ"O I덩[&��r�G�5_p���"O���d�35��hU0ku:���"O�M��[q��Dڐ��svu�"O���I�-.�z��Fg�\��"O*q���c��ܪ�G�)�`i �'I.�qj׼] �Qa��+p����']J� u��@*4�"aOk��Y�'|�t��0Wv<�ē,]
����'d��d��/XxŠa��.h�ʸ��'�	jQd�-rr�Rr����	�'�0���G�0� x��^6
�����'A($�Y�'`� � c	tXQ�'D��fH�J�J��%�łs� �
�'jb5#���	7*�1(�?v�@�	�'��4	�i��d6
]5�$"��	�'��Ҳ��!+x%��Z�-,,]��'�5��G�)21jS�U�%��0�	�'��;�.X1|�2sm�>���`�'���"� �� �P����� ˇ��yRON8?���:�X�]�r\�v���y"��7�R$1�BL�O����u���y2��"$��(M u2TA)³�y2CC�Qg��:5
ڊs������M�yX�a�8��M��Z�Ā�b��yb/��S��yrf.Y�X�Q+)�
�yr��G��1W�V_W�1m9�yrjȗ4
h4� �T�V�M*�G��yZ�P ����[�h��2o�hɄȓ-��1Ud��:|�sǅG	j���ȓr~"���-<��}��O�)d�\��!��P#R��[��	{f$ v�ȓ1?��4eO4`�T�"U��|h&��ȓ�8]:�'�-f�\�t�ےj� Q��}��d!"!���Jg���F��+#�H	]B>T� #�:�ȓ:s������JEz�H�B��ȓKc������rr �rjP��6
���h��zj�!��#|S��ȓ
�'N�P7�-��{����&����J�uIv�(��<b�>Q�ȓ0d�����Zk���6���<�؝�ȓ�0���#��K�պ1�N�,F���ȓ
�����B� "$9'F��%�Ԇȓ"��1g�P�:�b�-<"49�ȓ|<��80$L�/2`�Wȏ��F��ȓE3Z`���ʆ'fQjF��:-*E��c��P��i�m ���[�m�����.�&q;���C�$ `U��g�B�ȓ�t�����8\�v�V0�¥��Om�Y�%�nl�A��i�i JB���R��H1u��h7hۚ^^��Y@"Oz������B��i�gO�?q�"O� oʍ�����׉XM��!�"O4H{g�1mF�#��\1��Qr"O���� :�Jp���)�,��"O� �yje/p�d��[���C"O����GJ��"�٘�
�"O�8��+��c[%�ۼ'j�U��"O��E��VF��R׏LEaj�"O(��U���8�0���$ײI4��R"ODЁiӥ5<%�#9|��Q�"O�Ek��
�t�TИ"�U�B�Z�9�*O�]�pe�%@�Eʐ�ɲ]�T���'ɐ�4�U�xB�api�+C�~ms�'�ԡ:����(�R؀��������'}T�$�O/6=�S}%����'�ICV�^<�^$s��2'EJI��'�Rd��A9.!jr���.�y�'�r0Sծ�Z��pȓ�L0
�'a�( lW0�Z��H�hT���'Ԥ�2A��Z�p2�Ƙc�$p��'x���B�K�Ȉ��Fպ&�a�'��ٺ� �@xe�F�F�%�b5��'S�	{��Đ+�Ƥ�!�ЏM�:}��'[�ܓ2[�pe,@aB�˛Ed���'���)u*�~����vI_'7��I��'}��'��=��ei%��+=b1�	�'��jf� ��F�	�g]39��e��'Ш��S��`M|q{6 Q1B@|��''����gG�[`�kc����jD
�'8 X�W�\��h�?z�h���'�Fa�7�JfԐ*�Í�E���'.�5�eZp��1Q(�s�A#�'��L��/'#޼�H �I=koҁ��'�B��S-�:i�Lcŀf5�p��'p�Dq��,1������,v�*�'��5�$D�6N�Yi�M�<N����'��왆�Ђ./�R�N�/3�uR�'�X��͛cZ�1b�Ql��{$)g��lڈvv�x	���?����?���:�.�Ow�D�*H(�d���]wv�'�:W���af
*G�М�ŋ�xy��r��J47���M?�' �����!��+G�Ҵ9�ptz�C��i�Oؾq����Q�
����ÈO�$1�N>	����;.hm�viX�:��b�B�[}+6�?��i�O����O��)��89baHj}̜i ��2��-�O��=�|��40�*#�,I�`@
�	�ϒ��|4�Imӆ5lZQ�	�?%�S]y"��;�:K�L�<�4E���� G���R�'���'8t�I��'%R�'
$aq�E�	4��X�JǛ`��������ĉ��z�thxS��b �`a!����(O��A�.�j�����L;x2$�$"D
U����Ɖv��R���M�6-�+�Q����o�O�d�M�8lpg�i��Ǆ�kvpnZǟ��'(B�T>Qa���7�uʧFC(E$�%�����Ɂ]��JdO��*�D��ƇM�0��ɖw�$P��4��$ݩ	�М�;�?9������$��@P�t��e�d6O>�Xª�埴�	��DYb��J���t͜�25�!�M1̞�Aanx�q-��n�0��_
Y?0�<7%�<sA���0*��5��aS�iX�����8��h�d؍���!>b�<��#��hܴW��O9��� Tp�h�$yy9�J$��$?�)���ۂ�O�J�<�sv�T(%��((}��i>�2ݴқ�iW2�05#�hy��Z "�b��'�0���zӦ���O��'(���2��?��4A�v�ٱ��m]�ى���[�i����'�~=��@�*���D�}A���-�~��U>Y���RM�yzu�t�� A����H�����D�3<��}R��֦��)�D#�#<JP�S���J0���X uV`�n�3<��zR�iz��H�j�<��c��M{��	+a"0(�ሒ��^�`(��G���'��'����S._�d� ��z�.l;4�=���bٴ=�F�|r]?y�pDR�6��؃H;�F�ud��?	��u�')ˣ�?I���?��	��S֦9:E�C���:ph��9n�h� ?���y��7/��I�� ��%�82�'C� pS�Lo�I�%�d��'͛7�|
��9S�<bQ�K�>@�̩SAǥ#>��6�~�@>T��O�Ҵn�c���J��P$��'���!FM���X8�Jp��<����DU�d:2�で�+!�D�PASBn!�$#7�9��~ Z��ԯW�kW͹ڴqH��U���I�?	�Jy2BZ6k��DHQ�H� ���"�V�t�`����m��'��'ŲtH��'�r�'���%*$T��'á~v>�լI&%R����3��FBOk�P܋�!�(O��f� .� !��<20��7 P!0���Q ]&�V���%�I��K`�%��X��I�'�(�HB'��X�����Ex)k�����?������	;o���S��]4rmf�T�T����I�'��>a���ֲW�������5?���dɮ�$Qݴ9��|"�'r�x2(" \  ���ڴ���������M��* >  �H�r"\r��Z�Kf�y�{r�'�ay�/ͣ8r!����E�h���~��I��M+��i��'i��8�B��z�pK4e�!`�[��?���䓲�O����  �E_��[��i1��'�r�J��Z��'���'�R��ސh�̓�	 �����,n�"s�G��Y��ǟ�UP��擯x��Oq�$k���\x��;�Dm�=?: � �/�1/���@-�P*iʠ�B�z8��M���O\�Y�F`�i"���I����AW�y�`�ဌ�&p��vt�`��ܩXu���Y�Xm*���S�cy�e�FMF=U���	���>�<�2׃ �*���S{�r�SD��L����4�����'����3,p�xaG��kf���) ��!�OAQf�  ����7K���Hr�4sꛦ]��o[3�M���?���.�0o
�@%!7��.��5��B<k��!�	џ�	7W��t�f�P�>��� g&[��u3�N�_���׉�!e��4#�ʗ{��aIq�#�2��(�&Oک\�$�jG�I���A/O�|�>�!�.�,��@���f�u�D+.ʓL������M���i�X?a��C��	x��q�	��Q�ZM���6�?	����'�}����-�P�hҷ$5;v�XLܓ�hO�|nک�MS�4-^��˗+j>��c�0�0Y�O���O��Ofb���n   ���ՠ*���ԮӰ@v�>�o�-,/�N�
K���e�#'*�mȔ���4�6�'��|B����b�T����q�Z1���<���O�Gy��)�S|[��h�Md
�U�!���'7&6X�%��S@jT�?I�'��}b�bˁ;7���u/��[�QRv(�\b�9q���O����O���ú����?q�Lg��;S!ņWL4����7(�*Ĕ�=JT��L>~^d���䕼$�mz�G�N�',L��h\:�p����C��!�A�ۉ<�X���ٖ-n��IRn_;�p	Q�n�a�'�┠Ы!� 1�BL�L�WDT�n�d 榥�M<!��?��}r�ڂ%)}z��)��x5l�*�p>�O<I��R���H��CWjx���ˢT_�'�26MVצ}�'y
`9�(b�n�o�b�����.:δ��6eS0b$0�%Fǟ���)6>5�I�������\	cQ�^�Pn�6���
DRP *l�4��G��yc��hӀx
�@��(O��QD	�:c�]SE��xmJ�҉��f�@��S�����{��ԍ ����ݴQ���P��O��oڈ�~�/�7�V�S�Nª3��X��Ba}2�'������1�͊p❅l~ґ(���0I���8h�cgY�"���b��L48�J2�Ʀ�'5����>�����I��6-�����V�4�6�ԗ=����ǟD�W.O����P(�	0�X��@>a����I�W��C�����
V �0����ē=۞��b� "2���b'ĕ�b��}Q�lʸ*��'T -!����Ⱈ��ľx��$��i1��O���	�����v�'F�dq81��Gz���돿M���=����<��G���
�#�HPT�;2��n�'���l�>YmW⓿�ҝ�wb�8e@����Z�.�pr�i�2�'%�R(��03�'��' ���$ Q�e����i]���E��(Dd�eY�o'j��ѻ��[�� �O��DON�^���{�E�>�V�M^�$����E�|b���\�|�V��y�t�S!�O�r�#�I}�q�6���5���jOxӨ�G�i[ 7�]�	�hU"��,O�7-Yŏ��̄
f2�2���1$x�݅�	i��КUC�!�/h�# �]�>���'�@6�Φ�%���S�?��'up�1�'�,��9(BCE�[��Y��'�arˆ/   ���5N"����?!�vؤye�&�D�$kD�(����=)��B��ml�ԓ���o�% ��ՃB�\q`K�~����'�A��?��'L�l�Q�;�?����?���q����O67MY1D��L���Z�m�O�E�H�ⷌ��EoP9��+�,z<(4YtO�?Ir ��Z�.�O�JQ`B�FXh���ԅFPl[�ɐ!&v&TՁG�xy^�`�"�(a��0=Ylų�|�Ė4&P�*[��y�3 8u�L�ă�:�F��Hצ�^?˓�?��O���d�"C6��`3/��~p0��3�'���xX3)Q�cftA �����Pö�J��v�m��O������O�6-ȇe �  ���G.+Y�lt�h3�S�Ocx�3��Ї���!���6$x�4��a�z7M%���O��d4�ĥ>!�h  &  �AK̇b
�<0"�(1�e(��?)� AiD��O�6MR�NS
iHA�]@��YЧ�Y�$��ɂ2k ���Qm�n͙��y2�1��]�t�]�O���=o(� ��g߹$�X���Ad��	�	���p� �c� {e�� ސ��I �	%?1ђ��ji`a&Y%.4�$��-�>IGK�֟0�ٴ����'�>͓�M;}�F	�5A���Ӭ>}B�'��@��Z$�-X��(�N�B��J�J}�'�L6����'�<�AnƵ'�Z<3�L�RB�S�L�2yf|�	ٟ��	�z���k�8��֟��	6y�N�2_�Н�^.',���Հ�E����	-
9c�ܪ_Tq:wן��	W�!��YsC\�� ����`�zL�xؔ��K��:��:oXU3�$�UbPU�Û�co�O�
433�ly��8Y�2Т�#�:PJ���OJ))j���'�D)��	�����'��i�(��P #!�H%��/P��r	�'�xA�G�f�d3��!$(���K�O��n���M�O>A+�r�Z"dr�d��k�z�H٬e���0�$F�����?����?�"�����O.��*;�j����Y5cM�r�NX��I����N�R��i8r@h��i72`�U�N]�'<p�͙�uXf�� I���ڕ�!e�!�c����7�,m�*�o�%�(OPrP�i1��3�)����s��n@�����e�L<����?1��'X��l�!C��b )��JT�4�@ͅ�/�jA�D��f���	ăh?"إODo2�M�+O|3��Dv}2�'כ�P� �'Ć�1�x�k�Η&3`����#CON���O��$��k�2;Bȉ��@�I��B�pV
߫Snf��!��+'����%'�C�I�_o�T�V�ͻF�y��ץ�X�J5�ɟ:u���6%ʝ%=�(�A���0JX� �	R�$ܟ�lZ�Ԭ;�B�R�K��ا��4N�`���?�������|P~��^�i(���UK&�|��'��6͘=(�D� A ��$;�H����7Lr��jG��<��	(q֛��'��_>�P�ώџ�nZ����)�c۝{m43�������rt	��F��W� �����&�B������A�:.���]�f�{6N�3}L�݊U��."��WvYb3)Z$3+j�XH׆��T`U"&����E�EӁ_��2��4#<����S�����O�m:�M����H�4��ⓒ)�U���J�3�@��>9����=aA��)=���(g��Aʰ�*�ў�PݴD�V�|B�� ���mʋth���xy��G	Bݟ�&�l��
I�v �   ���;S��A��[�`�s�2��5hĬj�����cM�7�#���d��G�*�y6&��Ȑ��HӘ��D��1�f�O6��O
#}�rAF�Z5 }K���Oپ��Eh�b�d�O$���*` 
@��iǣX��I�$�w�Q���ɕ�M���i��O��F�-gV!�U"D�/�Xt��s�j`�I䟰�	�D�JP�A/Fԟ��IƟ��	w����'1��`r������a�ׄƮ&�T���?}��.�IL#�؟2�i�G�h�ksV���I�f�.)��ǂ���
���L�H4`��2S ��P�� �6�d�y0���Ċ�9��#eL,\�KO�>���y۴�?I��K8�?	��3�Y���	��Y�����+��M��@K�LN\���#\O�c��ڄ�͉Of Q�`�)�]�pï����4�v�|��O����xh\� ஬��%��(�(�2Gbȝ/��C��g��    ��,���!�!�<8h��O��oڻ�M#O>Q��?i�OH�	$`@�?V$Dp���zL�����>�j�J`�O��d�O��$ۺ���?���.�8X��JP9
�6��6b�:l ��c痐��a�3�Ϸ^#���}�&D��(�(O�#��ڸ_�����[�8�,��4@�#ꍻ��V�O�b-� m^�M#���R���(O�5zv�T
��4a%�SQ^$[� ˸g���jӤ�n�՟h�'?�$�'� 0����N�� �qJ޿�Q��G{*�|8��Q%�����`�50�5����R�ɇ�Mヽi��'��������! 6  ����T:T��N����0t��1�M+ �x��'8�_� ��	�	<Tt��e�"]R�hF�)��o��Q�"�"!Z�I5C��9@	�b�i<X6�%�d�|z+O�]ȵ��B⎔��� �h(�"��O���f��O�$�Or���\��D�O@�U{�v P�h�Lz�}�0��-J�`����x���`�i}z�ƿib����|�'��eR���F��h��=�N�ѳ�D	��F ��Z�UZ��ʜ,�m��(OԵ�$�'����bJ�V;~a+g��7:5"�d79�O���O��ʧێ=2 F��3|ƍHr��)]�����h��P�Py�=�d*�<.���#���y��˓G�|pZ�Z����C���mUzb4��lC���j�Pm�����O���Od��& �*`6��C7��[1 �L6-˞�A��٭C��܁D�R�R���U -�~eGyb��zζ`�Rk��A1�"�9=���z7�B�r���3 @�v����!9��HDy"슄�?�C�'����'b��.H� $��H (�:����8������������#�#�ItA۰�*"Fy
ד�?�i��6�r�L��/J>U� �3�-���*�O(��Fݦ�����O�P"��'�¼i��l��d�$� ��A�h.z�Y�i�i��H�o��@�ք�dˇ!�����HS�&�'�R[c\@��E�v;f���Z��]��4%	�L�P�҆[�.u��m�9yj��0� 3�>�>�F���e�3�ʁYF(G-F�7m��b"NӞ`n��`F��4I�����7C^h#ЋZ�$�m���?Q	ߓ�MsĊG;��(	"��!�d���	|�'��6��ͦ�&�`�S����)\5�D(��b��i�O�\��'�a{��Ǫ   ���������4�?���dF��TɺT��-Ee)�)p!��"��'�r�'n��I���)����D)Q�^b
`�'�ўp��4H�Ƙx��e��`;E� :@��@���O�O~"?���
   �nZ�����e�To�H]Z}(�JM�JG�U�v(��
���'�b�'���s,�o1��IFL�)}P��C�ϟ���e����5+��45d�pшD�s��
1��!��T�_}��Js�[�t�$��)3j��DTJV�0�G0Y~����(G�On%�r�'�T7-�Ȧ�	n��Z�+���`Ǐ>���BA3�	П�'��'Ȥ�B�n�fh����19>`�f���w�0�1%$� 1�ߎ6��Y�ɒ�v�c �#��%h��'�2���f�0���'�R�� ���c�M�:����&X)șڵF��.nd �uO^�y:,���3Lj��`��L���O���;l�v��E���(�2(iW�n�Yz�
�M�z�+C�E��uٕ�W>l��$����,�M[�� ւ��kHES���(�4�?��if�7m�O����Y����͸&���GH��p��F/�?�(O �=%?��jՏ�Jm���ʜ/E�TX�?�	(�M[Ǻi��'r�Ԩ��O���^�P4tp�"�M=*�j���^D`�͈ ���j���O����O��N������?�ߴAþ	�*�u��4.)aB��p�=Z����M)m7ح��ɷ&����]�d�,�?T��[@�cEA/GX��H�@��rU^<����VP$3�cGi�\�;'h��(�m8�	
V���V��~�Yb�Gz`6�
64r�Ӧ�&��I���$�Xq�m��Pc��[t�>m��'�O��"F�Ct#�=*�[5e�79`r!�%t�d�O�q2�Or�ɺl����4�MC5z�c�D�b-�a������`�B��'s��'fP�;��'�"�',D�:6 �'��1c�4ev:�����abO��h�.��t�K��M����#0�<��$�/u����k H��!U8�F�j�Fc�(ui�(F
kR1��z��eEy®_�?iƺim<��v(W�!.٪��W�v@˶Ag�$�Of��<�)��h�j�p�G(4������o�!�$��8�3��k���ҭ�r��4ta�FQ���3 ٳ����OBʧXDqb@��'
.X�$�Y�4Tfm@2nB��?!��?���2����b��+c�$�U;�mࡈ�?�uKVm�j)&��7^�6Q:�����'���;'�7j5p52&}ߦ�e�̺>}�\�3_9�4����fhqrg' $Db�����Ol���ڦ���=U�#"�E�Gh��J���J�.�������	�`���RS=<d-ے`�~����O�l�>�M��O� 2�O>^��QQ���,;U��<Ps��!��ßp�i>�A�F��I�@lr'�Hh0�ݶz�@e��	M0At�O2*݊D��=�8�xQ�BHNb�a(������y�I݀^]�Y��	�L���j�@^�
����CX�R�ƽb��yb -τ�H�����n�9��ڧ�
�rVÐ�7��5������?�ԾiJR6-�O����Y��aJ�dQ�₦O���!��?����$ʨ&nP�x�T�5i\0a�KϤ�qOfEmژ�M3M>��'�Rٴ	��l���P_��p�(�N.��O���D)  (��Tt�pQ��\c�P��&�ĐX�'N�=�Lpݴv�$��	2�M`T���"�禵�7 ��o��<	�|�P5K�����X���ց�k�����]	Gq���d/4�	⟠��4C�&�|r\?��)�N���@O�� �yˢ�S�?i��V�v�����m�ڟ`�I�|`Xw]b�i� : �Z� fxhJ )>Y�0y�G�7@��00�Ŵ�`t�i**��5!h$V0-��'��i�b'�D���gي|*XZoӯv #��F�O4H5�F�ϼ���T��M���|Bf�Ԑ���u6�̸�����<&�BNf���%����Ɵ\�'M��ʔD�Æ�k�+)([�D�#"O�� v�_.GxP��)V�XJ �jc�϶�MǸit�'���O;�I:{?��@v�ӛ.��q�X�G��=���9f&��Iڟd��ן���џ���O��;5��>����M�/g�0|��"R�")H��������$]'�`|�'jE
h�dEEyr���FF\:�nثkr� RC^� �$5���Y=E�9#���v1:��i��-t@IFyb'�$�?a��5�����>\�9���"V;h7�o�*���<9�����'�]S@��E��C�gU�6C!�� ��X����B@9��gr^�*wCHΟ8�ٴx���\�P�I4�M���?���V�� �U�����h<+pR�Y�`��f���	؟D��o�)ivʑa�h����=R�qF�R�����NR�d���g�; �|̰��%ʓmk���^]����ᘻ�|L��&�6z��AXt@)�X��τ��(OHlK��'�6�B��y�Iy�dW�_�����"�#A���8�M̗i�,�)��d� �	0vV�)`�	"f��P�d=��C�'�6MCЦQl��[\��a�ۂNn �I�i��>���'���'��'��O�i��  ��HJƧǉ)2<5���ޡS�^1bB=Sz �!ɺ+ܴr�ƹ�?	��B�?���k6%��D-�� C��,��3�'�6��릕�	By��'!�'�R�Y�-[�g�(1rF���@��$9,O@Qk�ɲ8�
��;�eZw��McN>Y"����*O|�2
����޴Hm��h �.J�j��J�|�µ�t�'%��'u*p���'WB�'���ց�j�1('Îh	jD�G��@���s�@۲݂�ʮER
aǌT#�(O����)������,�V �D.ep�2�v.P(��{�u{5@�3�(O�1Cb�'nn6�1$Ā�-��}��i1V�D,	{z��O�������?%?Q����M��#9Xdp��*��ȟ&���-���u���4O �heҷ�M¿i.�ɥkI4E�ڴ�?I����i� \�X� WIX�0��V�0j$���O���OJ��BJ�D��A�i�
	���)
]�S+TȺ�����`�!��o�~�@���o�vD�d���&\((rĉfz���	[��u-��8�Y6g^>ig:!!em6&#Z�0���I�[2NyӢa'>��OH�܃�	
�f�b]���
\Z����2����"|�'}�Ÿ%��g����B
�R,��x�����t���N����@�If2��
C�n�n,�D��5��?���|z�䕧�?����?��4C�`-�1�<^�n���O��>.l�K��+6�Y���s��H`��:C����"U>���1��.Z
i��+�/$U+SĔ�r|m��B�"2L�Ѥ��2*�	�6AT�8>�>ْ�wL-zs+ƹ|p<�ړ���
��D���Or��	�Q�I�IQ�>�trA�b��P:��pl�8m��@��'�a��źА�0U#�7'�%��"����܁۴2������O��t�i}�i�c�$/�~)���
z.j�����O�m;���*�"�D�O�$�OB	���?����MS��rC�r��Qx��ZE��e{0<���S>�Xx�a�b�	lZ�P�^�3 ��]�u�v��b1j����Di�e:�j�!��;�4dT�h���L)s6釓��'���R��!!�f��� ,2p�7,�%����V�I ٴ�?�/O
�$�dA�8��Z�oL&}sNp%�)X�Q�xD�t�
� �n� �%�4���lߓuN	m�l���M��'���?�N�.�  ��G�%�`���[�k��ND�]���8ƄU�FO ��d��4�,QJ�H�~Y�T�-ʓgm�'�V/?���c�j,�~���cݥ)V���6\�z�l_�*X��ug���(OdAZE�'�^7�\|�S�mcU/Q)M.�Ӕ�'YbA
�Ѷ�?)����'��% �JF3}���N�S@bEA�*k��nj��7-T?#<@r��5iM���eF �4��DX5R�i�''�T>)�t�����Iæe1W&Ʊ�X�9� �<~�h�h�#X�{1��Rଉ1jJL{EmKT=@����˱)�80(����~��QA��>xc���`
B+r�5�rHs�L�$���aw�a�F�9ջ��F�D��Z��\c��� 6g��.�3c�@g���4��t�ɇ�?iٴ�?q���i/��$�=!<Ȁ��,Z �0�'�R�' ~M4��rP"��_�K`�P�{��'��7����'?u���[����SJpɢ�#,�΅Jr��U�2�'�]�e�&N��'vr�'��םП�nZ6Os� �D��)+���9��"S���w����	�,'� y�
�S|d���M�LHӑ�J�I9e��؊go\E��ٛ��R&τ�h�� 9UƑ�1jF9��i�~�%��2���O�Xh�� K�8-�z����G!ğP�tN͟@��4Z�(�gy"�'���eJ����I:�ҽ:��/����+ғ�.�*�n	>>y�=���T�Q�
��qBu�2m_���?��|���)qf   ��Q�X��i)	��M��J9���^>!�S�C��E�zA8��4i�!z`�@��ʦ�!���facf;}���"Uq�dpZ@���6P"P�Z�����.�	�iY[�^�&�b���0��E�!c��t�h��e� ���!��Ix���l�3x���a%��TBh�]�V��<�"�i �7-5�D���݄R�`�VlX���JG�M�M>�ۓ��� �  @�?�� ��'�6m٦	�I9�M���2���Mӳ���b^z�1%��D�vHH�-P5=%r��>�z@"D�'���'��$}ݡ�����l�1��Л�e�%O-�U"�bY��ɦjA�����^c��a�1�Bl
�bu�g�"�y�P�_�<g �6�CŮԛ:���f�&FT ��f�纛f ˚w�>�Q��d�&S�Q���O���&�6�Vq"u.�̟���4[��V�'��I�l&��1 %.hf��g	�=pw�ڔ�/ʓİ<�@G+Q$Вu��SA��{R.۞pd7�"�� �$����<� � ��o��!(�"L�쀣�b�)~ P�X���ȟ��	��L蕧�ϟ���󟄛$��j
�9� ѕ}$�⋉-x�B̈�J۴Trp�Tņ�r ��	��h�<A��)fR�m������ !�A�r�i���:b��D�5hX7�[�װ�<qP��ٴo� � D�z%�B l�Ԭ�%kU��ɇ�>9��?9�J~�SU}ácȲ1�`�k�X�'x�?�!�^�-� ���Tض�����Gg�&`}�B�O��d�OȓO�7��&' �  �^���`��mqXe�R�JY��Y�oW8R�d���?����䓒HO�����  �}��K �D*g�f A�eK�2���GX�c�8[%lF�C-��+s��0/]F9b�i���0�!g��kG�V�y����j�ڃÏg�V��O����O4⟒�6=���y< �Kt�25��T���>aN>I���O,4QЫ�=O����!]�^�*-�7aڦы�4�?�u�i��M� l�����<����uㆸԘ�  B��B_�p���.�����y��Hg��X����) ��WhE�9}PL�����Ѣ����@V̄�{�޹���&LΨ��B�ȗEyȠ� �T�!"Ib�Iڻ��@�όQxLh`���,d�1"c��[�b����	*�M��im�D�+ 3�X@���/��A�I�[d@�4�i>=EzB�H	)m���gE�;V������p=)��in�6ͪ>I�͐u�ft�4$Z tPL�  ��$HJ�plǦHN��'n�O�u���'��'Λ�\�;;�ГD(fs�e#Qȅ N�Ȱa�$Y����U�ҭ"1P�0 BU�ʧ�
Rm�jT��5F*�mp�*X'P�L� *L�~p��Z�eZ�C�L�zVN�)=�H�CGg�,qY�O��݆_��A��Q=;�j�*���V��mH�p�F/�<馟~z˟�Ʌ�d����(�E�?-�5���şT���ė��ɁP��O" ӏ�$GY҅(դűs(*��������޴�?�V�i5���?eoڈk�,TP-�u�6��Q #��� rE������?i���?���z��n�O ��zӞX��?Lt�X��)��T���@n����Äǆ1���J�ǁ>�\�B�إx��xk�
@N\����=|�~�wkܮ�
�����M�����F���>6h�6��e<ur4��������(h!S�3F�@�s	eӾ�x��'$47mX���� ��i�	?ty�B`N?0���hP�ϬIm#=����~2�nD�Y���LƸ3E�(z��'#f6�3��릡��ty��L#�N7M}ӲhT V�VL���68��+K͟L�I���u(R͟������2�N�2f��U��F�VG\t挫?���T�~}���i�A&�P�tj��<QU��I��À���AD��6��Qh���BR�ְ{ ��q�lh�faZ�0+�U���d�
~�"�aӈcTlF+>
��8�
̸d���k���
�`���<������'"��0�AB�i2�#aY&CǦ� "O�r���;O����Bk������Q�K�ިsܴ��2��n�OΓO�6ɪO� �  ���sl�=X�f�:�׆b6�(8���؍�0|Z �.T�:dYKJ�e�<�*�ϝSܓO�t������DnξT�����Մyv�Q�e�G���	��X����t
�*e$qH����qLvy�u�9���
E���3���]���C��H�'`�aR%"96mS8|	�"2C�4SD�b�@�rq�,SFß�3�1O����e>�E��>"�z��Q�@*[���0��OV��U�O.�+���
��9�@@��""
�:4�E6e���ϓ�~B(�����?1z\��L�7F�4�w΄�sb7��xk�''&��3���Pt�r;+d��b�J_2IΓ)�´�R�>�i�	X)8�ʧm:{��Br�| Ŧ��$���ȓX�H���hN�SM�_�&܅ȓ3,>�k���jH���󏃋\�=��M�`�cp#\Q�I�f�>�q��S2��0�O/qd>�R�IEeа�ȓ }B1����b�C�4&lb��F�<�1"2�0��O� uІ�@�<���|�ܙ	ׅ�(y-�Q�DEd�<ɖ�U>{���2�F"��m�D��b�<A��� a�E���C�O0T�U�<��k%~�C3�G�~����N�<I�R#.sHu�I'�:�u/^I�<��c�jU�Q'	�6@lhQ�aGZ�<�/�m[�՛��/ ������_�<�7(�8.@��Q�,";�5��N�Q�<�@ܟ,�r�h&�O%|�p�J�ɘO�<�7�]�p`Ԋ� �|�Y2�l�L�<AU%GL��ŻŌ�4@�B��t(c�<q��"G�9�1��4{�����f_�<��U�i��)���7p8ADIY�<�����D�l���/@<�\�7��@�<y��֤ ��:F'J� ��U�N{�<� �@;��F+Kgr�H!͟ju���V"O&,2U$�5"��I��mt�e0�"O�-�3B�q>F��EhC�(d����"Of ����3��l�a�P,Sb�u� "O�3*�]���jS���vH��Õ"O(U@�Q�o���jӏ��u4���"O�H1��T�Y�.��ŀ6uEt�q"O�� ��H6�b�pQ��?0N�#�"OJ<`�A:#P�բ���~��"O�-�0!�70j(���9�R��"O���#�қd���0�B=|z4�a"O��D��m0u�r����\�`1"OP�AVN;��JiB�8ߘ�Q"O���Ɇ���`�g2kÀ�s�"OT)ْnôM|����E�?�U��"O�����,90���]�w"Od�W��e��Aȶ?f,���"O~dʖW�N�f0��A�MO8���"O��;�
��p�,t�ê]�[DN���"O��h$(�q]p�P�J��2(^-�"Or���`�u�6)BCd��F�hA"O�;��"�4K#"Q�4X��"O��'ꞷS˞8㶯�s���E%D�x:'ԵJ�~4b�HA�B�Ρ��B0D�$2g�c��|5$�]�Q���/D�����^���ak-Bq�����-D����OQ���XQ*�)t�l�2w*(D�2�k�6`1&�´��3u렼"D4D��*�M�1c~E���D�\32�>D�@H��RGNt��ć�>t�>D�$`��vL���3~jU o8D�l�f`^  �6E�FO�+D8D�A��5D�`��(µ8�a,�;-�`�Bj6D�pB�	�S�TM;c֕WT]+�5D����>hA�m���#$qA.4D�@ �j؇<jV)�*,�X5شB0D� �i�p̢\��)�.d�V�#�.D� '�W���1�M���Ʉ�7D��ڱ��q�Q��¿\B�bT�6D��qW�����EΟ�'�`�6D����Q&N\\	+���Q��8�(D��zeh�K7&�3egP�2Lr���$D�(:�(�0T��f��b�T�B��%D��[#ƈ"���H�[�׌��./D�|i�-B�{�x	�F�;S�LI9��2D�����(>Y %�J�44LNq�(0D��;�)��Оd�3�_�Q�:��`@;D�QbLwx��1a��(!��9D��� %Q2��i!F'MR��2�8D�0C'غe+8��*�j�PK6�!D��	F��=����6b<"�<(�(3D�PX�k�2���JR�5r�h+D�P��Z*�����F2<�V�q�)D��RE��"�p�h����"-�5�-D��X�L۩#9��iB�ۑ��0AbK-D�yӪ	�*�rt�çە"��e��C/D����.�*lX�hmSpMa2ȞR�<Q �f��t	�,��qP`�r�<�vI�QeV�)B���X���p�<��P�)@\݀��2�9TBl��D{J�26@�҇fP(G�D5��J��y�G�*�ZU�+�iΤ��� Ò�y2��<�b5(��\V�ؠѬ3�y��9|��kšPL,��A���y
� �YA���b9́���
��"O���c�ٴ%g�ĩ ��!򀔉�"O�9����)��%���4��B�"O�Hc(��0,@cV¶Y�����"OĐC��D��-�cm�d�L!��"O&�і�2��P��KTq�)g"O��sV�S�k4��؆��++m��"OtM($�^6W�J�� ��/.e�!"Oʭ��ŕ"K� �a�b���:2"O<�d�!P2�x�1�I&[S@�ڃ"O�hh��ߐu�f,�W/�;!N���a"O❀VBFQz�@����7I>$�t"Otdg.Y�g�rv�|E�4�&"O���PɃ��@�Ti�;.Zt��"O��0��	?w{�N��dL y!�"O�x��ս�Vd`��ĖH�,���"O����n��,��$�s��

����"O��(��Q?��ICA�A�(����"O�����Z6t�F@��Jǅ΀uK�"OFD"�����ʩDi��}�!�"O�4K�ƓT)�]�E�ɂ$.�r""Ol1��O�� ���xd���"O�����]�+?�xX%��om��"O��8�m��q�4��jE�C� �1"ODacJ�:�̍��Rm�$,�"O�Ȱb�LOΘ�A��8�N00T"O6�	��U+D���rEg�x���"O������(!%�@�*�Zp�"O8ѓE��Wr�I F@�f�64:p"O�M��K�0@zV%s�d�N�d"OF�bU�ױW]bx���6���C�"O�\b����,r�F�.���"O��� /���b�D;gФ1"O �+P��$:�у�o
��qa"O��8���0f䐻<��9�"O��1�B�
R���{�`��T:��"O4Iɦ�3	Ly;����S'$��#"O3��Ȣ7|4���L?]�uxT"O&P'�b�b�Jv�ɫ/TU�a"O�DQrH��]7�T�E"=t�b�"O�	S�OJ=ߍk'��7��P#9D��� �بuJKa#
' "����%:D�da�ʵKs�ġv9R|21B!j3D��x6#�GM�D�.H$*E×�/D�؁�C52�a�e#��IK�"/D���S��,;?�"邌=��#u�,D�(U�ۃ8�\-٠A�t~�rv�%D�\Cv�J9#C@=I�dD�������!D�,��j� E$Z��4�ë�+`�2D���AU�y���2���|\(��6D� ���M-đh��������4D��I�iY"�`��"(���rP�1D��ꁣ�r1:�*Ç'g�qCB-:D�|Ó����ĥZ�j�.[b��D8D�`hu���&]��DP��Nŉ"
+D���i�.���8���Yh\e
�A-D�x�!f g���.�8W��ё% D�,��Ő54qXf�@��|��w�?D�$��"	eW�I��w�lL3�*>D��B�ѡ/���\�N�����;D��26�ʝJ�8ɒ`�6WT5�8D��	���'��-���H�B"���	3D���r�+B{�Y�A<4�Ti>D�x���',.]6N^�E�tҰ;D�� ĉ�*L<
�Aj�΃�e��a	�"O��0�h�'!�:�z�L�6\�lyr"O��QV&ۗU�&�R���	qZP�{#"Od,"dk�>B�l��7�4iQ��"OL]{�ɏ�y���K�dZ�;>LH5"O�*e�
f��5�ˍM2Д:`"O|]���@�;s�Q�f��R"�5T"O�lӡ͔4e�����̦�d#�"O~����D<Aać��'"O<}ӱ��0���;3�Z<>��=2P"O摡�B_�<�-b�D�s����"OT�q��M�Dj���^h[�"O.Q�ѯՆ@ZE�vCˏb�c7"O&��g�¬��V�ǹ$���2�"Ol-�$���������[��d�T"O*�AKB����a��!jcX�Q�"O�����sy���I UR��br"O���K
�(�u��?hX~Q�"O^�2�J� SXr�1u�AT����"OB�A���J����G���>  �"O�X��,��*\�@R�V����"O��
S�G�D�H�Ѡ���@hY�"OT,#��7`����Ň�7O��	8"O�0��E��̸�"A�6�����"O\��Q$Ôt��%��k�)*�0&"O��p��8�83�*} ��Z5"O:�J�l��� �7ʍ�
t�yQ"OZm0B�P�)X��I�I�� �H �3"OUY��G6`4d�S�����Xy�"O4�0E�gfr1c6g#(�>��!"O�$
6M��+e�yS�_�S"O����S"%b������"O��SP�Z�x��)�O��:�G"Oµb�h�!Vm�i�Ѓ����0��"O��0%��h�z�"��f��8D��Yo�銔;H&/�.��$	#D����B�l-��B��@�
��]�h=D�L���Y��p�I`_4Q�9�9D���Ǧ]�H>z��7i
��T��D5D�᧠��~*rTA4d�4n�rT��,8D�ؙ��Y��(m�a�?� ��/;D��S̞���`���:j۾HHT�-D��)@Ҽ��C� @�Tg�,1ա+D��$�Y�c��+�`�|X���-D���v�*[\`��\7f�}cu-D��ċEt��9ƃ��/2fu��l�<G��)��L�����R��*ŏ�W�T�ɝ]����Ÿi����l����'�/Q@R��FJѿR�>��>(J|�V"[����r'Ş[���r���DH| @�Ǿ'��$P䯅�S4����gI\�'>NP�sC˧7�6���&c]Hݙ��"����Q!h��t��ϝ},�H��=�Oհ��'(�7�
X?�QV��I��K���'^?Y��?yN>Q��ɂ�G��U1�",&Zdu���҆'ҡ��̢��g�	�H6�QB��!v\��lϦ�'��O��M����?y,�����&�I#��	&����L�]솘�o۟��ɸHK"�������`p�)T>4�]w1�jqV?53A%ʔԹ��`ƀW_|�xRf:�$��9�n\;����_Kv����2-��L�LG�"�j�DF�h���a��Z'>�H0�UgA k���*%�Ô6f�o�	g�<�dئ��+O�D����܇�.�C@I��I�C ׸'���$0�$��8m	�gA�����Q
v�"8E{�OR�6-ܦ��I�Mk�4B���z���$)�lqc��%B��1�zӐ���<�����Z����>6������^�t`jud5ZX��q`aг$!j��	�HAHKua/Z��L�^00o�]��Y�V����":��j�Bέ������n�X��a˨\*���}��X�!��
�$&%ݺD��P���^��;شp����'�$|�������e��#w�ʃHY�����L�33*q��.O��XD{��IM50���uj�PSR1iq ��-��-���-fӀ�O����韴�S�? T�2��L[ҲHc�C�%`�V�F���SC������	�����u��'���'/��a�K����d�`e�+�^8�p*��Xs�G>&3��,Ȼ1���M��(Or5R����25��[	ܱS�C,� Q�P�[&z�`}�d3U��Q+��8+^㟐�ٝ<ْI��чe��}ʰ\���$D��QP���!�IYӬ9AN�A�	�NïZ�6T����?!g�i�OH�=��B�"�x �c�4y�nI�� �\���`Ӥ�$릉�ش���+�~�n�ʟ(o�
��$ѠE�k��թ��
{�(��?����?����?�С��aA���>{d�p�S�X��$M����c/qb�qK�4n�GyBf�'w�	+���CBr��M|`lA0�ʨz��x�˓�E�� �M��I�!,j��'�@���OT@oژJ��$�C�`Ye�d�B�*�	f��$�O ��;�)��$j�p��!��R��9"g�	"���<r�	џ�(��A&��)�
�<.��FP�
іqXݴ��$W��ftl�ǟl��L�/�c����[|��Z1#ƻWa੓$��W�b��O@�:� �*��ƌ��z��Rr	�`a�D�p�~���A�vp
C ��gF�B�P�ɰl�f0� �ʐ��0�'L�yH����O4<�B��O��=����5Y�!"�o�8IҥiI<QT���X�46+���'�����{w�R5[��a�] �(A���O�ʓ�HOvi��K��P��CL�r����'�T6_̦I&���׎/<x���BA�&����8l�\�������O,�Z�
�  �	!�dVC��G�	���˄MՋ|�!�d�"\���[Gϙm�x�[��[!�!�� ��{AO��F�"(;�\3@,+P"O��R&9f�p��+�B@���""O��2��!u	��2�� #r�i3"O���P�>T/ ���X�gZP�"O� �S��h~��'IٹMsb���"O��׼j��be�"l�U��"O���c�/U�x�؜b�$QY�"O�Y�,a�DSG�C#1��̹6"O��d#O?=0��>OD��"O4a�V��)�x�j�N�w4��q$"O�m��C�F�Pu�� ��^ :���"O,-��EJ�-��q����7"��Q�e"O�� �����`TjԺ<��Ѡ"Orq�g%J�e3�i��_��M�7"O�Q{$iB�jxXm;��'t�ƴ�F"O�=���قO��l��̬GgF��w"O����_B4�gG�!;X�!�R"OX� 2c	�EXn����ŝ.<���"O�$��	�|�Q�e�҄2�̓�"O�mk�Y�Q��T�C	��2Q"O*��# Vo�V'9ji��9g"O�`:U��>��*�Ł_����"O�`^(�QC��zI@x��	
!�*_�
��DN�iL�t���t !�Y�h�N�{�&�5Tu�t	��5A!�$��G�"ׅ��А2	݇�!�L�Ab,��@G֡I!"�#�đQ}!��I�-:�лp�ƾT&�*"�ʹc!�$C�Ec�D����-'>�&=DJ!����U��I�%C�C��Ie��T�!�Dٔt��@3C\�p�G�@�[!���7M�z,�poʒG�%���E�7�!�D]�o���ˣ�R�@�<Q:��1�!�PŐy�F-	�1��>f�!�$^<?�L3�ЕR��X���P�!�Ğ98L��I���/�n��0�Lg!��j\��5Z�N��M�.~!��"�^�kf����;�.�6zh!��+4��Z�g�z����6NV�v�!��Z% �ti����W�V�� �K�n�!���s8`����6�T��"��a~��'�ɑ�bV.���S�E�?I�ZM /��5ZEm�x���	 +i�d����m�����̢i-��bG��HH��mʑ|���+[Ov�@rI)��^� �k.[��Pb.	�JY����Z�J��3wm���4�Wc�0+�jaç�f�'���ߴI��Qĭ]>���f�;B���dEr�.�$��Iǟp'���O�P���j��CX�%�l��\M�dh�'�T��A@��UI�"�a�hM��Rݴij��W����$�M����?�ٴzvY�H��a�,����ޤj�V)t��' ��k�cd�S$�&8��V8*�Y��� *N^�Q�G߂,=zUBW�ǝ=�����)A.F���A��P��C�˕���1��ob9q`�7�b���)]�(������9��Z�j��m��X�����-O��Ю�Mx֭���f:�H�Oo��	����?E�D-6n��g'(m*T��%?*��OX�=ͧٛ���z���XW�M�=R l��J��
���7�'��6��XXD�m�����'W���O��IG��q�M^�D���9�cUi�~�y���4	�g�CL���p���8#�S�~�`�Ͽ��� �2��(�08�=�e/�t}��Y-TfJA�7�ߴI�N)8�	X�����G�S���5���M!�Fu[���ib�o:��ɍ�Ms�i52��56V��F��	�@A�&��R��'$��'ў�'j���s�E�[�H��V�3ℙE}��|Ӓ9o�z�ɡy�aY��
s���9��#h"�޴�?!��?ѐ�J�x���?���?y�����Q�J:�^e���Y�q�%I�0�H�0k[&/F�R�阉w���쟰�2�ظx��=��=Q7H�j�`�����h���OӛB��!�կN�6��y���,�	S�D�a���&�Q�B�p����D�l�(%'W ��ɖA���Iܦm�����9y���Q$4��iDh%���Vb��?A(O��$�O޸&>���5áI��<=�2�A�&7U���챟`1�4b���'I�7��|:����IN� �-3�o�`��9��B��$FhEYAhQ��Y�I��|�IПTsXwZ��'>�ͺ��l���U�F��8�Iz�F�`E�>�!�w�Q7��� ��V�h\��̾�L����Жi�6쀅Z��P�-�Ge���f�U��X��	̑r��Ə����,yK<����C��N�Z��%� ��8X1�1ƛ��a��O���3���|�U�H�y��y[�L�G���P��xb�	v�'/���ऋ �����*�4��ORumڡ�M�-O����\զ�	�0n�0!����؞)h�)�`шX��q�������?��0rj0��i�2�Y�"S�Z�B�d����頢,ׅ�dܘwC��V�@(�CLU�'����S�ۍ>��`	tF2m����"k��O�F�9��IJ_F��s��?A��l�cp~b�0 �O��(��7��O�ם+q��ӤO�{m���E:F����l�?�|R�OZ���R�l!�B�?�Vi{C�'%�6���k��I�Fʌ `=��P���wpT�*O��F�sf���9�I �D�v� �  ���͈�	
�Cі�*��	X0d��;�Ld�+�UXJ\�>��U��Nc�4�� �7R5b8���U�N-�3���F�Ħ<Q�����P�ʑ�S(T���	"�ś4�luON(��R�_Z���7w e �Ċ-�*�x�4��[�.�OȓOj6M��9^ �  ���
  �y#���	>X"��׺i���uA���X��E�8v8>�%H^5nd�O�S��U�S&�dY��ig� �W$E5��mӂ�Ez���U�2�n�9}�V�9t�yiZ!�	⟨�ߴ��'���$ٵ��,�hPB�;M1���J�?As�i^r�j�(-n�H����J	�6��O�7� c��� H�~�`u��� >������X�WԟD�����b�FQ�:x�!�L��2�,1�6�����&>�f5�����c��dk�i�/��<y�ӻ��������s�"���.xj1�ef�L��0�K�h�G����
���d�On���'I�6M�/�yү��q��̣�%1b���GA��~��'����i�_���Y�X�t�j0��d�Q��#��D�O���lXU���0��C~���Nғʚ�m�@yR�8d܎6��O��d�|��ӱ�M[�%߇w�\���dw
>�hEDG�eWr�'[`P�gM�w$�8%#[@�\3��w~�8VT?���s�����O:POr�sv+�D�O�@|����D�P4j��$	�Qp��G�LΜ�̧؞5��OW�!s��B��
뤡%���ce�O
@o���M����OනY)R/� !Qc)��tT[�{��'*��`�'*��ҐJK7\2BL@�D��4*d}jǓRěVb`�JO^�#!n:f�,Y� �W����v�6�F��Iq�	z�'��	�� ����
��eO�'p��T�Wޟ�� 	�ٟL�	ȟ����;�P��vɎ=pw=�WE�MѶÏ3f�QrM�[���!��Q�YT �<�#��T<6�P3J^�K�}P�	]�o=���B�Y!�� K�?J�>������!,D-'s�O�m��'�6V��)�.�̈q�����e���}3���՟�?E�$
	0v"�w	�_�@���'��"=�e�v,}Ӭ�[t��1�P䀗s46Ѐ�<�@��$V���'b�[>-R&�ş@m�_�hU�pd08�h4�1#-1� `��������+GZa;@K�T���*��0ᶌ�)��ם86���r�L)O8D�N�0y���j
����'N�D�Zr���H3>�	�@X<4~�J�?�9��K�R���!��bR���À�>����柬�ڴ{(�F�'�>����z��qh&��~R~���:}�'��	Y��Z`d�k9��Ѷ��#o
Qqe�u�'��6�G�%�`��n9v�tin4Ar�L[pk��7���t�	tX� ��� 	  � �2�Bɷ*�pT(�8h��2�I�O����ʦ]k���y\i��8ny���֩�1r�j��?Q��?����O�PY����il\d��瑊���
Fa�TX�<ܴ&:������*U���@�=ڠ
v�
?=��R��0G�6��Op�$�O`��%v�d�O��t��PA1"��R�,���N�Q����� @"�K�ML�-:�!F�4iPĀ���o��O�z��;���{�,iD� ہ
�+h̥���6@��B
))�L���B�H�뎓)i0x��[?�*�w��rRE�G�m�R��%R:��r���OD�oZ0mZ��,��"|���� �|LY );L��Bb��A��������c�^X4\T(����\��@R� !���?�v�i��6M �D���i��`�'�`��ӉK*j�{k�џ�CW�_���	�������Y[w#R�'Y�vE���#�M��{:)`�↶)#���W�]�E�(d%�
A�h�qe�K�0"�����5��13��
k�ӲJX���b�ޠ}��q�� %-9~Ȁķ�R���.�&D\~��<y����ᖣS�+嶴)&�l�=pci�%�?�s�iݒ6��O���?�O<q��Ӽ1�<#�/^�x�l�E�'zay�e��V�j$0��\jTެ�6DE2[�l�L��2h>����ny��'�1̻9
�� @�?GF1�O��&iPw^v<J�o�O�.���I;f��iBda������St���2Rr2� �U�}��Ha��yr&L|9�}��S�u�>lP+�9�?ɧ�X�$�*99��H����	�#?8(L�`r���,ʼSXC�I4�pE���o���Dǯ4�T�aSN�O
�ۆA�+ZE`�c��|Fy2N!f�&M��B 9?G ؛�l �0?Y���!*x��@]���c��$���f'�����- �O�H�U��53W$�F��=rt������J%=ŀܢW�~j!B�:�x��d��)@��!PF]�<���şM��g�ҥ<`j])��g?aB���A�KW�XT�앧h�THS�\,U��ad��;te[T"O�<�N
;9�6Ṑ��+��`B').}ba�	V	��٤2��d�
\OjUi'n?�<���Q�|�!�D�
]M|���
^''RZ� Ȍ�� 8��	�Px�G�<�2i�oD2B\�%j5���y���� g�)!�E<DE��y���1�y
� ������ .:��BR�3�����"OҴa�`аj��'ܼ���p�"O�MCG�	�UAbaco�^��A2�"O���
|hh�֩�#�`aB�"O�م��cD<�H���Mo$��B"Od�3 Oʾ+欙#�H !C��""O��Q�Akr���Q2ZȩW"Od�����2* �$���_�$�94"O��� ʡ%�ZT�bҖ"<@AP#"O`��v�/n�q�!$�$O8��F"Ob��#M:<& �z�d
(9��,�"OPaW[-4�P��̩.*��"OHsӂ�/M�$� ȝ#���#�"OJ	g7u�@���g�/S�"O.�XC닾%ђ�&��1���c`"OdL�Q��*z 8Ղ7��'.Й��"OP�S�h �$W�H22��2BZ�ʖ"O��#�M�=#��bm��$z]�"OL@;�i�SX�Q��!��M��"O$�c�fk��Y��M�&��Y�"O�Y�IX�j�,*��ِy�l�"U"Ox�3����Z�x@�8	j1ٶ"O�Z5ǒj-�hF D{��]�"O���V���u�H�7/ޖ(��Ir�"O.�;����\���.0�R]3 "OLP[Eb�,��@�/�c��)�"ON�3�N�G�5INJ�I��� �"O�H2!��N ��#���Ybrq�`"ON��H�����aĝo����"O�!��G�%��E#�kτ���C"O����� `�����	�&��)��"OrRf�̞=�<�T��X��A; "Ohm	�dBn�(��A��n�zY:d"O�(�dI�8�f0��$p͊�h�"O�	ĥ�sd�8 ��"O��[��&F�`�)5,� }�(�"O^-��HN�?��xRc�ڶ��r�"Od\
Oŉ<�\PH��0Z�b�"O�hJ֮�	O>�m��	�gB�q�u"OJQ׌�,=���y���	ySԀ��"O��D��td2�c���zU\��"O���CfE-@������QV��`[&"O��RD*�b�*c�[�%�2���"O}���R&H���l��\��F"O�tcA�$�RQ��a�+��#"OX����C�p��Y!��is�U��"Ov�'�@�o��@���Ƈm$�@�"OtX�e`��0pj�`�M�"a�X���"O��;���=R�J����?��]�b"O�u�` :s����&�Ř3����!"O��d�@<+�F9A'퓣����"O<4 ��L�ưiq�I�n�z�Rt"O�i!�D�ZG4Rs���Z���"O p�BcR!H�����f�$lY"O$)%�٣N���dVi�њ�"O�,�A�DD<LI� (]BUꨳE"O
�A�D<����(�6TY�ػD"O 	*Rl�`��9pe�έ ���"O��D/�� qЈ�R:�"Oru��M��=:�`I<n�P�"O�H��Ս8#!'o�5_aX�I�"O�A�T)�3�*@�v�`g�%cE"Od�A�-ݠp�L4;���w�e�"O���$�9syPu��$ݳ����"O� � 	���{=T�c2�Lu��"O�5Q���2Xi�	�bW8'ޔ��'��$�qOb���Y�8����P�y,U�H!n�{�c<D���+�A���W����z�#���?y��u3dHIx��(:I�ȕ:vΙ��r�8��0<Oʝ.Y?�x�0�O�P2b)ϐ��PC6�φ���"O� �d	n6<�r�d�<v�2(zv�|��=r�& :�p�O04e�1FN3�q�l�,A����'	B��`�}r�D1�Y�n�콡V�Ź|��'��+���>��"�8r�-uuh��&Suh<�]\~p	�삗���(�޸�V$�[SfX1��"�O����07ʃ�w�|��-<O"u��A��}�h�O���E�P2N��eaBm��t84D�V"O��y7o�1<΀c�0�P$�|2�	4�xRDc�\�O�b�0"�4n)P���H)7@�œ�'�J��\�0�m1�-�Y��8IR�I-vk��'��A���>Q%mѯv,�c�
�OfB,AԾ��ȓ���JGa�0r���GF	i&(�q�J+v +�8^�V�^�.��|c�/�'o�M��00��Ԙ����	�h}d��uҘ�΄�(:D������~e�n�S�*��։�yR�V5ณ�)ՉJ��k�#݈O���ꆜ�(��������l��v(�R=��I�'<�A�DG[�+o `�� ͉�
��Hv�A����6��S�O��@��@ES�������p���"O�E�ѯ� X�8T�D�3F����Y��j�a�,#�%e�'܈L{&�	�Z~���1OL�*��=��u
���j�F%PcX$-�0Z��[�G�Hx��-44�p��Q?0�cEշT.�0�7ғ�
%إ�O*��?i�l.],ѫ`#
�аI2D��2#�YM�����k\X��#�qӠ)##��'l�AL�"~nڎR��Z���=<p�1�f�$utC�	7|D���L6%�.��6�����`����]7
s*��? �� ���I�q���P��%�E��MV<,���A��@iX�xs��U�d0�"ŀ.8f�k`mr4�RゞV+�#�:Ӽ 1��-1*��S�O�8�`A♶;4�ᐃ��}��Ҍ�ԧE�x�@Q����O�LQ0ā:p{�\�� э/�fY��K��?	��H�:�����DA�!�ߝ*�&C>d|���Cdp� X�q�X����j:Vm��L�J��i�&(�zcj�(H����X8)|:�p���#���1d�-[����җ|"$��Y��c?7-
x� %S�+26pV��E� (�����%��9[s�E>_1 �����}�8�˚�3{L��5�'
��6ip�A7y�ȉItc�}��d�8��$��"�hOn���[o�"Dj� [���r�̜ \x�%E�$�UJ�/A��!���Ad�����Y����>S$�#a�`-zSdA�:���e%n��I�Dm�<��g��g��H��$"���S>�Q��tU�L8d�H(DD�	�gg
p+���F8��rP`�V4��Ot(i�w'�q#hbuF��%����!�,O��!UC���
xS��3��h�]jq J�،��F	���!U&!���m�Mc�e9D]�fV�'�̤��Ɖy��d�p��6-�`���#�(���Br��$
�nʓA�~�kҊ,�,ē����h� JG=�?ɚwXH݊�KԨJ��������d�:�'�LIJ�4y��DR�˨^�:48#C�0?�bY� oO��3#B�5>��C�֤K�Hڦd +�~�؞��$H[�����p�6X̬�D���%0�B�c�H�D�f�y`P�7��S=�0.R��ÆOIU�8rr�F�Ge��*OV]c��I��clK>��[J�4:�7����CL8l�8���@8>8u��V�����? F��Є��Z>��I�iv�E��d'v�I�ol� A`dm��
Ӗ�O?7��V26�ёiT�^���0&.H�G��iM��!�
6���(������d�8sQ�-(���y���L����>O��"�'��Mq���RkΜ@�M�5n�нh�36|z�;����ks���eh��$��v�QVS,�n���l�?oN�h�"Oޝ��%ɸXoLP��U ~eڼi�(i\����>q�&1�gy�H"5t*�J�%��QtX}{6��,�y�J	�K��K��%jB3u%
�����jQ�Q�T]A
�bf�X��LZ�%Y�n�"?�h@���hNB�{d�ι��p�< s�X�~$��Z��@�4�� �Lx���%LO����O�xbp:�I�h �mI��d�ή���l���OŲ��,M�~�2��T�3��s�%��=�O� ̀ ���7[����&�X��5IF���a��>y�L����+�����ܼcQ*F�~Ep�Yf��H7%F��a�<��dС%��h!�\; ~��J�e�
I:b)�s�إ#��>	4R(�ؑ{O~
�˓�� �	�J
�vAdt�����p=��ݑ"HI|�<�a�P-@Q="�W/<��L�<y�h�Xm�|�TD:,O�1�1kO�ƴ��K!
�:����B�L�����&�S&L������8���H�>qa&m
G�(�*D�O��%��4�����U� ��r�#L�^0���=�aH-c����5}�3���R��.V8$�R�#���"O4�p�������:S��#,�H�1r�'z T���7s�4�O?�a�����r�	j�m��\�'qB��"�Y�U�.-��K�JЀ�&�t�'A*���UA�X���[Ȫ4��0�V�Q�/b(�Y�0�Q�j���S�Sc"	�`@�-�����%�tr� �腊i�Q�Ɠs9`����U	2`d*�C.8�^q;�C�[�Z� Ơv6��s�Uw���O����BU�} &[��	K�^0�ӓ ��h��a-��BU�וW�ʴH�oK����IS���J�:U(�K<�*A�={pb��֝����\��ځ��k�+��BԨа ,��|���&y2>�!��1�ؑ��i@�<I��nn&S�E�#��ْ��q��p��Ƃ1 -@Dkr�-���O؍���;P�䉨'�.���X�O��Sdh׫I��(��L��SF�n��T���#(r	�����>������!z L�yT�9*�d�����~~�yr'�8/�z��r�|x�4�����P��S兄\���C� ̰B>p[�O�H�J��>���R���P)���|r�R��H��M	� �X��C�Q�)T1�����+��>��,0�B�8����"OZtPU�JOH�r�cܑ�H�V��QC�|�����<�q��lO��x���)%t'ʱ8f@�)P����Ɠ3�n�8��}U���#%p�*$��IV
 ���w��;Y7�",O�P��)�c�OA�5�$��'`�!�� ΛE�	-9���R� �x5޽z嫏?)�8C䉔b?$�󡞨^k�R��^$m��㞬�Bo6W�a��'Z8�V�cak�6�Yy���,�y�j��yf
]9a�4QW@P32G���y��\�&�r��S2ICFq����y��V>2�cS�M?8�X��±�y����G��U5�T�gmD	�o��yR�
On��aʂ�b�jYX� �)�yD�V8<|Q�뚈e|`)АN���y�_��9j�*�3�P�'���yBH*O�l��C`�:]�v���yr��?#�3�� oŔA�F(�yRk�����p�֭]H쐠����y�!�-"=��jE�T�$<�	��yRFδ2��Cq&�yBz=w�P1�y�ʹ O"̫�Kդy�nt�F��,�y�s�}����pdc�-1�!�� �F 0$��6zS��P�A&{�	��Ei�Ñ��S�O�Fy�rᓣ8� ����2�R���'Yp��P��71: 8@�} ���E7? �@��JF���}NL�'��`y�H��Ȟ���!�̰?�i]�QH��2DnXLvF,���_3w:B�K�Θ�F�م�ɑx?��y�G�?(QCD��b�#?��2Ɓ��ic�ӯ3�65
�H9 �R�aBiC<[]>B��1.H�I3�k�?w�J��D�Y�^�\t����<P-���H����[�i��)��j[�]�0�D"O�E��(�g�"�˂�g�|L���D~2�WB������1��$+V�H|KW&
X���w��i���تU����앬=	����g�4.�Ld����Z��$��`l:q��1�|�A�W���4��OC0c�D�p��/�iF�S�b�T��D�'D����BO wE>PaM�����3�&T�h"6��@FR����7�2xat"OtB��C�bp01@=T�,@q�"O� 2���@����/�)"��
U"OFX���D�u��� �.��,r��"Ot��؛
*��� ,Y(x`P�"O؁���@�Τ�D��Zf�0�e"O����E�`޼���wed4��"OL�0"l��O̸ܲ��8({dT��"OܽY�l�%dP�Q���n� �2"On5zeL!>�̪g&J8Y8X}zg"O��v�D;N� 2�
;B��A[""O�|�hF>oj���"�tmA%"O�q��</�L����[��qX""OXI{�@0u$��0�b�8͒"O�RW!�w��
�hY�PL��"O$e+�遰*AF�b�&@�R�X)�"Ol1��*�9m��E{v�8X8���"O���V�?Qt�<ã�ޑZ*�p	"O�#��G�$��肀��py�3�"O�z�ʅ�D��Ti�j"I�!"O<|z�h�>�!�����3g"�@"O���M� �DȲ@'�uM���"Od���ʭg��&��<�B��f"Oe��%f�B	�`�#�V�X�"O�\y�Iߦ�ZUP O>)E΁��"O� (���� EnԀ��]�f"O�)2�E0���!���k3,Ls�"O*0k1/
�8�Y��#�"Q%F��3"O�IڲB�M�����NT$�YB"On:�OH�H���5!(5a�"O���`��A�9y\����"�PpVJɑDp����U�<�1�M�g��^���ú��T?)t�d�"�vS�dhGG�/ �H�RW�H��]��a��C��z�����4+j��'ɣj>V��M[� E�qIQ��ӟ�Ɓ�Gk�!�~��fɉ%mk�����u�ɇn��\�.O�>�p��
Rm��$�I;�Ь?5�:�qЎ�T��06a2?E���׃w=�""��J.��	1�����CEf���9����w;�@c`��!%n�)�� 8n�LC�CI���$O�@q�����O�&�S�!N�X�!*��/�V�3�O$PKD*I�_���w�O��5;pNH$\����QBN�S�:�)�'曖�5H��a�'*�a�e�� DlA��� /"������D<O6%�@lN�I/�����B~|�K3�a}`�?h�$�O���|D�B���z�ɉP�K��y�᧟�Kl���S	!�U2Q����E�ա�
* �����l���ty
�'Y��ԩٺU�,(��L?< �Ul�A���S-O�0��O$�E��� ���R�A�l �	SB4A�	����p,�&�f*U�rN!����А[4D�<1�Hvx�KSN�P>���l��ID,G,��A���p�$���D�p0�r]))#~2S	E O�2�B$h�1@�Фf�L���tS�D��=9 #��Mk�T����X>t�Q- 24|��/S�,�꧅0@��
2c��8��:�-~[���i�P�� ��I�CU�`��J(Ĥ�*I�P���1DM6Y�<���?9�bw�9j	��5�ԓsp�r�
M�v6B��� @�[�L91� W�w��PD��҂>&$�g� |CN�0�'�29�(��C�}'	�'�ČSx�(���O�8c�zg��x��^:a�̥���0d��g&��u�_>��e�5@.�a���b "��!"R,YQ�Y�'��Ύ�ɧ�O֘P��DEk�)#0��Hh��C,O
������S� �OQ>��S�|Uj��f�>���n4cx!�6>�qa�o�+�l)YD�Fb!���%�ʥ��-�9�lh��}�!򄙇8&��z�*٢^ƌ��A(E!򤇞!�d��g+�C�(uȑ?!�d�f��p�D$�A��,�&+Y��!�^WfY
ph����� "��>5|!�Էk��� �4�R�#�M�<r!�D
�
� �굀�4��@��8v�!򤊓�Zq�0!E�L7�d��V@B!�$�l���A4ʑص"�)P#!�� Ty!ԁ^�x�x�@A�z'0q�b"OND0��ԇ9J��w!L�`	6\�4"O��f��?e�:��/�P����"O�E�Pc_��$������$i�6"O\�r��^
f!�덥`�:�j�"O�!�B^1�L�X�($d���"O����G�0Bv�$%�1���X�"O,t�F�0�k4�%�¤Q"O���L��?����3"S1",��"OzY��!F���@	�bj,��"O�aȂ�J�7[0e�v���(l�ٺ�"O�cSK�-o�Dċ'�qL��%"OZ���V�5��Mb$H�9�|X�%"OBs�͡���Q�'��f�r���"O�E��ΐ�3�,�z��_QM:=Ys"O^8���n���Vc� "\�p"OjԳ�� =s��b�GW4|�f��a"O��p	��0 y�4ƛ'o�⸘�"OV�hbD1���E�� �H�`�"O *�FЌy����%��!��#�"O,�I�蒫/4 �¤_*\� "O�����~�@(�G��%��	�"OtD9�� <�� �C]�	`��R"O�E2���$(Wl��%%K�"O�,(��	+{2�IBN7B-��h�"O��e�K�6������K!^}��"Or�;RM] K>$`C �4#};�"O��Q��ҡ�j`za 7� ��"O�	hU䎭�<��7/A�^(P"O�`07$.ۅ���(x�2�� �!�ѝ~<�jK�M�����m��!�[�W�Td2��t��I����"�!���U��=��
���`�J6U�!�ę �3ŨA�3|��9 � �!��4c�f�:c�<q�����Y�y�!��n��V �Yd	@�$�+:�!�d�[0Tp��?�VܺFc�Ry!�$��B�S$�,H��,���{9!򤄬q"�RR�V^�X����ɀE!��_I�vts\�v,���:[
!�Ć�U�~�9��0���Zveă'�!�D��Wդы�nتeLH����%f!�\�<����će����5d!򤞔o hXX�"�K'��20mU?C�!��-��X���h&Ɲk���9�!򤏑H#�����b���M�Ne!��Z*(���Ò.Ԃl_ܴ;� #S!�$X�/-8����E@be�!H��8!�D�1_Tx��"���T���3T�ŀ!�ą"�fY��nܤ�N�ZCk]��!��
�I���G�5+n>|`L�pp!�d��ne�I� /�.5d�X��.I�!�$�F�� ��dC:^�Q�cТr�!��ȣL�4��Љ��)ox�s1�Ng�!�$pˀ@��ĕ<PK,�Ys*�{!��ߺ ��h�dȫ��i����yv!�$�'N��@gG,e�\����^�tk!�Q�����G�o��%	!g� _�!���{�l�KǥK�u �G�s�!�ċ��hAb��&x���#f��!��"~1���k��e�ծ�v�!�$Ȃu���8�`R
wn(�.2l�!�ĝ(5T�QD$H�ŢʥF|!�Dܝ*s&��Ə�dg�Ab��yT!�� 8��D�&8��\����X���"O��y�H��:Z@�CD�~�V�
E"OV�)Tb�a��\�?x�*6"O�����S�dM�"L�
p0�1�"O�i��a�ipx���ߥmZJ�Ab"O"��3C�"yu(-���i  ���"OL��A�n�Q���ɼP1zP"O���-�7˔�+`LA�	Yb��"O2�KVGB�r��<qKÎ.r���G"O�("�Đ�[8�A���K#rʔ��"O�)rDq�,���%޿@m�B�"Ob�����nCxx2��J�mF�P3"O�5����36��	�%Y]���"O�es�"xB���߃ ����"Ot��AMו/�L� �"ʾ'$ˑ"O$��DEL5T��|j��9T���"O�U��ċ4,&���Lۓ|H�q"O�t�bL�𕨕aX�phD�V"O*��aiҜ~FF�b���VT&�`�"O~��c��*3���Ȧ�A�rv"O@�j��ǖa�ʌ��׉X�P� "O��`��_��ɡ��ʒY
� T"O&5A�Ñ{1ru� A<+VɊ�"O�Ł�c�.����a�A��b�"OR��.�4Z_����`E�y82�"O�$r�A�11@�����3n���X7"Oعa3
��PW\a�a�D��H�9�"O:� �K�s�P���LS�-�SS"O�}���!����	�R"O,�Q6���j+2)+�B�*Z$�e"O�� $0C�Hԩ!'I.K��S6"O�����;vn:t��
1 V��G"O�|���ԚG��k���]�Q�"O�q��j��I����tJ�x�&��p"O(L ��4��XK�dC�玁9B"O�ts�X0
�\R�$�6N�ҍY$"O�tr�GΆ!�x��@�zܖiS'"O�pā�'�<��D  o%B�s�"O�J傽}	��T�X�)�W"O�0���#>$����&c��Y$"O�
$�΋%\\ ���0'6�L�'"O�=��^0w����H�~]"OLN*H�!�: �����"OL4�"���AB���paLU��"O����JF�iJ$�'9:�H��"OvIC�A�pT��� ��k��I`P"O"4��P�;�����`X�o��E;`"O|)����UA@8c�o߰ˠ�u"O|J��&nӜ	f._#�腀�"O�1q ������/�`G�lӴ"O�ycU��:*,P)S��)3��[�"Oԍ���G=.f����3�UY "Ov�i���6a��q��O�X(v�@�"O
Xqw��9zMQ�B: 68xU"O\ؚw��b�h�ꋣp*��[F"O����39g��"�)�F�x�y�"O�|"b�Ӝ�՘P�[�Orlt�t"O޽pw�QD�Dk�D��A��C6"O���eB5���c�D�\���W"O 	��ѯC ���G��B���"O0�R���7��1Po�?h�F��'"O�U3o
e����_�.�j�p"O9����*36�8c����8RG"OF��E�@6/`*� 7|��AF"O� �TS�OЁ8mz��b)W�e�<�"O��#�-��K��8{�摈M� ��"O��G��6��@�s�ب��8�"O�9��.fd���OJ�p��5"O|�1��~|���7��9c�>�x1"O����ҕv�r�w��*A��1�"O@�!���ƅ3��I"O*8J��9�BظP&��R�~3U"O��a҈�U�D�S�	��bD��"O�@��!X���Yv��#j�,yP�"O
`����@HfU�&��"4�^T&"O\���H��CL4��w��A�xY� "O~�"�ӢD{�=K��R�2g)rc"O�aS`٠(��S.�9Qx�	�"O�	���� �0T��ҌBP��iS*O���̅p���N��f±��'���"���x�\�S���QƠA�'���31I�SŤ(Y,��:(�'}zm����vt���e��:ԑ��'X�qT�!q�{�+��~}��'�>5�N,J�P���*��{�Q(�'O��GMbX+�|	�'�6��a��5Z�$��O˸��'lxurу�&c�1��IOJ��r�'�qt��u�H�4�@�JQ8��'N^�h��Uu��X���9@�1Y�'�"Y�� "�>�R��iZ8���"O������l�V��o�s�$��"O6TBニ%<P=��͚���b�"O�AXV�B�	5��1뚙p�^��"O����O.���?���"O�yH�MƲ��M����|�Ҁ
s"O��Z��G�M�t��F��_����"O�\ SlXW|�SKڦ��x+"O�"��n���ʖ�nD�V"O��Vb���jE�4�7a�-��"ODAҫQ4H,F9C��A�FL�t3�"OH4��]@j��D�"��$��"Ov8�ҮW�9+�q�gn��/�ZA� "OD�ᠩ�p��̠�'@�Q�����"O��%���bq�@fX���""O�\
d}�x2ф�I�0�i�"O��B�L�n�&d^la{�"O��#�]5AYI�3��VXyY�"O��'��L�^��Ç� Q\��#@"O��#�ʚ
f�b0i��^�T"O@�h�C�mE����PC,!d"O*�#'eP�`�QA�˴:���*�"O e���2�`��nZ����"OrT�u��x�,ѕ���G���Z�"O�Q6)�?�z-�TkL�	���A�"Oq�tk�l3-H%нL/��3"OvL�a�T<k^�Bp�
z(�e�"O�t �5<�F��tЅ/���"O�	���(E��� �*��Q��"O]bBF�o$����3��q��'`ԈA�M��R���ѝ;��!�
�'@Hq��"��ް!��7^j=�	�'�>��  ����	/5��8�r*:%���>��'�\����%rH|ʉ���A�X�ۃb�*z:�sciĺ���?�J>����?�+O�j�F�kݘ�ZP���~�bı$Ko�';���e�p���ئ5�	:JֱC�Xž %!B�&�(٨�4�?�(O��8������O���<i�LԊv( 	���.�n���P
��- �$�;ZJ��e��d@kQW>�j��c_�+R���`['UV�b��6wH<uy��ۡoEtq �0#��z��t�˰���L?hH���DC&$��hѣx��6��ey�`�?�����?Y�	(dig�#����g[��T��J>���IC�8��3�&
��e�@NIC��>�M��i��'��4�O��	�-X&��p@�
3�� �G8�!�f#H�M3���?a����d�|j�O���@�	b��ha�V�F�bq�i0.d^�ca�0��j$�'%�`� Z���=q���8rɂa¢O?R�]��՛P��E*�
U>9:�ۊ��ʼkxj�7N���7�Y�_!�?9��i�V#=���d�&Y8���6e��z���r U3V��|B�'E��im(�pF 5y�đ�Rs*Y`�'�6��Ot%m��M#.��QҦ����<�#dU8zn���,��5�>�+�������'���'��IĄl��t������E�q�b��� V ��ީ^�<�:��<I/.:��'��MK�X0v����1 H�x�T�"7�Ԓfo��h��@�]�|������DƖZ���bӈ��'#R�[S��d6J�c�k�%t8t(L>���D+��xm�,x���P�*1��&@�����Ǧ��JZ
k���ʧ�}S��22$J&�M�-O����n�Ѧa�IKyRS>U�	�cr��K�|a�M���;T����	�R%��)�:r��V$Qa�������f�;��Y+I���&M^-:ׄ@�b��xjP���lTp��!A��F�L��&鍫�Bc>�*��΀=p�c3�Y�_ߒ�:��8?��f���h�O�gĄv�����[�f0�K_)2�!���X�n%@�Z;T���L�.%�џ�@���E�Tlj� *��S
����1<��'��,�~��Iߟ��I؟��'m���!��iCL�8FO�'fHIBǄ�9�m��"Y��$ҲG�1����`ɋ�~�nPx�x��MI�Fk��q���-�FũT�"G�����N?A����c')(H����C_�4�kBiř6���'r�	2mb�d�O��=��HIƅi���F�fH+�G҄�yҤ� b�a��L3pF�4/ݵ����P����'��	�2O>x��ˣS��ԫ�Ǽ/���Y���{�������	ޟh�Xw�2�'��	߄5���ӰF�1��O�'&YT)�1�I��YPm�<�,�SBՊ��O��a��Q(Y*2a�/RR��h6Ą�SL�5�T��K����Ř`"��?!�L=0���4�V>${H�O��$�	�4�	s���rU��.(Z����4 ,P��"O$dZ���2��@�>X��*T�|kd�,���<QT�"�O��0)4�OC�����/�MK�����O�$�O��pd�0���ff_�ڀ��2���%M��ش|�ܙU6�l�?)�x�<	0�Y�G]���!��"�,lb��'M>����ȆZ6X1W"��T�ܳߴ%�n�DyF
�?�����޿kM��x��@.C����aDZ>%��'��'Bl��7c�� �.��'fa5��I���oβ~�9���ɠt�����D��?1/O ��v��Ҧ��I���Oo9��'�
�A�Kǲ	 DA�Ɖ%n�rE�'���"�j$Y�$J�q��!@G��O�I�d��i�r�$��x��1����Ā9	�е�Ԥʡ�еA�KV�P�\��#�)BK��T�K+8����� |��	�Tp����s�)�'*��X(�3�� �T��b}���a���5$C�!�L�jQFZ�RDbd(ڧv��h)�E�u��x4��cJ�Hiݴ��)�.|���?����?*O�L��F�< 8����Ó7.x)(G�K�/C�|b`%ߤX���q�%r�`b>} ��Z�E�����nA� �^g��9j��r|�=a3�[�4w0��e�ߣ��<Q5�iR��`� �'�Lj�*۷F�T�g�Y��"�p����$��\ b�'�ў�3�@�@}ji93O�>"�`��OQW�<�3�4\ʒ�j�K6H�r!E\y�E&��|����_�?`��q�63I�����z����$����	�����ty��$, .�l2���c-��*#�[0W�����=$�s�$���r���JT�����+�(�`iU#TG�)���#�$� F�+;ℭ�vdQ:[�>#>Y�a�$�4ͫ�눚~�R�
��#��O.�d�O�8D�d�AuJqB1�F>hd@S�CG��y��*q����ϛm�a�������'+剡J��@����$��������iD�� ��V
�4�$�O��Õ��OJ�Do>A��@%kiL!<�(��I"h�����*K�
����ф��?����$�m0��9D�C��6M(&�4S(�Av�U�z�(x�TĄrL`�+Td����To�O��D%?�5/`.j����؋C�^���,�n�	K�(a�����3%� I� ��3�O���	�4��`����.J��(��ŝl 
�d�<�Tb�Vv�F�'0�X>�&��������jgN8qjdK��џ���^� jD@R�gqȌ�$���?�O���/L1`�	��G
|�A�B�K��<�bǄҞu���F���h��!`� ��5̂ԋ�5!�`y!U����O���,�'�y�N�K��E�ĳ,'�""!^�yr��J�.�J#n�-�)��כ��O��D��n�N�Z�!��[	[���O�y���'2�'v���a���'rb�'��Nڬfk|�*�	D������hM� �r}�eY�9`����y���6��8�M_a�9���;l�]�$)�>��J�/wb�=�|�<���ۭJIZ���,C�Ȃ��ß�'^�8���?����V75�T��ЀI�a񢐋��3MZB�3_�}�����"|��0����<�q�i>��My�J^��r�3�0.mjݳ�'˯��u��U���'	�'����')�6�4��΁#n��Ԋ#�X	$�<���C=���G%CR�A'E2N�?���a�? �q�����Y��
r���x*�'_7����/�� gV��)a�@�%�ɥXR๘��.AȬ��C�[�
]�G�OJ�*��O2�9�FJ�f�j\em]8,_�Y�0"O�1�0��.fR�@ұC�tRbh2ŝ|B�|Ӧ���<q#�^I��'�2m�O �Fr�V���cߟ��'[)HG�'4��'N��q��g���0d��;Ը0�D�/�}P5�W�$�3ca��@ax�Hϲ#,B<�o��<�l!	A�Ǐ�XY���E82�Dէ݅ka*�q�L��>���Ey��?�Ƿi��6��O�ذeꌫf}� �f��[�BA���<���?IL>E��g	/��k0f�is�uc�/Z7Ԙ'rў�'U_�Fb�y��IB��Ƥq��5e���k�6��O"�l�8�+����Iџx���2
�Y�I9p��I��Q�\��u���W+�i��̟��gI�"j�@K��ԏ@�bq)�	U�f�\]��N�o�T�%6Yi�5��/g����e����d�e����"� *���'�ǡ��%��˚��S
I'�a1�I1iǚ=ZDʂ�jh�aю��	ɟD�t3O^�����8�^��,�2� � T"O�TAa(ôvRfE3�i[<<�x��I�h�R���� 	����� |���Uu����O��d>z���a�G�O6���O��$|ޭWDK�P�쁺d��5aW��j%eӿB)~Cvk�4E��k�C,a4vc>A&������xݤ��g��eր�z�
��;��$�4�2Ih ��( �pc>�%�`[��9
u�2R��H5&���r�ɁJ5*��"�3�X�fX{� 8��z�K2�ZB�	<%\���&-��h�IU�',�\g���B�	���͠�C�	W����'��]�(ER.0n"$�	��H�	ğ��_w���'2��rD4�)"�W�$^R��C0\,J��G�Ü]��ٰc؅z��bVDY3zP�p(��Ĝ4�Yq��֋RA���A�DI�c�`Ť=XBfo$L���!K�p���W�X��� �\�" ���r���`s�'w"�	|�'�Z=�ץE�+�ݠF/��1�&p��'��!qB�O�mp��)�'S���	K>�p�i�S���������Oج��&!eX�g�	��m�Ƌ�O:���I�v�$�O��Ӳ�h������UMӟ@;�K߼P�|IKS(�Qs��	��*O@	��W�R>�ڡ�@;c;n��	��&ܓ��X�lQ:����C�mFaxB����?����
2�����d]�� �mͫ	+�'H��'�$×D	%1���{A��k�6e2	��l�Bo�82���`�D�&���QGŕ3�?�)O�p1�B�O���ʧ�?)���3�p Ct?#Z�S��ԍ�?9�L7~!zqgذB��q�@F�4�����B�N��&�"^/p	�/���I�rȌ����'qG��Np�O��qq�/��IzbD��AK r:zX#�O�Ȉ�'�b���<) �&A��@i� �`\�"�@�<�5���� Y�/G�@E��:r`]q�'���}���c"�QY��N1_��(H����M����?��O*½P��ؾ�?����?y��y7��6f��� �%͉m� z�aS��z$J��A�B2L�e
=Cp�U�����'���*������ߤM+����9+]�1; ��$a�$�{'䎭�n$�#�	v��1c����H\C@l��Oh���1?��ޟ��	y�'�����-]�.���jA�<m�Ů�yb�����dD�=��!bdQ����Ln�����'�ɓ��K�'Ňo����uL\�=j@Q��@#Hl��ٟH�	៴C]w��'2R)1�*i
�IW?d��I�F(��;/H4:��`ˬq��W�Ό��-A�~�C�ֹ(��tjfi�5���o�&$��q�Q��q�W�c��">��$�4�� )���(�BaRD)�)|����	��MC��x��'����>oE�Pڡ%�0B�Љe�Ԏ&'p��D8�ɖ)����g 7_�v4h�,�V6^�O�yl�Mc+O ����Ǧ��	ݟ��VN���b(�@��}����Å�����zj���I���Χ?ӊ<�D�^�N�(a� �I�Z�)�/Ԣz1 +�`�!']�!pb\^����'�20�ҡ�ӫ�&�.����;@cɒf�� 1���I��߃7R��V4{���'��	$.������ C���'�[�}`�O���$?�5��Z>	h�ةS,�]p����O�ժ�"G�X�J���n�7�]a��'0�ɢ:�Z|��4�?A����)Ca���)WԪ��	}�����៧=:��$�O�Шl��)>"��r'���T>��ORL����[��2��Jm�xZ�O����,8�����R�O�U��Z�NIj���"V:���h�O���w�'(����<��m��`����
�7acH�S�<��X�E��|��)
�Mz�d�"fS�'��}���2�e`2�5Y��bWđ��M����?I�Z�*Œ�eW��?���?!��y�/��J��AZ+]Z�(H���2�W�
X|RD�� ��I ���yr���b$2�(W`*`Rj['��;� U��EbRA[�pZ��y
� �8X'�Ռ7��4x.ۅ\����bE(��ۄ\�r����5��Y�V���{���0�M�#8�!�d��6� � [1+���ڇ�K�P�剽�HO�)7���6�HtJ�W	F�νI�֕��}	�,�Z���O����OJ���OJ��r>=p��ɗv�)���;1ΐ�C&�� �����JE�	:CE��a���/�B��D�:i�6�H>-�t���)�v�S�A;`�!�<{�9���I2(�8�+��!`���@��xp
$�O:��;ړ�O�t9��	�L_6�P�쁨8ɸ5(�"O\��Լi�� oά56�)��/�DӦi�IYy�L�
��6�O`�-RN1�#gʈ ���m�y��퟼1gg�⟐���|Z��s����&[����w^��p����TC�� w���u�����OH!����ì9&H5�'�J$�Tl<GM�	�0k5��a��!����-$�G�D�J�X���!�~�ȓp���˒��69�%z�-�?	E�����?q�K'e���5)N�uа���A�{�	>
h���4�?����C8���5U��X -�#6V���1�.bg��D�O�y D�.�\t#�.c��()3+Z8Vz,��.(�7�Ӭ?��R ����T�@+A\~R@�=p$��C���>��g&�:��0cgRH��ځ5� (p�a�Eq����E8zk�	)�~��'��>�͓i#*8��>qe�Ak?�\T��C�ܱ�v��)+q��!�0�޼D2I%�'oP�%	��P�e0i�扔@�ti��4�?��?Q�̇=�~�����?���?��w0p�cSL�q.�9��B�R��H�gC���a�B���<���j�̘O���bV��\?�!�-��{��\f��Rլ6i1�s��M"U�pe1��+V����|B��Ŷb�
�I�g�΀ГL��y�@S%G���$>?�(A��IY�'gl}�C���d��i����L��"O*a5��9C#��Ѩ�?J���R�p��4��Ŀ<� ʗ�}K�#��Ҍ/`X\1��X��Xѧ����?����?��J��O��$~>�{#�.,9 HcS���Q�VT@P���;QFX���-&��z��\x�����pjE�7F�J�t#�"6j Yi�Bۭh+��3�.6�ؠf>�(�\lPG��bٜ���Ɋ%k�5`P���0���P�?ю�iCZE:�a�,A�ps���'&Ү!�!��B�+9��c�9I��Q.M^��'s67��O��Uh e���i���'	�b�lK�X7���&��+=8p���'�2�ޫoa�'��l�og u�7!(G8����7 �$��I�JE�8(�̨1��	�'�*���N6�aGf	p`��ӵ��W`���@��0	�Ӄ2�ta@�@�'V	0�)��֬c����اBV�s��:�U	�������?)���S�O<*��f�H�UN�Ug.}�T��yr�|��i�v4C��
��l���� � ��!g�����æ��ɽAM�}�	�@�Iڟ8�0"Zş�C��&	�ܹ�vʄ�'4YQ��ğ��	Aφ��Pǟ�!�@�E�i��[?]�O��@���.y��\Q�@_�����O�����Ț.��e
��N�#&��lR���G�U��Ԝ��×�
b��I���¹��	�f��̦�3O|����B�O.Q�j�3����N�"�<�O>���0=9#�e�����
9MelE���Cs�'���>)�����S�܉p�GQ�!5|u(�	�?TX�f�'�B�'��TK�*��v�B�'#�'��N�Qd�0�Ǽm@�u)��<R�㣈sO�zb��{Od-����6�D��+Y�K6��/T$x���}�`C�t�4�VF�Q�� �+�d�.>��A�M�%���L#��� (�)�O����ON��"��ĀI!��H���&`l���n�A�<����QYdE2�x���̙gy��.��|J����$�&r��c	�#Kג�p��4q(�I`�!�J�D�O8�d�O����?�����C�pl�$�f�əM�UqS�4`8H@G
Z��̠WGR�N!���ɔ,[��I�m��NJ��ha#�33��U+��b�h!��P�!b����k�'���5N7�eQ׌���"�M�?q���?�"�S!8G�h�&�R�)���i���C�	�k���3O�R�q�Vf�� ��O4�m�Ɵ<�'=��J�A�~���=0����48v�-�F���y��Y��?�c)���?�����Ī���ʙ�%���Hnzi��E��4D������<�<Q�W�B߂�D�B�&���'KZ�=N����e�N��b��[ ~Tx�E+���0��U�I�o����O��A8Vq�����@X�cA����L>��0=y!�!}�f8)�-^H����Bb��؁�w �i1��ĥK]��zC�4&�ҭ��Ay�R�`Ԛ6M�O*��|�Ɗ��?�b�C�N�8p1��T��0�ƠR1�?��Li0n�\jjE�FN�!~���R?Y�O��X��Dޯ9NN�"���dȐБ�O:��!q�\��A�{"H Z&A$�ӂI���z�̥;q"e"���H��Ht�@��џ`F�T�'|� V��p���6)������8"O�`3��D�@ͩ��R�r}^�'�	��h�i��U�N�P�����}����cpӈ���O��M�<�����O�$�O��dgޭ�pcE�7l����0�`��>[�ر��X�0��#�O�!w8b>=$�Lx D��")LMp��3��p'�5,�Vݑa`�|�� �1��D��t�|"�R.f@.	�c�{�r� _+Z2�'�z����Ϙ'@�B#��#r���7���N��y�',��S���7�`��@�2����/O�9Dz�O{�'��}`��M�z�lQ჌IR��x�� TB����W�'���'��mݥ�	����'q�Ut�^�`^і`R
"���Ƣ��P�&eK�M�Yg���d�%~�>s1��;R��="A��=�8i��+$��)*�*Q��p=��
I1 ���fbQ��4���Љ^Eְ����M�C�in�O���b��@1?Q.���+K�p	q��dg����?��#ɺ6{t�3��źN�d��7�c�	�MK���.e��m�h�$*6&���[�mț���6I��0<���c�'���'�]�z	��rq'�_�0��
Ó*�"EFxr�>T#� �Ո��
a�l�0�0<!1����<YVM��u����c�>�.P`u�t�<I�lV.BHZ�E��@���G������O8(�K���ir�}x �;"�Z$$��v����sl=?�(�2�i^�l��3�@�Djq�`_�dP���O �0Ǉی
!(MI��	�Z�5�)§*��)�Fnz��zS�����(�'�*p�`E�DY��xCcN���>U1 ��*�z�[b���Lq��x��>?������	q�O���3Q��E�'�Djr�� �ˍ�j�!���=cRZYI�%�#^,iSm<�џ�����͛ju��`P.E�H�0� ެ'���ղy���5C.���I�?��	ʟ�'u�y��f�*��X�B�@���eZ��[�j�O��hн%�1�1Ob(#χ����#��R�x�����2�qRi�O-VSA;���y���g������-^&���A��?��O�@"�'}��ɳ'ɘ��S+�h*|l�1+ �G#�Y�ȓ�vI�ua�-�j ��J
5��'I�#=�O�ɣW�*�SW��|�q�gļ?z���Ҹ|��$1@p{d48�aR�&�(�m�	 )��GG�F	���;//��W�I�@+8�A&��F3�=�� (����	ٟ(��@��I��s�H�+9�?�'[�u*a���$�V�V�/�fDE|b.�<zj�츐F��|��S>� ���@;���A$�ȸpDa=��Q�	��l�|�BI�)P4�����5����)�xy��'�r�V_HF�`�U�����y^�ɛTFdE��R���Z�^7$RP�I�P!���?q����i�@m����O��H�oڳn6�m*s���G�����O�}�%D�'`z5�̡b0I�i�Y6.�S��+��6#����H�%S)Z�JG�^�^�	�v�C�@ȵd�4�F(/#�m���ԿdGq�\�'��,A��	E�^�h��0:O���'b������>��{1�@�e�T�'�ݷ�r���.��xR f��j߾�� �CupZXF{�f4�O������/N���5�@'�������?I��?7r��Խ�?���?y�����e��ڱE^��8��L�1�:��F ŷ*<4��v�><n�b��׬��i;�I�[�V�c���f
����,gF�!�V�X$��"êz� Ys�`5��46�4��O~��e�0M���R��*\pq������OZ�$?��y�Ie���g&�&;���yЍW%�yB�\�Dtp����,3tp��=�?��i>��	Py� � ;�f���-�)J�fm����y�	���'�B�'��V�b>�զP5.��b!��!&��4A�΄��P���j�*���⚍O�M᥅P����Gy��U a%8Ub�A��J�p�x�"7g���q4I~�؃G���`MҤ�E,}� �Fy�h��?��S<)P�ӣDM3K��1�TJ��?��,�+IBlr7�S�AI�)"3�P �Fh�ȓ7@�l�FHϭH��b��#"��'H�6M�O(˓,�����IK
{������>�U@ 	Z�8˓�?���?aTdσWԢ��EC��}'��a0�V#}p�h���[l�r�؆ZxDe�+O��1Dy���og�m���h��cqc�6t�
�����m���ӴPx���A�
2JF�9Dy$��?i��ɘO��i�IƼ�j���$��4�-O2���	�X�i)Dkt������}�!�<	g&�(����S�18�Q#�őfy���z�R�'��Ij�T�'�2$�/q_�@7 �9%��4��@�<��dNj,$R�jG�H��Ԃ@ψ/G&z�Aw"��O�&����:��spJ�"/����'`�����Ʒ0�dۑ,�v�&��垶 {nD�}��� &��5�D�sf�EA5K��<Y�M\�x��X~J~��O� ,��bAz��u�&%�$?��6"O��z�	�..ʐ��T�7V`d$P!�I7�ȟ:�;���M�q�Z(
�8����OL˓x�4I���?9��?�(O�	�� �d�[���6���:V$B�0w�iC3��O����s*�tJ!�?#<Q���L�JS�eDj��b
���
���}3��%�1u�M��O&�1���+ɰ|���u��]{џ�|ᐯ�O8��9ړ�yB��=��i`6�B�.x`��)
��yB(_�lp�@0�G'wȭ���O �?1��i>���}y2��Eɔ��A�ӓ�X0��><I\tZu�'D��'��U�b>!�#R�<�Pa�ڧ_����6>�^�w�,&�8�2c]���<q�����xU2u/ږ�R	ʃ�}���0S#�&`�2���;��<	c#��0`Ǫ �΁q��9j� �����D{"�I��r(�E�Y^b=��nXV�C��yގK&��P/@�'����ʓɛ�'��	�x�L@����f>����K-5pȀkS�(�Bd!���OfTЧ�O`�$�O����B��7]6jҢ�0)�^��i>��#�]\���F���t_P��'�>�5C��l�d�RȆ����Z7�!)�f�xg��c�X/�D�!�O���*擟a����_j���4�țp�0ʓ�0?�s�tu1�=W��VH�Cx�)O �i���}�2��ƣ\�7�Y�rR�l��Ο���Z�'��DۼQ;��b�A���'ȹax���-5��$QRd����/M'⟰mZz��d
�O�Ҽ{姉4���3#�1&��9�}�Z���9"�d�ɽ�l��ON�)�O��	�v��5��J��?"��E�<H+����ܦ����6��E���<�U}nz�M�͟k����:5M��t���͝�H�K��?QG����y"��,�$�Or���Oz�I������
P��ZAO޶S�h� С�OT��/����v���
�?7��B������Y�@4@Q�J$fw��[��gL�	ԟHbǸ����O��$�����͊Ft����`�u�o�.`?ry���	�B�$�O��.�t�Dd�8H�k�?7�� ��;>W��Cc✤KZq�㟣%`�nZ�<�ԉ�۟���Zv�'�?������_�dҨ�2� Ρ��Уs�2=	�@�'�����?I�����h��r���?im�i,�A�G��%����33�&ii��ԟD�@���ID��/&���?��AbE�����2)t����%�BZ�v�H0k��DN44��'����'S�d�?)��}8���_T�� ��͚B�|6m͗]���Ĵ<���O~��D�����?��B����jY�bO]�::T|��)�*�y�M�|�ܐ�D��6s�1�c
�$�M+���?Y���?����?�+O��$�Ok씰�Ȱ V;HVL�8��K?�	H�	��'&�h�	� K�ɹ�A4(�b�X�!��W���'Ā}"`� AĔ��OB��%O�����!�pRׂ@�8@ "O6���催)��<�5a�1+$���"O����j�b}���R�|'���"O���E-�lJ��$ ʵB+L��t"O��l�"0d3�Z<�|yQ"O�}�w�,i�0����
k���	g"O������l8�)�m��G]��a"O��6�"v��U��K�j��њ�"O \"����s0K��L����I�T�Iß��I��Ԃ�l� �x|�F�@^h��0+��M��?����?	���?���?����?���mL���HV(Ci|��S ���&�'��'~��'���'�R�'V�	-u�r=�fV�L�T�'����6��O����O����O��$�O��$�O���].��x#�WY?��[5 J+0�jEo�Ο�����X�I��X�I����̟H�	*�IKF揠a ��Y��A�[�V��ݴ�?���?���?���?a��?i��X�0i����>po!:���01��Q�p�i9R�'�r�'!B�'���'\B�'����M 3�=ⵆɲZ4��bj�6�D�O����On���Oz�$�O��D�O�b��v&���h�@���JNҦ��	՟��I�$�I����	��x�	��N"Y4^�Z֍�%$�R�[��M���?���?���?����?����?�$+X$.R��ӺM���X:f��V�'��'1r�'��'%��'����,a�6F_-'h��S)�9��7��O���O ���O�$�Oz�d�OT����RN��v��PJAGG�)ioZ�� ��������P��ϟ|�	���ɤA�Jx�4���0�/=$���	޴����O��Ɉ�m��鉎~UiN F��0!'�v�Z=1P�D ���M�'R�(9����x� N^����7�'ۛ�0O�S�SMIjDl}?��b� 
dE"Ⱥl������OƟ��O �R"(�놌�o����1Ol0�o.�i:U�Q�c�l��'0�	m�I��M���h̓�� |� �?|
�V�j���Q���syb�'�8O�˓q�Ra���.	|��q%��Q_JY�'�$�jg��I�L�!�O�i�&�H���y��6g?�S'#T%$�<�1Î��d�<9���h����0[�t:�g�9� �t�����oӘ�cu�����4�������*��$mZT���bf�H�z���O�7�O��(
b���I]�,� d�]02�ݠjJ�Hy�ԇ\#*��FLZMF��=����"�
y�l��������C1�ةNzʓ͛�L���'��1ps�@8S��h���P�q�%ːEy��'k�V<O("}J"\�Z�P6(G��H�����'�&q��Zp~��7@b|���fNd��*%�X�M��ᓵ�+���%j8����E�<	�eD�f02\`���%W����aCJ�V���ӡ��$URX	��N����"�/5����|o�L���~������
�+,�`�gϱVRd @�+�>Y"v`��E�H��f�B�jY2e��2C�9!4a�+f%Jx1�bgm)�� �7�p`���?3���F �3�ΙH<<`�Q�����({s.�1��}0�d+"Gzࣵ�$a�@%+Ec+^��5�B/6D��H�m�P�VݣLG��XPw� ?�TcX���म��q���q!��H!@�D�R`0�����Y�D��L
B�F`V�+���r��_�I�g�ISp�5[ϖ6-�`A�4C��pr����f[��D9����Nq���CI�/$��	�&Ǜ��j��ƚ6�@#��#TX}�i�|XU��O2�PYݴ�?)��)��J�ሂ/��%f	BvXy1��?yJ>9���?��i��?�O��I3O��r+�K��F��?����?�-O��8�bNt��ßx�Ӣ#f�Żf,��~�l$�4l�&��%� ��؟�����$%���>���_�NP�=�dM�����ĳ<y��X�]śW>����?1.OT�� �6]���5��-,g�u"��'1��'m.��P�'�ɧ�O>�)w�� 3�1���N$-^|h��7��I�i�����S���$�O�ܚ]��M�Qoш(����qȠ\��d�.y�>���O���1�SПD�	�2�(#��1yͰpT)ˁVj֌1�4�?I���?�W���J����I�O牦f��eU2~}����	X�k����OH��O.T���|B���?a�����C$N�<�w ˑ�����O$�č#H�l�ş��O2Y�<�I�zC�|��L���ޟ)��+��ݟ��	����	����I����	V���'��i���ݯ8Nd�����Utu �j�O���O�O��$�O �p�eY�4�j�@`�G?I-����%��U��Ķ<���?�����$ʎQb���`ɒE/!��àB�=����?Q����?Y����b�%0(���N0=��PP��P�lk/O��$�On���<1C�[	q&�O����d�G,�,�E�� E��r�'G|b�'F��>P2���X#ϝ!Y�L#'�H0W�P4���O��$�O��$�O`d���@�u�	ҟ��	�?�&��	��k0��},�mx�GScy��'9��'��'	b�'�Ӳ2v�EXIT!
����%6�d���O@�D�S^�Un��L�������?��z�\�3mD�A� $��FR�vw����՟����P"5��ڟd��k��*.�)��T$l?Z�iQW�{<�t��UI�y�ói�Iԟ������O���9����d�+D��k���%kvl��S�cP��$�O���$�����Ɏ�Hq�� 1�}�����a� ���4�?i���?�'J�5�����'
�G�B��8���D
�a�֪D����'���'�,��f_>a�O��=O8��ō"m�0h4��	<�.iU�'I��A�����$�=P�f(��ݣH^���,�D,����OܲSc<��ϟ<�'�_���(ȱhڮG���"�-(�ԡA]��	����?���?Y��?5�4Rs A	W�:d�vH��4�LqFx��'F���t�� �|�Q�� |����O�n@����N֟��	ʟ��?I��?��+�F?I�E�X�D�@��� �@hAW��̟ȗ'eg���џ��4��t�{�,
� s,`ע�ҟ�?Q���?iV�J̓�@�Q,Q93,���C��z��	����?�*O��d�x5h�'�?���y���>a�h9�/^�l�$�FLI>���?���R���<�Οެ��a�F줸1�[e۶���'��e�֦��O"�OŶʓ.q ��ZШ�G��K����%������Ѓ�F�P&?u�o��'_s�t G$�?XL���2[r�W�uc��'�"�'��$V��'���U�<)j@!�ƍU����?�F�>���h�0�d�+��S��� �0FÖQ��n�ܟ���՟X�!O�9���|���?���$`;�Q�7N�S�0��ʑ�?i��?���>�4��+���'}Xq*sgQ�I�hM���Ù#$P��������&ԱC�&�A�c�1 "�s�iMm>ze�4�'��'��3Oz�:tDF�n�����[�R��Iۅ�|��'�2�'tB�'B�К'2�W=Xx����:_�.$��J"�'џ���ןx̓���֮S*wâ)f�0��G~R�'��$�O��d|>	9�E��k��� "ˑ��nl��c;��O�la��8*��)���O"������S�&-��D�s<��J�͜�C�I�:A�MaW囂�j9�F��V�Rc�pX�:V��$i��\iD#�A�odtу��M�lP"��4���;mz�R���(8F��ħǭG�ryX'�*O�f=�B�3s�,�������'��6>\H�G�|�� v*e�?��X�7�t���͂�]�f�#�k��O�d�wi�3��`+v��)<�*��HV-:���u���e�Չ��F&r����/J�I��T��?i���.؁��	H�L���PG��q(�?��O���:�F� ;r1"p�A7O�\Q'�+ .}�ޱJ �S�3ĝ�BFZ=\���\>��≟?2㤕� 
0&�!kT�.�D@`�2�nӼ�n�؟��~z�	��hLњB@Px)�q[��ߕ'��'42�'�P���	ԟ��� �t�g )i�0\�G�x�!|��LmZ�� ܴ�Mk���/,@HŸ���7����W�E?'A�7-�Oj���O�̉�b��hU��d�O0�$�O��X�n�P%�S������ nd���f"6f��Vȑ2F8�9�!��O~�6����?�G�V#��dy�	�DC h�_.h{�5x�	�
g�L� �Bǘ/D����D�i0(UϻH(��Q+��(ܐA�ꈓ4���Gz���'@��	��|����'�8�
�o���I�+�&Š�`
�'� �"�\ i�� �H� I�D�����զ���~}B�;g� �p�%j!4��0��]DBp��. <�Z���O6�$�O*�;�?)������K\��]�%c$�V��!*�>N����^�iE���K�-��!┆'�c��#.Ѳ{�(4��L�g��� .�88�t:[�����E0>����1&���Z��¢g2Ew���GH#T���-�O�Z	b�T����
�o�&E�� �y�!��<ṱB�*5���	��[�¸'c��PdV�M����Mk�C^.7�>�fb�: ���$��F{��'��*��'D��'��<hU��5)Bt����΂u:�[��Vap�l)9_��RҦ�TX��S�Ԑ{`8��F�9�R�*a��&!߮xi�
�z<f�7+�$�����v�Q��h���O�	nZ?�M��4LX��pp̄>!��!�3HR�K��$U�Drߴ��D+r��4֧tch���.h�Ѐ���x�*�l�F�+U��3!O�A�#�)�V����i�ªi����@I�Zg��$�O
����T�F~�ƼySO:mh�Mx��Ё*�@���iLٟ �� �ԍ�R�� O���蠩����3P?��O���Ѕ��) ҭc�m�h�t��K<a5��1l�X}[ aT(nD���Z,_��S�|I����?�P�9�O!�t�'2��O���t�fm�C�����U/�h��"O<ea��P�d�Z�ٳH�9R��=X��V���d�&ʓ|3$� mۙL�q5�W�)x�g#rӬ���O��OPЀ�O �d�O ��wc8�����i���R�"'$�H1�p �6����U�aӲh"��,t�t$?�CN������^����1�	89N���t��fa��MW�M�4��)-�6�`����i�k3�f8�"C=2�pd^6)��:�j���M�WW�X!`��O���=�����mڼs,������h܋a���u%�̫�'(�����)=�L��G�R�ԭ�~��'�X���?���h}bE�8��@)�%V�S�=b5��:6��6�%7T`�$�O&���O�D���?Y��������%Cw�T7�4x���� �@��n��`��`	�(�]���P%2��bw�S�b^��>\���k@N,LO��(���K�0���R��^������R���'L-2�l�;���Ƨ��B�Y��'y�E���S&R鐠��!��_
(�{b�,�	0 gr@"۴�?qߴt��Q6 �-���j�d��(�qJ��'�Z5 Ab�'��)U3B�"Fi q$�MY�S%A�P3��cw��0=�I��	:Ⱦ�:���-����� "i�ј�U ��h��19��Q�A"@Y��ß<�'�:,(Ї
��!޺�� ����~��'�2��I�,���R�I6���A?2����)F�<m3��T���K�2p����'���V�����4�?9�����&}�&7M�]��T�G,]�sw�� U�Bnz$��Iݟ�X%af��@��Od󄈀��P���	�~r�	��ZT�!i%F����  @�	���aHf��" �xeA�m�%$�ĸ�}P�
�NZ���"
%p�ȡ(Oy�!J���ަ�J|�K|*�*x�=�ѫ��MҼ�Ct�%�qO���6�d$���LTvE�ԏ��d��"��c(�����!��4��ah����R�bݢIq�!0�T��h�N�D�O&�$T�j�����O����Ob��w�H;���`2�qg�(���	��Ťz�D� ĉA
�(�o�b����']����D9��X�F��#7Yr�c!�T0:���؄Q�̐yg�J�ym^�>=�@Ê!�y'C��N`�&��8b��Q0L*N2��$Ty����?�}�I��n�B�@�KT��!a2�[D�8z���^eqO�X���P�	�T�D�1ෝ>��i�7�!��?��'��Ipr	�&�b�±kI�fb2�*�)ݺ�đ�O��d�O��ďݺ����?Y�t����%�/��C��DT&E�ÀȷB^jH��(6-���"C=,O&P9 oJ��p}����S�����2����-;����nPsX��Y��ҁ�j�k, ܅���^�X���O��n��� �'-���t��j��"t-A4�ʸH����	�$��R؞�K �̓i�N-"�[��&m��	>��s��&�w�˓"�u�%�iVұ� 8��wX�{��Qu�Ũ�՟����.!���	ϟ��I�Qm� ��ÖxL9�k��
����5K��	H��6G�#Y�����'^R�k���W�αh��#A��y#�ߢTB�W);9B�q��."�4�K���
�4��eh�P�oZѦ!Z��X�e#�%�rh�q��Xql
�����-�?���)�~���¡A�)tYd��7��$TC��d�J�=ZPk˙d�aȥ�uf&��'E�u�'�>6-�OP�$+�Y���t�^�Ix�����}�zA�SI$D�d�B��7ӒpH�,ԉK�rUҡO4�	�u�4ը���3�ʀ�fd�c�P�Ol� w��(y��]*rHH�7���8�"OFX����&ܺ�WFƽw�h�8"OHVeթ1�rR��B4}�&��"O��
����>M�.4e�8���'ے@B��?~�����P�Թ�	�'<��a0�O;1�tڰ�IP�
�'d��Yt�@%�R����Q�L�6xq
�'�H�p��<�8�)��޷E㚀0	�'���� �נ`7N�rW✔�j`	�'��|1���)ST�y��K����'`B�AAm����F�XF����'��lZN���,���N�~��	�'�HI�1�	�a��<�Iʼi;����'e.�#3B[�7�<B�E�k�����'��(E)(4���#��[c֎�;�'�Ν
�뇳GX����? f�Q#�'ְ=��K�*��V�%ނ���'r��*��w�x�e�3�6m#
�' R���l
2t1`&�y1��:�'�I1'g��O���Ce-<b��9�'�Rl��*��>��ܲBEb����'�x�EM�@���$�� �$�h�'��D��M)i\�Bg�����'{P��S���:��B�
���'�
�����0*��1�$J���v���'�1���*<��4i40�
�'��qj'B�}ޠ���F�yB�	�'�>50�C�!dm�m�S͕&Mo^�*	�'�BD��	^x�l ����o�-��':,Y�0�<D."���@��s�����'��h;��[yP��c�0L�	�'@�Ș֯���6H6R	�'������P�"�"в]ߨ�0�'��}J�HN;̎ PMJIW��
�'2�����_����7ǗY^h�
�'�&���
���H�;��Gn�.M*�'m�5�%D�q��X��'a�m��'ܡ�g+/	��\C#�"h�v�9�'��$X��Xj ���HX%k~��*�'����.��^�D����fh�a"�'(yZ�JP�#�8�"q.�S0X��'>��ҋ�6���)�C�7UH�
�'�HBd���Xֳ0�DdÜ�y���,�|e�R,]*��B%mڷ�yr��5|�`K��I$^ ��2���.�yB��X�&�CULӓM-*��#G&�y�IӖBG>�i&L��C�J	�d+�y$�9~j�V�(=��ȳE/˂M!�C�I��d��㋊]��@ZY��!�'SyY��_&�D4Pr���5��'Jܑ�Dճ?�Vā��8x��{�'kr���*��'}l4J�$�
LZ�x�'���R)�-&�:%
��k88��'�>H�e*�^j��įO2Kd��
�'9�%���ډ]��h��Ȯ)���
�'<DBcO�4)_� @�� >;�pq��� ���!oD�Y��)QM��k�=OD����2�p>����2f���p/M�*��}Y�X؞�q��<.�����'��L��O�.~��d@O8�� �'I�<�օ!6�;��S?:/T1:�y��ӿ;,\!�D�k_�F��!)�y!"C��$غBG �yZ(��a�]@7FT�*L�,ُ�!aa`D�?Y!�4����I�����H�i{t��S��C�It]P`h��*S�<$sSN�:EyX��E�o�
35Ⴌ��ɭ��l3���#��y��@Z�?�R��S+F~}��〶wT���➞c�H�4	ɺ)��q+�HƹB1�0�'����L��!D�&؝��aPI<�C�B�84��� ���=s@`$�ӈ
D��Vn?�a�$N(`:B�.���c@Y1'�α��mgV*�b !Y�=�	C���;.�0�@�#�SW�	�n���%c�-������H�
��$��{�B�r1҉q,�E�uf
�/�(�'�D�y6�x"ٶ^o�D�o*,O�ajt�R�8�@��sL�*Q7���'��h*�FN��^�0�㖺}��0V�E��lY�T,{Ԛ ����b�!��|���p��D P#n.��I;?�T��Rl-2�\���T�� t�ͩ焃4V�ޜ��$�
�y"dϣxeP����W��,�5�X�HI�����
dR��R�j
Z����L~r�J*�DIor�[�	쮙�d*�5�a��Z���TA���+%�	�di�/.�*%��~�
�M�#H�����/r��򄛉n��|�F�.+�Ͳ^�\]�����7lx�drCɖ�ru�#��'}�@`����I���N��9��	�J�B≓� 9�-k(�:��J8l���fbA�0��A]��Ã�
a�Q��6�S�Y[��Z-O�*�n��EJ��C�2�bX�5��
�0�g�s���`�+�7^��H��a��Pv�aw�*��C���Q���;��k�R""��>y���	�=r��z��)2�x�{ؑ�(E	]V�B@R�Q�'a��\�T��牐,W`��j7�n��0·�Y��">�e��OwH;#��{��h�˚�"_�0���D"���!���L���g�]O!�D@�i��뇪޹+q����X����޹|���g�MӘ	m�������=��OtBe��Ku8���,�m�P�+�'���y�ڧ~���Ũ-(	�	��PѸQ�G��=)@��"gS���>(BO�Y!���Ft�Z�EF'HIP�F�'��x O��h|q�惐$���""���C�<�rDpf#���b� /|R�8�2�P�<+�	�+����&!��P�D�-��	�� �!Tq�mä�$����'��4@�Q0E�b��N�R-&�2c W�� s�dP�z��!��d�D�6���dI!p��1�朶M��D��
K�J'܁{k�E���էA�&���	a�'T�:蒧lM�BlZ��Ư..~i�G�B�|�.��d�)��8���:C;8ı�1.y���@��'fP��c�OI�8�W>�A1�Qu�'eV�8d	)��(���ͨN��r��y�Ԁi�йhZ��pFP�li�1�K�&����&�H-m H�nV&��{�{�ӌ\�˧!�8L��h�jZ��*�+�lCRE}r�[��9���+Q�r!����#�>DQ�oJ�0�bAЃ��q�(��2N�%�?�`Fim�?���"1Rn\	�@ɠp��HB�JM}b�� N�k�'�)RdP����+4�"|
c����I��
�$jw�XطZD�<Q�&\KVX<�%啧\���j�l�7h�a�4%�"^QZy��˨tˎ $?}�<i���?.5��e�O>�J��p<a���$Y{H�*���R�d[6hܡE�����/snB
�/ְd����dȵ8zz}˄�:%�E/ay�)W"u$R2kJ� Z�II^��/��$|"Ү�:U�0B� JR�;'ײ{�2��Ճ"<q�CC���~�UCV�pcp��%"ʿ4�*�:D�|�<�bC�S�b|{��;6X�+S �G�<�=rYZ���Q�n�bpJ	K�<��ͦ#n$$@S�8B79s���N�<ɀO�3<J92G��2�4M0ČO�<a��<�~d;T�5\�]C5)�I�<a�kx�f=(a�ܲ%�vTSbE�F�<�D"�]�Ta���סq&pKA	JB�<qR'��BH0�)��6[�Z���d�B�<�v�Q,P�]�q�_�"@�kA'�~�<!�`�;?����G',0Ti�a�]A�<� �2d�LQva��HB2PA��"O�y��Es�@��D�&YJ�bR"Op�3$�C��U��%��Z�.Uh�"O@��$��C�Fщ�.M�$���""O`ِ��B�-$0�b-��P0L�u"Oxг��V4Sn��1��Ǩ-<fx��"O�� E������p�閍+ uQ2"O�� cg�j��Q(�(�>7�d��"O8���"�-̚�ز��[�*u{a"ON�֢�T��[�A֌����d"O�P'�]�����*��H)"O�e����9?�kV�� Q�j���"O���g�9KQL��7`�>H�Αi�"O@�a��F'H�tT���>˖ *�"O �b2 �6���M��i
\��u"O�DsD�S�	9���w�Kk����"O���#�F�c^
}RE�ӷc���"O����.���s�Ƣ}���5"O�-[S�b���z�lˠn�&��C"O�E�W�r?����KK$0���2"Ot��kU�@ư�he���`^ڲ"O0Ls&O��H�n�+x$���"ObT�jr���Y���& �I�"O@�w V����V,Ҥ7��kQ"O��9p�ø:�\y[ua�J(P���"O&`Z��_P�Qp�N���=)@"Oe13��*M�R��'/'x�0U"O�e8��m�<CR��9ep-k0"OB���摦m+@}P͗�lz�c�"O���#�\fؕ���I�q��(��"OD��!S�H�r�c ��Z��)�"O� 镅l6���;�pI�"Ob�uF �����ÇC�N\��"Oj�y��+*?�ѡ�!̬Ժ	 @"O��9ˊ0&Mk��_�U�2��w"O(ݫ��E('��GOP�`�ڼBQ"O�5j��D�=u�� �Oޕou��5"O�ܛG�ޢ)/�|��c�-8S�P�"O��i�i\�`\�P�3�Q8	B��P�"Oe�Ռ Fs iѫ�;���a"O@�Q�GׅpDf�Jb� &S_
A��"O0� ��F�.���$k3��"O����j�*D������o?���"O��`F@S�j�# k�m�ʰ"O�͢��[!**@ϊ5�#�"O"RцY�L�UZ���G:��2"O�ɔdZ  P�7&%L��1"O� x��ޯg�x1t�J=�Y�a"OĔ���G1jѬ� E����A"O�����g�TTQPᙩVT�ah�"O�]���b��,eQ�S����yB!�	�^�0�C��m��qDL�(�y�b�,p��v_/XfqR�
�y҈�&Yq���#�I���U E$Q�yn�,+2�%bļac�Tbn��yȑ0�8��GeL��Q�A�A?�yb# �:o�i�a!]O�Z�
���y�)�1+�i�	O��-z�j���y�dO$|Ҡ��9?�x�����y򬐊���0�ͼ$�5A)�:�y�GҳRv.�k�� UF��1!�M�<�F�9X ���֤"Z���Nd�<��J�xfn	�
O&S��e���Hk�<A��1����#vL�xC���<� h(��Kޗ����'N�M(,B"O��r-�MC��C�������"Ot}��F2S��ŉ$u0���"O`���eٗR2�s�OV�`�<��"O��2��0H�A�C��$Z6\K�"Ob�s�� h��sa�ǹW�ָ�"O��6�T�,bLC4@&����"O�|C�ơ?�B<ye`U�E��y��"O�PA1���0��PB���Bd��"Oz@x��x�
YSӊ&K���+C"O �)��ǅ|�>j���G��|p�"O�Xӂ2y��)q#A�V��ڇ�d�(@�bѻ�����#U�H��'��4�'jD�dr���E�Y-��9{	�'�ٙ��O�`´H��0{���c
�'(����(	Z�8�)���"~ ����'5�+d$����4�
}U���']�#�i
aJ����a��}�'�,܊!,�C��$@p+��`����'J"L-){
L1w�Ѻx3�Lsv#�y�<�v`_�U{Τ �'W�;�l�:���z�<	�#�gp�:���-�RV�Gb�<���3C�>�1��O<u3�q�Z�<���6خHQ
¡kL2pQsa�X�<� �6>4��nC�Jo
ݠ@��U�<a�D1s���#�{U�x`ӊ�k�<�1��1�6I��A1E�^��]�<��EB.m��k#��):4S6U�<�PbQg�&���(x��0���E�<9��N�Vx�,�lPv�.�:��}�<a���![Cqqp*��/h��"��E�<!RF 8���P`W�"�.�AG{�<�@�-Y&�kw�XUX<�F
O�<���*eH��(q�	����t�<!E	1I����5C�<O�v���DGm�<1t��)08͓� C�]�vQ�B[D�<�R�OfH�u����	b�L2С�K�<��J&jB`"և��t�q;��1T����(\�[��`�A錤&�A[c D��ʄ�˺x ��1�� �L<,X��=D��Х�%�ށ0��-��D���'D�$��剕)��Xj7��:~��
�1D�гB��0���Ţ�2��s�./D�U�&q'�٩��ȥb��)�8D�a�Ą�Pv���C��,D0�,��
K07�3S�RAG�4� '&(1��E����ݤb!�D�6q���͐
w�~,i�i��W�hQo�9`^�r��OT����Y��XG�]Pl�#'�R3[1T�˗�8D�D���G�8��d�wm��Q��%�W$\|5�FY�=W���/LO�C�nS�H��q�I�}�Hذ&�'��}��IR��1��wV���&������	�3�t�ȓ9dBb�� �oL� ��-@���=A�� ��#� L��#|rq���|�ɈN/��8�gIY�<Q��\*q�d���'8L:tY��/J7�̤�F�X���?Ѻ�|�'�J��D��sZ�2�`��@���!DpЉ�}��h�DzA�&�1�Drԁ�8F���j�L
z��\
��ɕU�P)2u�=}� j��5\OL�qK_?w��bq!�2f`.�����=���i��,�bi 
�'\�hE�J�Kɼ�	'�]TX�=Z�{�&
lt����P֊\D��"�t�$�&b�9}�\��%Lݪ�yB@@1a8<�� @�(i���A*X�h��˃�O�4���'A�EE�,O��"h�?q���H�+!">�s�"O6�ZŅJk��8�Ө:5�]0�i+�Q�g�1'��@��'U�ي$��p^�
�����#�x��P�V�p���FJ�*Qt�{�L!�i�QO>D�� t��Q��V�Z���@N�A1u�	4Wt��U��O*�3`O; �`�:`���]��HC��Cv�����x'$=�B�ֲ^҆�����Q*��sJ�3h�n">Y�C�0p���＼���Y!5A��Zހ[5K�:�y"���fՠ�n�_K2����1��'�2����<�Q�Κ9�~b>�(c?u��2��
P
�l<�O*D!̒�yR��*�}����H0�P�e@5$�>�S� ���J�AU����')��[�	:
�-����~u����OuY�e���M�&Z�-h6e?�gy���xU��c� �b�̠�wN��I+ZЊSM*�O��H%/�5,~P�#ң/\��c/�r\�������]~��O�q3����k�;��x:�H�����^o�����cr��֏�^ L�RrI�6lڂ!����~¨��y�NP�x(� �M;��$� C>��үG8=��`�'P�s�џ�6LZ�^a�U�c��� �� H ���.A�={d/�1Pt9���:k��lڒ'��'h�h�G�[p�'���	��'���W*��Bu0+O`�B�O� �h��ɜ"�BlcZ��O!����@ 9_vD�'Oڃƕ`Ĥ�){���I�0�0��`��}���`��h�h%w�*L��ۓW�(�)��>0<��G���oU%J������ēX�I���!�3��7@��C!^�,��\��J¦�����'��<Jq
d���Z/"��I&����1��(�4�wKW7T�?�2�׌{� �rH���Q3��T.�ΨZ��9p��8aP���laO>aT�������9����O~1�'��0 c�ƥ:��D)�h֩]�:�A�O&��VBɜ3{t��N�>F��ԺP?O�g?Y�$t�d��G'/��Q�a�?�#�����D�1Z|V��-�[�Ҵ:��L#IND�j��Ynt��%U�3��5��LT!F����^�?�$���1ϩ>�G�:*����&Y5<f0��);d����a����|�.��E{��@́:ސ$�'@�<q�2�[�#D�a{"�O&=Kv��W�]9i�D��.~��L3P,<O���PM0V��>�px>Z����藼B��Es��;�A��㧭	�h~�)�GIg�p�I�(dI�k�6ָ@�,PTH�e�R�49�$_0 �C�L��~��;+ܠ��j$�IT�KnP�r�G��բ�ꋄqd�ɷ;��j�%�$�!'�ׅJ�(#=A4��,l��	)%n�H�<�sd$3���4o��@8�)�3 s� �Ӓ~�<�h="�+V��5b�0TN�2Y���(R�"5Q��Y'�K e-� 5T��6��7s�>�"�ϣ|(�1QAMӸ}2��;<O�0SE	�9��:��\5�l��W�݁o�|�?9���9�qK�j�2ػ�Ћc�1+w�8�����#h�@5sd��"}�Y�c��>@���#����Ƃ<�|6-�,[�*�K�L��$�j��Ğ32Ͱq�Z�
��K$���&���6'�;W*�I�DЩd��h��Ծ��t!B� k����ݢ��H+S���0-�I� l���NJ�z��k�D�u��"=�e9�ʃ䟱4bٓ�

 M����+�~JQ$�n �O��I<[���jYV��&eW�0o��K���
&��E��mՊ(�v�����|�c��Jj֬S���*���ચ�AJx�����|��4cI+*�*�O:�IK��ߓY��tL�=r��Klf}�+�Ƶa�
���2�F�#����W�D" ������]P�x��K�C9$������Q^N�KW3���6�N�IS��d�A���ʔG����O��IҞm��`]/*��M{0A�� z�(�"�"�)[ч�K���E�<�H|��*#F�x��.qXT[�K̽X)B0@�i���>yT戦U\��Jb���`�"�"O�'�iY�iE�dV�y��^<bor���N"��ɣ(S��ٲ��f��U�K�#���dÓH�TiᠫN�K�����F����.zjź` ^��	�_���'h��2�$�V}�"ľ.�^���㙛VLV�!��� ��O:y�B����'��t{@H]"��y֯�([�zTb�$�ɦ��Gl-}R�ų�D~��	�[�� �nOԞ��'���ċm��Px��/}b��7��y��~�u(�_�D��sgB9{þ��c��pR��A4�O�- Q��H�hl`s�A1>�T5*A�>���@�B<^�kV��<i@�Ox�P�T�L�`�Y�_��lЩjL��+�L�f��M��|D�91�X����#<�L�Д�ೆ7Ox��L<��z��a@�lcP�.e>���g��}H8<�ȓ<V|@�C��. ��2T��8E �g�D��@���?�':�@�&�F6_�<8�.%H5i�'Q���n̥h������N�c8*�ہ'�|l�]����9��@D�QE:%��`I����DT��:$�H<��'D!Rt� �v�آR�hE���Y�<fŁ:h;0l�-������	z̓Co�豍��Ă�W�|�Q����j�*D��y�"�0�n$A�-?�P1��I�y�ě?���Ơ$y�(5q� �y
� �X��g�ε�b'�
?�����"O&$�U2T��U�`fS�Ĕ�+�"O�-� EϘ$��9��<B��̪�"O���t�"{n�y�RM�&�py1"O��C�BF�]TR�:E�K���"O��@��'E���@r�S�4��eX7"OZ7��͙��I���w"O��k�7`��`�w��'Ϻ��"O<�L�<��A�F&qm� �"O"�ϓ� E���ĦOi��Q�"Oz����'j�S�4M�فu"Oj@{����N]#f�0(� � "O=�����@�&M&�ɷ/n.!�
*��)3�fFT�Z�M^�]'!�䛪su�@E�F�q0�cW�$,!�� .��0TmM#z�ޠ��_�}�!����� �5�Ġ��K1�!򄒷 uH�9TjK*��l��D�T�!�$�k!2ujt�R>G�"h��C	�y�!��D��A2���s�,y&�Py�!���yX�ka�t�V������:�!�D�<�A��#۾��ѥ0�!�d
�mR�銊~�Yq���$�!��ҿ B�ծ[���%c�?+!�T5 �����ٱv؄�)��({*!�d0 4���ڃϐ�BՊݪ!�DI������m�.��\���_"!�\d�T�9$cB�7D�5�t�'�!�ċ�a�^H�S'���7��)d�!�$Ŧm~m�P�;��o�/h�!��W�$��q
��|	�H27�&^e!�dQ��	�!��{�ج�㉮l>!�$��k6U2��P>�L�Q�� i�!�SH���N_+sǞ�JZ�����'����}w�g���>r���'`L(�UI,�yq���@9Fl��'�l�9u����U�1lL1�p�
�'Ⱦx�aM[���Q�d*#h�h�'\�z���(�ǀ��%�\��"OB�B����<Fj�J�G�r���x"O���B���_l-�1��X�J "O�s�G��0Na�D��B�����"Oɒ�Z>s���+K/q��Y�2"O> 3�0��z�i��q� ��4"O��Q>���wB�3h��1b�"O
��5�3�e�eAQ�,�"�i�"Oр�ҜJOԳ$���($�3"O���f^8;��q�6��(f��z�"O��.��1RV�5S�A��"O�X�s����\2L	f#X���"O20ؖ�˗�)����"#02V"O0��������%i��8u�Έ�yr��1685HPM��2z��/U��y��E���ɨe��
f.�6B��yb���dyޜ	`��{]����y��z�NDBkAd�  ���M�y¬�VL��T�\!�P �y��N$Q�4(�&��Y���u�%�y��PM`	PeA k�)����y�`CWm�ٺ4��+�h��M�8�y��Ԥ$z6؃$�!2��P�;�y-L�1C�=��̂	���+���y�d ����%�L���6gX�y���#^|�e��.1:�T����y
�  
�W�or��Ĉ$>��"O�$�2_/�d%�z���g"O��+�`�0�C�Y��zc"OU�E*�L[4�(�Yl�F�xb"Oj���%��Y(�'K<j�~��"O.��`ʹ,�`K�EW� ��4�"O�,`Ǌ���7�O6��"OԩY@�B:YK<���ϰz��}A6"OrŹ���׊Brn�x����3"O��yp���?*4�1���Q���"O��	a�Z-���a��'�P<�"O�QD [��HAB {�� �P"O�A�kE9hQ���Wj�n\4(ȑ"Oj��
R�:j
����k���"O����,�F��8r'����ģ�"O~ [��s8%���Ԍj@p�(�"O>�8D�g��p;�A7[*.��w"O�8�s���g|�Gc�,>.��"O��0���	��D�S���%Ѥ"O&����E�4�J�``��*F%�ģ�"O��{"�-r��u��X4~B�ؠ"O4]�2��L�q�Ñ5�n3�"O& %9E���Bc�0�J�+�"Of����  ���ѩ{*�1��"OL�p ��U��؆�̩g7�X�"O��9& ��iHd�`�E� �����"OЉ��0l�n��ĎR5��9��"O���PV��e�#g�N,cU"OȁI�i�2�x���jvnp��"O���� ��1g�Q޸j&����)D����MX�3w��ߌ$����`;D�Y-�e�$|���"d��aV�%D�@�FE��]Z� zAf �;���z�"D��y�n�:a�e(h��e# D������a�Ш�"��?���	>D���Q�C":�@��'�tQ�E&D��)fh΄]��u
�Ď7x�����b#D��s�m�c���tD��d��%���?D�L�W�.<랑3�#4ٜ�i#c<D��A����Kva
mк9}��3�h6D�l���2K�$����oM�A�6D�0��
�qIf��H��~o�M��i3D��æ	��oڸ��v��c����1D�PS�IR�ը��`l�0�t=�Ҋ1D��$M2|�B��d�=XV�����/D�P	�c� 2G�¢Iɠ���5+D���C�(
h��#jG�9j��T�%D�lZ���J4t����}B1�+$D�$+���Q�<�SC�S�^i|y�>D�tRT�G��-���Y�1D�8U鉋	I@I�%P�e�Y��/D�p@���N!�:R�� (�̰Z2-D�@���< ](4��$��B�ɓ	�
9��&���K�掲H�B�	�vL��1&�B�HD�ArE�E5 B�	<D�D9�'���T�� $�B�	����]�R	T�⢌�:N`NB�ɑP� Xb�1B @�`�\Z2JB䉘yT�����I0d��-� n\0:H�C�I�^K��p��̱S��APMA��C�ɛI#6틷��<��'F�Zy�B��o�|*�BK�m�nX@�E�v��B�	�[ �m2��
�ud
����%ZjB䉽g�.ݙԪՁ�}���;g�LB�)� ��U�pˊ)X� �64!va*6"O uX#�C��E05N��G
�J�"O��2��א�(�*��FO*5"O��x�����ū�0NJ���b"O�=#S)N�f��cpØ.VBQ"OT=jc(λ.�ZL�q(
gCyCS"Oء�#.P%*�>m�SI�	^��p�"Ob,�'�ݔ%�v!�Ce�Db�0z"OB	#�CB�V������I�bx�P""O�(@b��j�2)�HU3Cv��B"O��1"��|Y�a[H�(WF�Q�"OZ��F(Y;����f�5۔�q�"O�\�Ή6B�	��&χa��p"Oz�j�����j���*:�RG"O�4ڳa��a,�*����n 
v"OB`I���T�H�"7+у<����B"O�:��Ȃ6�Z�r)�/G���0"O�GN��yx��kN ?X+�)+Q"O��Ãē�s�	&�+*��KR"O��F4l{t�jo569�"OL�Y��,��gor����ÿ�y�˓�9l�8'M �n�z�Æn˰�y�J)_Į�ƍ�a;y6-Һ�y@  ��Yj�G�D�N�s�����y��)��̛��Ŧ;�đʗH9�y�KY�S�N�I�IBt�0� ��y2">'`$�� ��f��E�gP��y��=R�����Q�ZA�Y� ���y�M��Jՠ�lO�	<�i#SE���yR+��)���� �{f�
3�D �y�c@4 ��pM͋x7*�S��(�y��*aX�I�hz����B� �yr�O�H�p��@�Ŧ�>�
sEA�<�rDl�t� (H:��8��Ef�<��*V_�	P���m��1�Śc�<��P�Rv���b�	^��r.�c�<���k[��ɡEE�w���qB�v�<�`J��z�=�$��@%���J�<a�`O+*p����1|$����NG�<���: ��G�zs���e�E�<�7OK�l��GF6pPx��#�V�<�$i��%�6��B��z�>}��^P�'�����*nz��a�k��Yf�`�Jպ![!��K2�كf��?Oj�ys(N;qX!�$�6k3��J�@On�fļU6!��M�{@d#���6l r�*aē�W�!�DA�{����^�4��1��8N�!�P�zD��:b�;LH1a��}�!��3���ZDnϭkSRa�E 	U�!򄈿�B�bʉ~��`��b�7i!��7��X)v� �V ��!Ϩ<�!�DLh���G��N�9�Fށ_!��\�8�ر�O�0:�j������b�!�38��a[��ռ !|с�9
!�dU����h�X�$Nuj�B^�!��Q���kb���i�P�a �ͨS!�$�@��(��P'о��G�N}.!��9z��c�E;z�8��e�.O!�$	�M^�@�蒩�2	��$�c1!�Ě8<�L��e�A�s��$�3�!�DV�U��՘D�!q�@�A�w�!�d�R����OU�DWtih�A��x�!�dZ�S�����Gv5�a�$<j!�.t��Hh!�ȉTֱЀ�\� K!�� �\3go�5V�4q�� ,a�nX5"O�1`���D�� ;,	��"Ot$ڥ�W_:��"�!k.84�s"O��cw�2P�6y�G�N�zL�P"O:�ش��6y�8�� ��p����U"O(鳥cĂ8�f��d/Ν��@�"O.Xe�_�K ec'͢Ag2{F"O ����8��Ѡ%ԉb�^, t"O�h�@dU����ADǑ7�Q
�"O���ntlE/dXM���G.&!�d).]�i�H��/��5rr'��z��VH�
VNאy_��U���y�i��b`\�#�\��T�;b/ݗr�*U�ȓZ�q�C	���Cf�s�p����dA��>����2<p�ȓ��"�� ]#p#F
����ȓ#��I����/yj��I.U�NɄ�E�	Ӆ`��fd�eC� -��8rEX� 
rږD��l
�?2���Z��Ԋ��zA��8��9(X<)��}���Z��]�{�4h0CP,L�NՇ�Li���5��/vXD�C!_��RԇȓV%�brmҩ%n�ͱ�H,xOJ��l0h�%ؙ3W�!P��$���ȓe�������r��%��B�=��(�N��U�\x|�k��$V��5��@��!��І���' ӻU�ʑ��A&q	�&̘ ;��3`(�r���ȓCI�)�s&Ŏ��LR��'uY��ȓ+~�k���?m�*I� @M)x�d���i�9rb��J1н�-�,c���j�c#�&\Mʼ�o�~4I��]1@xa5�@q��!g!8b�x��/劈�B�J�d�F 	8[[��ȓ|�D� ��'0]L�:u��6tC�Y��w�X�Af��.���P.�X}ʝ��q�x �lG��<����1t4������YI�
;`^$P&bU�Lv��ȓ]g.���5�n��0Z��0��ȓS+��ЕKνp��%Q�L�OC���6<�)2u\>fc��� �Ŋ����X��u��Qt%�ā1FJ���2�9s�
�*|��0KϬO�}�ȓ"�Ș��d�c���KDEc�� �'����`ʴ=�8AԌC� X��'wP%���B!B!@�cSl�)7͚��'U��A�{9�RB�,��8��'�2��LPRg�hY�g���Ɉ�'��i�m�6�n� r'� ��u��'5�z�Z�����S�
�NШ�'�D%C�.��k-�`h2��NH��
�'̪��n �ij��^����H
�'Z�)H�&�: ��\{�� ��-��'ax�a�4: �fn�*b�<P��'����C�9&Gt��@A��.6RՋ�'�N���h�N<�@���'OZș
�'8��і'ѫOb�����30ChI
�'z�$l�9ED�W],�d	:�'���Zb��:I��m���	W``���'6��6I�P2#��]D���'Հx��+"�DҒ�S
gd|��'|H-c%H%u�x!@Rb�&Z� ܚ�'w���v���Ҡ��(��a�'�<3@`�Y� ��V#n�
��� �6��^�`�jT����"O�yc���K�X���&�9���z�"O,H��#�	�e�<Gu���E"OȰ�G�	\�I�F��l
e�W"O���� �Hj�Ѳ%	�|��"O$Dr*jT�3�J�"�~�P"O����Ć �%�t
˾}Fq��"O���=l�:x�J�k��$�"O4�:��OӾ��Gd�ex�
�"O��s��S"�RyG$�D&�`�"O��*V֝M'���7d&K�"O��9P��h&�`B3��'%�h���"O��x��	l�����~��<�"O�	;���x.�Z ��6��	��"O��$޿-� �2��e��@A"OXͻ&
?.�Z��ªr��l��"Od�1�Y%�:�R��N7�T9 B"O&�w�����*�^�<hG"O�%S�Kҋ���q��X1�\H9�"OI�A�E!+�񡴋͋q�Z	3�"O����ӽ\�ѻqjI#3�܌�"O��ٰ.W�xr�x���\�4}1�"O���iB�9��U�L�D��9j�"O5�v"ѽ5���� ,�2D�()�"O���/N�]��$)'�Ġ���Q"O"d�¡ߜZHx8A�.�F�R9AW"O��"�O� ���s�ګ!�Ԕ�"OTQ0�$�Y��JF�u�8Is"O�����Ϫ+^hQ�C�I���"O@I�Q�Z>N��V%[�e��EbQ"O1��ǌ�Ak���Ɔ?>���"O� �a��%hn,�B�I"���"OƄ�`�$y8�ԙ���S9���A"O��)� P,D�x ��F;�Ƞ`�"O�z�(V�b��#�(S|�P0�"O�*@�P(n� ��%Z6!���2�"O��Y�G���BEʇw\�|�p"O�cङ�$p���	�m
�K�"O��`Ë[z�Y�����.���"O�iB`�	V�@�pBa�3�̀�3"O&�P�Ǉ1���
T7e
6%�2"O�K3
D���y��ɳ�FD"O�9�cW�h�բ��U C���E"Ob ���9=±�c�ل|"O`��G�I>`i���R���{#"O���@�;_�V
�l�1�T}H�"Ox0�0�2}����&!Ŵ���F"On��2�B##+|8(�H�E���2"OTH�gE
D��m�7�ԻR���R"O�LJ����J1lZ�ud�"OPEbRK�"tU��]�EEr Z�"O�(ǈ��l����j]<0���"O����)H�ęF
�>�Ԁ!c"Or�KC���"5�Qj���ҍa�"O80P�M381F�3�8�Π�s"O�̱S�A���JY$h�b��"O:��aHɽ:�xLb1�W6o�)�V"OliA�;��A���!n�Ό�A"O�Q�W%�GP�,�7Ş]���c"O�Dy3m��2�xM9���詁�"O��KǡC9{�|!3bE1h2��"O�as��U�()zƀ�H��$JU"O�yj�$C�`׮��&-��"O:�q���&��"ޠ#���( �'�1O� ����6�T�˙'k���Qg"OR8��jk����c���Gt �0�"OL�2��L�lQ����5xe����"O���v��4(�@qx�η0Z��z�"O�9��&K���#�=#=�lЂ"O�pq�����+ k,���q!�$��`bX|#Ć�<_�)!CŞ�_m�}2���Zccߚ1����c�w�R�E(/D�L���A�����,O�6�pU�g�+D���w���h"H��F���o+2YY��6D�8"�-�:F�źb&��@���c�5LO��d	�'�'%��W�V�9��c�!�]'E4nԙ�$�-Lٰ��дj���M��(��8S'"_�Q耕�6���M@�9D��:�O@(�Vd�w�\����v�5D������+�l���Kݽyj�\�7$5�O��I��|\QAAD�Q�I��L���`C�I�^�Z�#��[�Xj�FC�	5 z�˥�̪=`�az�S09NB��Q�ƼPG=�v�(�
E=4B�	0k�df�Տ.�AS����zNC�	�a���A-	 L�M(�B�	 J! �kT�=Onu�ը�@�B䉜i��YYg�кp�La���$~(C�		!�����@�8wB0�r ��`C��Eˮ���N�0�
��5@
;xR�C�I4��jUd֑=���;���P��C�Ɉ����f�UhA�� ƅW����'�	�>�vD
$%�1���Q�.�G,~B�I"*7����F��P��2��
�C��7P!@I�a�8)6Ԥ��.�4A�C�I*�<�p΋�M
b��M�%ɢC�I�!'����ܮ|:��Xp��6�8B��7D�6���۩Ma��*���JYJC��(3�H�HcO�o������YB��gsh��'�थ���+y�B�	#0o�� �A7WI�E�"���D��C�I(K�D�B��Q%g�ɀ�J�	g0��h��p(��եL�L��؀B��'0D����k��T�l#�%W�|��P�C;D��a�t>&T��e3�a��.5D�X"uc��?Q~��S�qw&��^p�<��T>u�f��X��m�K�	V*l0��1D��ӆ�R�
��B�!,B��1��hO?��&����F ��A.�!��Bi!�Əo����A�C;g�$4H�Ywh!��_P۶\�W��E��21?HS�|"�x(�EO.��%�
v+T�3�L�	ϸ'�<#=%?�H�ڶ#�,�spd�0 Ԏ̣ե.D������/g"�D˥n�e�v<�#�1D�hh�*@�M:�,����P�(#�g0D�8ڴ�%���ٶ�K:z�F�أ�1D��BA��P(����F�T)/D�X�F'��\{B��p���Bܙf3D�(�i��$�{g#M�l�
3D�,q�fC�>���Վth�]�6b-D�4:p�^�iY��7W{����)D�\ԭK�X�u+�i�\pt`0��3D�,�-
�K(ā����h=N�W�-D��m�<��T8T@q��VD)D�P8b*
~��B�-y�JJ�*"D���uI�ު�{g�I�3� �`�&"D��0��U�/�Ex"�ǈ{���Ж�>D��ʷ�1mY*؂wFح=n%��� D�� h-��`�=d����0#�PS6"O6����I2�M�+��A��"O��z�FN�@ �"�m�<tﮑ�F"O�`�n�4��H���ֹ� �RG"O*��c"^8�Qq,I�� �$"O\	JP���%!��j+W'��L�P"O2$��;Z���Ћ֓ ��P�"O�1&�M&*����@� 1!"O�U#"���j�	G.k�ș!�"O�d{%�R�w��8�sct�"O������4b��v�ŤnRn�""O�ɪ�.�_����m� GX] "O��k5+O�i_�P�e��4,��"O��q�eE%�����e�,ol�YC�"O
�g�LZ�𺆆<o�d��"Oб�Q��' u94��)O�9�A"O�p)CDU�q`������0;�"O�1��>Z� �����a6&Y
�"O~m�3C^%���dUtyF��V"O�[B"N��L��$��r�93�"O �Ӕc��+���c�
��5�"O�2@eN�#���`Ç7��L��"O��[�C��Es���Vl�g� i��"O�Kb��$y>1PT�+_����"O�,1�HV"*�ʸ���҈@��A�E"O^0�.��j�ˇk�lg�I��"O���DN�\(�I�JR�+Pe��"O��-(D��X�Q&{�-8�"O�]9u�B�0�����]<:����q"O�X��
	'�h�wH̴?L���"O*���hN�N.��Ð�`/��qT"O\y�8({��;�$X�"O"u�t�M�9#�űx�  p"O��9&+¼}�ԑX��Nވir"O�eiVlN�)��<��d������"Ob�p���h��r����M�g"O,�a��<B�<`�������B"O8Q Ԥ�(���bC6X�B)�7"O|�6l�--��p�D�ܶ)�}f"O
��t�تSI�R#�� ��!���>������C��	�.��%�!�$��/��賃m���v0�%K_�L�!�d�k���Cf'�^�h��S(H��!��'ot��@ ޘg�
��5'�a{!��	9*j �JP)�-_�Ε�@f%_!���<|�Ha�fȡ?¾D3$���MM!���!t|A��(�0�T,"ę+$,!�$B!�4�I��ѺU��@C���N!��8$�z�zq��,O渨���3!�$�)Q�x��&��k/J��p��=xj!�$K�G�I23C�����IV� �KV!�䖻z�ָ��L:N�x�k�%r�!�D�M��ⴍQg���-�Q�!��V�ƥ�n[=ae�u"��@�C�!�$��$�-��F��bF&���D�x�!��,B�^-a�: H�9p�+|H!�d�[�zA�^TcRQ���C4!��>vm�!�ա[Gx���/!���3uM\)���#м͸���;^!�$6.���5D2G��С��_!򄌍5��1L��^���@�+L!򄃺V����2
�1RH\���Q
�!��A���j�圶f�*�붭f�!�d�Y��h�2���n�Ҁ[w��# �!�� ��`���QӼ5���_B���*O�Q#�ėh�N�v),�3�'l
l���x���yU����PyJ�'�F�AUDV=�Ș��V�nʹ��'ނx:�J�'R��u9�-�$}����'�����rz��%�P���a�'�N�h��E8u2� �R/��C�]��'a��*�O�,M��X��B�Cc^���'D¨{�#U�AB��Q�-A�x0�	�'ռ��Т�A�jL�Qi�
JO����'���:GI^,7�np��6H�J�3�'W��XON�n,�������>�&ٹ�'l��C!e
�"v�`肯�.�v6"O�IZ �\&�Ne��C�9d q�r*O ���U�{;�Y�&L� ,Ո�S�'�����̄Hq��0�@�	W���p
�'�M�#�[���qb�8&|��'�l�w,� J,RD�q`(<��'`��A��~ڌ �C���L�b�'�Ȅ`�|֮�A���@��'}8����I/��U����^z��
�'����]>Z���c��U�&Y>��
�'��`#-Q����&�=��'� �X
��m°��)u*� �'�2$�S�O���j����4�'ڤ�a%�1!|h8�iVo��dr	�'ݒ-pl��
�d�Yr�N�c�FY �'趈�0�֑W5�JcZA��'�,<��-�r�1v	�U�:���']��2���a�T�U�`��4��'�h� CJ�U��!�@S���h
�'� �bO�Ѵ�`�K�L  
�'!9�����8(jK��ٓ�X��'�����]���ɢH���Xh�'�t�����Q�j(3�l��}���
�'vi�tBO*��M�bW���PQ�'�����	�x�Re�T�Z7j� �
�'�N�����,�X������p����
�'�fXKaZ�@4DEᓇn�~0��"OH�a�#Ģyhp<���P�B����"O�XsFS+.�� :���jOD��P"O�8Z�7�(���C�f1�"O������n�BP����%(�Q�"O: Fh_8" �{cb��3�,ʡ"O����g�P;���!B-lU�]x�"O4����92��c'�8<�P�Yr"O �
et������P1���S"O���!!P�J�А�#Ȇ H�{4"O&��$>挃s  ��)�"O`8PЋ_17�d�!t�׾�>eF"O��c%��]������_��q��"ODdӅb��9������N$�� "Ox�J��W�ОH�! PZ�a�"O�Q�A+��K���1dY�V"O��Ɓ�9tn����ƾO��m��"OI�v��!���FMzH��"Oj`X�D�	hY��FXNJ��s"O>|�d�P>�h�W%^�B=h�"O��%#�����1%�V�#y2�"O���M˾r2���C-8r�"O��S��*Y����B_�#' ��"O�K߀}V�QFL9,?>��"O�X:+��_pAf�'+6XF"O�D�T��B�SPE��@
��s�"O� �%�RČ�jW�4�!D�p�$�2�"O*0��Y%v���C�P/G�e�T"OZ��%B	P�B ص!Q��G*O�	!E�O^z\��E��C"� ��'�B�t�n!EZ�H����'�*A	��� 0�����#�1����'��q�NB�$��@	ՃY�0�|��'�j�
b�ʳMiX ���.�ը
�'����@�O���"o2!���'���Y	D�7��leD/&Â��'��8�p�\�!ʴQ4�R�
�P���'L�����X0De6��T�~����'^&��sF9Oe�3�% A&��'�V��_� ?p��'�5�X�'��RC��E'�eP�g�*�.��
�'w��k�[�F�LE �^�nzpI
�'Y�ɲR���x���8o�9P	�'L�(�LS�KĒ͊Ua��7
h0	�'IR�Bb�S)��C$��Y�p*	�'J�$a#��^?J`I��z2�	�',�`
Z&G���i�c�m�
��	�'��e���G�NVܙڕ�R�bxdP	�'�t%ѣ����V�`��/]��mJ�'�$��e��VFDx`Uʇ�B���'���w�P��@;V�� KN�ti�'֤��%�MuJL��5ݔ@��k
�'��-Z��Į?��Ju�^�14��	�'�\�ѩ܅%-���o�9%\ u��'�:q���
	" a�#�43Hmq�'2x�d�?-m2C�
9�`)�'���Y⫓��ܠb��2͈H+�'�:+ �1�����GŨ�$qK�'���7�҃.8���_�q�Ȋ�'��1�sP�����&b�+g (���'��9��ׅK䈁���Rd�Ѐ
�'�c"�!Gz�L�UlI�O����	�'�ڡ�k5�NY4k
I憤��'隘RB⏡o��,�D�Ƨ:���'�0�!���
�4I��5:D����'%F�3��"�J�!��4UtY��'�dE��ET�+D�T!�>jk	�'���5�;bF��0�M(3��	�'D� Y����C�Tp"-ז2�8�'��!�CJ�:!z�x��U)�fp�
�'��� Mt�t��֢Ũ �P�'N����)�3 �Jɣ��D��'-^iǧ�Q$�RF(� ���x�'��	G���y�������
��'���!��Z�~QS��v���'�xL��ҽQS����Q�jN���'�N1�a�V�t(qe��f4�x�	�'p����.�""����X������'hDA�6!��0��6�ԧ��p0�'-L�@���W����  ����'^�T*���j��b��d�'J�m(UD�.e����WX.Z�x	�'3�bu ��y�V�~�����'I�܉6��9� ���A9.�N���'��@(�׃M&�T ߗ(�6��' 
���LN����&O
x\�"�'�"��Ϟ�InVȩP� �����'�z	���c8������B��P�'�񠑧�u��C-��?Z�`
�'DԘ��U,
@LB�2fn�
��� R� '�g�>`��
�� ��"Ot�z�ϑ�G�V�Ѱ��S�^�"O��X�X,���	7�� �p�"Op9�)��a`�!ч	("����"O�̓с�\W�`���"jj$)
P"O���El�9��Ţql	4fF�z�"O���E*[?�����F39X�1"O�����2h¶Al:� bD"O�\��٦A�2 r�3�T��"Odc#&�"�(����	�I����"O��H�!�N��8%�!d't���"Ova��΃?w���8|2�"O�f�1j�NPc4J jt�q"O�\�m�7z�p�Qo�]��"O^X)r+L�p�Rq�&��8S��1�1"O��RDC��G�ԡz��̶�ł�"O�lyG/��7�Z�Mݹ"꜀K�"OR��r�J3B\yy��J?�M�@"O��*�k�%���i��<��"O209D��1����j3����"O�+��]��܈R6�ɬ* ��d"O>���Yj��,��$M�-���S"OP�V�ðZHn$�Q���Հ�"O� �f�ڃF�(p��ܝ_�x���"OF�S�~�>A���H����"O24K
�R��,��6�Ax6"O��Be(��pȩ�SMPId�$y�"O��EgD�5�����v?� AT"O��:�k�>f��@D�>pa�"Ot�B�(X*���yI�BR��Y"O9фb�B�~�9��h�xٛ4"OҵC�;F"�7n�{�*A'"O���\*#^�m�C�G/jt��1"Oy��x�Y�v�5Gh�h"O������EG�̀�jÜB`8�ڤ"O�drd� z�.\Y6�q5"O
ЙJn4<iR���>���"O؅��n�^A�Q0X�l�0a"O؂R��$��  �n\��ݠ"O��`@���8At4��l��(
�"O�`X0�8sf<Ys��~K<��6"O��b6�	�bW�p�0�^�"1�)�D"O"�r�B��DNإ�5���8(��"OP0B,Bj#��Y@��D"O�a)�>H���2��~��+"OI�үϊW�8�!$�4Y��)��"Ol�p���5H�D!Se�Zk~�9�"O��4L6&O~�񗊊�=�TG"O8�x�C�:�eℯL�gQb��@"O$��qE�)I��b�C�"OPA8wl(Z.�#�� 2f��\#u"OI�P�ų4%�%��<�8���"O�A�"�ō7o��u�E�0�ę��"O	�d���(Q�6���ݶD�S"O�@�&�@�f����%���?�*�k�"O��ӱ� (dm��,��E��"O¹��Dv���򦕦%�z��A"O\%�vF�(/��Ѐ7#E�u�z��!"O���N�m��1ip"�7)V�k�"Oʀ.��q1SM�>L!��$���U`��d��xv-�(!�-G��y�)Ϧs��u�C9|����cM���y2Z18��,	�b��t�$]�ӊM�yr�]焥��%ߒ{,@*�"�1�y
� �x��:�]Y1.�2�h�S"O�y���\��AZu♚_�2i�"Ob=�A��`��6!�z�|YkV"O(u ��@�<G$�X5��10�rՑ7"O�m������-ʶ/F�^؆�bS"O���t=�Y��nհt�>AZ�"OB� -�rX�b�G��
�E"O�=I ��R�P��gM4��i"O�TuE�!mo�\
�L	�wT|`"O���D�V
/1*�i0�
@�=�"OV౔Ș�AqZ��⅒K�0�""Ov�B��*Fy>L�u���E�\��"O<�U8It�i#�ۻ("�\�T"O�2؎�_��2`�-���"O:�wFA�PEb�H���.��u�%"O`$���
����R�t� ]H�"OT�����5L���H�� �0U"O�<���E�]SJP��h��T�$m� "O�B�8��QI!�i�θR"OTQ��/=�R���U	7�¬W"O6�kP�Ai��RQ�ʢj��u��"O~y�sm�
%�z��������J�"O�l:Q�G�<
ȼ�S�Y��(��"O8Q�Wf[�5��`�p��u����"O���9_�*)ࠫ'S�uy�"Or�!�Aϴkm��K�q���c"O�9�M�V��	B�k�	wn�u�"O��X�f�yv��U*Q*AP�[s"O�0p̄{�Ż葷tiF�5"O"m�Q�ɭ.�N��e��GW��b�"O@����x��̫@B$�u"O�S���Q�&1�%K�&P5��G"O~����&
ހ}q��΍�\H��"O����.Q�c�!�ǒ����W"O6�������c(�?r���A"OR��P�	 x�2zC�ʤ05����"O6�#�I%Z���;% �>  �l��"Ol 2Fn��L1� A�ao`%i�"O0�CA���^�N��o��m=�Q!"O���GF^V�6Hs��
LI�Dc7"O��@�+�RH=	�`�/72�l9�"O8dX���O�|�놡��uL�""O扛�!�]�rT1��7�l�I�"O��b�F�m�JZW �0~H��%"OPQ⣮Ȃz�P����Ԟ@���f"O>��ψxa>��4��4��` a"O��{���#'։���%l�� 2"O�̙��*:��*���&h}�"OHD)�Qe�� ���[�4�<jt"O�V�)mR�ᐥ�Q~4I!"O��CC�N�M
*E1P(U�|�8a��"O���mڇoN2$h�'*f�x��D"OR��1�E9R��'È;�yD"OF	�f��I�|�YS��
�J��G"O����h�:TT�:���t��A3b"O�Z�ߌ6��uX�KӁM��1"O�Xy��:��@7�޽=��a�"O.y���٫c�>��7o�%�����"O����g�0!idl��֣4��|�"O,��Eԭ����$ݧH�6uh"OƄ8��Ոa98�)�MͻgT��T"O�eP�n�	#�xC3��4O�-�"O�JR�U1K\�5aت�Ҕ"O q�&�[�
��2-ҳ\��\(�"O� j-8��Ԙf��$QE�	D�ޔ@p"O(1 ���)X5�G�\����"O�I Wj	8L@d�bΡmOpK"O�e���ٜi�|a��D��r��Q"OT�)��"�"���M�4���8�"O����ҭg��� l�^e!��"OT����>C�݂p \pcl5z "OH��2	� ��9��"jƨ*�"O � G��O����#C�z9�"O��0$� {QD�)bH�-�&�Q!"O6t��M]�E��3�`1�2"O���M�*�݈�ܩw� i�F8D�8��!=1�$M
 ̕�-�+&�5D�|�Ɛ�K�f���	XXĨ�g/D��9AKĮ3�z3(��-�ā�g+D��p���p>5c�C��=�!�Dȧ:<L�W+�$z��(V�
/!��H�9	��֖!z�!Æ�.)!�D�����&JEC�|��Κ-]!��P�Urc�Z�iDt�Sr'�7�!�$�BTT�Z���o=��Q���s�!�	
��4#���\�����-�!���c1�X7ď�XڬZ����)!� )�,;��F,HUkTAV�
�!�$)vVx8��f�_L:��d/L�Kg!�d�%n�ʡ9''Z���+�)g!�dB8�p�E�{�����/Z3!���eaD�[�J�@a$�(	̽-%!��#�p��D#�"%0䋴�֕F!!�$��P�ꑘ��8#�؈���9U�!�$N�o���S�HV����A�;!��
&���:��I�5�ڹK�嘈'!��ҹ0�� ��	�2XSCKL�!�d��Z�Ty�j�d�X�0 ���V�!�$�x�|�yA-��D���E�_{!�E� H4{g#��n�f�+Q�!�D��n�H���L�;}k�m�E����!�d�?UN�Pg��\M(����Y#!��ڗ"�����.�����s!��&ud����Ǝ�E����v�O�5�!���s*�`���R1Q8��b.�.�!�d�	U�E��JW���s-۔K�!�A6V4T}�dܦiBNԒ��Ysi!�D��/>8K� ٬r��y#A���fM!�d�*at2P� @�7?i|�ئHؽc�!�D��cC:����
Q8�d`D���!�̦]���S�B#2��P� Q�!�$��d-���5��<�5E�nX!�d��H[���c2�9*�N.W�!��N��@�����r4r�#߸�!��%2�.���I6z��l�vCb�!�r�,m�q�_=>��T��U�V�!�D�+{FPe!	Q+�t=�g�εu!�D�1O����J>���:�*�Lm!�$�$��H�6lZ' �>�a�H�r`!�D6ْ����>8���֘I!��N�fW��T���>�2<�VL��o5!�䚐l�^��nX<e�,���Jψ5!�D��v�R�3�b\�2a�@׋Fw!��;.ιJ�)Ǽ4�6H�Cf�c�!�ĝGk�����co��9��R�a�!�IY0�%�`KwӜ���� %DC䉉c'���M�,�x!�3G�<O��B�	)} �\{DG���L�z�m
�^TB�)� �%�M��*<�)�9DN�: "Oڜ`��]�{��ؓ�� 9<.��"O�cK˻ry�<�6�bE�);u"O�(F�5}��rQ�K�H&2��"O�)S	5�*=Z�d�F1��4"OTH��D�:8bL8����YD��0�"Or �V��U`ؙ	R/�xU���"O���$�J��d���ŮBXU2�"O�q��L�&Y=��ӄ@�*8ld�"O��pׄ������ԋM+��Y""O,���,�&��%:�.�5W�<5"O��(�f�/\L�W�ńW$�"OZ8)�ՠ|�`�a��h��\ �"O���R�8Ω� �@�s�Bŋ�"Oh�Q��P�x�`D�}�� �"O����ț�	��Z �	~�$�k�"O0�0pӜ6pЙ��<Rą�0"O�Le��"]��h4�	�_�0�"O
���j1��
�gE-2P�"O��â�5Qt�y���T��W"O
�@�o�$���h$�.��j�"OPɪ@��1G͂��4�ʄ��"O~�(g��!BѴ��
��p�ۀ"OE�%��61��Ɏ��@59�"O@9�	<C6��1G�\3S��蓔"O" 	�OU3q�TI�;����P"Oʉ7$Ry�,��U�D��"O~}z1lZ�"~����)43*�5"O��R0�߫oN9�0%߳*d���"OFt�שհ=����cѸb �#3"OYA��0/}����Z8I�R"O� ��T?0<*��Gˎ�8��0�"O�,�$Ī(Eje��ʂ�6@0r"O4R����?�^Ahr �����"O^������A�.މn�\��a"ODR�8:���-V��f%� "Oڵi��E�4z
r�	D�
4��"O0��c��mvʴB����jʌq`"O�q��N�>�0OH��jt�"O<�d�±+���)��(�����"O
|���$۾1��%�d�lE��"OY`q&��%k>��#�/N��8�T"O�K�(�8Ѿ�[7�Sd���"O��HG��*$eDk5J��*>X�"O�	��+�3s��[¨[�-60���"Oy#���g��p鶧���8��"O1��Z"��@B�aC�/"L��"OP%#�ځ1V��Y��=���K#"O$�S����Q�q�_�CV�p�"O���7�B����@F�C��X�"Ot�@F�B%�XU��T�oݒ�"O�  ��JW�x\1�qXĀP"Ot�Ro�$W�*da�ㄤB��%�w"Oڈp'�J�j��) %t�X`1�"OtY2թV*Wt�ș1BƖslli�"O0#*_�Osf�� ��O��J'"OjE�"a^�e����W�s�!��"O�٤/[36���%�`��2�"Oƨ�#ʂ�+Z��ٱ
�i/n�"O��w	3����ɺn!�"O��P
A!,�v�Р��6!�dp"O� � 	x0H���	$D�e"O�]�2kӶ:?*y9�O���Qc�"OT�X"��>��
G"wЄ��"O� ��;W�ڿ:T��s�HB;MЀAd"O���-q���J�Όfì���'�0H��Jr�3��!Y�l�C�'>v�q@�W�Jh���\���0�'Xٹ����r���A�B�)�r��'�n���+�R��q��L�N�P�'_�D��Q�WOx��#�Dd��y�'�Рk��N*�E�2�ȳ;���	�'�8\ط��	h ��P��/G�ꀢ�'�6<�����~đ񧛆F���'b@��H�@�Q����G�l|��'��0З`�6�����A�H@��'���@(�*b�)�B�ê,�Z���'ZM�� 5��}��C n���
�'�F��-�m: #A�ތk��4[
�'����D��ڲ%� ���d�r�{�'�A�!�ٺZd�uh��+A�p��'�Z�]dN��6B�"�)�'.�!���L�
L��&NS�l��l��'C$�`d�\a��؀��N��U3�'3���hL2�5@0�� |���
�'�z��� �
���,�)���ʓ������
U ��$��-9�ȓ8ZE[����T�*   �>.�̈́�z����I>��c$I6 #���e0�U�q(�R�z��w��$��(�j��R'[�_���1ӡK�$�ȓD�t�iv�
g�i���Ϳ�B��ȓ'��2�W�$��� �ȿ{<\q��&��0�S�ء5>�%�g��:"�HՇȓ`�H�����H����GS4_@LՅȓ(XQ����d`�۲�h]�ȓ~Z�&�"fx[RϜ-����ȓ�����H,��F'�t�����td&����<,B�dK�1��&5�b�K�}�0�H#���^h��ȓ��h��Ѡ�21�oG�N�p ��qdJL[�� �t�S�&��犸�ȓl(�#LOݼ,(l�.3Aj���=�����8 x����)IpЅ�[�l�7H���V�p��+4~5��*T�n�~����["o_,�ȓXx��_7�j ڕGW��=��#%|���#E�8���斎uఄȓ6��P1H��[���ɶ�U�2&�-�����ӧ�-R��ˠ�t	�%�ȓV}����ݛY��|s���f��X�ȓo�$��L�9l5c%��!1��ćȓK.�A0'�(5���0� �9`���ȓ"��l��9;��p8V
 0.�*%�ȓ�إ��Nٚ*UT顷░/��ȓ{N%�� �4/�ly� �9�r��$ޜ�7jnA(I��1O���D¤}���'��EP��.*��y�ȓl���@��_t0 �bN�"m�ȓD#l�� �qF���ŏ6h���ȓ\��l�ª�4IvP��Ā�]���LZ�s�/ķh�&挌I��܄�%�T(Ӄ�*RN*deB]rxԄ�+�ʐ5(�;k��!%N��f������э?C�D8CeG|_����&|��r��R5?s�a
�@	�I&|�ȓ[$�%F���p�Ɲ�4�
a�ȓS�8`�藞'X� ��Z5(l�P��S�? �i �«'㌕x&!ߙ!��Pj""Ov!V���Й�Ҁ 4q�\�B"OZًUdP/�b{����wh8kc"O�	J�ƙ&B"2l����)W⩊P"O���Pl�3���;�H*6$�F"O\AJ"��f�@���#�*���"ON 3A�X0B��+�bQlߠH��"O*H�Ib�f@B���$?�b�I�"O$�#�%ڱE�z��qK-��}r�"O��)g��&�v3ri�!�41�"O0-�Q��# � ��1�M�K���"O�X���-�dibGf����-=D���BLJ<��(a�i���1-=D�xᒟ/o��)P%&!���U�.D�d�3�K��*�J���|�l1�E.D�dQ�
��!MB��H@�k>f	�eE8D�@����.���61�i3+D����M�Y��]�0��K��%D�j�A,cX�S��ژT���u%D�����=��Qڒ��_��`a�&D���Bb��9Ϫ-�$ ��!Ph��h7D���P@������R��7<rx���8D�̣bFV.wF�h���	q �)��6D�ؘU"��I����(�[��,Cpc1D�d��� :��l�ċG.%$�fK-D��#G� (xHه��o4��,,D��P�{Q�d2f傝s�Tq��f+D�PX!�/q�q�U9_)H�:tg4D�9�����`L�w��O�N��g%D����B��ԙ�`-�dmdõ
$D�d6䕍SK��@ @3���A�"D��P�[�g���xL��_�0Q�<D�8z�� +�|�v�]
r"
1��G'D�0� )�#**����n/���h��&D��jGk{����R�1+@�5 ��(D�Lԇ�(�����&��PJ1G<D���o�4pW�(�u�X�
��8�#;D�42��Q�J��f֜U:��O7D�Ȓ��������A��,��1�8D�D�Q ~U��A��|k0@T`7D�8ѱ�l< hq�@��A�SE5D�!�G�-_�" ��&1'<�=��F'D�����V tԂ���>Ԥq��.0D�c$nM��,Ds���3fyx���0D���f�1���Tj߾O�f�+.D�D{���5f���'�A�Tm���+D��8�"Z�4p�HǸQP��`B7D��3e��<+��kN�SĈ��d5D��(�� �Tx,E"̎A�$H��G2D�Tc�
G�d�¥	���Sb�O;D��c�.�j�(�lؽ^b\�D%;D��㚵N��$�ӊ�Hkf��P$D�p:'��&�R8⑫��Z@z<�F� D�Hi�͉� ��	�1��\��y%�)D�8�F[�9��E�&e��0F(D�;"OX:^�����-�)>,����K&D�hI�n�9���kˎI����%D��k��G;����
 u��iBP�-D�`Jg�i�
�J��j�΄y�E-D���ǃC� }���	DO���E�+D��y��gF`q�w�@V~�)��6D�������%M��M�t4	��]z!��;�^� ��u���!ʼ^_!�DL�s�f4*���+tcP9�rmӨS!�� Ni�!�A. ��sT
w�z� �"OPY���ª�0
�bԚc�<�` "O���C�(%Uܸc�]�|��1j�"O��k���~���`�Ab?0�
�"O�pc��@�{G0�/]>3\(��"O����Ә
��EQ"E9F\�5"O �0���6M������O��҂"O�� 6 
2���t��\��ba"Ob[`��'p�RI�B��*S�8=��"O
ݺ�*�j��E��X�$��0ӕ"OP��p��^�Ū3��5r� �[0"O~P���O�?|���GU��J�ǒE�<A���z�x)l�z���f��<f�C�g	�	AfkĽ|ڜ`I�
�{�<1��@:t��AQ�94�T)�L�w�<�^.��d���f�꼳���q�<AT�:uY+�LFb����j�<Q��$��\��L%d�2�s�"Z�<��D��ej��٠Q>�hS��l�<�w�2�
 Nm��V�j�<�����-y�\ږd\_1�Y�lL[�<��솕<^,��m��%TaF�]K�<���	H�ȲaK��iKh�҂Ga�<���_�qìbt�F�j��񐥱�!��V'�&;�L�	4�Er#`J�o8!�D�8"�
I�E����0-_ ]"!�!n�:9���-l�`d�nK� !��7qD��'�+�*��0�K�Y�!�y��9DB ����7�A��!�dϝ?�v$+́�6����Al�&Y�!�)7�4hF �*�֌�ҪǬt!�$�[}b�Ĝ�G�&MaR�8�!�D�k	�T��
"�B��ɽtS!�D+o^�Q3#jK S�h�!�N.I!�Ĕ ���#7A����}�ƏE/O�!�I z~5`�"������\��!�$M5Qε���.�G	֞�!�D׺vI�@ �#R�>�ۡ�ϡ*�!�D��j�8���NJ�m�z��F��`�!�dR7Q��$q/D"p�k� ]{�!��^fLi���ܲF����2��p!�$��GWPyq��1[� 8�ƠS!�S�Iȕr�A��~�@5sQ-�>O!�d͋0t�M����I�\Ȣ�ʪ<!�ˊjD�easj��HpaC/�A?!�8������Ύ{e*'_3?!�$�(B(���c��l,!g�}�!���/�6���)]�H¦L�!���ky:��!�('�=�CѦ=
!�'P����́�bs���!:eN!�d� 7Z��;CB�L�f�����>!�0g� ���Ǔ�:\u�F��&!� uk��@�ՖR���3��_� �!�$�,�L@k&��D^H�͋�f�!�D��o���m�^aZи"A�S�!���.�U �!߲4(ȼ:b�ɇy!򤅆Q�0r�bY�8��`�&��+b!�7�ŨAaZ7S�РZ����N!��B�v ���F�%4�i�/�?(=!�D{�<y��I<"Ѻ��g�n!�䖉@/du  �mb�(J4��N!�Dٓ3��PV�ӵw]\I�е|���'�f�Ja�?\�N�[V#6TL��'���p���:RY��o3��0	��� p�K��ɒA�z�ENL��`(��"OE����*�h���SU���b"O�8�Ƃ	Ԡ=J�B�
o>,�"Oh �0K4?֍ِbσ-;� �b"O�c@a�Qߴh u�Q.G��11"OPU�'f�=;|r��T�j�`2"O|��N�Q��j�$�'9��e�"O���悟�<���B�@�_�<�{�"O`��SNU4KLJF�öo��$��"Oƕ
'�;^�8c�єx���&"O
��1HCk/�DX�-X�G���@�"O؝P��Z��у#��><`)�"O�x��%Ȧ1�d"t$H	hش �a"O ���!�|U�f�Y�y�\�w"O��"� #)=V��p�V(jhv�S"O��F-�7l\��H�=��ݘ�"O ��5.�%��B�%_�|}��A"O�i
3�߰q�ڤ�!d�9j��?�y�mXd	I"M����
S+��yR��<^�)�@�(=����y�9�L��Տ�?kr!⑆�(�y� H7B��HV�+CT
����  �y��Dh���{e��>b�i�sb$�y��"����Y�6T�+�%���y�H$\\��ui��y,�Y�g�-�yb%��w�^|��j�xY�=S`ႁ�y҂E�_l�ZB�D\�v0*p��*�y��ӍaV�#C�'�:쁔g���yb(�9B㚱 ��2&���rBW��y�ܹXr�P�A?��0Bh�7�y�"C'��Ȕ�~���s�?�yRֻT�n�d�@�z�F�k�n]��y�/�Q�\��R��G04��bZ�y"�	I�Y�2g%D�չ�nF1�yBo��c���+6��/ 4�b����ybOT�s��\�@��n$�y��Ug�����3��8����y�dYӶ����5�xY�e�*�y� �*ӂ��ǌ]&1���qF(��y"�Խq3-� �ځz�Y�Ę-�yR��1��<���SkΤ9 ছ+�y��'DJ��q#؏k�yzg̜��y"��9��	���2!V!tDV��y"��g�0�s��7�Zı�̃��y�.�|�(� �"�>Z�H� �T(�y����8k�TP@�g�n�K����yR��HxL��A;g�D3���yR�<	F֭��JƣK�@��"C��y&Գ?�h��kT#p.^�RB����y�<i��0`�gֽ|�R 9�䐺�y�ݖ޶�q"J>���(#F�8�y�\fw"UCA�'�������yB�aKf(�L,9vL��m�yb �;dl�R`� �|{�bM��yRJA�	Q�|��[�EJ��j��
��y�@�zڐA��ɚ$2��قѡ���y2ꐫW�9ASI�(�y1`&�yrk�'5b<Ѐ����%GX�PdԾ�yB�חM�ҵ�áy\HH3Ɋ��yR�O����.ԼC#r]����y���|[��!���-�N����<�yb-��� � �t�����h��y≟�'H��1�S�l\�p�Rg���y$
"|(�@om���/��y
� ^M���)G�x)0w͘����"Or`�@⺌��O�V����"O ����F)�`��G�g°��b"O
đF�	�Ng�����^)5Lj��6"O�´,��Zw��L=j�o|�<yQ�7P�ՐS+W$����`JN�<���
&1,ԫ�( V��G�G�<�L��m��%F�4Kg��<� T�V��|qV�6.l�+�b�z�<)��G�;�
�[ӥک °�9�c(D�Ļ�Io�H���:���` 'D�$�Vd�����To��X�~%i�j?D��jQ$̔����hΠ;�͐��9D��K�l�<D<�ʇe��D�6D�LZ�G��2�|��e�Z�W��� 3D��C4n:~h$}���˗|�Ƥp�O>D�� ��X�܀�S��7(�����<D��Ye��1����rh�Hx��&;D� �'N�K�ܐĊ��@�v��u4D�(æ�\;E=�	P�
�'FX=y3�7D�x�`�W2����cʉ>��*��'D��0��w�X��)>�ɲd%D�x��� \yz�"	6I��|��5D��dM� �UP�ҭ�L����
�y�%H, �"u��¾8����Ď�	�yR�\=~�ш��FZ ��	��y���I"��3��ݺB+x����5�y�Ʉ8u�ĵ��ʲ6YT�!Ņ�-�y��$p�� 6�G�+
��H�Q��yb��"}�5-��s�:����#�y��Z�vi>2�ʔ�p��ir�\'�y҃R�R�eM�#\fv��&�
5�y2G]1�tB��@3K��\���ƌ�y�MC#V��h�ʦ=?Ј������yB�U�z�8�KV�i�r�҉�y��͟t9�}��^�="��h�oV4�yb�Sxa��Q�� =1GD��T�Z��yBo�� 7�P��J�$f�ZUhҩ�yR��1!~�3�W��6,$���yr�ݺ,�6, � �&8{����y"h��]���Zt�ƣ�֬��Ë.�yr M�fg�I3P��2�3Ѓ���y�i[�r�0�oϻ<�^ 17�8�y�oho8�D���.a0R����y2�J�4��p�%�T(ʗN�1�y2lM4R��u��^'",v؁f��y�@�cM �`IΓL�	K$�y��@-X�s�g��+;H2u�D��y"m���T)�"B�Y�jdXt-[��yr��4�~5��PYj��c���y�iF'm!(�آ͚�@
���͚�y��Ҟw� ��cKS83����@���y�K�K>ֵ�G �99X�hv�]��yr�,L�2a��i�5/Fĸ����5�y�cL�W�AH��,,���ŮJ��y��P�p1jQ{`�[,*	f���NB��y�#<%���# ]�nR@�2�K�y�l7 V�)WÑ/(�|�/]��y"�ؼ�*�;Ca�\��+�����yr&�d��������Z����y��:��!X��(Bj�$r�M
3�y��C�;|.��%�l������y�f�6TGr��,G�yԬx�N�y��@��@���Ei��
d� �y
� >-bፒ��09�L��~v>�SG"O��HTO�;)H���d��Yy�Q��"O�A��CD�(К�8���Lr� "O|D�b��%z�����8� �+P"O�8sr�B<f(��x�g�{�L���"Oj�� MP�<��'��>6�8\� "O�<�c���xD��S"C��|y�@��"O�I�ϒ+Q�*\`'aN':_p-K"Ov9`��R�1]�,hQ���l��U "O�CB��kU$ٵ��.R��'"Oh�闊E�y�Ɂ�g�T���"Oư*5�0ᄼh��܂Y��+"OB���HF�2j�.Ak�|���"O�����:I�\�t�To��� "O$�'N/&�$8����BI�g"O�*2G�7W���r�j�=�0my�"O�M�p�[T����×%?����"O:�b֠�+}N�l
`HA�@�M�"On�J��C�B��5۴A�|�NP W"OH�a5�}D�`�K]�`����v"Ou��'��z�F@3R*ΛO�*��"O�8�%F@�l��t.
�/��uW"O��Q�ćF캗��>��q3"O�{��Z�1�@�E�C�αB�"O$Iy)�#%B�Hwˊ�b1kg"O�p�AƼ8:n0Jw*[�'��q�"O���&Ϣsΐsc�:�K#"O|��AW��bQlx5��"Od��N/3րz�A�c����"O�q��BN��k0O�5j`4Z�"O�Y��A�l�^�򤎖9dT�R�"OtQ���@��:� �[�1�E"O4\q�)p  ��!��,=V@	�"O�Ia��ЋdE�tdߎm�h�8�"O�a�BB˴ 1N qg�G�@��Q�"O��)釂6������gG�Y�"OH�a����ه%�3�F�m�,B䉴�P����ޓN�E��o�& B�'E{�����K�	�B,ܻA��C�ɈHm�$�9w�#Q��a��C�7��2e䁕ư�P�
V5g�C䉧�XA�tl ����a�q�C�	m�>��W0�����ԉu~<B�	�L��	��_� 8�1@T���B��C��0i�H����%�dX��D�
�C�I�
U�ˢD�/^�^X{�`�SR�C�I�RL0��O<V��eU.��p�\B�Ɏ+��k���j�6E@@bőg�B�I=g�"d��h��i"�QFOF0��B䉆t8�
E`�bw��He� �\�jC�I"
8`��υ7���ڠH��+�C�;hG,uy$	O�l���o�e�\C䉦4�EH�h^�A�AF:�B�ɐ������Vx��v��9?�C�I7����Q'>5�$1�#c@'u�B�	Dv� ��<-N��� �jY�C��(dS��o�K��y�/�t�C�	�q@��R��<0s����-g�C�ɧF��@��˓R���)UM�=��C䉱P�\��ѷ7�fM�-̑s��C��31��[*m���(�rC�I�[�1��c����Ce�,C�	>�F��S/U�i��!���&��C�	�$ox$�d�"lάHF�D�!��C�)� �10�`R�x��Q۶g���S"O�{�Ȉ8�J�Z�A��T��	�g"O��H�ӏcr��p���m޺���"OPHAq�WG�� w��Fي8��"O��#�)V.Aرo�B�x��"O(j.v�0-P����k��#7"OxU3�/�){dyc����)�b"O\�gBF1ݐ��� K���Ti"OPp�� ��<�@�[*�csz�:�"Oz�R�G�
m;|M���[2J��Ƀ"O@ȱ�J^�}��qq��/X�ȃ"O��:��[g����F�7)�ʠXS"O����*@"y�$'�'�m*�"O�ԡgG<IE��d%ԁY||�ٰ"OFm�C�#$m2<2ծ
:q&ȡ"O$��FKT.T-�J��ǰUp�p;R"O*��b��Y��վ<^� +b"O�1*���% `6��2-�""ON4�0ECq
u@B�W�!�>}B�"O����Lޠn��А"�����}Y�"O\(�GML�j�:���IтW�8���"OR���d1U���[�!FEZ"O����X=C��;A��S�y�"O��lE#fz��IR]��	zF"O�4!t���r������Q} �� "O�<`�%M���BD\D<y�"O���N�0NK��� ��/LUI�"O
$��BK���u��"�ͨ"O���f��lW���,O@����"O<�!7gV�B��!A�C?.�Z!��"O�9���Q/yz6�ص�V�4��	��"O&9sO�y3�x�qΌw��0D"O (��M/u�`R#��0q�AF"O�Q�SmI��q�L��?�^I�Q"OF��LEL�\�KT����	!"O�-R�J$���&�{EĹ��"O�q�`%כO�>�sR���>(&���"O��I�	ɳt� �Q��K�'zi	�"Oj��EbZ����v��	T�*!�"O������a��p4���h��T"O24C�σe����d��L\RA"O�a
6l�*�����Gn�H�2"O$��q�9  P������]}����"O����-|�hy� sjD���"O�7�I�m!L���hA�9��H�"O����ӨQ8EAF/|�4�;R"O6�8-�EE001�&҅ =��!$"O�� ��,R�x�zq�'h��0"O�]	�
�D�l!R'��x
Y��"O�, ��'�4	� !�*p�"O���3�Ѫ4 ��A��2X��z@"O<�Q��q��Yّ�ʝpnhD+�"ODU�C$O-$�b�U�օ4g���"O.u�Ǫ�:�fXďhZ���"O����T�%5Xt�q�� N��"OޘөF�.����!�;��J�"O���oQ�9�цkǠg���"O���J��V������	{U�M�"O�h��nжj�(��
Q�K:f�J6"O�"�I�p���C�ʗ�?��{�"O4�s�,�3����vv�"�"O�d1�W�,�z��/$u�"O�P[u-
T��*�`0 �"O@���@.
�� ����R"O�  �³�Fk��F��`���;6"O�8��'y����եT<k��P��"O�Ȗo�� ���k�䁅n�p��"Ob@��EJ�n���4�U�C�8�
�"Ox�b7��D�|8����"d����#"O|��B�$fr5��E	+z����"O���������N	�	��+�"O*]���������R:��څ"O�EdN"�D-9@�Ya�N̓�"Ojp�fN�D$�D��8W7� 1f"O���CW�z;�tr��C/��ZC"O4��S�ܱ]zZ�f��;"I<L%"O��s�H�Nq�K�M8�Y�O���7m�I�D�J��& �@^C�<Q��s��!�E��#{:1S@��e�<en�%6��i�'������J)|�<Ye���vn�I	ņ[�Z(��ץK��hO?�{;�0i�EJ�dgBQqf��rF�C�	�,�r���X	)x��S�T��RC�IG�~uj��=*9~�
`'��b�b���/��$��E�d� }	f5���0!򄆭�YQ7!�	<��|7:kYax��I'[�4<9E��g�ҙ煌R�\C�I�1�tdq�ʗT"��8`!O�"�^����Y�L�"�b52�ʃ9q.L@�"O��vNU$a��k�i��>XFᐧ"OޥTi��2���R�H_$oF�d�G"O `��@����7�Y�a�NIR"O�@ê[��d�1���S��u���	�0|Jb�	h�輐ш�D������s�<I&N˂A�q�T]�raD��V����>�G��2��9�n�IT�ARA��O�<�E� -_������Q8��2�r�d/�S��)�JUy��w�Yx橑�\�0��V��0���<:p�˰�e�ra�ȓ+t0�"���� �3g!�D��4�ȓF=���1��0W�vM��#�2v��-q�'/Э�jҠ;��4��N(_�t\����)�t���2S�A���	?N6H̹E���Px�iK��Xա�4kxcT
^�jD~�"�'_J�K6��6i
����G a~|��.���3U^F�J���>����U�C�I�Z�]��c$��REeQ(=�#>a���[J@��WeH+$��-���
K�!��O��	RU��:��9�ǆ��i��z��%�/�.ypvl�>2~��#�UN;tB�ɮ4f��2EG�K;L=�-��O�>x�ƓfU�䛒/�d�nY
��X�T���� �M��y��ӊ ' %��+�s�b�3�b̉�yR�*bQs7M�;6�\x��b�
�0<���$��H�TlK�a\fxT$��y~!�J�$���b���)$���5� �HaxB�ɵr(e��J�Y�x��ݖt�"C�I�aIQ!o��v�B�X���1;F C�8AV�b1���Mml���hs��B䉫{����@M/��H�Ն�+C-*�D�>y�Z��%>���~��˴A�z	����+ �|��n ߰?��'�*<0�Mnľ�ᇪ�4H��q����M�'�%,O5i��4i(�a�{��!q�ə&�Q?y�@,\�f���GLX��� �#�O��eX^xkQf�&HT�#�c$Lh�m���y?q��d�~څMV�%kv�' T�g��i�Vd�@�'�"�i�Q>���c�FXj�C��<}2ŠcM ��-�O8xPP��/*� 0h�M3^d�b�'W�������j� x��oخt�l*��D0t��F"O�u�IMJ/ք8q.��z5TQ��xB�{��hO"��1���zJ��y���M�M B"O�]�i̖E+`i�Ul,);�|�>Ƀ˄Xwp��)g��'Πl�Gi&;@���J6�v�ד!̶�O0��@bQ�p��dbU�S��+��. ���DǕ�C2A
L�fg��60F���O����#K�S;�ybf%�#^n4mK(<iu��a�6욵Q�}�@�s�
�M��8k�{��\�d�0��g�>�`��C�yBʚ�T���۷�`�C��=��'ў�Oܼ���,?fx�3c
]�:�r�#��HO8��dg�1`�����a˔���i��$���L�p��aF�+�넠*�!�Ě-G�z���7)�YIlms�C䉮lv-���!�8@H���v1�C�<�d���G=�$٥�Z$*�B�	�nL�s���4��$2p�2o��C�ɏH��U �p
��"��$xpC�Iv��h �7/&�<r6F`C��N��PR�׋ko|�Z���+l�8C䉇`Vީ0D��#2�Vt��$�OF:B�ɥ}O�[s��W��\��A!n�C�漴�K7_ζ��@K����C�I�N���'�Y�0���*�C��M=��� L*6-NAٕDF�x�C�I�p��ݙ��F, 	baä0I�B��4����� B ��"����dB�	���Uj� �U <1: _P~C�	���p��W,&� =`���) �xC�I?���$��\ �f��`;:C䉵s��4A͝x4���ŏknC�	IԪ����O��"l���C! �B��$@��mѮ5ȍ�����B�I�� ;%#L��Y�g ,]"B�	C�b��� ��(@]:  )(�BC䉗;��`�V
�H^y��@�%vB�I$ks@`��R�y`�(�ڋoC�C��,w3�u	��r�x�HvMV�(܊C�IJߎ��h�$f�\Hd��YVC�ə=j�4�f�
����$�ҭB�@C��5Qi�d�pC7u:�f���E�C�	�|�P��ҙe�9h��	"��C�IE�<���"V�,��0��A�>B�I�YC��p���"����p\x�B䉞O��nP0�F��S�D�B�ɻ8ĉ�e��h1Vp�B-i�C�
��yQ�F�/�j�*��x��C�	-}�<��j��P>$D�s�:"��C��6�dDUm�<M�d�6��2W^C䉯iT�l{1�׾RH o;yRC�ɛ;�B�0E��~�^e[SLÈw�C�ɛˠ)���$�PA�p*���B�	�mx�����s�6티� \�C�ɟC�B��𾐊wh�UW�!HW	0T���6��h�V��ĆAZ�t��"OFt��G�9:l�1�q�۰W�jA�G"O� �f��*���y��Y���bA"O�T���\!����#Js��"O�P�%��8�`�P�-k��)f"O�	QBG^���Q!�Y�Rr���1"O�!8�\�?��Q��\�)]b̢"O:�8�Ȏ:#[F
3��<JW��*�"O��3��2���K�,�� ��P"O� �-�#\-��(�F߀P�t<��"O��x��\+�8UJ�&��+�"�"O��I^'p�d�[�E\�Sp��ht"O�m��$��	����D�IV���"O�A�ԡ���<śdٞ7���Z�"OX��ѪڻTհ9�@+@�R�,I�`"Of�a�ĝ�)cR��q���!�h�%"O@����*N��)���3H�6 ڔ"O��
�KL�b�\\:@���~��X�"O�X����iC�в4�G�!��D�p"O]cNi��9[��ٴ{�1qc"O�4�Gk,�|H�eM"�B8��"O*� U�ð`��)�����#k����"O�(�gViȮ|����Ji�ԑ"O�	�� ��g�}�P�B9Kr�$"OV1��U�Y�	��`�k���@"O=�`�6B�,�F�-��=��"O� ��a)��1+�m��\�a"OVU8u˜\?܁�u��}�h��"O|!�1嗆ʦ���B��\p��"Oj}��CJ62@~�{�a@�T�p�"O�Tj�Ė���ړ���PDR"O�Q+6��?�|�2�#
�X�H��"O��9�*ݑ2I���!��B��9�S"OUf�{$�L���9��;�"O����*η'���aUKݾc�$U"O�ѳ�/k�=[��@�"�:ݠw"OX�RE�җB�t5��˙"2�]��"Ǒb#�ۢK�A��K:X~�Q�G"OR�낄Ƈ$2���ұn~T`��"O@0C�	�|b���i��hvU�"O�Q(T���}��X��Z�[��a�"O@ڵOG.~g,�yҰt�\x*a"Or�s�욁nz`�Q k��`��a%"O8HYb�۝KF՘��ظ;�,��"O4���lã�E�#��f���"O�:�ǋ�8���5u��r�"O0s��=,\h$��+��7�2#"O�ի%�!��ajS��=)lLp"O�x0�޺pAr��BO%o=��@�"O�a���E����'.�U��@�`"O88iA �$��\˳mS�F-$`�"O�!s���&T�u����t�C��+�x�u�C7n7<�(֎�C�I�y�"���Ņ:�.	�c��>X~C�8�|E��R�j�:��͏-C$C��q��8���ō&�{q��J�C䉊,�ĩ"$��[/�؉�-֓L
�B�I�z1�`��)�p�r���CE�C�ɵ]e���{���6�׾C�	�oo������T�P�4�Z(T8�C�	�"���+e/��1%�԰Gi�%D��C�ɝ�vP���C��-`df�uͬC��h �<!��M6�d��eŉBB�ɂE���C��Qиx(�%ЌYB�I���j�"=Xz��� ��C䉵m��Ѕʃ�Lj���0W�B��1�ʥ����g��$��>nRB�I��Z(�7�]�K��T�`��i��C��W�
%�b,�9��"f!�!V.B�ɦAh��@�(3_*�BQm� B�I�WZ-z���4�PP�WP�b��C䉬)��k2dP�6c�ka/�&I}nC�	:��e�ᅛ�L��a(�"͑d0�B�)� 2�!VB��,��ճ��إw�V�+�"O`iP�BV��(<��+���e"O:JCKK�?�8�b*U�}� t�"O�`1��'����c(]FH����"O�ɘ�-û:<����'I���Q8"O��@&��x$X�q-�=,q�KP"O4]�"*Xݠ��V�@�SY<�C"O���
K����I��nMx���"O.-Su�G*B+j=�P!D� I6��'"OT]B��40��U�G�P�k=�`aW"O} S�̪O>p�B+�Q.��"F"Or��2�D6E̺y��C����A�"O�|C�.�2#f<�`�E��rlw"OH�@gڛ<��d �
��zǮ�r"O�4cI���� �*]�F���"O����u�bA�j�g4��W"O6c�N_0�\�R�Ϯ:��M��"Or�E�,dH�ƈ/�� iP"O�Ѡd@��4�F�U Q"�#@"O��;p $eWJ@��+�H�Q8�"Oиc4�ÙcN�	r*�5R%�Y��"O��#H�6i�Z<���֩;C�$ؕ"OlT&��!�V�BiĹD,�Z7"O�D�C�//�l�*p��/��9�"O2}(��(TY�5j�ŉ��R�"OX��D�SA��B*lx۱�$;�$;�'/r��"��L�O����Xo��a�ȓ V��#��p.�����]wH��Rb���4�ɫ2i�H*��̈́ȓW���XR�`��Y���s��Ʉȓ��U�V��=x����Z�g�($�����.ҬH�����
m�Іȓp�Pd�C����D�Q���ȓ;��Tص�?�(�S ��ec ��ȓޔ3������G!�d��ȓ!��@�E�Y$?�Zm�K	 !o)�ȓq��q�S��$`<)"K�SkU��)��9X��@�&%��c���4C��Є�d� �X���;b���rۯ��@$����I����o���\��e�i� (�ȓ)��tK��2%�r��W�*	�����O���O���󒅑q9�Ԡd�|R�)�SJ�^QI�H�����
�%U�C�	�4E��A$��P'|T�"ON���
2���x�k��o
́��'sў�Z��: P ��OT�#�Qs�L5D����K9X��U�-����)7D��ǯU�SF܌0�Ǖ8��5�9D�p�E��l����#Hv��9D���d	�
����/ĕ������"D��Ӥǈ�^��{��]!�p�ٗ�>�	m��ħxy�`	�-c*��%��.x�.	��X���rD��D?���F�r�v���M9�#�_�h��uP����KRPF{r�O��� t�,bXQ� �^����'4t@R�R�?��xI��F E]� ��'�,p��R�)�l�qP�E�~l��'�و \ |H�	�GgY���0!K>1�'4qOq�n�[0��9uv�m����4ܜ�
p"O�)�Acb��ȍ�cl�2� D������cVi8"C��%�b4Ȥ!D�V�^���X�� �<�8�2�*,D�|c�A!U?����^�y9ق�k�����+��1�cD�J�����	��C�)� (���՗l�Q{wF�t�t�V"O�T�5#΅��@c�ꟹ�v�0�"O����y��D����u����R"Od��F��� �vhX����b)�S��?��iQ>[zL��ό/9�8��t�R�~"�'5`U3V�Q�z���0Sl��w���x�����ofyqm(2��z$���0>�K>1ԇӂJ�Xh�!G�3m�\T#ZJyr�'7�H�i�\6��q%�#<�1���hO�h�r�	�W�&��� +)�,p0�i-��dD%�[�H�(�Z�C�S=!��0�9� �a��E"կ.t��
O�-��@ωA��u��^�\�*uK�"ODX�ӁP
V8���$P��9�"O�`Y#�ͪ
4]�ǧH�� A�"OΕ����Bok�<UZ�I2"O\`�e�<!����%�+,���b�"O>\��nC��=R�V%���A�"O��2�M��Ā,��.a��홑"O��*6�A�[�D�r�^',�jH��'��O�(I�(
�}��]�6�]�sɼ�@"Onp�ņ��QA&����,Ģ�I`"O
M`��*)T�&��2"BM��"O��&l�*���	��Ѱ,ν˅"O�I��Ɯ�����dْ��A�E"O6l�P(�*d^��
F�O�� Q�"O���.	�BT�q;��ސ!�z�w"O�@ � 5e	@E9�� �H	8�*Od�0֤[n�L�W �>i��2�'�F���!� ܮ4���2f����'j(x��F�����4$8�C�'��2��Nh��Z�^��A��'Y�����&�r��(��^F��(�'�����'��'���BӌєL�Z%b
�'�t��1�CR�D�I�
98�'�`��c�W�,���DL�������'��eʄ���y%^-���zF ��'��I���,*JQ���Q�w��is�'q����\�n~����X�|�	�')v	��O�C*�T�DA�2M�0��'҄�bG� �0��9�+ɛ=��=��'^�Y�X ^~���Í�-��U�
�'��-��Oexv5��d��&�:]I
�'����U"�����lO`��'��
1Ņ\�l�bX�f�\��
�'61�c�\�UHn����.R},Q�'������}�aS��?B�Ra�	�'l%���UӴň$�V�:��-0	�'�:�Q(	a�t�sK� aDށ��']t	� �٤T���s�U\rԱ
�'N�|���"6	�o͜Xڸ,��'��i�݃=DY�b�C9X�h�'׸H�"��*Cfr�48���9	�'I>ܸqB��4 ���1��&����'��{N�#@����Ȓ ��h{�'C�}S#�ۖ�䫵υ'�@2�'����+�400�õA�Z(k�'r�L�`�C�bE��8ROZK����'@��G� ,��`a�E.@/�<��'^�"��S#NsHH�N�8p )��'�P!J�4b����D�$J�'�����´Y�l�ם?���'GX5�WƎ,.d&=P��4K���)�'*䌙�%6�&�Y�-�F����� �$�W��v8�P)��&R)�"Om��O�p�L���k�##O�})S"O`�����vmR����ÖCD���"O\�jW�O�tdL�h�"�%��qq"Or�&jͫl@I:�ɘ~ژS"OV��<})�4�,�1|��	&"OUJq�O�9x���M�=i�"���"O�Z�k��Jޖ@�eɜd����C"O�<�� S29uf���G�xD�B"O � �t*.$9�a�~.��V"O<������<$�Qf[�
_(��"O���"'�{ɘ�;s%�)R�V�'"OH	��V"�>e9�i )s�"l�w"O�m�T��Tf�kwȀ�W\�Cb"O���)�j�����gSB�y@�"O:tÃ��IiN1i���:}�&!Y�"Olx�"�(|�1��ҋ]]^�a�"OȽ�%]S��� �CI$��"O��p��ծ����1b�oFj��%"O84C�
��"���:3� 1�,}�"O�9î[�b�� -D0������yr��1$�z,��A���q��b�.�y�h�j�=ʧ���%#U-���y�gN����X�>��Hd�N��y�S�Zf�$��T&l014�
7�y ��N�rggY�@�� S�yB�Ш �4KP��wW$@"����y�O��k�����[5i1��
����y�L˾{�x̘�NT�:I����y�#/�Vh:��T��*Qc5����y��%qp�����/"ql�Y�+�yB-7s.��/�|^
G
�yY+�
86��J���5ߤ�y�m���\ 'Ö���\�4o��yr�� ]���jG�eTk�
��y���K�l p���{ TY���R�y���3%��i$�J�(D`,Q0�	�y��^�:��E��͜O��C�� �yr�>��ܸ���(:��zF�ݡ�y����9�ށɅ�b&��0���y�AŻd�L�3�M�Y,��8P��,�y�A� �|�p��AΊ�)��R�y�Ã�]Պ�`��*1��
��D$�y2����42!@ߧ>���W/��y�,���(*#g��5����(�yb�ԯSe$l��hB�:B ���G�y���8 6)sb&
�hyl��$A*�yb��;"��'�b��H2t�݌Ǹ'k:%B��t����8v,L>��^�O�(@h@��-X�d�A���I�<�@�%f�,���ue^(���Mi�<6S ,�mi@M@�IG��k�<���	�=e��ǃ;>����P�����V�HU�)#��<[����D�� ��"B >[��J� �|��n:� Q��3W������;O@.���ɀ��a�����HY2Y�B��ȓ�F��0��z��!�JȰ?X4�ȓ'oܕ#�*H�y,����'��g��m�ȓ\%)��'B#@ƖY!
A��ȓ)=6�*kǄl]�]��aC�
h�]�ȓ8�|Sਕ�;�5Ȑe،�� ���ŧ���uY�
"�*h�ȓRZ�p4m�%b ��O[g5D���O��&�I��>�6ǀA{�Յ�S�? �\�;�<�Q�F>-�y�'"O�53$�(�)f��4�y��UB��6�����i�% ��ȓ^��ٓ��q�p@����-�v���J�h,�E-�H���+Q;@��f��)�F-��jζ���χ�m�m��E�f�A� R��lzt��X�D���ڼ� t���4T2��ۺr:��K��!��:a��)���¶/=R��ȓ}vT|�b�I4g��AV	I�d���q����D�ɴD��b�B�*~���Q�Ik%�³:�|�h[>x���ȓ
V�f���06��` �-o�$؄����JG�I�E��e���Rm
~��ȓx�`�m^+6��pIdk�'i�@��3D�X�6^����"@�8�ч�q]��뵏�*��
`͟��(��ȓ_�|���ȁH�P��S$/=���k�u1���(�<#����X��/3�œ��a�XS'�b�� -�P��N^"5�*��cLX�k�`x�ȓnÎ� ��c�ȣbbK>��Ņȓf<43K�[���p�˅C:���eZ�;������ӡ'�	s��ȓ%rJma��:��1"�P�Zp��c��#6iO�6�Ƥ�.%��B�+�hA*�(߰W����3�?aynB䉲/��85ɕ>l%�\r�o�[JB䉙K�z���H/NΈ�Q�z^B�	xH�-�Ɵ�F;ɑ!�!dB䉳D��D��޾n��  ��M�n`B��!׮ep�Q�'������
�C�ɊYf�|:5�='���+�NơS�C�	&x� %e�6Y�(2��y��C�ɒ Ov��LW�O��e�ѭ ��C��%0�(�cC�#H�q��N���C�ɪ)f����9gW,a	v&�-n*C��6�6#���"���'`@-.��B䉂\a�|ꔃ�0o�f�y��O�C䉳7V�ӳh�z6R4�Eϛ�[MC䉞d��t1S��$*}�c�h����	�3�H���'�*�c3Ƒ�h���d��5��5`��(0��`��n\��Պ ��� =.�:����O�nZ!���;(��	��J1�X�����E=1OZ��䡄G9��2��0�(�ꔫ��,i>(�go���"OB(���Ɂ<��z��,I�y����#Yؔ�soˬV��DX�*.��6]Ry����)x¤��$Ȍ�6/��Ɠ�Q`7��hĜ�����
�"�ju��tR��&�L�	��5��1��{c Ь
��h���<]O`��I�X\�����|���tfP�2^�����F�p"��Űww���3O8d�Æ�-iȨS�u�zXд�x�Ԩ9��� )�r֨
�E�Y�'3'd�P����Y2��/=��]�ȓ"i�h�d�	$���q6(�>S��!b2�s@��x��Zf����`�'��MT&1�)D����E˚0O��*��$D&&v]J7@�*L��G�J�M�RL
���&q	�ؑ�A��<�2�
M񾸲FB�e� y���BS8���j�Yj���	��G�*�"կ8��a$F�Y9�FV�T���N�]�0�3��}��DQ(A����'+<�۲k��U�XŃ'	�N��Q��3��k�Z�9��(jD�M B䉂n���Csȍ�3�q2�S�J T��hO=2��[� �$I@���yJ<YW��8 ����00r�H� *Ma؟V� Q�=�r�H�wL��&Η>0A�)�葢.?�� 7G��o�n�3C�\2�<�w��y�$�y�٤!�\�m_�'�:ݹ'�R�Dx�mRҮ�[����L�@Y�6�gx�p��,mvn$�O� �8b%ǌ�Hla�Ǩ�'�l!W�O~Hb0˛�E%�@��Gi��fG���!�$�(X.pM���	� ����u"O�YB�H$jjp	��Ժ+A@��2̙%L�d��!�� ~@���$ը)��/��&����ʌ+oP�� ǩO�H��S
#�O~�	��P]�R�o��j�t�-J�x)
uX5�Z�0����jޮ0���0<O&��CG�!��T�E���#*~m���I�6y����,��� �$�hV�QB��N�_�]×n6E�Dr�h�c�m2	�'5*���� J_>C�W8^�i:�'�&���R34(`]�#Ŝ�e9<����H\<c?�zE%
 ��8���#���G-D����=�	B7P�(J�0��K�L��a"v�%��J�.���
!�J<A�`�v�<i҇��9d;�8I$��i��,
ԣ�v�b��[�`�H5e�;T͖ ���_�/��-Е��RX��C��ܸ'�νB��u}���*z6�s��U�2$�t�a�P6��O>�z/�!y�ā*���h?V ���*W�詨ш�]������
'��CSJ�Z��vo%�m)@�i�l@.m&����	`�\A�f�����#G��Q&N'k"T�)��@�l'q��0h�B�	A����ϟX�X�f��s&�0�egh�#���t�ʍ1�,��x�P4��W�'5bYz�m� �b��WMq��靵vm0'���գC�*!|@��0i~b+c�9�O��P6�<��F/1�����P�(��	{E�P�xi����L�
�R�=��&D�zH�-�V�9��RqJY�m��y���ɛB�8�؇�߫��5�O��*�\�!� nֱ��cڏ_�*����I�-�6�4�YF�'�1Xˈ�aq��p#D�lc��O����Ě#Nt+S(�&e�8�%��p�O0�S�"ېR��L��K��V�q�'�T�w�L�����(��G�4°�E�s"T�jH�}�v$0DH"��'��'C�i��}F���mߕ|[1����Q�wJ��n��:7�4PS���lY��k�D\(Z�Θ�3#����b?\O̕(��ݝ^PrVO͘FۘĚ��'&6����0��=�E���db@m�!q>��V圮&���A�a4D��S��E9#������U�=��"0�g\ B�*!�H����GR�<#�P�1��8-����KTB�p�N� X�B�$7��|�ȓa��c! ��*}
L��.
/L�6��ȓ]��,����6�TE�w�[/u+�ɄȓP���c�fߵ23�Ƞk�*3��̄�C�݊SN��d���ۜ-�>��ȓ2:-:�ER�;g Y2%�#)h䴄�U�ܩ#G͚3E�  dрB7 ���[/$����O����J��x��?�� �C�\4Ix�	a�:����ȓ1Sҁ��L�7��|Ab��x@�\�ȓ9��Q�Ƃ? |6���J<y��p���%��<ѻ0+��j�>��fبW/��\*�L�V��DS�ɇȓ`�� rb�jp���処I�Z���&%���T�d����H%LU�A�ȓ&����F]#k��T����-��ȓd�H!e ��r&@虂�ԍf�ph�����j0枠S+Y�ĉ�B�5�ȓu�x�t��
�@e��e�2�v��ȓf/�icpg� c�l�ː��j]fa�����E�ʹ�~�K&£uq�5��|oN�T�X�2��ࣂ��pGȓ~Hb͑U C0"C���W�B�K�A�ȓC���$Ύ������G�P̄�ڊE�t`�g�$s�c�7s�`ņȓi:�+1l�<�l}�#��	oP}�ȓm���eߝ7�8h�7H������ȓz*h|�Bfm��]���w(I�ȓ)obl��%֢$�"DH��a���ȓ@�č;d턗O_�ݓf�	%B�p��N���T+I���6&]&����'�h���I�+��l	�J�p��ub�'�Ġp�S).۶<�S�I?i�&�*�'���a�	�R�����̗=�M���� ��X�8z^8��d]��h�T"O��Q�@�7E<I��$��w!�"Onx�Q�ޅWs64�$I��'p�qc'"O�%"$�<B��=*u�1AZ��c�"OF�CW�D���)GBC�M�� "O �JQ6U9
�p��#v��"O�0��ǂ�o����t�Ȝp�V"O��Z��^'���7�G>�D��"O�AxƤ�u5�4�A��Z���2"O浂�hV
1�Α���%(d,�"O����"�*��[FF���xe�4"OL�
T(S�V�ic�GZt �Z�"O}���`�|y��@�+cl~ �v"Oְ���*z6���G/��B��f"O�l3�K����g��!�Dћ@"OX-⑁N�:�+EkI>}���S"O��!*+�t�*aE�)���"OHP8��۶W���g#ɥ�hЀ�"Ob�т��?/���:�Ǩ��A�"O"-i3���E���@��ʜ$����"O8� 2Ջ"��(���"ȐT �"O�8(�,G!q\�4� %úFZ�h8�"O��H��ң��i��'?{(�CS"O}X���R��q�#DRzu"O�����>qL�����)9v���"O���Fɼr��]��c�8la�E�"O����C�P��1�sa�0��"O�ܠ���\� �;«K@���9%"O�"�f�2_!b�(�`��L�"OJ(�Ū_)1ehh�͕�ޅ+�"O�y{2䀾��]��
+o���"O����ɖ����̕��"X��"O6���`���YQE#;%`�s"Ot %�^	$��YRE�,:b"O��)UD1�kG�j���"Oj�a7�L�W��p����.��y"ON���NM��=
5C�f��xC"OLY	��Eh���2FDL5t�2l�F"OX- G�B����LB�"�܈Zt"O���s$�N`ZH��ּe��=��"O^�W�P�5XD��M��e��u�"O��h��ùm���l
G�ԕ! "O��Q���*$���4L�(V���"O9�*
�>�"��ۣ �"�b�"OLHP&�Q�-~��Q�KN�V���"O�FK'/L� 0T
T�^>�]�';��Cl�k2j�";��U�	�'Rȡ���9P�E�SI��e&��	�'.-[��L�b��4+Ģ^^E̱j	�'jd��޼2u,p9c�S�Oo�xx	�' f�h��*u���˲jP����'�U��)�&-/pH򂔦Q���`�'���:�*ك08��s1��A�vD��'mPyJ����E^��Q�IFh(�X�'"��f�3{���2K3Iw���
�'x�၁CP0K�F�(5�e�
�'"��r#��"My�|�V�� {��٫�'�H��W�Z+8'�峥Țzư"�'z*��Qc�1���һbd��"D�$StǄ�i��P�2a���T�a� D�(�^�
� a`R�F�-"6��� D� ��bǲ���ô��Sd�-z�?D� r�	#xt9���¢r����Q#;D�P�U�#`͈U\?R�X���<D�� `��7�UK�!3w���`����B"O*Tg6N���d�&Bf�6D��&����|@tE�3�Bq+�7D���t	��\P�'�)��yC�5D����i��!v��C�N ��f�1D�0 ��(s�|�X�*L�U��X��=D� )E�_,6L!���1%���n;D�P�a�,q��mq���>b=�1:��<D�ؙ��4|��Zfς�)Α�d�!D�Pc6���O
)����(�� D��K��Dl|�j鍡*V����,D�x������@C
D$̨��6D�܀�($HB�|!0���x'�A� !D��p�*N"vEt����%��A[��8D�����,�%�1ͬu�&�!�C&g���bִkζ] 4*ûC�!�$�� Ğ=PM9��!PW#ÓP�!�I�4nȹ�c�ۍA��(c�#��!��i�DX���f���!ղue!��7F����Zz�lQ�II�Tp!���~�v`��`7B5#��S!�DG�$�0S�N<9
�����	 {�!�^�r�ҩ��N���1rƛ��!�$�S�*���ܵf�:�y �U�!���y�,a&P~В'�O��!�$�
_���$��x13�[�s�!��-"g��q�ŎPjf8��HOX!��B��r$����%�F��r�!�dA�f�ܽ�����`l��!�$�JK���"NE�\��\p�g�N!�D+E��%9�#��2��JtgY�4!�$��EM����R�wPM���	!�d�	����e�>X��\y���8~�!�18����qh�`x��(-^)<�!�$�'��!PwnI�R�Z��$�Q.d�!��"f��X�g�f|�x����&!�_�i|�� ��dV޴���P�!�d	�y�T��dR'y�F �F�	�!�I$���`�$=`Z���+�*�!��&=N�K�%�1l��@K�#a!�d_;[6��{�&�J#*	�lǋVb!�D�.^�T�0��L�y"PS��T!��[�
m�U	��C��HS�J:!���	���фIٝ3��MP�ޔ+!�Ā�;*ͱWmA�w�H�P��>\!� Z�Dq�3eQ�ϔȚs��e\!�$��-���'ه�h@S�/݈v�!�DB�h� Tؓ��.��`�.�2a�!�$ΆPꤘ�@�Ȏ\�.��" �)<�!���H�f��?����� �J�!���<���ƙ J�t��!�
P�!򤋿y�Z|��D�euT�)Ʈ�1
�!�ѭHR*)��V����nʔp�!��<<�FT9���<5�y�w�,<D!�$ܧ<��b������	�f,!�d��]�� ��0n9�mZ�G]�!�$��T�Y
Q 9���Ð�V	V�!�d�b����Ҍ�g�� J<P�!�$5�0LF+y����,��?�!�$tP�2d��tٚUhx�!�d��$}ܘ16�X�FQ�7�S/j�C�I/G�$�e�^Z���"5��
��C�I�fJ���[�t0���6��C�I�?��yG�;]
�W��x#@C�)� >�٣nͻ[�0Q���_'A���"O���*B6�-����weA��"O��y�J��4U^������p<�� 1"O`A��]+!Ϻ�I7��<�Q�"O2����9Z=$��A�g��� "O�b0�4Vyf��B�0l��a"O�@Ғ���Ud�,��L��PQd"O���p�P�E��h�DJ�>ud�m
�"OLQ���Ӯ@�r�
��W�h�"O8�Ƀ	g.��j6�B�B�`R�"Oh��퍓e��8c�KQ���3"O$�ӠGɢG��"n���J$��"O�	y��ڮ���@AB}eNܰ�"Or�8 ף<�`;Q��"=^� "OJPt�p����Jz 4�@"O�����/0O��r��Q�N����"O0$��d+�4,J2�L�v'~<2�"O����0B�l�Ǯ,�\ ��"O��;�FŬ�0�!�S9Oި�"Ov4*5.������Q�g�4��"O��G"Λuq��CWɓ'~��!��"ONe㡪�;#tբ`"�V��[�"O(��,�Rx�a�¢?M�0!ل"O�����"P�F0��kH�2���0�"O�u�o��"�ri��1U�%J�"Ox���K���.[u� �y�d@�A"Oj�-@5r�>�"��*v�R	�"O���(�:*��Z�*��l��Aa�"O�eҁ�H2,"Ш�4Aޙ���;D�`C"�3#�&H���E�RYY0�7D�TǣP!e�X�����a#�+'D���p�V�4���$� v04X�8D�ܙUEE�Z#+̈B\�)(��>o�!�S:t-�9Z��8"Sj[� -�!򤅙:R��4��8���.�C�!����e�Ǣ���X9ǕF]!�dr�.����͈]�"�iu�%D�!�d�%�8� ��Ur"�ʱe�
C�!��֐�R)J�i�:)��Z�!Y�!�^���PP4��#�q	�'d0����,l��x�&*'�A�'R-�6KFx���%��E����'��\p'�]�a��a;o�5?BA�'��0�Ǉ�G�����a�!.�H���'�|�	W̓,'�VX�O��Tp�'���1�/�(i( �C#�] �'�4Xqe�R�B�~��3�l��'Gb��
 (@��� U�,(�2`�
�' $�� �F(��Q��²*����	�'2�1�'��7B�������R�p
�'ξ�ic��J~�dq4�ϑ����	�'���P`���qk��#�	*�4u��'��+c$X);��h�-ӏ�8�!�'w8�J!�K�fњ�ȗᕽN8	�	�'3��� 8>{ʉ1�Ǐ8�b��	�'6|8G�KwP�ɜ' ��Y��'lx3f�H @p��W���8+	�'7J��C�׿ �2d���_8Dd�)��'(�ػ� M�89
��A"��C��@��'5v5�r�
is�<���%>@\���'�\(��)S�+��X� 4Q����'^V�����G$@|9�Kڹ!D�T�'�
x��؂)Ԩ4� $+���'8�\�d��2CF��\�a������� \��f�B��8����΂�Q�"O^�X�H�!;\��@ӊ=֘A�A"O�xp�E\#6����&��7�>D�DxF��;q�x3ag�-
��9�t(3D�h�2K��V~Y�U�؀�޷�$1D�`@��$N���;�M;����,D�`
�@�.x�c�Fɉ�@���o*D�HP�!�s*F�z�n��dvXq���<D�\#Ў[�.3$��2I�b�.-;D��!KE�X��d�]y�#�"D�SEM��
t������Y�ѡf�"D�d���O>MBFy����.'���%k>D�<mޣS;�����
|7�t�S�Re�<y+��4$�e�FB���dh;�M3D�$�.�:vn���Ñ �*�`�.D�t�k/.|<)�V���a,�§� D�@A��:�^��l˟NH����"D�Ġc�~b��x
�N߶-�b�?D�H�́�Q ���@�� ����:D�SRM��Nn�U*�m��<�52B';D�xh�I��eZh�5��+j��@�D4D�L�$�5� bDR�^dy��)D�4)�ᓦ��"�"ԒMyN�b8D�@���xC�tq��U�Km���,D�@g�����uÒ�r?�˲�*D��@!g@2Y����ïD*u��$���&D��t
ػP��%B�	3��P!ԧ>D���G��Sp�d8���%Fiلa=D����*P�87�a���#G�H�ˣA.D�8�׆�>��� R!�,'v�A�*D�\8��=�8���tRV0�Ɗ(D�X�VdT=fԚu�a a� ,��($D��b4�Ȃ
�F�3�ݒE��顫%D�D�VA�Pzޕ(@N5J5�!�ah5D�<�W�M"c4���G�;M�^�I��,D���%Q�4����b��:>��ٷ�&D��!�j�piܼ����(W�(!@G1D�,蔠	�)��!ɇ�C-6hI���5D��ae�V�6 b����Nшw(4D�p9V._<EX�A����$b4���`2D�l�U`�`徭����V|��E*D��g��%�Dq[�g��S��XCф>D��'��H�8��^1�x�Vk:D�h#�M
>�r�!���$Xx}��;D���-��j-<�z�_ q��`A��*D����g�]8ͳ�j�(F�*�1�B&D�P�J�M��xs-��!��"%D������.�V�X0o�<8&���+$D����O&k'�=�B(�Z x�D	$D�h�/�F�����
qP�i:gi'D��ʿ,��*rgS.6�\S�%D�tS���=Ϝ���B��PY�/%D�� ��=8�^a�U�� ]��f�#D�,J���m:|�RdJ��N!J(r��%D��9`�C���HE3�b !D�4��kCԑj��#11X�aF5�I#j�HSj�=Pc�`kBN� aw �!�B����2\$�\Фf��
�R�j�I��%�M>Y�JYi>QH�'J
]�L�l��?�&-*��QE��<?�$)"��1���S�ݠt4|�V��?n��LPB��l���L9�ZQ%�"|z@�K�NZ�(6��
�������<�%ϲ`�h���KJ��qP�c�O���h�ŤP�VUB�O׽A�����4Lإ��'�v���'���(F�(��|B�I+�����w��I{�G��t������X(am��p�}���:9V�����}z�[`	�4�6��sE� }.�L�	?��9I#Oc>	��M�s���A-)3&(Vg���JX;qk�8К"C����'9"~z�g�? YEKѢ�B��M�b��	I���X��(O�O��)�ǀ׷t5��!w5&��O<aF�#�S�'6��A�%̈́3p�<U1Pd= �jt�''��Gy��� M��[�k�O=r��$��ԛ��7��<�}篑�j������BZp���KĎ��|����џ@	�J�?D�j�·J<���ħ<X�31( �u'&a��ʕ��v�p��� �DR:�^M��N�O=Z�ې��?^��\#�锂.zZ\�qoJJ�k?�IA	�':D�����5YU����mי �豆ȓ"H.,����K3J\-aB�d���2=���Ώ!�Dd�!
�jp=�ȓ̎)r-��=��Cb���[V����oq0-rViL��DN� J��B�	��T����f�t
s��@��"?Ɉ����p��p�%H�EQ���4F�X!�J��`�X��ͭy<�$p��%�!�ǥO�`(�Q+�-A�h֊��$N!�ď$m̩3��è?����X�KC!�$	��H��fE0E�)�a�C>C!�$I�hD�
�o�$I�a��ްq)!���m�mcE$M�j �Ig^@!򄓵R�|�B7AٷJ�$tzD��?u�!�%A?LKr�� :H�<¦�."�!�D��0�2t(�Q�^B����Y�G�!�d1M M�u��m�J��%�,�!�E�%w:�[�[
뒤�W�T�e�!�Ď�n�lQ�'ID6T�,�!�Ȋs�!�$�
�\��ܩA����Y�!�$H�b{j�*E+�&!�A`ڪ�!��� ]���I!� X�!�߃U�!�8�]Ӗ@�&v�( ���ԗG�!�$�,iE�Dpf@ݘyb���
�!�$[�? I�PfÎ�~)��B�-�!��/!�Q��Fؐ��C��Ts!��^��v���D�K!`��$\Z!�1����V��#4	�=���)2�!��ާ��S4�Oe^5b�ډ
�!��P,v����H"7��q1Ѐ�L�!�dK0�QV��5�jɷa�Gs!�i�VA��mU'z� ���!^�2i!�dS�(	�-�C �cŞE9���f!򤛷�f��%+��i0�ƁY=!�ř9T`��Ğ�G�聛d`-</!��K vE6I��&T�QӪ�!�سPˡ�䂢��12��k&��C��y���=I�"�k��R��NX�&lф�yR�  
H�9V�C��>��� ���y��������<�n�� ���y�N�Q/��y��8N���TNG"�y�\�Va�$��&��)�HJ��yB-�v��H ��ϘpN��'L4�y҉�� ���A�y�jU��dД�yh�&s�������8C�mc�`�;�y��=�l�����m�(���K�y_(W�z����-j^p���I��y%ż8�����gU%g�l ����yB�˝`��[em�vWȵDGK�y�#H����ě�|�4�brL�%�y2�R�?�����mƉ��`M�y�\->���JaPr���Gթ�y�oR�$�XwG�m)Z�	F��yֱ҆H�6�+�Iە16	r���y��U�_7T�`e�� ����"�-�yr"��%�hB0��.n���t,-�yr!E�rS�T)�oɅa`z�� X��y
� ��Ju ճi>|�%K�9!F\17"O򽘕	Li�iH�gň,bR�"O�����=HH9�&��D�p���"O�0"� �)أ��F�!"Ob��2�\[�\���_N|̠�"O��q �rn s��Z+NVQ��"Of�sb�P|��:�⃾k��
�"O^hHa�W67�P��W�[�fS&Q"O� 2�c�!<%���û?�<�U"O�d��mD� )��P��G*�"O6թq��;��`S���)}"�)r"OI�TL�lL( ��J&W��S#"O
��ƤUnP`�����\��8"�"Oj�Kf��l�R���ύG�r���*O��0q" ;j�"�b`˜TŢ���'���R���
4˴�p���^ۦ�9�'�^U����)�؈z�l�U P��
�'6��ϟ8=�	Z�e�|�t��
�'����$)�2�z�����,� e�	�'����P���|u�(di�	�'����jZ�g�8�S�̿��y�'�@p��r�v`h��X�Mv��'R�� _7�|=S�ϟ��F��'x��5'2g��J�BT�)��Z�'`��ǌ�X9xA�L��n�r��	�'�)��e��<憐�7(O3��ܢ	�'���UmST�!�"U�2�d̚	�'�>�f���e�h��v�6�		�'���1�S
y���Ï^�s��k�'S���CMͯH}���HA1dv~��'�d�@�l��WK"ɹ��O�`vb�'z ���74r�"�o^6�s�'a�����Mi:����լ`î���'g�Ճ��>#�j0F�B��I2�'��}�:��L"J��Z&�܃WW!��X�ȝ+���w* ���ޛF�!򄀧l�~��߀@�y80��/G�!�"e3B�З.�?RM>ٺwa�4P^!�T�)��8�`�-I4|(d�ͷ�!�D�7J������J=.-�ABH&�!��l`*lp'��(G�������P�!�$A�\���:KY97@��Q���!�D�"M(�@��胎-���/\��!�΂P�@����#��ӭ
�!��;�����X��:��0� �}�!�݁�Jh��#	��x���~�!���yF��@5��<��ۧC@�[\!�$a�`���D)  �9	7@ʛq!��F��z�F�x�뢎�%V!�DE�%�X��s!����j�*t��"O����'�s4pA�B`��M�Q�v"ODxz�.BK�N4�Vn9)�"�C�"ONܙ
M�[~��؂�� +6���"O�8ۅ4B���K�#艊�"O���3fY'P��,��X�4 �P�"O䘢 o m����g� �i"OMٖ(�wt~�s��LM�$ہ"O�UXB�)� XKW�4Q�P1j�"O�a��"��z&|A���ʻG���"O�Z�&��U�ĵ��G�<� ]� "O�	o	3L���ƶ���AG"O(�Y�E�\O]��f^�]���"O>�`$MN�g'�H�!%f[��]�"O�Yʑ�β�$8zw
y�N��"O� ��R��8(�0ɦ���JwЩ��"O`�y��H�9�z��oP�G�n�
!"O4�!勆�*밑��N��{�Z��"O��;u���$)@e���}H"Oƍ2��N:>���#c�����pt"O9��$]-�\���4o "O�[�)��z#L4�䀀�Qh�!�"O�[�Q�s�1`��!��%�"O�=�r/�$,�n��훃z�ؼ��"O�0�+K!0��|	%�)(��!p"O�="t�J��}�1���&OtH��"Oh��c�#S�
���c֟o6�5�"O�����p3��	���yNՉ�"O��T�)c�1a#�Lܑ"O���I�Z��m�&E�o��]�'"O�hf/�=TأBIM�O�$�""O�\��⓴#�����'�)"�"O�A��
�X�vǜ��\�6"O h�� ��H�aWH^���y!"Ol�˔�H�3�t"6A$plbu��"O��R�9JP�	db��yU"O��">*r���%ƌ&Hj�b"O.q�sF�KD4�вD�n0�h��"O�x�!ë@}��e��\��q��"O���Sa�3wdm�F��1��6"O���A~�Jr$�ף/�J���"O�A�ɐ�"Ȏ	� G��y���"O�קۍg��E2���#|�H�"OZ�kS)���R���aBƨ�%"O�Q�W�À�:$NF.;��!�"O��B�F&} �JV�ض[:v�r�"Od�J�C�D� �ڥ��8�(��"O���2<�|����M%����"OR�C����A�%�TW��q"OESDK֟_�4����VJ��(��"O.�3�Ԕ^���Ru��)d.
!�"O �Cը�`Z��C��V&�)�`"Op@Q3A@�v�5�]�Bk�:�'l��D�O4F݃ f�,�h���'{T����� ��,�B#�)@���'���� ���VCJ-)�����'5��{�#�)c�#�,��1�h�:�'%@����_�9�x
[%-`Q��'-*�4n� �.�3��M3��MQ�')� #夗�i�d���L�|^�j�'&���-ƇA�(��ŏy�PX�'B�|�� dMp�����wb0%"
�'�ȁr���w&����,2<q��H�'���WݮI�p]�P�]�94	@�'?�l��mJ����``G�8W\�'/����(C!�4�8���t��',���D �C"6AzĲ
��%��'���0�l%C���q���I�',`-x3G�4$����Q@5h����'qĠ�TL�	r�TjRG،]����	�'~�2�`$��H"�_�ִ0	�'���z�Ǭoe��;���1�+�G�<��<���C�6��#�@]�<Q�&S4<�@Wl���0��\�<y'O9��K��>8��T�QoDW�<	��4~�|�1����]$(h:pg\�<�"`�-<Tu2�ؔ&�fJ��T�<�� ��f���#�G��r���J�<��*	�?�y��P�k�pe�JV|�<� 25��h0k��#���70ƺ��q"Ob�Ɩ��՘���i�T8��"O*|��h�8���Z(.j)�!"OJ����]=W��� <i.�j�"OT�1"�HPp�1��J p� �e"Op|ɐ�I_J���Ӎ>,��ڀ"O��1��<&�@iR�B���!���`>.}[@�7X��K4!�%J�!�W:�D16�V�rH�c�N$T]!��D8���(w�3S�()�.;{!�$Yv۸�S��O"��S�lE�JY!�d7;Ú`���'v���q�M�.�!��]��Rƽ�����.Y, !"OީjaǤt*x��/I�Z���"O��뒤 �}c|��b���+ۖ8�"O�Ԋw�\qKp�qlFe�~)rW"O0e��ˋ1E���������"Ox����{��H3uKW�QwX]"O�ܑ��φZ��]j0+�!*b�t�p"O4�d;�
e�"햼IL�+�"O�T�CϏv 0jVL��X�$�1�	ş���E��F�i z[�M�c�/����6�T��qOl��u�� �CK(���)@Z-q�p1i��N'ת���L�
?.aCj޿nࠌi��I1��m3���3Y��ЌS�n�D@�-T�`�����$a��x%ASe|(A0�剄Sx*�$��MI�4�?ᬟ������=_�:�*�O�!V -��ƚǟ �?�O��Oƴ	q��!�"�c�
g� ���'�Z6�զ�mڳ%��X�DkFP�AGIe	����k�dS��Οh���`m�pO��#��Ѫ0�x6�W�z����X;T��1��]�e��Q�jPfZ��7������_�!�F� �v=���iJ6-I�ĞA�u�7p" !���Ĕ{`	�T���"�
l �@V.`=�\{ҥ���Ca�Oz�m��M��䈟���џ���E�� )Ν	O�~2�'U��Z���ɗ~��Q����s:����*FhQ�\��4f�6�|b��"\wlĨǋiR`A��Ur�4�0!�<!P��Xe�&�'BT�pgU�B����1�@-S���A�ɑ��B�m�:`�pSV��&BV�I�2s�N,���|��v"ą*"��3�,{��+$<$"�&�`a��(eX-[��ؑ�&B̓+�6%�� ��d�ө �U
���'�8x��0�&�:��O��ķ>�%匱�hmc C���y�f�
E���3'�?�$�t���{���+ �^�h1��
C�"�g�d�mh�	�?���{y��Pj6�}�"�J@zR�IևK�(�h�S/��y��')���_��bT)�I=E�Y!Ӭع,g^x���BZL ⇇��T%�2�H��(Ox�B���{5���HΓJ٠�`��@3Lx@��D<
����*i����4�HOH�AC�')� ��I�BГ��ܘ2j@�i�H�8RQ�6��O�ʓ�?+O�b?�j�l[4|I���ՠ兏Bs�B��?	����i+Z��h��IРD���I	�MD�i�剞d�40۴�?�I|"���6x���Μ��ա��R��?���ML>��P��+w�aG�([�L�Yt�.Ba�Sj
%�v��@B&Rp5Ey2B�.��0l8$�6T�bL&Bڡx!�\��!\�B��C"J*j�����鉽.]�����xK|��4c�(z��	R�H\pE���Z�2��'�O?��KwR �#�l�1q�p��`���E��|��f�T$n��A3�lҐ.h�����66L�h�δ��+�ٞ�M���4����-�dN�@� ��R�я`�)(׮�<�� ���&6�uoa���@ܥ�@`�6�����	O�"�˓�5 D���@���M�3o\�J�]��m��l)1AS�+���]G��+�*X��SV���`�A�ܦ�b��O*�nZ������?7��'8�&���XS�Z+�g�6n�~r��`I0랸!ob�����>61�(S7.(ʓ
��ևrӐ�?!��u�pDA�(�	�0���Xg�|��'KTP�� ���   �  �    �  �*  �2  |=  �C  J  �P  �V  ]  Lc  �i  �o  v  V|  ��  ݈   �  b�  ��  �  '�  ��  �  G�  Z�  *�  l�  ��  ��  ��  ��  ��  �  �   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d�O�=�:j_�[����q��Z�|Ӂ��H�<� ���.�:�$Β,�^���\D�<�$��
c�
�sa
��A
#nC����<)��7Q�D�u$8]h�����P}�<���� U��\+ OT�%2��ŋu�<���^ʤ��H�K��U��ASr�<�7.D�(�3��5o��Ձs�I�'�ax��ӊU�$c�H��xF���"��y�Ì�I�4 #1m%��u�������0>i�/.f��4�s��4D��`	�x���'��p;E,PS�U�B��D��<�'��8�I�)NX��a��u��y�`
�&F���4'�ZpbeaX,�y� ��"�f���S�iJ����y����h`h�v�L����D1�B�ȓt�V}*vL�TD@i̯t$h�q��~�	�:zxnt125��1�y� Y`)�щ�nl�5��ޗ�O���4H�Z�F��O$B�jv^��!�d�O2�HWJ�*9]x�ꁷ����@��y/�'(c�,����:�.��r-��yr�ǲl����"6$<z@�%�y"H�I�����V�����?���hOq�XX��g
-Ph@�ݱX&"\#W"OLl;�`B�dxh�o�1^#���i�����H�S�A�4�ę�#� �aL��I���� ���2���,�tlV��s1"O^�`�퐰l��H(2"�|S�"q�'�H#=E��-�>G] }ض�^"DZ0XR���!�$	 k���4��~]&u���y�e���Z�F�:&Q�sȓ���`�(.D�h���G2� %k0iΈX���6�7�Y�ayb�QI(���*پ#�\p������hOq��l���H2����,NRZ,(d"Or�i�P��r�ʣk��
S�D�Ӧ��D-�bO�J����S#��P���D/1XZTi�x��M�rX�'Ka|�m�(f�m�H�?�P���E�y"
BQ����-�gj5��(���0>!��9E���)]�M�ҙ���t�<Ic���X(LȆ�J���v��n�<�-E
Cl �X ,��%k�uې�q�'2����O�R�1w�>'�~A+��U�ghz��1%2D�,��%�.E���*�=t��!˴���'�F=O~��h�'D(�@��nY�	�eB�.�BB剕m��H�a	Nac(-�2f�1Z�,ʓIe���ͮ}�D@8�,�#M�j�!PiGb�����j�'v������Ï�9��`��`O"R�
˓�0?gH��NPr`Ƒ��0"V��\}B�'ӛ�W��E{�'k�m(����`�(TnX�>le��I�<�emaӼ\�'J)q�>��qbR�>+�Q"O��3FA=��)�s�	%6��x��I?�XD�ԩ2S������
[���v)����0>��1V��U�z�u�v2��O�7M<�&
�&X��$/6� ��w���e��� wȞ5��x"F-}����h�1�S�̐��ē�~�b�r~2�=��'�Iٓ%^N*V!�NC�%	�|��'�<I!��Q���%���ی{B�)�I���mIb�~fp��B��i�!��C�2���b7�̦T
\T�qL]K��<�c_i�"����q�s^�$���ȓ��́F��v	hiڱ����n�s(<)�@�1P߬9�5�ыe{ح�ʗc̓�ў����c�a��L��`A"h9�"O؁�7�\��i�b-���"O��@�ܿ_LhK�!��f+@�Y�"O|�K�r.PlΛY�0�s��'�y�C�Sn����� 	���CW	�y"���,�<��4p~���Nм�y"g(g��|2�AObA�AC5^-�yBb�"��L��ȂP������
��yrNٕ h@d����*N1R<b# T��y�ߧW�b���G^�HI�)$$�y�X�A���р�8E�-��L�y�bL�GG��H���B�d<�q����y��T+@����b�Q�(���y�ḽ3�|��t�ĚL#�(E�P��yB�R���C�́)/t��dM>�y"��,���`�����=����y�({Ɇq`�g�'����K��yGֲ4��=�EB��%|�U�q�P3�y��U�yW&�3�Y����O��y" m��eh���~���LY��yr��yf��:c���4����'�y�[�+T�8��K9�*U ��_��yB�V2�8|�҃�Ho@���jJ2�yN�h^��z�o�=�:	X�˅8�y���4KǮa!�돾-މ;��W5�y�� 0��2��Z�)�&tR�]<�y��
�e�������(4������	�y
� �4+�
��T�p�b �X�?3���"O��!ҥ;MN<\`�Œ�zJ��h�"O�5㱫�|l��!��)M��R�"O�i���7���TC	.�hl��"Ot���۶4<C��(�m�*O2�1d�F\X9�Ǥ�po~lK�'�^�#U�B�R)����t6���'� �I�kJ	Nr�a�M�]���[�'�R�VL�'ᐡZ��Ԑ]����	�'#���h=�m 6�5P��'y~�rPـ�BX���y�����'�|!�ȑ�Y���νb�X���'��I�%�^-:%��H1P���j�'xՁ�`���Z���O�C)�'�&3!�G ���YQE	P�(�2�'�*칣�b�4y(���V��Ś�'B��c� 9�h�#�N/Pu���'���p��4M�ZLi��U1L/��z	�'�e�s�� cap�R`BL�)�'�\0`��(mB�Y���F6�X�'8�(����;�\I���>,���k�'Jb4����r2FX�*�e��'`�0P#�L
t_⌰��,%+����'D����V�&��4$��&P�l�'�N18��A���A�B=���	�'پ���퐴C4�!�cgK�4���'�8l Å� �l����^E��'��0�.^7?_��k��֟{ᾡ��'�V��tD�_^&]Kq�K�l�����'�$|�&c�������ת]h20��'��)qiBQ���k��R�X�DXS�'��aA�Pq���S�yZ�'���I�].t)��p�N#�^���'8���Mˇ}�l=B ��&�xx�'���F�N�\�5��������
�'����Vi JJ��BF(\����'ݪED�rɖZ��I:|A���'=��i�ƕW70���#w�"���'H�Z�@�m-@y�Z�%�J<k
�' ��� /zZqp�+]�q5��j�'�X�re��c:	�r��q�� ��':�ЇeԊe�x�b�S��c�''�ᠤ�ǣ�vX2ѯ?Wv�[�'ڹ!tO�+��!;c"�0U�j���'��̊�oα\�؁�"��Jk(��'���� �YKt����G����'�6���Ş?�h�8a�[�3�\P	
�'�Π���S���b0��!{8��	�'���,=b���)\�נ�	�'^���G�I�/�:��g��H}�l��'� [d�R
9i�����܍T@<( 
�'�a!�ە3q�0(pLz �J	�'8�H��E�v-±�nY�H�<��'�`|)�	�D�N8�ש��A�����'`���uPx��ȒP�B�+�'�nH���q$|�c��7(��'�2�K0
���*����w��d �'1��ҕCK�Nor�C� ��Y�Q��'�F}z�>��y���*S1�#�'E�Yi�8>p �R Q5~\�Ԓ�'N-�r�U�7g�`��]�I�~��'�����b�~���A
@���h�'Vy"O&�hQ�ᆗ%*Uf�k�'<�|&.��h��h�p���.�|T���� .�U(
�7�l�+�K8Gj-� "O2L�Wt`��l��6���"OL�"䇸#�b�Z�+ƕR�L(��"OH�d�O�"!	�
��|i�I�"O�<H�IAc��i�C(Z�^Y���a�'���'���'V�'�2�'c�'���c#mʊ ���h��!MlE:��'���'�2�'���'���'T��'�H	B-Ȅ��KZ�B/�����'���'��'�"�'���'��'����+/!$�٘4�	�� �'�"�'���'���'*B�'��'�<8$U��q����+T�ܥc2�'#��'x��'���'���'���'!Ti�`�;YjDi�'S�	�0�'O��'gr�'���'$��'���'A��Z�RSV-�̓d�Vш��'0��'`r�'�R�''��'�b�'>��S�;H�j�( J�"4�'
��'��'���'��'��'*w�-N��Ã��
u/N��P�'�2�'���'���'���'%��'�:��	r'�y��[9."d��'���'���'�b�'1r�'$�'�L1�P�Q�n��dX��VI�t5c�'2�'$r�'���'���'���'��2o�>��K��� �0,{��'�R�'%��'���'��'�r�'��������OW���l\��줡�'��'��'�"�'��G|�j��O��bB��E�ĸ!5.J��H�3�&�oy��'��)�3?ag�i����e�s��"hE��9�*�����ͦ��?�g?��4pC���6R_P0�� ݼ��'�i�"�ݛ���h����-.2�y��~��aB�*�[���&	8�I�r��?	+Oh�}��	�j��}�e �4�&UawC�S��F�����'�񟠭lzޥʡ&@8Cؒ�R��
+S�� @*�?9ܴ�yBZ���jM�B�vӸ�	�$Z��IdHv�Kw�&Y��I�DT���M�v�`hF{�O�B�\
B�F� �&	�3޼5y�I���yr\�|'�TJ�4,Ih��<)Į�)����!E#��cb�&��'Htʓ�?�ش�y�S��4O�2Z���m�{1nm��-;?I� v�^�r5�]a̧\�R�S]w�@��	;�>��fR�yOv!�PO�.0w����d�O?�		D���T8F�1��Jܽ=��I�M��hu~��r�(��ӵxoН���[�\`r�m�h����П�nZ��"�G٦��'��9`Q�ڱ��qA��#�bx�ℝ�	;ʄ9,��9�p�C�o�+!�e��F]Z��L>��F�z�|��L>j�Z�Z6.�W�<�VjU�{P�����
L�w�ͨo�@����R�\���!£u���Z��V"krX1��L�� Z����Ȧs�0uJR
!z�X��O l�Sgɸ)X������X�P� A�65i���7)"D8*tJ*,<���e̶( C�TaȂ	� �B�I�T Z4�Y�N����%K��0,�	&j��U������	�?m �O6�F�a��p4*A�KW.4� �i���'NAXf�'ɧ�OwTPb����b�` ;T��
$0�(�۴F��`�i���'L�O�O���@�̴�~�\=y�)Ӑwв`m�9%��X�Ik�)§�?�Ң�:nJ�٤�O�N���yeI PM�V�'���'K�yp��)��OT���x��꘍��q�u�����W6{3���|�j�I�f�f���O���ձ;��A1S��4�
�.�f���l��0��E����D�O����O�Ok�
h�r|!3��7=�x��S����'�d���'d�'���'MRV�)�w��ǃ�6xaP�l�0|n���d�%�M���?a���?1,O.���O��$�3B�nrO�t-J���d�b�X{q��O��$�O��O4˧�?��վU՛�РM�L�׹��b�eV4�q�q�i#2�'��W�p���0��'dX��I7S���G���<���xc�{�Pmjܴ�?!��?Y��?a��NG�];Ɣ������.��vl�&JP���Lv��7M�O��O�d�O�5��)�O��'U��R�X�Fuqfhϥj���H�4�?����䖿v��%>Q���?�R��Q.��=�4�nUh�뵋Ԣ�ē�?���8�A����S�TiXq�����K�.0 )5���M�)O ��`��1J����������'����-R�>��PD�H�"e�ش�?���EA����S��(�T�(0��� ��%��l%�4<�4�?���?�������)@�,��]�#��+��,�E�f*lZ
Y�q��ٟ������O��'߮qPB��+�zIy����3�D{��~�"�d�OL�d��O�&�oğ�O*2�O&	�Al�``� /R.�,��i�r�'�a�$���?����?��O�r9�f��/u�^�A%5%��x �4�?��a(<>��ǟ<��ܟ�%��X�)IX�r�Bԍo�@\�T�E�v6-�O��C,�O����O��$�Ob�D�ON��X�2�414��� �f4�  t�l���S�Iş�����'b�'���hp�.g����Ñx3pɃ�	�^���I쟌�'bcפ��)�K��=���W0�HLA0�\�4���'����OL���:���3.���QRH�uI�	,��O��d�<����ă*�R�dB���;��GZ���i���4.��=m�q��?�@ �-�<1V�S�Zd �:C���sv��+.0��'K�	ş`��m���'���5����.�~p���#���u��9���?��#L�!�N>�O?� �-�uM5gQ L(�bX�{팸RFY�<�I�O��!�	����I��SryZw(r�Ҧ����X�
^�m1b�"�4�?q�!(�<Y�� �@�Vջ��#<4y#��b��V(�>}���'>R�'��4]��'@�B�cp�M�!����E/�8���ɱ�i��ɑ$�|�c!ҧ�?�pf�1�]��P� Ң�Q'8����'p2�'�|���?�4���D�O:� �>�,0�Nٳ@;(|��%M��5��ş,�I�|����.ʧ�?��'�j�S��U��a���w�.Upߴ�?��a\����{�T��GK��D	��_�+�\9`��Bd��o�۟���:�I۟�	ΟD�'�`����*;uk:Ԣ�2�%�<JO����O*��<����?a2�Ҙ-�r�Q�U!BT <
��M�IN������K6���x��%�ʓ��4&\f��D��̬#�O9�B�	�M����b��-�̔cT%ڌv����2F�[\�L��ϔE`v-9E�& �H�[d�!Wڴ��e ���"]��!I'
h� �Ǟ�Uhx�0�рa�4aKz����6��yu&Fr�$A���azl���;5P��{E��
�۔$�4�ؓ��N:\,�C�� u:�8�$��6TT2�a�<t�8t��O��ړ�8uT�ֆ��2[$�	qi�O��dW�\�+�aM���a��U Bpt���O�S�u�\���Q�#/ֈ�EA	;i5�'�0(B��V�����ќRP�S������O�B�b2�ؾn�pت�n���m�N��U��O�doZ��M�����OT����#:5�H#c"�(7LM���|��'r�'9�	Ο|�i�EjAh�u� ؇��db�;Z �������ߴ�?���i��a
D�<�j��ߧFnX�@OC( �6-�O(��OjiE�$#��D�O���O��0X���{B�7u�a�&Y�(n�����է@�����B�w����%��Ϧ�*��i�h#LA�ONܙI�Ɵ�Eh�(��Y-q����P.峵 AOS�>aoZ�{<��I4�N���Ei{�}aChߙ�$��4<��ɚC���4�j��)�	��+�#	�&��� NH�M*�B�	���%�s!O�`�`��(��i��k>����޴�?�.O�0	���:���i�N(x�*���_�Ƚ����OL�d�O�����c��?�O����
�3!�|" Ȓ9 O(S�h� O��0
cE˼0��!*ÃL.U��#?Yw \5H7�r��l�dT{�CY�F��łtᖻ,��u�,NTr�w�ɥ	��h�1�&Qr��3c^�vҮ�0d�O����NM�Pݨ�\Z�����:)!�)�����mт\�r��p/,r�1O�d�>aʒ? ��'�b��y��Y�7�?W�h͙2�ѥTT��'��I��'NB�'� �*X0j��]�b��mZ�7-�*-��T�ߋ]���ش��x����H�1�4Ô�W�N K�Γ5�TH%Ɔ)@�.	��G�Nr��G�e�PGyb�
5�?ᐷi�6��O��e�:������(_����'�<IW�i��Ib�T��Z�AZ���*� ��M����V��Ӱ�p-��i�(z6�W�f�ʰ��O�������MKQi�>mt����?���:�*�?���N�\&�Yҵ���un���Β�?��U���{�fW�{�"���	���M��~�,��:��J�3~�3�62	<�a�>����8m
��c��k�Z�l�o��nެg�� �c��W<�ȓ��]�<0�'�ph���z<ɧ�O	��qGY�3�8���ڡ!�T���'`�}@#e�	t �Qo�$�!�i>�"��@F������ʐ(C0�_rmZ՟��	ߟ��	.ir�|����������݀Z��8���^� �Se<�М���ZDD�oڟqNzx�v���'A"�'� i:]�����Oȥ�@At���f��j�故�M����������i�$IМ'���r$*�,j�ݰ!����i'.y�P!�'�������͟"�'��	��� i�����y��H�g����˒X�.�Y�^6RΨ{�ND>5����O��'#�)2����A
\��(*�hY4!� �D$;\���ɏ'���D�O��d�O�,���?����t�N?P
&�BՄ��l�0���Wtr�"���u��4ɴ�	L���"Dm�zں�-�B��g�O4q��d+&LO	s~�CS�г"���W	ڰg*�ȡ�'���!��;7&i�6Yâc���yb��	�@t0RAW�
R���d����'�Hc�t�ƪ�M3��?iC�S+6�t��&�)CN%Ӥ��"�?��������?��O���2�K\?����8ӛ6�,�v�+��U����%�p<Q��	'2��
ac�9#��M��40��pn�P����A9�a��	�<3B�d�O��a��z��^�U>B����O/ET|x��?��������̉�o�R>�Ċ`]+M�\m0�O1nں < p�ΐ9u�*�AүV���Yy��
�E�X7��O���|�@\<�?�D��,-f�����IV�ArR��?��eRZ�;�Ð�7d���g�Τ6|HX&W?=�O�Fm��'M�b�b���K@0>E��J��S0KӐYTp�s"��&l蕪Ww�'chH(�eMFȘ`�C1f��O�1C�'�"6MZ[�C��{����v��t浨S�V*Tvc����I��T�S�? >뇧[�T�������=��dۆ�'�<7�ʦ�%��Z�$G�dJ2�\�0�,��΄=�M���?i��&���a�.��?y���?��Ӽ�ŏ'h%���.��=��U���S�V���pᢌ�mT��	H~�<�&�ɧL̠P�f��]l�`4�]�p���NG=^��%�B���}B,ʸX f�	0%�����j��U̮�r���:j[H!������v`����?I��C*b�U=��9uD7qu���}�O�R���4{
��A�}oh�ӛ�|�4_�v�|ʟʓ]��J�c�\�:�
�=�
��@
���p��?!��?�պ��d�O��C�Q<YBD�w�]K ��`��d�l�%rdN)x	��3�2��˓m��R���F�*a;�^�B���� �W0%aa�w>:J5'�'K�B�@3T� �pn�,��5��nת�?q��
����'������?9d蝌��lSb`� �?��?)	ߓ{�A{�E�I�LU��UV
E�O>�Q�i��6��<���U�6����'������m���'N��bPl�t�b�'���"�'���'��s���cUk�k�%C�7�L5�Z\H%a¯P:� a��Z6S��x�Y;��qA�{��պP�O�0���`B�F�@��,E����퍴ȈOHb��'-J7����I�z�0d)r# �2mS^,�|�'\@6�1�	��O_��A�ޞ,&�P�ϊ*C���
�'�x7�O�}A��*�FS;�JP��T� W"n�z�	�@��[�'�@EXf[�f%����rUk�'].�q�肊_)'*��K���yB�BJ���������� ��yB�A�4@^��D�� by�� �y���GD�Ʌ�P;]䁓g�H��y�%�R����bӴ,
i�iCf�<�ʶ?��x� B� �ݳ�Nb�<��JT�t7B�	U���J��!u��a�<�$��h�)�&&a����LC�<��%	�`�dܡ���?,��0�|�<�UE�M_z�B��0W�  �DL�<��ʕ������J/ �9����F�<iD�ؖ&%:����ձ6N¤�%�F�<q�#čc@mH��_�B0����k�<f� � #�*:=��T��y"b�>XNz5�C!_.����p����yR`�##J�����<=Z<990g �y��Հ[,lI���3#�V�Q��L�y�`$�,��4�F��
�����y2��l�h�
�2z��N�y���,��3�A�\��d��y"/�Eʀy�
��Ѡ�[�N�"�y���v<���A��2}ĴAi�ٖ�y�c�od���c�"o��X�1��y��\�&r�(�S���B��y����	�H`R��чL?Ԝ{�o���yF�d�D����$DB�CCJ�'�yr�ڤ��E�g �9{�oϕ�y�g	�5�ba��O�]�^�u�P"�yR/R ��8����`Φ�*�ۄ�y�-ف����V��D�8q����y�*�%s�❓�hZ1m���;Dh�1��'�� ��4y,�9� |l�4�F�N5a*�ͻ��O�(!6B�	�R~�bqE�)�B��֪��2Q+��G
V�$����O�����3?1��³V��qb�6��Ъ�E�D�<�B�u���v�|e$ #��hT ��U��>-G(=�SN2\O����!��9�lJ3>��t�v�'V�k2�	?7�H��h��fr�{V���
�)s+ٰi�<d8
�'�\hx�'ַvۖd�AA��_�6���yBI��6��@���W�b|E������R�Ý����� ��y�- &� L�7obE�f*c[ 2e
��O@�}�pPE��O*�����V!���"���hI'"O����n8B/r\�w?l�|J����?o��!�*ץ<�p��
��~塤j�!�K��X�lY
�鉰@Ҥ�w�A�l�����#�&oN,�P���3��у�(��Z׺C�)� ��!��,&b��d���1wƴjV󄜇q�ƵhR�	;��Î�)áx��(�q���?�v��R ׅ?!�DA>z���q��ˡ�EIE�S���,�\!�v����
tO,�g~��LKaSC�,(�J}����y(� l 0�ڒ�[=�����4��Èmh��k>lO��84F�e�l2#�J.����'�r��DHE?�ME(1�nԳ��\t�ҁ� �Mu�<� ��Ci�萄/ͅ?����l�'�p��	�W�g?��,�Cېي�ύ�6��Q	ȞM���3�Ov��N<&�ܭ燊�~�P �Aca$�a�����c�Q��yg@�6�I��@ܧ1�:��շ�y�i�1/FE(��L,ʠ0l�	��lJ�2T�T��s�q��|��dU>;>d@h�͟�i��D9$�'~Lqb.�A?��Gڇ�^pq����#��E�������'S��UH!ϣ^��3�+�2��ɉ�?�l���"ފa���'��!���F�iaf�5������<��bK�E8 |��GR9cY���D��P���X��'$�1�D��"��"��A��2DJ#]�4��A �<)�����Tl�i�AB�D�k��,"�k�5��%z�0�O� ��֩�Nت$FI�zp��������vAi�㔭��Ħ�T��u��SV�<f�> c".�<�`�/�V-�T��&F�6���&�e�'�y��b�461���%v�,Aܴ���� �:�x��퉤.�j����/���3	�>�h7�ɸG���	�R��DU%S�Q�t�bt�#J��j�� �k̃*d􅔧�s�l�WmV1b(B�Ǻ��L��V�1Uf����r�=�%��a
��"2�K%�ܰ�$�"ތ�'P����D�A��	�<�$c�`R�-<ՠ�`
�H���#4�{ŁD,ty*􆜸Z�;C��W�H�ÆH'��K}��;2bj��P,	n�$��<�Dh፞�l�x%J���&Z���[�-R+/t�d��#A�]D1Ӗ�d��Ӓ/�?�H���$�T�"�0ěx��Y,h�$Eze�ǽ5���ORH�'�`hc�ƀ�L����fK׾0�*	�,O2D�sË{�� D�XZ�3��O��>ɀ��Wk�hZt�ם�
�ZQA\�<q�n����DƪJ"2eBem4�k�$l����؍�a,t?�p��C�Lϊ��C�͸A��@�Ǻ'�d��<���Ы.=dO�.rrĹ�E��j{����O �p>)�.�~o�	�%N&�^aȀ��ay�C�:x�ÒSf�
�z���<;l���4GR��ܘ��ƈ
%>���d��,�<�3#!�1U�|��c��0x~A��KS+sEN�+�E.\��'�
�SU��0|��` ��hPxhha��	5%�	���6"����<�"����-u��h�`�l���&r���Vo��V ���'��i:�}r��J�5ruk8:�-1gF��WN0�F%M7���"����v��
�ўP���ۂ_L|�r��ɁW,j�y�C���C/ax�G �*>��A�Í5�@���e͌JC��?{t��[u�l�'��ͪ0�^� a`��C��<8�r���"���K�.A2A,"?�����Ŗ��W�VUI�fi>\
 ��B�rƝ{Ć�`j����$��-C.- �ۦKI6�s�;.\�'�j�	��1�^Y4�+s
��z�O��#�lw�� Z�JVtB��5�b� saF�o��䈘^/���*�*f�=��B�鎉���?!��`b(�#!(*����4B���ئ��K2i�0]�+A3d�H��eJ �:%���%?p�5D{�e	5#ш"��#O	 �� Ɋ
dܖ�O ����*�(�����f8"��IK~(�a�yB!�`�B_ճ���"1��њ#�1"��8ò
$IȪ ��+T��&Л�@l��A�����TtI_�K2�_������
�Lm�pۮi�D�"��'��S�@�+@�*�0U O�%��l�J<y2��)@&�)��R�{�I
RӤ ���6ϦAӅ��6/���aZ�c4u� ��s#fm�!��d5NCK28�33������<5z��ʘ�A��S ��C���!U����0?���[oƑ���Za�p�TN�~Yp���n�zH�I%���<	��GyR�˩Y`BIa��[\l����ȵ��?�r���3�|H �z��ju���'�Hy{�Lʗ1 1�C&NJy����I�[��<�AR�DCFq�H�k�Ԥ��'��@�1C
N���I�MC���)$a��+����|�!548��@N� ��AS,*�џ�J�b�'v�J��0��@���C�m�>�SBŦ	���H�|`+O�V[ᗀ��� �	RC��p� 0>�(��DN�|~�òɢ`=ۓE�&c5�	���d�Qy�m��<ٗM�<Ѳ(�d�0(�q��h0+�i�N���Ҷ ��Q��Z�O�N��EZWn��%T�ѕ�ԉ�6OJ��K<�S��f�M�*���PM=�5��.2[��'�Q�PM�|�"�D�$\*d��{R*R2n��b?O|Pk�j+��A��D{�]qqO��� n�P/i��|�����X�se��KuR���Ž/��u��遺N��h%B	�ay��#5L�'�� U(͢b��Py� Ԭ1#��4�;D��C�ċBnD=2�^%p�u�@�8��N0����>�����%T�P��
I�XM��9�!D�pA�6:��j�<n����2D���Ф*����@�W�`���N2D���\�l#�8��LD
8����`�.D���a@'� ��֬� ,F���+D�0�k[�vsf�	�J�%m�B)�V�3D�@)U�ݻ|���C-ێO��[P�2D��)֍{5�	�En�0�~�j"2D��9��Dtvp�V"�BpS4�.D�d@��[4-؜��Q�I3S� ��g�(D��CU+�<1H1�VN��3��] Dk&D�4�rlI 5(��5�1�µ��#D�4X��M�b��AcnFeLU� �!D����M	B�@t[��+�ܨxe*!D����I����bG@���H%, D������tuVL�P��g��H1r�>D�tcaˉCe,}Q6�KI��S.'D����&�`�еqVa^'Crv�H2b$D�LѢiݎ^���LZ�)]N��k#D���ԃ�Aw��	"AZ.'�)���"D�\C�1^�
hH�#ͨF;�9aB�;D�xCgDdxI"H��<\A�vj:D��(Q��U�����e�-|�t�Y��9D��Zj���e�4>���� E��!�"�D�� �L���ْ!��>k�!�ĚR���Qw����Č/���Ұ"O����Q��B�#bC,��H��"On�	��Ū��i����j��	��"O���27�ᦀO8 ����"O��j�h\�X�8��M �SR��p"O�@:s�
</�@��k�,_D�r"O�XU��7��;S�ן�6�1�"Oح����c���B�v�.\��"Ov}��fm���R�?�)s"Ox�QBHˢ.��tP�����"O*���H[������)xx�<�"O��Ұ�_�r&�4���˂\��`"Oހ�n�+�� ��J*?D$ ��"O����<Sa���_.9� �"O@@%�L�3dl�A�"R�>��C"O� IbF��Z �L �MbFH��"O>�y� ����XS�_xX�1j"O*<zs%��,r��W�<F���ӷ"O$q���$P��1# �7�� $"O��eֆgZ�(q/S�*���X�"O�94��K���" lŚUZ<=z�"OvY1;�5��`I���A��y�f�\�@��R��g=�����R��y��T�`\�E��,�9��Ê�y��Q9W�4�r.�$"�労��y2��8H˸�@*��ȽУgܯ�y2h��B� t[�'�+� �(���'�y�Ċ�|<�ш@�&��dcR���yb��g�J�b��N�{b�ŋ�y⡘�d��aZ�6&t�qo_�y�+ko�8�愀Q_���E�W��yeGNv��׏�Mq(	[5���y��.�he�ܿK�ո���y¤��nVpٹc+��B�� �U��y��� ���d�n��2�H�6�y
� Nđ¯ۈ7��z��ՠw�}S�"Oޅ�j��[mR�(�$	vh��"Op��e"��A�H��a�K=cb�JP"O|�k�"�)!���i��Гp�`���"O���)�s����P/"�)9�"Oİ��?$�Hsԋݤ$X���%"O�<
0��i�$�	�J�&~:����"OPl��ď�*5�P��L�"*8���"O�c��ћ�0]3èG�	�ڱڥ"O0�1㒴bdP��M��P	�"OJ�Hf�l�,��2~ࠣW"O���(��l�z�n�Ã\k���"Ov4!��
B�c`�;<f��"O�%��a"t9Hu/ґW��M��"Of@�� U$�D�FV{:�X%"O��K�a��y��8�֭AUq���f"O>�{���u����,فa�� �a"O ��5OΕ7�Y�	�&WN$!	�"O�{B�
5h������!0�D���"O�e����	G��a�"���*�"O�h�wm�"s��t`BHƦP��"O��*�˕0��|w��(~�BT"O�����}��(��4J$ Ȋ�"O ec���B=��K�-z�,*�"Oܥ�6���w���Q͜�Co�PA"O�%�B��۬� լ�37���02"O�<P��\\�������)6~�aC"O�p�*TTMBPʡ*�vlD#"O�9Bf�ƿ.�P#rI18vFL��"OL�s��R���E)���u@�"O�� ��)�P�� Q��$q*�"O8�#�L�`jL�HegHz2�S�"O� �D���<�P���(N]�$;�"OF|!J?bu�I!G5S�Lx�"O*D �*�:Og����O�K�b�C�"O�hc'��?d�Ȉ���D/J�&�s�"O �j�G	;.�E���=V��@�"O��+�I��XQ.�sR�/<�%�p"O.��VÌ�F���a�̷���ʷ"O��� R��t��e׊U�$PC�"O,��a�72�0��jN�}��"O�a1@�DZ\ak'�X�H⬝*�"O�S G�@�@H
�E�v�<��"O2p�u�i��)B���"O�m�\�2�i���fm�d"Od� �;ގMS`��
��t"O�8U��>&��P��{����"O��aQ���[����hA){�1�6*O�T�c.�$8U�����$u+����'SH� �X �������a��'H~(��I�Dfv "SÞ����'l�!�gƟn�ѐ��MZ�px	�'_���g�Z�'�<a �`Z'���	�'�qp����O�d�W��6}B�Ъ�'"��Uk�;q8��7ƞ�*ld���'��Z#�ň)��ңE3u�
5�'vbDy��4=�����!� �i
�'9콣��ƝB��X�b�މ+�U�	�'l.�r����E��3	 ���'~���(Q
=݆�`Ҩٳ(�ʜA�'�����5EB���ʿIxZ�9	�'FX� ��O��bլR6=e�d��'��Ԑ�L�����I�"L��ة
�'�\U�QB1fH=�$�Ɨ=�H}�
��� ��-[�pԈ�h�H=�Ԙp"O�[�ƙ�v�j��e�* .9P'"OMr�hՉ><`�;!+utAC��'QqONL;0N��qX^q��*Цlp�F"O~4;��Ȕ�C�*\P��@"O䱸v�ñ>��� в]H(�ɳ"O �"R�JM�t�@�$\+�i.�!��g��ˢ��'q�� a'�B�FL!�$E�t�\��h�C�r���΋�!�$�"'Fxhkʷ�`����=z�a}R�>�T�o�6L�-Zuਢ�.�[�<��ȗ�N�h�*�P.���oH|�<���ܖ�\P��N@  ��%��@�<	g�H:'��C��ي*�X(�'�@yx�$Fxr�Z�o����i�
��Q�Q���y���zw����ۻ18~�r������"�S�Oq�@���_?i&��``�4�xC�'J�dp K�66�^�X�	�.�	�'�p�8�jM�*u�v���uD�	���~rkMp�Ƀ�H
g�&��V�ī�y2L LPfyه!�_�<pXF�Y��yR�2R��1��Z�����iY&�y��H�c\¨:���J�vq���F�yB놽2i�� ��E <G��8$F�J�<q��$c�<0z��ב&S�I� ��o�<�uN���Rӂ��qy��P��E�<ق�ӓc�.��
��f���i�!�C�<i���v�H�h��X,ku�y��W�<i����`����86E9@�O�<���
.fe�t�&}���$��M�<)c#[�zc�q�.Z7w宵`Ј�Kx��DxB
_�W��+��^_�T��n%�y�	0HET����Xn�|�`���y"�R�r#P����1V�,Ey@�N��y򥀣`�iBS���RlT�!���y2�Q�R�Aq�m�`���Wl	��y�M	�x-xU;-��^Ԅ�� ��y"ʌ)Vn�y���W4�����yB@ʳV�����OR�fU�E�ߵ�yB	כ&�V�ؖ&�D,j��H�y�'Y��"ܹ�b'C}Z0q�n	�?q�'�^ r�˗I�xd���ط&�Z�S�'@6$yF䂜t/�aK�IU"<m1	�'s�e����X�0=(D�^@'����'����_�]0$4Г�>��=ˎ�$>�S�$�<p�܂C�7e
�$���I��yR@:��{E�5c�bmS`i��+vў"~Γ/,F�+���	�:3�@�tF��ȓ+r� � �*U�P � ��:�PY��6�37�� 8y�k�M|,��I^�I��%z�"��R�L�M��bb��x��󩀎?<~�P�m7����N��?%!�d�8-��E:��:$���Ƥap!�F*t��ĳ��O��9u�!o!�Q�D'.[�O�>6@iF'˽cP!�D��3�6��ԏ�_%6�yf��:\!�dȩ0�v� l��T�9Z�!�X�}"��g�ؓNvh�	�	@�!򄌇1hH䧗�ewQ�('*�!��\Np ��ܛ^��*��C�b(!��9r��h��z[N��u�Ӭwj!�D:[e`��T�&%{�\���9"�!򄘾[X��aw�Y�ft����l��!�߁+��и�˅�>iQ�&ɌV�!�� H1�q�^^�LT�hʑ-�)�"O��K��(g�N���G�'�T �B"O�����Ť he F��!"Н�S"O"�XL�z�t49�E't��"O�c�E�0l��3�MV�|�l�3"O6��
�v2��MЦG��|�"O.�a�ؒEd��� -@�Q����!"O�`H�&�$=΅qū嘜�"O2�KŇ�,j����*P���T�P"O��!"�
��33�J$O��Ѳ�"O�q ��.
Z��r�5�ڵ��"OPh�b�߰Z�! ѶY��)@�F?D�tƣ�0"�2�ʶ���*�y�E<D��8�	ک ��1�% �@A%D�����;l� ir�A�=��l�cm?D����$�r� ��M�:Qc�*2D�X!���7T�B��s�NCB	S!1D����cƷq���P��]���P�1D���ܻ�`E[5��i��YP��2D��"�!;��ڶ�X�	���r�>D��!���9�H�bu����0D�̹D���.�+�
��δce	;D��3�Ȟ�pgX�`�&Z�%+T1jt�+D��a`��N�01�,�YL@;!4D�x!G+
5DM�QJڏO�R=
��<D�ܚ�ˌTTmR�Y0�j���-D�d�dCͳښ� UǗ!f�z��&>D�X! ?!\��C�F�m۴�KC+9D�,�E �++
r��$#�� ���J7D����"K�n�e��W�"$���3D������`�r&�W9���k1D��9�$�##���IRA��/R�B�"%D��! ��<*3���7��<��ȃ "D�`�� 9W�uq����se#D��k k� M��źTA��4����6�"D�|9Q�N���(��J�~2�!)E�>D��Ì�u@���Ћ�3���L=D�x  ��p��h�D˖%n���R�;D����j#9aƝ� �T�Np��)�B;D������~t�ff:{UXU�7-=D� 
u�	�=�1[S*ڴ2��x�1K=D��Q��q�<�8�f֑O � �e�;D���J�yw�u� ZwOڈb�:D�ȱ��>��{�v�t�#��9D�t ���:VWBq�a%�]�\���5D��1k��T()��T# $j1Ѳ'5D�$�F'8nR�9�Q�&����=D�+���u����"fU�$��+8D�@�"Y�O�TD�#�J7 f܂%�4D���NiÆuȥ#ʞS���ä1D�X�У��V�2	�g�ܐ,�$�!qk.D�$��LYgDd����t���
TC.D�h�bJ�u�+&J�>���RF?D��1�
U��X��%3^P�8��<D�;�ÿ;(�m�/C�J��K��&D�H�ځ02:���ʞ�Z� !�7D��S��i^ġ��"�,�k�`7D�D�b���p�H���=~�a2b'*D�X�Dm֞"UHă'ܚ^te�`a5D��I��Y� 0�Lڵ/q^�r��%D���0-�
	�`W�L�f�j�q�5D�T����9R iS��Sh8�3O5D�l�f�]�옉!���!� !D���`˞��24'ƹP���uc4D�� �E!g芌5�m3��U!u].Mkb"O<�"���f��p)YT=p=��"Ox��.��aٶ(��C�n5�b"O�����90fR�a�g˪3:��"O|���S�������%��j�"O6E�%IE}���cD]�s2"OJŊg+í���	m����ƫ	'�yr%�W���ʂ*�)iژ\���
��y2L0Y�f�1���hC��׈�y�I�XWy��^�]����`N��y��ɬwT�E�Wâcaj�b�R��yR��/d�\3 BAEa� c���y��J�L�r	�)K����b�V��y���*g=�0�F�L�~����E��y��ʉlm8�9uMĚ}� ���΀�y�̊���ʠ��	�Z�S�6�ybiwr���	���������y2�\0/�n�����>&���צ�yR�Y�H���%"�4����V+�yR��f�9uG"��I��L��y��u`�}��H��e�y��W�'��h��/�.+fP9fb֍�yb�B�m��@+R�v(x"�)�y�,F#�X[���2��<Be���yr
̎r�J�8gS�$T�<`"�˅�yb��0qXt��F2"���y2�L!�dɻ�ԧ���s���y���h�Xu�"g�%A�Y*����ye�61&����(w��kU%C�y�K�"kL�� f��P86����y���9%& /$؝蠀�T�L�	�'B���&��$�\X`1�M?J���'���
�'ӵ$ڡ���=�\I�'�ԙ�D��n���c!��/��!�'��E�T>Gp��3@����ph�'x��-D��"�0�bР����'��1%�S� �u�îU�rD,|p�'�L��d�H�A��`�e���%�v�<Q��ֆ1,Xغ�o�:u}���#��M�<�r��9,W���&fL�< �,A���@�<�%^C�x�XL/_��l0&M~�<yvoR�1�p��`U�3)hI�R�y�<�(Ο]����T�ϮQj���`Cu�<1�ꄛbށ��A�h��Ɋ2�7D����a�>l��X4��?�b13r"7D�h
E@�-3������*8\�2�#0D����/�
}9��b!�O�,%0��8D��*SK�6j��SW͒)4v�r0�4D��&����ĨZ��V<k�<s��3D�(3�ES7V
���g�*b�lH��3D�`���0�F� =�B�ǀ{�
C�	 >���{���`q�8�`F�N�B��} nM+���� �|���� ��B�I0�� 8c�$;`���[-�tB�	�w� �8Dhօ,Y2m�TC�)O�tB�IˎIS�$K�Z�B}P�	E�o|�C�ɫFu����A[�@z}1�X�0��C�I��I��a06�Z�`s��@�HC�I� ;�M-w�|X锆%vTC�-<�^Ԫ�k��]-�Tb�
�"g�@C�	� �����)TnD���n4C�
A����]'�>��#��y#�B��3h��ȘCB�O����D�P98�C䉡��� �I�#x�U���!X�.C�)� �[=)kj)�G�3k��(��"OX��Rt8jl�`�E8,)�"O��T&NE�PE�կN|IJ8��"O��ՀB�H���`���"OPy��S�eG�$�l�#]R<�f"O\R�S��jz��BVF̵�a"O<�B�"��7`�P��d��E+�"Oʝ����+N�,��co��'�p!� "O@P;,ٓ[���VoI�F�8��q"O�A���Dh ��A�,ǜa��"O>����/ZN�P��$D�|Lâ"O¬��� #��p������"O^� �A�;�|ͳwl�4uf5`�"O�@aF� �l<���Ń`��Q�"O��F�֑a���/T�|���w"O*L��-^�������S�bԲ�"O^�Ebw9�-�W��*6��M�@"O5����b��U�A��}z1"OH���,��@3TE+���I�"Oa ��ĳa�t���F�w����"O~L��"��>\�9����-0B  "O͛��	�BW��"B����RaI6"O�t��BC�,7Z�QQn���[R"O��ný���1���4���ZA"O`�ٶJQ�^8
m��b�[D��Ё"O�C!�	���x���R/-�D4jv"O<[�%��J��V@X�.�V�Zr"O�5L?lX� k'AO��
�h0"OY�r�� �h��v��F��x�"O:X3X�¦���`�HLu!�DR�X	FM�)6���se_$lb!�$�fk�@r3ϸglj��d��L\!�=$(`���@!	1Z,(p��2jK!�@0��7LR�t��{�c�(U@!�Y�n���d@[���uHS�\)!��?l�Q�b�G�����NH�!�$ׅ�,%�w�.~���Ҡ*Ҵ@�!��ȼ"(�ٷ�]z��8a�̉t1!�9S}#�ˏ�0�@��&�!�d>e��A�A��,�����U�!��%Q��E3W�]�K������j-!�d6�v�aa���8�N�aC2!���pX�L&��
N�8(�"]�O)!��w"V�#(���``�(
!�Dݐr1,U���k�t	���"�!��W��	�&ő�>S���;�!�Dǲ8�"�E≯R�6x��ʗ$]�!�$N�1����b�=2�\��� �-�!���"�h[�ڦ:h�C�b֓4�!��yZȘ��K�SHμ:e�ј{!���;�D�U��S�8I ���-0v!�[)-�&��0��7K��E� H t�!�$�3e����[<��d:3��j�!��7#���!�%� �FCҋ#�!�$D�q/ĭ�d�(�ذ�b��-N!򤊼/�(a��Ԫ�Ul�{0!���(�(�h���l+$��AL�/8�!�DZ-*PPx��,Y�(E����lΣo!�Z�^AҲ�3
,�8ȶ��k!�2@�t|���)+����-%�!�1EЉ)���*�h��On!�$�*k�Q�S#{�$�:��ىia!�U&�}����f�%���ЋU!�DH86��X���Y;���ѕk��+N!�� ��#��q�:��C*T#X	�t"O�����߅A�d��a( �&�)�v"O��@��z�>�: �R�U���"OKǈп(�rHh'�=�pe�p"O��Z���Q�֬8!k2(��{E"OD�9qR\ A��ɛ�1#T�� "O���Ĩy��c����R�z�"O$��:XX�Tر ��zɈ�"O�����}�H�he@̴8��0��"OJe9s��)�,�zB��'>�lՓE"OHS�畭����mO%
��!�"O�-�Slܴr�"܊��I��� ��"O�ԁ��)eR�J!*v|2�"O� �tC�%E>��r��ɠ@�*t��"O�5eG�H���)'nQ:Eg��"Oa�A�^l�˂ `. a"Op�W�+r1�Egj]m���"Oڕ�@d՝M�(�"�o���"O��PENƱz��9[t)��$� ���"O֙	�KG�H���R� �0,��"ODx!�*��Lv �� L�M���� "OV��6��
�����@�4�k�"O����BȤS�V��0ś\�����"O��[��,1��t	��LPu"O�{���Z��+�A n��5"O���c&�=��iQ�`��?ȮMjs"Ot��3�?�0�I�3Z6�[�"O�p�A�z�Fm�H�LA6Ո�"O"��N.������D7���1"OZ Ԁ�H�.� I�4��4"ON`!�
2'?0�Qs��:N-(t"O�x�WJ�j\x���OU�?�D�%"OT��Fmâ@���r��M(=�\�D"O���2@�=0eK���e>��"OĜ`�N�vdXrc�k�0�K�"O�բ���."�YPI��66M��"OQ��k[	r������x.�0�*OR��Tc�=5ΰ��B�B��Hu��'��vD޼58�s/� |M��'�j�RL���&�2&�fzؓ�'���� +ϥ$	����@D<m�d�{�'s�m@g��%\>Pd�'O��Th�$��'X��E�h�a��툲>�Je �'s� �@l�[�Dxh!�K</��0��'x�[�p�И�S�$�
���'F�<��ګ�$�0�&��d�P�9�'� |J3��vU�����)��j�'�z 0��V����htT.l�8qi�']�%)��D"I9�)(�L�r�,#�')��ȶm�d�|�bcY.��-h�'�l��3�^-f^-0�o��P
|�z�'��	9 C��,��!�M�V��
�'Ҍ�0�LŶ^��h���>> =`�'j���BԼI�l�P��9�6�s�'*Zxb�hؑ?����	NV�M*�'��<c��ɝA�b1x�#ȄӚd��'l̠���$l\�Ц��%b�*�[�'��@�Q�q$x�+G�R�"��	�'v>���'�@\[v��v�� �'�j���I����кb��<��'9�h	�+;,H��A�'Z���'#�3��Ӗ?�P�k�Â
MP8Y�'톙���کX�聸s�IБ9�'�v�� �]�1p��9FK�@���� T�s����:����ƈ�
�8�t"OR�sD���7����$ߘhlr�(d"O� "����T�0YbuDBR�$+r"OzȊ�GK������57.��1"Od)x��G�+H�Q��
�0,�~E"�"O �����3f�ph�����-p"O�p[�
	f�]H1��o�z"O~50��J�f���zcM�lr^ͨ""O�}��o6x���T�A6�1d"O �{��D��yw@��0�"O��"�ţ@ � &����x�1b"O�ХI 60�h����Z����B"O(t[��ܶ|*�3%���nq��E"O��`�W�B���E��Q[�t3`"O��x��A�c�B"Ӓ]U�  R"O�mqEb��r�X��Dk 2Ra��k"Oƥڄ�V/`:ƥH�I�V��)�"O�9n�c%��#d.�'^
 ��"O�x�d�ơ��!���Y��	�"O�� �"�||�S�׻:��Q�"O�ᐕiU:ZE��.�
r�8�v"OV�����>��1�8^�a) "Oȁ�H²r9��I��ҟw,$)�T"O�	��� 0�D�҂X7˂ �"O4� ���05��BE�=��}KQ"O��"���YU�衂!K�l�(���"OxD	�_�#������8~R�{g"O
QaD�Ño����><�&�y�G��M^��P���ub!�梃�y���!�^i�2˓*r��M ���y��C(j�6DXvHI_n�|����y�N.e_�8V�DP�P��퇜�y��J�C��$�@(M)�-��,̲�yb�D�J���A�87\DX�I@��y�d�!V^�M*FB)3l�Pu�H.�y���O�QS6l[�*-�1	U��y��,/�F�� 
Z��J^��y�)�J�c���
X����E��y���;�đ{ġ��	�H`�ȑ8�y"%Ϩ_��a��X�1�6���y˟%�>,��Z�.`F��U�\-�yRD��'�p9��٫%��9%�Q�y"+��n��<��H�
ٔ�:#F�3�y2���g;>���
�)���yҭ���yB�ޱ<`�����J�����d߼�y2�ʁ��Hƭm�d�b��/�y��&4��IC�ÒP��+'Û�yK
S;���Ǣ��!x�',��y��@:VH�@ � �|ܾt#�*���y�"��H�t� &u.�R��-�yҩ�'>��!���]	R@s�����y��9wK�<���0H�z�v���y�(���"�õ�F��P����y�6/��q��Ռ�R0([A�'��:&iU�KD��`��آ#,�8�'���� I ��tj��' ���'�nT���ݶwlN�@ڼ9N���"O�m�w��e���	g�+] �M�"OR�)v]>Ernd��	��P�`A"O�(gi��q֐��b�7Ԧ\y�"Om��H�I����aͪWi�"OʐkSm r�C� ���pq"O�᜙a?�\���	S���"O��s�
JxP8��'�4��a"O� :qq��L|�	����d���"O���5�r�b����G�i����"O�-���ʄR Iz&�Z/QP^1��"O�� Tk^�C�X���W�TI��"O���P�K�8�8�a%��!ڴq"O���@@(7����W�<��!�"O~�س*WF�p�	6��d��L�E"O~A��$��?�����!l��X��"O�|j!g��0�yc��g(� h�"O��
d��ke&)��`�<B}��"O��S �#����G`E-I�t"O�l�ӇW��d�ʍ?I�0m��"O(q�&�)q�Ԥ��)D�X�b���"Oz�jӦZ�9>DP�'X� ��d��"O�Y�qdn�R�8��ApT��@"O�AqC Z��cRu����1"O��)�3!0�̲� ��r֮�Kb"O���gG4��D��òu�Ո�"O8\Q�%�>(o�8ӑ�Tj�Y "O�I
����v��(�y�׍�!���hTkЍ�!j�:M9P ���!�´5�X �Ձ"�^1�@	
vD!�?h��c���;B*%���Q�!�d��>�9��Jؚ+%:��%m��!���.�����{!�q3E��4�!����|�P�Tl,�"�HT.�!�D�1�U�DƏ
LΨ��gLR����l��}1e^�s��A��B��h��|t�w�4T��5�
�i(j��ȓ ��bQ�z;8�d�$Ae ��ȓp_Ʃ��EL���ՙ�m	���	��pʐ���ۂ^�Q��jX*�����e������25���u�����lt�s��M070���V�D��؆ȓ~Є���a��!�(T�#炇��ȓD�<B�Al�B!�W5P�MV*,D�����V�zS���`kW�}�XA�*D�h����-���l�/K̤q�vk'D�0V�>,�d��q�H�%�@�R�b%D� �@J'o��᱔��<����� D���cgc��d���J�lj�>D�P�� �2�X�+R�n pЁ=D�,#t&�$��3@�M�m��:D�"���*1ZX�zi� /,�Z�g<D����&Fʽ07��>�"��F�;D� �J���(9�`oM� � L���:D���d,�"G�d�	�>����$D����MJ#.�Hd��*f�*I�$�'D��H�`�5�z�XbN�0)K�pj&D������-�$��l�����D:D���g�\'�t�8t���<�t�;D��J�j�
,�r���z7��j 9D���i6T�Q#H�U~z�a�	-D�Ȳ`�DZ��YQED�t|z�C>D��!�G�^�	&��s͔<�'m8D�P���������C�zT�1 +D��j��]��]�b U	7L��q�<D��·g��p5�8���!�DXQF�:D�@��_�	������ $�8Ԁ�%D��+b,+	GU�錍<��e��e$D�����HX����ǶN̖It�%D��bv�/D��I�i;n��9hơ#D�����V,zx���Vǁ�/T�%��!D��`��N�t�	��F��V\H�� ++D�� �yKP@�7Tal�8�o��k����3"Of��7��/�@dS�LD2|�T�("O�Y#��@Z�E�#b(d*�"O���W�CJ��J#�E[���"O���VE_#F<) +�� �["O��K���4f`9 1�C���I�#"O*1��/B�
����j\�L��'�|�b���.�x�J��\4Ut81{�'����
�A��=�!�*K+�}r�'ҵaѪպM���!i�w�B%��'�Aܢ<����@�7aԴ��
�'U�Q��n:�ȇAU�G�x1
�'g�h	1�¾1
|:d��E�($�	�'CN�2�.M��ïA�Йq	�'p��3��Fh5�b�Ԃ?첈3	�'�.���
�37V
%RC�2<Bl���'Oވ�Ebr$����LM�1D1��'�H����N]���Ѓ	�-���q�'�:�A��1�5�/&�*$��']�x�!-�R_���ↂ�-�N��
�'����H�E�� �`�y�ĸ	�'dU�w�2J���腡���`��	�'��h���ˠ�!5i�$�\9	�'��$�A)V�:d>tH���3�\P�'`�h"�Ŗ!ho�G�D�e"O�p@��,?�ZL�#N��?�� �"Oހ�%�ATp�# 
FXp7"O��A`E��F��@��'��HU��"O�l�4��:-�~���&J�Z4��1"O��2si���UB�8�dR"Or`�#U�;{�p��G��"��r"OL�f�C�mŨq�䖼h�hS"O��PE͑8�	;�,͛7�R���"O������a�.A��6 ۖ�y�"OF��0�̏V�.�paa �"�5"O���"��.}�T[� ܛ~��C�"O�����')�$�h��m���yT"O�����'��v��-�~���"O�rYu�Sv�F���9i"O�LȳB�5�R��2�O ǚ�[�"OP}�C�;]>D�b��I-��ዣ"O"�b"��vj����W͂ B"O(�����&�����B-�`�"O��@�(�r��CC�F>�E"O���5�խ G\ʃ�G!V��yQF"O�p�a��=��hF�,t
b"O�\�G��tk8�X��F�m�<��"Oؽb�O��n�X$kF�ܣm�U#�"O��X�׵d���G%ʸ&���R"O:����#^�@jq���:c��ad"O�RPA�8O�>��C86���c"O,��������c�#ġy*��"O����#�7�|�q��W!G���!s"O�U;��Ǆ,���f!S�	�d\�@"O�J��,�n�*�`��dtk"Ovܙ��b�qʰO�oSP�aC"OLH�b��Ď�8�]��"O �2��=�6���&��]#P��"O�\ō���1[S((D����"O�tcR@\",��S!�χ?H%��"O�j�Rhr���A֏�A�"OXd����w�^���i��F@�""OZY��kJ�RPq���:T�'"ORt
 �F�x�x��'T�[?� q�"O� <���o��1Jf$�Մ��{Ԡ��"Or�J�Ϡ6��`G�A|xN�� "OZ��� l�m�e��?Sd�QC"O���(?UpH���83J�R�"O蔡!���<)b�JY�2�U�Q"O����P��)q��'��Ӡ"O@f��S]^�wBJ�$��"Oΐy�ŏ�yX��o��`g0�ɂ"O�Y���$=�]���Ö/G�ȈU"O6@ W�I ;���� ��l��"O�+s���v��f��
$\�0"O�3˂ .@~0@��TW�T�@"O|��`�ƾvR8�����j��M�"Ony��ѾaG��R%B�*)�y�"O��`+��Uz$�
��l��`"O���oƭ&�vEuj7���	�"OP�� ��n&�ʃ)`�,�y�)D�4U��aI�J#�YO�h�E&D��Y���r (<�H/b<��Y'�%D�re#�	&,�A �&v�P�vn1D�da��63<I f�џODQ��3D��)p�V�w`�q�5�\'7_�c�-2D�\�g�"_�$�����6l�`8�&D� K��ȑ�X � FG�pB��:� D�L���ùq��ق-F�5�h��Q�(D��J2�Y��D�� �čc\h�i%D��Yw$�&Fɂ������c$�P�B?D�`#���M��y1b]�<���-<D��;t�W�_v�̪�J�#�"�G�8D����	˞`r�t �X� !b8D��#�HC�*�a�K�%�Ш�6D� ���H�!`"�⃯�C&��i%�2D�t�\-Xut���!��Ev��i�+D��i��F�P&,Z%�ϝ:(l-���'D���!���A2�-U�j�#b$D��x�HF�?�q8�.�8bch-�H/D�h��KŢX�ꁀ�e��?$r��'D�ܰ���4"�����o���;#k D�����)�v`��\.
�!3�>D�X⤤�/,!����7z�[�$>D��B�e��Uy'�	05D�yd-'D������>!1,0���_<���bm#D�H`gI�X@���V? ��Ao"D�T�1��u䞵��
*k�F���$D���fԡr�"T �9$�6�2��!D��	p+U;I����I*.�)�o?D��b��L�́�enܾV ���1D�0��\1��L�� U�^�yφc�<Qd!��TY�{�Y�elX�Y7�b�<q��DØd+�
�>�2-9��HG�<і���[�q!��G} &�8�ϓJ�<��)3~eåE;kU>��.G�<����%s�N�r����o�F��c��B�<� -s�`C�"G�h8��I���D�<���}���A��(!v0�&�h�<y��E*8 �a�Ŋ%:�d�)�#~�<9�d�V1����CƤb?��р�I@�<�s��}k2Y��E�q+�YYw�{�<A�.�2��M�A��
X�p�GkRl�<����d0��0-ˈG]&��e�d�<Q�ǔ00A8��@-�=d,��T^�<ia�]�g��22��*g0�j%��u�<���,�R�kF(B�jdH���Jo�<A���	���0�E�#Z.�s$Rk�<� *ȳ0	�(-�y�@��e�R��"Ofa�ҡ�����+�]8���"OH���M������/�zK�"OFum�h��qF�V��N�Z "O����A�q��B�J��3�"O�s$��9a���a/�<��Sb"Oh�e#�2n ��2t
���"OE���5a��}����4+�.���"Ol���I\
b���8�j�./�>�#�"O|8��g�H�Xe���
�@"O�L#��-$����F�0��"O`4q��֒sF�mC��[�H�ԭ��"OJ����Ů ifʎdG�D	�"O�u��`���"��2y!��)W"Ol)(E���39Ia�%�!:�@�"ON�2�!��=�I�0�
!���"O$]�k�dF�g/(�.�:�"O�]��+�?����dA�5*��*�"O��C0Nٕc�$q�C�t(���3"O�[$[7Db4�:p�O#�h�"Od5c�g�n����A`V��"O��P�� DL��F,Ԛ����E"O@��tL	h1��bfA�'Ϊa�e"O��K�B3���B�12�"Op��f�՗��AE!F�H�\]�@"OS /ьbҒ�ytO�o���"O����	LKl@�2�˂p�@�V"O�h��nʼ�4�߱k��Bd"O$,QuÊ�:��(b�޿glN�s�"O�����5��1�ʀ4����"On�C�� �j��u�O�^>���6"O8r�6l������ɩ6���(�"OH�kܧ�$���E�w0L��"OK�E�0p�E��\�Ac"O�1`����5]�k����C�����"OŁ�S�Y
������O�$4@�"O�5��M�
-5 ������-�^Y�"O"p��ҳ|�de#�.R�2��� "O�����X7^����2$V�)J���"O���G�lT ��$``jc"Oj%9�NÏr�����+���"Ox�x��V7�����gB�:��9�6"O��z!�h\D��E�j��,k�"O� Z�g��D������̊u{(xh�"OL���~MZ��A\w5s�"O�a;���u>�J��՘]�3"O(%pc�X?8�
a�&  &� 4;�"Oj��fh@�s�Dqb�	�A���B�"O��R`� [�� 'ψ\�� Z�"O ����Vh���5��RA�Q�D"Oj�G�(r�B�*�dS�J�z���"O���AO�f��b7���a%^UYs"OfE��	�!Y` t�W-�<:9��Q"O����N��I�[87#���C"O� 0%%˵q�<�:���	?*�h"O�=����@C��1�EQ�!�T"OFx����:&�D��'˃
�쑂"O��A�j�9A�\P�հx�`���"OnqKe�ݐc��Р��9�f@�F"O�0)�ʑ+t>L�1��;�|Q1�"O^ [�Iȅ�D3B�αqt�`V"O� �E�<���$-�0mjH`(�"O�����ǥo��ȸS��&��a8�"O��B�DR����	S����5"O� e��MX�J�LTQ��T����"O Q�d- 2�FD�e�D��ش�"OqrQD�	Y$])2I0!�:�Ã"OL����]�L֚�ҥ�M� ���"O�\; _�=�T�Ԧ,��'"O��8
_��Ud�)N FB�"O!�F��_�s�b��E	@�5"Oz���&N>�
���	��"O������(�-S2��*�j��f"O�D�d�K+K���P�ܩ�2Q��"O���JF�%o^=$�q�5�T��y��	�2:��	u�.���#5#à�yb��%K=���ԋW�7% c4���y"Ǔ�~��4�0���/7���i���ybF�!X�d��T��S~�Pc2���ybM_�SN���f��?<&u��&���yO�z�hP��%�+h��E���
��yr��o��zPAT�U�4�pO��y2�C*��*�@֊=њ�w.���y�*T�CPX�T��4�Y�I^��y򡓔zy�Lq��ׇ,J�;'�ߖ�y�
�#>C6�r���*�����
�y�˂	[,� (�#���t#�Y=�ybm��/X5i�$X�5�,m���ߧ�yrIWbɡ�IZ舁(Q��y�&�r����.Nx��%��yB�n��I��n�YUa���y��B�2�F۝�V�ڥi�(�y2(V?lfd(	@D��~i���㜔�yr��q�,:�!�q���`5&�,�yBi0<*��Ga%!���s&��y���d F,��$L�&����)�y�DS<�j-�WmN(}��E02E�"�y�� +q���7eW�E��ы!i�)�yd��
T*��
E�Ha�̀�y�{Kh`i��[ Sx:Td�<�y���	r.e��o��I�7�S6j�!�$L8!�l:@/޸;|�U�F���B1!�$� >��*ԬcqFm[2�ǟ;!�$S�4����v�\ ## B�R�!��ɶ���3��+d:��d��$�!�ǄG6���M�a��0A���!�Dşc�4� K�=1~��sD���!�dΧCp��Q���qL@z�`
.J!���-S]6�ڗc��; �X��Z�G>!���{J��c@��	&$mr�F�J+!�C�~a\����3  �S��!�D�4\H|(�M݇s�B�@r3u !��R�s�xJ7	=,Q�Sb��n�!��D,�qx�	�V@|)ag'C� ~!�S��d��W�E_VT%[���>v!�dH���xS@�׀s84�[��_�!�D� <l��hʞ=�	p�!�B�!�@��"K޶|Y�����!�D�
K۲@c�F��C��{�'V�3�!��1j�������4y�aD���!�DN�J����L�%E��!b�"Z�s�!�^>�d����$�R��Q���!��E�/�(�(>r=�A���H�!��	�y������'5�(� jP9�!�dT�u�
hjq��� ��J�!�ɸDO2!㇫
F�9�O�B�!�@��Hs�	EGR�K7��X!򤀤 P��hA�]묜��KC!�� �� �ک(,�ܪM��x���#"Op=�m�H�Ų���V��Ѓ"O<).�"L9`d
ݚ(��UP�"O�U���<|�
)��#�@�dY��"O����	@r2����M�|�g"O\m&<wz,��kF�r"O|h�%Җy��� h�| T�"O�D�Յؙ}i�H`(�4A�H"O>@0C� ��d+2턶=�	:�"Oj�b�H t�p��^�*v�j�"OL@�aDO�:��|cf��n>��iR"Oܵ"��<L�^@0s�пIL�D�"O.ȡ��L��8��B;oA�횲"O>��*����Z���=Àa"Oرa�Dm2$Q2��f��lc�"O��H)~� ��sI�
�RP�"O̬)�NY�@>�-�ȓ�d܌qʢ"Op�;��QF��B���~��"O�1c����s@p�G�]�8�Ɛ	�"O���r_��Q�-�;
�mcS"Ol��$@�  N��9Q-Ӱ	V�mف"O�pw��k�vx;�N+6�d��"O:��pR�`Q�e,�N��P"O~�c�&D&}M��!��5i�� �"O����Bf�ƐX,I�wr�,"�"Oy�։�7r�+�%oU��r�@Ku�<@���9C�=�t�ۦ�l�g�<���; j>���l@�Sy��*�.�y�<��H�!� S:e3�H�"�J�<� �P�Z�b�z1̃+';��kG��D�<`/~���d�ɱ�x�)��L@�<a�� �9Q��(��"A�ȓ'����X�!Ȝh��K�-@��͆ȓ.��$��B�6�J�ZE��.%�<Ԅ�mœeB*(�!�r��T�.��`�ά�f,��t
� ��G�]��ȓ*q�|�&k�Zʾ8��k��7,Єȓt>�r`l�h�ꠂC�ڨ�d�������RGP�b�0��GLO,��܅ȓ)���� n�w��pr��%"d
D�ȓtR,㵩K*,x��b��1m�`��:�݋�f׾|�������eĂم�.j0�x�&�/	��`��<z�ڬ�ȓ��US��'�j� ��y��E��A��|�2�:{|���(�3~��Q�ȓ��r^,S�n�Jᅔ�,��H�ȓ6m8����=�J92W/�: ��U�,��aZ5�@|�%��$����ȓր������7�r��#Y�\*%�ȓ^��Xۖ��2�v4�gB!~�A��Cc*�質A�_�Y� ������ȓY�F�K2��~�hrDC��J�\��u���靼S�ųw��_ݶ�ȓp�|��$U��1��D����ȓw����[-+���
bĸ1��cx|���_B�V�&oL,G��ȓ70��G�Vl:𣧮^K(���ȓS�BmCѣ
W�Ybe	m�v���Ff�=�5HԳ[*�T:Ĭ��N16���uaR`QD"ϚE���[!rE���:=�"��6H�AvZ�
,D�ȓ L&����?TŤ	iF��2��4��+n���ș�-8�X���Q!�$�/�F|z'���5��s&e�.O!�� Ru4�W�-2�q���T�sPzH�"O�y���ZHl�	T,�4>F��"O�h�A������0S�9G���"O��櫓�"kT!�rʝ���P"O�1 �LVC��#�"
���`�"O(43b�[T�`��@M=T8@� �"OB���@�a�ҵe��v.(���"OH�H��éc�)[焞4PMd}�e"O�4��Ě:{�\�� �(�r$�b"Of�zs��J�t	0EJ	
r�6�"O>i;�\�@����Vh�E�&Y+d"O� d�U����CV��]��)B"O&���7�&�/9ή9�%���y��D0���R�ό6Soh<sD@��y���6�P(Z�aT c�򡪣�1�y�nE�h 7�V]*#BͱQ��C䉝 S�)�B�4���qh�(q�bB�I�'b>�Z�7���wDH%]�C�ɡ��A�p!�.t���S���<k�C��t wF�6�>=y�(D�K�XC�I�-�������I,M%X�C�	�5� ������M�������%��C�)d���te��vfr���
�NB�I>�2���Zk>8��HM+C�C�I%ls�(`J-8W�Y5��
  C�I�F0C�Q�v�*&^��/D�� 
մI���R�J�p�ZȺ 9D��!FQ�B�v�J6�
�O���5D� �E55�ہIM�_3>�u�5D��ؕmơ��`ݛx�aD#?D��h�D�(2�D�iG��K��Q��=D�lgq�!�q�ʄ)D�U�Ӆ�~�<áG"� z"oX�-h��QW�}�<���9B]���:u �AE	Wq�<!��<-��[�m�A�q�Ҭ�C�<QNX;.��VlS�O�t�5��@�<�TjA�$��rr&�	��@����}�<�u�E�;.<�S.�<ETD�#u�O{�<9�c�/'Y��`œ1~�beG�s�<���]9�z3��l\B쉵k�k�<)V�bqI;r���*�0{���r�<I�(�+J؜�qeN[a�����c�<YL�
�x�N"��J7�]a�<��#_�<k(1�,��)���h�A�<I`�K�W�
��&i�?T��,a��UU�<��g@4�����	>4W�����G�<�e(z�.��t#X�=_J$�D�<���~x��%߫�^����y�<)ဇ/X�"��2L+GBx�Cu�<D��>� �Ώ���S"EY�<���ϨN�^|��" �ќ�[��}�<��8p�L��pKG�<�t,�E(�x�<��&Y	PL�e�
yE �(6H��<q��ۛ 
�Q�a�A��d�QnF�<��c�?�b���)��L16 �"m�L�<� ���`���*ΰe�p)��a�<�!O�)3lڱ"� �_
xU�G��`�<�D��3 �&��$(c���U��w�<�!��8j��Q� *
:_z��P��x�<y�DOD4d���8FQ��귣�K�<��� �Y#4LȌ@wh�X�D�<�R���{��3EJ�[��5�ǈ�@�<��)g�UA�
W8[������T�<��Ŧ	����	�������i�<� j��5�	�c+��K�KN�n�z��G"O�� v��<�1B5��*l�l�h�"O��B�f�;J��(;VF�f����"O�L�P!G�y`trs�Π����"O��F* �//�|[�TSo���B"O��)���q���᝕�0�!"OLPqGHT6u��o�~�h��"O��iT��M¦��-Y�J���9P"O1�'��������8*�4( 2"O��㜙	�(��-��h0��"O�`�2��P��MѦJ���"O�Ɉ$��X����MR|m@�S3"O ���-7(�ȱ�l�`v pc"O�)Z',���3"���y+,���"OT�2c�X&1@�2��6"F�KV"O�{�JW� oց�C�G
9���"Or�������XH�&I=0�t�X�"Ov�1�ԋY	*�+�nU*�(��B"O��'�K�X�8)6�J��49""OT�7'=���7*�Fv�x0�"O���C�	-�@s�脪l2I�'"O&��aE]%��`	@�E�Ĝ��"O�%@áY�9��������Lq�B"O�# &��n[��ۢ�٧g�|}	�"O��	
�|�*Tjǅ�6 !��:"Ofd�pBιH͈�kU��9	���r"OhU�eK�)S�P�D"T�Ӂ"O>u��%,Zu���Ͳ'�8��"O&�d���)�����!�JC��b�"O�yb���G&��AϞ+,\�|"O�z#��02�H�S�,�i� �e"O"� �C�;�v`b�H��M/jY(�"O�4x��,� )4h�?P8�Ԛ$"O��Aqo�!]M��H^43F�"O^��c�y�D̫$l���D01"O�ի�X���h��.پ�1�"OH���ցw��2E��H��!�"O�}�-Ɛ�FQP.B�A�"OҀ�%�2=��B�Td�"Oj%����E�DI���H=D��m#"O�)�F"	P�`T+���E p"O��c��:)�AQ�,�\)D"O������r�A��5%�	�V"O��
��&��lA�&@U��"O����>#���X9xAR�"O�@��*�,����j�) *]�"Olx:��)
�kVd"�:LZ�"ON�@#�*�Є��̞N���Q"OT�6"�YP��С�I�u��I�c"O~��bI
%`|`p@���.$,� "O�|�t��,E�ZuA��ϣo���kb"Ob\����M�ZUu/�ⶐ�"O�IJ��C0o2"�@��� ����#"O@�ӑ/Vzt��c6��9UhB1�$"Ox�ӱ�!����vi��]_`"�"O8\{�e֚*�|0#P)�4mc`"OF�3�k\�[���%�Z�8��$"O0HÃA
4�!�ׇѻe>�[e"OE��jՋ	+f���& �hpq"O�]h�� `�0�z���@��@V"O�X�bf�DU�|��,ȁ�P"O��:�(��5,��9��s�`���"Oȥ9d
ư��	�M�B�"O��@��B]�3�"D�Vʲ�P�"O� �]P5獷!jj%��b�Z��4��"O\�cf�	4/�䌈��-L�$|"O�-A�l8�P��jS]�����"OBd�D$(Iµ3F��?n��uBs"O��Q�lL��J4b�.�'Rt�H��"O"���≐.,��XmL�h Mѵ"ONi�!�W���C $%��;�"O�ceI� $	����Y^}��"O��f	ͷ" �Y�Ϝ�	�P{�"O|�Fj)?
�A�H�-r�Z�A�"OR��3�Y)>�Z�)��*r�dmzw"O����ϕJ�<4I~�j6���yB'J>G�
<ʅ�Y?A���j�C��yB)փd��	Rs��l ��LC,�yᝍiv��@%��c^��%�׬�yb��H"pT�vJ��s_�*u�I5�y�j�! 6�|�$A\�g$�Z�����y�J�<���@X�I�Qz�ݽ�y��F�0��
%I7��p��I9�y�D���t�� �!_^�(p�^��yr��ffnE�Sj%Q���qb��y�)[N����"�4Wب:�ܭ�yb!ߴk�⌓եB�&a�0k�\��ygO$��̫Ů��!�H����yR�V #�ƕ�ʅ:!�nԐ0�ѻ�y�ԪlBls�-X�@)�P'�9�y��8#d68�c[
$�tC@nY�y�	�/!�|�*��˭�����)2�y�̤h�bI�0�ϐ#�4-b��Z��y2�E�bEX�d	ǋ?܄Ӄ���y"�m؈ݹ�A� ��1���U�y,]�m�<� �r��-��A��ybÒ"~���V�Za�2�+'J��y�e��\��e�O;�@pQ��R��y�&�>J�ٸ&+
iBx� ��y�]e* As��҃3-�ć�;�y�fݞI\-z �n�#2
��zRR��ȓմIQ�E�;�J���b�<X��"L��Fc�hH��,U�r:~���S=���-�3R����d'��h�ȓ;�VM����t�*y!��r���ȓ1Dȳ�ǎ7SVɣfe�� XЄȓCn��:0����K-p�>h�ȓ0t�H֠H>(���%Î�Q�0���P��]�Rf�?%�,��2,[#���3��k� ЄGS0�dg� �jɅ�+K�ېdC�e��\*�H=Xt�	��sOH�7!G�޲�)���5w�>�����X�@n ���յHђa��c����Fg������8�
���3����5l�%Qv<Z�b٘0�E�ȓ3:���t$��*Ĵ| �eR;`���ȓ[��j�B5{S8�d�ضJҀІ������ZB[�M��)�6W-���ȓ�psF�C��J�
&�U9A����ZU�PJCz��A� 3 �~B�ɕm� �a"6F�����c�C�I�dׁ�s�h��)�ex�C�ɠj�(� �	�rh�E� \���lLb�i!Lo�ܸ[�O�
nq��])��A� Q��m��AI1(�ȓVPmJw��4~u��a�Ԁfn�� ̴�eA˻VS���<,	U��7Zx
т %*���+J1�]��S�? �=�e��pa��Bn9Y��x	�"O�w��2�<xƯ�/$�F�Y�"Of=Ac�J�!���o�u��4ؗ"O�a�tL^2,"��� C���;C"OR�/W�y�Ȼ���(I�Dp1�"OBAء�^�<���; χ�F	����"O�\�6��J�Ƞ�쐠 �!`�"O��F�؄R�f�B�kN�Q��,S�"O�i���+=~+�*_!n� m�"O2����tg�=J�¦w���z�"O��RDĘ
�z�����k)^!� "O�|�پ��v�?����"O|93cMR8�x���ՓA�
h��"O��S (V;*ط�θR�Z9��"O�4 Q�V1rƨ�5�����@"O��� �I'g;�)aD\�{�4�´"ORm#B L�7��m�"�N�x(`�"O|�I��+|��hX�G�Whp(�"OP4���Z�XZx$	U'I�{{R�ZE"O���2+�"zY�,�@�Thb.Q�5"O�ȱ��& �j�e�G3n��P�"O� I�iD�+F@	�#/�'��S"O
�QdL�B��1G�\�P�"Ox��?�lH����'G�V�@C"O���'0����َY���.��+ҧ2�"���H��*���1.:���ȓ9ߴ���,��P@A�Z�ʔ�ȓ/��b�>��A�Vb��5�ɇ�[d6�i�D։Mʅ
a��o����ȓKdhƽ/��}��mJbʂц�t�Zm��[���K�aOT(���u��"Z<7@1[��dT��ȓRM���L� U�U��Y�@��ȓ �IrVmI!L�Bu�BcB�<Uh�ȓ��ᙤ�5N���r�GN����ȓ(�r ���ϑ�PкR�.R����k<n��&@Ɖ5x�����6v���ȓT�.}{��'$	�@v���y!�O���'t&ʕ;~q.��V�^�`!�D˾<#�D��ƚ	X��p�B�~INB�xVQB�Kv f���L�5i�nO��=�~2#�]�h������&Jl�v�S�<���'p��a0�D	��be���V�<a�E�,�������C�\u떉Nz�'N?��jw���%�RҸ�᧣;D����
=�!��A�'m~M0�$9D����
��E�@�N�|<�ɒ"o4D��b��Y�nIJ8a�ʋ�x;ru$h-D���p۵=Aԩ(VbJ)�L����'D������dYfA�"
6킹1QC*�	F���'����o�M�\�֧�&^ �ȓ ����	�4fY2��JΆr~ ��C��+dm��ꄙ��~��DzR�~�`��- 4�5ƒ�[��#��o�<�a��A�Ā+�gU&"Zs��k�<��H�=�4���S�1͎���L�f�<1���S��,zW�B5Up}�
_�IY?��{������+.�*��L$y`���ybZ�Bi�!���z��W��y��:�B���B�~]�!�G�Q�yB`�;��Uj��Ćx��IJ�	��yR��!b� ��WD
�C�0��%�?�?��',|�:`"r�^UJc�P<���'�0aY"*�y�vZ)[9Nڲ���� �p�@{t�D�!a/~�����"O�]�d)B<)����b%@<=�Z"O��Z�'�X6%�q��=ZjԐA�IC�'�� �1��4���`�g��o��A�`�L���5+t�QILT'I�]�.ǖ��c���I�:1���c,T�>`�q�,��J����)扦/7N�Ǆ�_�񲳃� VV�ꓐp?��%#�Jt��¦p� �#�b\�'??UCefùw�x�BF�Q�3��Qp�I5�x�!�63Ҡ��D&�*��\�揄�yB'���i@Y+|	I@��tB��	2�މc��S%r~�!6 A )0B�I�!(,�3A 
vX��]�m��C�I�?�T�4���^�|�Zb�kʬC�ɚa~E�Q�� ��٪«O�{�FB�	�a����vFY7$x�Q��C)8�>B䉂k��	Zq�AH4u!!��&�>B�	�#� 髠@W�B�����V):B�I�mw�$��(]� �4��9{P:���2�ɮ����"�KU��� dh���fC�ɚD�zdY�H.C��1Z���
ZC�I�>.�"AM�5z�ƅjြV(�C���<Mk��E�ԥ�©�;4.\C�I�^I��%K
�zL+u��	:jB�		5F�1��N�;n�0X��:B�	A�+p)Z�{R콘'+��B�ɪ{+D���-V1Q���(���<PB�	�a`��4 B�j�u�#']+��B��[�ك �ğ9�����Ϡ&mZB�I:(F�H�&��<a}��2�N��6�@B�	�J:� fΗ^{$m�ӄͿ+�NC�#I���pT���LR"����U�hC�	�E&�(�T�ݒJ�����W�>C�I'j��@�ï�r�)b�%RO�C��6?�6��ԂH@<ÁF*;��C�3�*(j������J������B�	�RM�S
�Kn���ө!pSdB��JT�'��Vh�I( `Q(HyzC�I�0&��)
.l�a�g� `�RC�	
9�U���Y��p���� H0C�	5_ݨ��āG�(Q8��H�+`C�I�?�@ I����ɩ�F�fW�C䉟4[����ɓ[̐��È|�C䉢Z��D2�(<@�H�G��#n�B��1�Q�R��6U��PC�@,X�C�	�F|сGX6|����Ǉ�&d��ȓ�Dxe���jL�x�D�?�z9�ȓMO����{�8`%fε*|$I�� D�j�0���c���&a��%�ȓ�&!���'���h��G">Dj���sƾ���N�(_��

>,���h�mʦ ��%2�U�\"�`�ȓ�>�"�MZp�6�\�F���A<)����l|�8A��	]�>Y�ȓ}��͛�b�2c��8S'�!Gډ�ȓl�&�R���z �A(M��7p: �ȓil\������,���BW̗�L-:5�ȓa��yq�_"9��i�YO�&0�ȓM"xڣ�D	 {��p��Cx&��ȓ7��TC��-.�����H�}q$���j(�{Tc��|�\rS�ԏ�0��ȓ�r�Ô'	|�������\��ȓE�x��P*Q�
�,�p#e�-=J��ȓ'.~�����=��=PA�?;:���S�? FĒ��2���@��'�R4�c"Ov���nI�oJ(�d.	#7l)B"O�����$p�=�'��m��"O��B��Zu��a��-q.��"O������R�3 F�5��5
a"Otͨ0$G;|��ԸFeΏL �C"Op�X3�-X��U���5R�F�*�"O���*ؒ�!Eb)+��4"OP!HqKҤ1&�JP"�,=#꼋$"O���4d��#m���߃f�f0"O�h �KˣŮ��E���F�*]�2"O����,3`�L�g[���h�"O��`DI�d�n-�G�?|�ȭb`"O:L{��,6���ɑ�<	|�mre"O�2���� pD���Z-Qm�x��"O����||DA�CJc�� B"Ov5�Q�Ӆ���$�!���'"OPA2"+
�0�B�"��U�1��Q��"O�ёc n��(�k̸$�8�[�"O�LxW̞;y#z�+3��;��1H0"O�Z�i�'7Y��B�C%}'XȻ"OzUW���0ݞ%�EJ�]2A{�"OP�7,��(p*�d�%H�0Q@"ONE��M���ۢ�y₰��"O���T�J�f~���0t��9�"O@li���6�T@��X6>p��R�"O�!J`�/0�1�t�q]x�#"Or�fJ�G�T˒��+SΝx�"O�
��MR�*���IP���v"O�eX�G�c𭫇j�c4>�S�'�6yK�C�7_+�"�Z��ViH�'X��ʞ
�Hy�k�<X�����'�	bV�Ӹ 
�����' �8�'3ҙ:�-	�������}���'���Qb��J��x��_�p���'+$x��[�}�tl�1�܇�
�`
�'63Q�]0M����N���D��'��գ�.�`�9У�����'��\��d"uÕ?��u��'�����N-;���${Ì���'2,p��@�44�N
����'����X���`F	܌�� ��'cʩ�㢀!@ny�r
[x�$���']X@R�<�����E't"����'Q=���$թք�H�模���`�<�0�Y�y� @I�l@ +$��0��E�<��ጣG.��K�OA��b�HN�9����<-�Iv���<�AE`	J�����
^HAь��<)$A_j�� �T� �K�]O�<�G0X`,*7	CF����$D��k�덉o��P���&2�+��(D����@���=aí���:Y1W�$D��)�1�^0 ��j�\=��N/D� :�m��/�,8�žOZQ��-D�`v��%R�B���.�}I�+D���cF6l��dc����f�T��#�&D�����:}\
傣��b�<:A3D�$0ɞ}�.y�6��>C�m
��4D� T�28�fЈ&c+�Y�F0D��hVAC�H�ݫ��
3|���i$D�����\�-;`�G5���6�0D��Pf�P0v�@X�E���D"D�����X�(P�Y�y�n���d%D��1�\�-�clZ�B��$!D�� ,u�0!��,0���3)�& ��"OЭ��M��T����i��^7:��"O�m�!)�b���� %�)9T"O�A�Q�S�r��!����"OV��	�\Ԝa�g/�h|��#0"O���w�E��zh�䖲c�h�#"OF`QRS.�QsBđf�ب��"O�͘��%:\ [�B�=2�̸3�"O����Tx�f����xI��"O�a��D�@�80F-6i�T!�"Othy�A�l2���#{xE�"O�h�
���c7o��q["O(�����c7Թk��Jy�M�3"O�t1�����,�欇I�| ��"OL��0�.���C���J�"O��Sa �)8�diFo� �d��"O\��Q,�,5%N�Y��U(3�M�c"O��9�B���� (4͜;�ʅ�a"OrI2+˼z��ԌB�%�&|�"O��� cؗNJD�bW���, ��"O2%���أ_��8���2�pؙ�"O���(O�/(*�Y��K�"�vH��"O	�'�P%{:|��Y 2��"O�X��`Õ's�e����G.�P�"O�� R,��5�h�7m��x�"O� {@�@7C��	J�Z	V����"OV5�l%lP��V�	"A:��"O�(��@�*�)[�+
�:R�9XV"O�tK��X�5Ț��7 ȓZ�=��"Ov@���ܶ`� tɣ���Y��(D"O�@��" �F��d�G�)<h��
�"O`�a��@=b2�����/���9"O6E07(؃�|�Ao��k���hE"O�ň0i��6ز!�MH�v����"Opi*���rJ�S�+��!��QR'"O����	+�@C$)3>}BHb"O6�:b`B1$��ԙ��ǬRi��"O�$*Q�
�v�|�P`��m�("O�mHЌ�r �0�d�D���ȓ%��}*�~�N0r୞��ڄ��I�~�L4z�x2)O�{B��*���vqF��^�y�D�3lhcăvІ�Th�����!5�PvBa�$�Gy�M0��i���#���y��0Xsڙ0c��#p���#�� �^�ݴg�S#0p��3@#�`��Gz�����c+��:��9R�M���<�CkH;��	)r��C���A�h�.DH࢓+�0Y~a��==�l�j�d �;��M��ɬ�,!˃W� $�$!��+a��' J�Qr� S�P���\%f}��:c`D�'�6�
X:�N݇i��"(N�x��4�!�W�<�b	�JE���P� �b�D�b)K�r,���d
�0b�&��,��!�"Ix�DL	Q&q�w�>��+ �\��z���3z\��'�8��1�֭j�"`� ǖ�e��a�r�fp٢�NB�ud�x&�޷(��H;fV,i�,xڈ���p������*O�m0�eѾn�џ(h���p8��6��F��Q2�%��]t4��.]�6)��gM��)`%��H��=�u���=�tfq��p@A�Y����ӆ�Ty�a e��:P�ϙ"Z.�qQ�/-F ́���A%�����8-j,Hkq �C�:$j�"O�X۔b^~��	��Aߖ�������ٵτ>b�`�Po�R��}�f�'��I�|^�"�B��KRHM�-�����VbJ�IG�	n؟<����ِe�&M���jE�%j���ġ�ͺ�ti�,�P���!��"!(A0�×H� e�?I�2p�X"�קO~8�F\�'Nrl��KE�4�$E���7�8W$S7|�I$(��u��ȋ���Y��X�c�A�R�s�K�|����?�Ddz�D�*�f�1/�>Y���$�B]�գ�z�Q�V(��q($b	�];h��'����Ex������hC!r$@�R�"O��BQ�ب#v����3u��
,Κ�"`��	v�	3�A�:bT��Zq̸?A�-Y;
��1��w�HIX�#�N�A��I�P��S؟xc"/��� bmx���2l�r�D_�w-p�4"V�qP�	�Af�"H��BW"I)pE g��f��ð�S�z��I�\�b��6�Ew��ꦃ�eC,�@vb՚L��uh$gV!F�\�ÉF�.0��@Q�Q�v5"d/4>�`x���'���*]Red@�V����O@�
c� 4"��z��N��\PՎ��1<<8�b�C�N�Sc>�$�B��
,�)�p#�"U"O.@AV"�5�(=K )q}�!F(Cb.V�b�3�Ґ�f�(HI.��c�\�bK�%λ�h|چ��13��;A��3p�q��	�O͸�-�/R)����
��f2�@r�J�M��Bu���p�BV@C�%Ӥ��tM�,U&�"=�pK�d�5��eA,A�-��w�'Y�4�p��*x1��{j�u���I�M���2��\1t1ԏ�0�����
.R����$�L�ģg-B2���I���N7�I�j0�)�掰�\�J�'qC�ջ�CVc����(�JO����w��P nժ�"O�%��g��L?��SR.R�
�\*�I��Zs�����
>%�$�HѠ���OKqO��C���_���ZfN�
��@���'���ka/��-Ix=�b�)�Ƅ����:�tu�2�V�-���.`F���82aڠ�0@��CјHxTFƙ �џ�y�JL)e#��b�S&����Q�F<z](ə���_4$�%"OT\Y���B�d�C	P�r��Ԝ�x��'ȓ#�����iً)\�G�DȚ�?Wf��a�
�%]R���>�y(w�f�9�aU�&��s��
�x$X���B"jްv+�th���yҊ�3
�В�ٻH�ho��Px�ə	.��u#��֐���L�0�Da��`Ҩ_3���A-z�ԙƮ�߼ �X<(Z�Z�(9<O����)^�R�O����!�1�!�b�ӛ�F��"O�9p�G�yj���ԩ�D�x�@B�$�A�|$)
�'#�X�₃�)�
�2�"|v*��c� 3�7x̑z /�1��9�ȓ{	�IX�C�1@*��vhğK2����|���B�SL�E��IO�q��p��e\�]Q��ƺ}�f��� ��$v��ȓ	ѰyY�L��b�X�"��L�����c�x(�$O4N�2� �E�1����
���{D�7,dUC��@�7��݄�n*��C��N�D��c�5I�����38�Л�K�.Dn�!%�	>!5��X��R�\�L��ȱ#%�D20��ȓr��h
T^5/�偕 0}t��ȓ��ͫ�]7-���	�͕(=pp���$���:6qCƟ~}.���8b���G�9�@	9pf��N2r\��A��JZ��8|�`g;.�ȇ�g��"��ϫtdP#Q͝�%�ja��e���cɡ82���2 �-{����X*�x�̯i�n��7��0[ ��?$��A�A�<�Z䟲_�La�ȓ%}<���C�	C�ʌ��/-��)��N��⃈Ј")�5���[*��e��O����r��WF�X)T��e�֭�ȓT/4q�S�����e
͝Oݲ��ȓ/�Z��/�B�a !��nst݇����H�&�r A���z��9�ȓ$�=���Q'I�P9R��='�bلȓY�l2bJ(r�LU�(����)�� t޴ˇ���#ʔ���L�쥆�,, x;��A�e5�pK#�=�La�ȓ�fd��_L�^���B����ȓs�"%��PGޠ�wB�.ͅȓUb�K���DO�tr���
(Җ��ȓz��ե��8N(2d��d��Շ�="��JK~��YdA·SS�)��WƦ����t���(��� -�ȓni@cDE���Etޅ�ȓ�(��E)�!f���Y ��7T_X��ȓP�LB���@��b��Y��Xq��S�? ���$#�pi@Oߵ��G"O< 1��� S�	JR.ؓF����"O� ���"٣�͋�q�h|"�"Ob�i�i�`��͒��.F�ze1�"O��;Qj��I��!���R�n�E"ObQ�1lY�Ye����9V a�"O�t�!�9/�漣S-\��\�Q"O��c�*�7n"�J�G��ԉ�F"O�(:�֣���H����5��H�"O` Y�d�P�l��m�1�X�x"O��Hs��(Q.��eke��"�� N�<)]�P�&H8��q��J���ȓK?Z�"ȂiklM�W�(B��ȓ*x�`�ƛ5r$�k�-͒ ߴe�ȓ1��P�$��X�AS�ᏓN�\�ȓ�j!6Ӟ j��Y1����l��Gk�,)��5��2w��ȓCM(\Xpf�/Х�B&G/njԆ�ya6䱡�B�}D�d�()𮠆ȓ:��Z�Ꞣ�0���o�3J��a�ȓl��p �Q/�3H���P�ȓyv|�ء!����@2�؅{v�4��a>V��!U�a~@j�)�=.���|���3g��H��	�G�.Ʌȓl��XD�4g��R�ȃ6 �X�ȓ	5�)x�ʒ{U�}Zu捸ub�}��4Q����	(޾UkCd�����U��!y�LP8l�"O�.0|����.ld0t�T.�����X*e���Bْ���&�6c^����(k�ԅ�!�H��սFB�a�B�&{Q$��ȓD�4�a 
� �v�R�D�C�IV��T�D�]yؐh�֬H0EcC�	�xe�o��y��Ƚpt0B�	�.��a���U4o�4h8�Bƚ�B�I� J� ��_�e��!1؎C�I"h�t�ȳᒄ/���⭍r�C�PC\tzFUr�A��,E/�C�	�XxD���`$|��8���7R�C�	 2�Ȧf�U[��a�OP�^C�I-�.=����G��u��L&�B��Yta�'+*(����$$K7��B�	G��92JL�z��صDK�P��B��)7���c�!�鱤
�s5�B�ɼY�pɛ �,>r����� q9�B�@�Sg��8^�.���*AxB�MK@�3��Mee�e#�
	�6	
B�!z�ͳ�n��6�|��/�+�C�I-Dۊ՘Bw<r(KG��&(�C�	�V�ۓ��F0)���k>B䉢T�"e��NG�u���-J�u.B�Io�L8h}|�8�	H'o��C�ɫϒ�s�m�0c�H�Q��I	L1�C�	"z�F�k҃,4\ଡ�E5�C�	�!O�(U��@�!��
��Aa(B�	�P"hY�ב>h���T��C�	�uΎ�b�� T=s��5+��C�I*��Ur�˝OO�CuJ���C䉻��2�˴��u�Q,�_�C�I3{���q�۵	�	�(�M�C䉰)�&�"v�N0���ivvC�	>GB�� ���*���&��,C��28��3��k��i�6�1�C�I.c�xj�MLf�*\�V�U�6�B�)� Fi��,�7��8S��!E�6��"ON���o\6־� vO֊Q��\��"OP���_�P�Ƚ����C�u0A"O@��'[ w��A����j�c"OZY@֧\�/l �1� �g�!�"O0��gbې?:J�H�J�"��� "O��)��3Fl9 BB;m ��"O@8z��@\�����Ț�d	S"O-㍳m�lD���2����"O0�a�l
�:z8�����#J
��""O���3��X�@�'�E�VP�p"O�
Q������-ˈU	R"O���c��q�-	p%�kf�Jb"Oڽ��g�3荑$܉p�s"O@�#E]m���]�?DF�b�"O譛�Cz��ё! �z=��3�"O��
#��>b��/\9mN���"O�	�邰q5�8xP���u"8��"O�u[!
�K4�mp� {:�<"�"O��ciN����!-d/�9�B"Ox����P�Ro`�B���� ;Xh*�"OD�〬Ph@�3��]�u.&݉�"Oh0��E�33w��h�1X,X@;�"O�\Q�̋q�Qr&�.�8J�"O4�@`	�6\�ل�;+隙:r"O ix��PK��%��R���F"O���M�/��Q`�����1@"OA�$�J ����T�a���`"O Y��(H n:t�� ������"O�@R���M���)T)ML �"O���>>�f�#��]V*fi�S"O޸Q��M+yJ\q���<N
�2�"OƉ��h�H{
����"wr���"Oܥ�&�� ^q9�i�G��4"O4-�6JI e:%�1�� "O��#�D�5Q:���)�#&&^}"f"Oн�K@}UjE%��pl�"O��b	�\���J
�R�"OTaC���y����iF7f���C"O,��gFS�%�d,����2�`��"O�q@�*��C�H�r�T�"Op�R�JP��GD�M�F"O\x[b#]7!�5��P�H�D�:�"O0��"+�!���@��ˢ,�li��"OX�0�f �0Jt��KӓlJ��R"OH�0��;�8a)��PU��"Oҁ���߭LX̜Bh�]�<PQ�"O�lS%b`�j����]�@��t"O�#e&����	"$Ғn�ƴA�"Op���NKư��
c�:@�"O]@���b%�Ĺ�#F~B�5a"O!`���PX܀��֡T�(U�"OX��D�	�J�zUj �[F"O2)ٖH)8�p��$�KBj��g"O�����%>���$��TX���t"O<ѳ�@��~�Xg�Ѕ%��$��"O\|�d��=�8���<��$j#"O��*�A��a�)+�$�A�+P�y��PE��� ��"���)s�C��y� 
xi<A����S̶D�%A#�yMM�'��5��8�� P�H\"�y�ε�d���4��#��y��^�CVi�L�q8`v���yB�^��8dK�&h���ڟ�y
� ���%ͷr+agM^�E|���c"O���4gU,YD.DQE��3b��"�"O�ݹ��z�i*
�>A8@�"Or���7��d���C�1OflR�"O~m���̹'->l�i�"O�����ϕLK�hxŁ�|/rh��"OΈZf�[�=�zDY�j�4C��"O��ΐv)P�P��6M��<
q"OR��� �X�˅+��E	"O����lҋm��� C���n�<�R�"O�a����+���4L�[��ۤ"O�=��-�,�x0"'�Z )�L��"O6dYSdGz�r쁣�L�"��1"O���ƌ5������y�JP*�"O�1�"V�lQ�pI_���x"Op��3]0}θ��7	�@aЈQD"O�#�N��8��M�/׭=c�e�"O��"���/� �Z�cO%^X�"O`!�2g
P��1fAY
w"@��Q"Of���k������X$:P�$"O`EP�Yz&@B�	m#�la�"O�l�F˓�HH0ErUA	�#� b"OHUy����*2��hq��>%��[�"OD-����
3�X*��E��i�"Oha�@�׋<�.���.Pd8��"O8a�5�!RN,:��G�F�-�W"O:8�mݧf0����aY��8�"OTd���Ou�" �M�=��"Oʤ�� ʐ;��� �C*"��Aۂ"O���T@ �B�O4����6"O0�
�L3j����3,�:5P���@"ON)0�Gl*@��i57K�8�"OR��6f�.�h���=R|�1!"ODB�f�	L ���șE� �e"O�}�3(X#}2�pM�V�:QY�"Ou��/��<]Xe�06�9�"O !ZG�
�B�>m)�ɓl���jg"O6M�u��1_�X+��"(�.%X�"O��	��+�1a�7�8zV"Ol���Ɯ	<Z�H��J�X�20"OH�&NL�'�:�z�l�.D�"O����K�N�Pq�!�D"O>@1g�_bD����R�*���R"O������V||{f�ܯ�.�[�"OZ��U��~�n �#OV)�* +�"O<���	M��Xⶏ��>Dj"O  ��*�� ����	V�l�+	�'/�����V˂4x�痄#� y��' �����l�a
�+�Y�	�'�:�Ş�E�Z��f��O��Q	�'#؀H�l�R���fO�p��M��'o�=p�=�����5h�a�
�'M>P���#N�\8c'Ui�R�
�'Sxa��DZ����B��k����	�'�4 	TL��4� ��VY�H��	�'ݎ�a��b(R�#��U�258�'Q�{�D�<�V�s#�M�'6� ��'2��G��� [�p�B�ܜ|�q��'��L�B��8t-^��%"cF �
�'��L��J*~kR�`�,, �1�'����w̓4"ߦ'��2�X��'��Q�g���i��'��<��<s
�'�P�	��x��̱u�4�P
�'ʮ���-�6môTH��۽7����	��� ��W˒x�v ��é����"O��SrG\����� G� ���"O���UeL�p� ��EN_�@��"O^��#��.I4��'+L�O�nU�"O6%��E[��X��
_�=���;"O��aP�ݵ4/��;&h"w�L��"Ol����ר8���ϭt�P]��"O��K�S=(Hej��S*]�
�IF"Ol�g �*�0�WI�b0T@��"OHm�G/|nl�;���MY���"O��R���<�|e���"V" \)�"On@YQ�m���L�=#pl�"OP3m�>i<�sw�I�]��5�q"O���7!^
�q�J��oF 5�b"Ony8��U3tXj�Y�+�A��|[1"O��I՘nq�]*&�΃ZR��"O81ee���m�v��
�Fɻ`"O���!�/p*(x�-X1bƜ�(�"O�0;T� T,�z�fT"UX���"O�	��ո4&<(c��	�읻�"O*Y�g�h
q�9���P�<Q��"@60��mY�6����ARZ�<��n�dh�������*k.��QT�<��b�26�"����#Ƅ�G�U�<7�*Ȑ5��,�D؂���P�<Q�@�a9�4q1/�N󄵢t!�P�<�r�H�st�TӀL=A�zћ.�v�<��L�~*�岆�Ҹt���I�O�<1P/�y\t(2q(��*<�{5�F�<��.�3xQ�$�K�r\n�#��A�<Ic� � ��2�#Ǯղũ����<)��
fpT�s� <&z�qK�"Mt�<ڲX{���e�̾d�,tC7Ev�<���!)�~H:v勡G�d8��y�<�B!�5��M×E���Y�i�y�<Q�.��s�����̀Z��	Ū�R�<i�߹'��P�ɇ�(�n��V�<��χ.I��McJ���%H@z�<�j��M:�-��.%.l���w�<��9T�(��'AT�@��c�
^D�<�El�,e����rBΰ�J�BUG�<ѥ�ڌZ팭Aa
�$h�BFZ�<مaшZΘ�����2���N[�<�pG��)3؄��	�{,2P{�ARo�<i�V&#�,ak�B�9������i�<�1hZ�֐�Sɐ
�R�B�a�<A�
� ;�j<�F�؀&V:58��K�<�jX.�l�I:B�pʄ.�j�<�@�0"v��r���$�:M3�ώC�<)F�p�Z�Aq/N�7A���R��z�<ɒ?��K��ކ�E$�t�<a5Ň�,@��x�b���<`㉉w�<�f�S��0P�C��L��qRțK�<��L��l�H� W9r7������\�<a���|����h:M�b��'��A̓J�|���,^A�08��O�-N�8��'	��hK�+�Q���0IA��*� ᡒ|R�څ*a��S�e2F��ԅ�y� IS��F���y�"M[���0|r�ٜ����gJN8?�z4���Juy�Kߩ9������|��	�pU�D�f
ҹ)����U7B�m�"����'1\qxC!��������TlU>���"l��$����_M�T���'����6�'�x�S<Fi��}�"��j�����H�h ̀�k��~*�=�v/H�1���I���M��;Q 
ً3���m	�|X��ʄ.�����=8��d�UڮH�����������I��<<DXc��9N�`�a��:�f]���O�˓u+��}ʞO<RӅ ͘D2�q�F������{��@K���g�? �-�T��oT>�0��8m"�[��>�q�9�S��^��)0�Ӈ<qT{&��>���	�<�<E�TIQ�	ꜽ�R`� d[�4Z�W�[��%�\���O�8����?a*�I	nS�m�f��&c�`S��v�>-��?-��Hz�D�l���&>���D�	R<� 8���?E�`�����?)�c�O���CDM��TP���F�,����(K�:bb����3$���$B	qj��l���$�!��CE/{�&܀R"O��WC�)t/���p����ȕ1"O�ȱ2�Q3 ���U
;-XQ"O�t��g@�IO6EqF�J�s P�A"O��b1�M�bj~0iD
�/L�a"O�e��	(3���c��1���1a�	F�OƢM���,4D��q�<p���P	�'(�pe"��4�4y0	S@n���'b��g�S�'>=s���:��=k�'r�l��ݶD_vѡ4a��)y �S�'-h,
�#� OO���Ĉ��&�F%��'
��8'K�<� @۴jֵ�ReH�'��]#G��#'�,�`�:��D[
�'z֡z��d*�]��Ѩ.+��(�'�(����<�ʝ�ժU,)�0$��'ȦqU#��N����)#���'��A����VФk�ԧH�:4�'
hx,��_����瞯K���k�'%����Ò�,8�[��υLeĪ�'�m�KK91�]�����=��'�:����3���n�x����'���c%�AN�HK2��\p�Y�'��]R&���2���[" �Hh(�'�<���=1b^�#&c�#c���	�')x}�oM�?�У���*N6:���'bV��wk�Ht�4��h>H���'�ⅈu�ÃBz���$��3��+�'��8I ���!Aq�ȣ-�N ��'�� �nØm���Q��Ǥ����
�'e�
A��$W�
\�R,C�[>͈
�'�h�gI�"&ƅB��ǥ����'����W��p�j|P�hg�ё�'מ}� ���h�̈�ʁ�jP����'��	`A��:�H;珁�5���'�����.�w��%��e��1Gzm{�'�U!�$�wߚ�a�+!\����'p�AE���4TD�_��!��'9n����K)�2���1w��(�'����ĤʅT�R���g^��5��'`�,�U ��PH�M�6��V %��'5��
a)��%b�Cz���'�JI�&)��(��ٷ|�.Y�'�6\QF�H=e�$i&�P�_�B53�'��%�BO�O�ʨ�Ԯ�1%'^)��'8��s@��R�x�J͇'J ��'@��93��k*��R�CJ�Mu(�y�'� d�H���3�C� t� ��'��-��-�;������$4��uI�'��\�5��#N��K$�
1F���	�'��LPO�-`!�D���� 	�'Q0=J&�ޯ;1�L����ސ�:�'A�d
[!:�0y�RxI�L��'����� �C��I��fSe|��Q�'��H"�Bٛ+_� qF�"]3����'Y�)bڮ+!vYǦ��O�N�;
�''L4[S�]���p�3*:L�<���'|��0��~���1Fh�&&Y��&��� �n�&dg�-�GD�5ID�p��S�? p O[!q<���-��l��\[�"O�)#c��$p�@��C��V�V�QS"OH�X�	�$���8i�bui�"OJ�಩�<:-L�k - +��{�"O�܋������0�W�8��D�3"OBЫR��%pHQb�J��|S5"O&����-4Bh�l��a�T�2"O��'�&B��Į/eٸ9�"OH�@�V�(&��r��r��`��"OPMCd'Z#���yu���k���2�"O (
��)�`�a�R�|l��v"Od�t%˂.����[�y�8��"O�TK�Ń�\�l1�����: ���&"O�@`�/�0(��� ` �n�2Y��"O��Y���ek5rD�_�>,��"O@ՙ�&-zȾQ���U$|�f��"O�|sr&�O�ʠ:W��8Z%"Of䁢N�
& D#DF�f8	�"OtU!$0T� ��#�->Y!�"O�I����b�|����Q�D��`P�"O�@��eS�9����̐��"O������DH!j 2�0�%"O����%�h.�v�����f"Oj�j�=%r,tX�M0s��lb�"Onl&�p�@��z��-�D"Bc�!�H=u��(�V3o��Ɂ���t�!�DܿZ  �T䓽_<�A�ˢ�!�_�n� 	OY\Jբdk�J�!�d�J����,Z���@�!�!򄔬q"����̌S@0(f*J �!�$9�b@aݸF��{�)�0hU!�d�0	��e Tk8s�.���/^!�Dʌ�RM Ϛ4�:��E!�dƚA�rl�� �"S❡A�G�=!�d�(&ą��Z~.���cbT�3!�I�Q�$N�)�ɧ`ܻ_(!�$��Pn�����X)�a�68!�D]=,RI��X-�~Qx�Q�!���ya Ey!���,{�( �i�!��J%]L�&�O�4�j[v���w�!�d�,+���EQt�$� �B(r�!�:#���JI��3�0 V �n�!�� O��m���W�5&�`cR Q�}�!���L5<�y�ɛ�O!>y#¯L�%1!�d���p��5��f�S
 !��Гp�T(��[��@��C!�dT�[��h�a�\.$�����	X�!���p��pˤѷ'����O"6�!�zɮ�Y"��&>�����d۶q!���i���Y&f̘ܨ|"�B\;!��1^X<8��|ӎ(�=x��;@����*̄R��¥Ln�DQ�ȓqY���0dL,8������=��X��2������N���e;Gi�2@>І�L���鳍��@� �퍯V����Bx�cըi2��gK�- f��ȓ� )�D%
�g�P�*��_�Eؕ��x��L�5滑�b퇸�$��ȓF��1ū�1@��̛��U3L���CM����^=4܋�P�JlnU�ȓ ������ۚh^$E(3Ŷt�68��^���в�ަwE�H�5)X���]X�0Pu���\�|�X�e4y�	�ȓ`۴� �`ˠ{: �CDѴ.��%��S�? l,����mHA����3_����"O.4�a�P<+~�уCG�0Y�h�"O~q0b�|p��3�G'=tb"O�P�ԅ�"��Q�el�2Xr�5�b"O����J&VP�%�&�V�P�"O )�بD�1R'�@.��C"O�4��.F���i�&: �$��"OB�7��%k�EQe��<5�PAu"O��9�n\�M���拵&��XD"O�a��=���"���0}y0"O8!K���YV E�%&�"|��"O6���(	�ld�`J���x��5"O��R��I����m� /���Z�"Oj�c��ڸ0�ٳCl����e"O�c��˴H0���D��'�ir"O�P&h�'/"�t+��U�L�@"O�5�d%��P����dCҘr�}�2"Ol���HF�M+F�s��в2�|�V"O�TA�ԕ�f�h�j�4)��,��"O�E2u�5 ���nۊ�*�"OV ����W�Bu����0%ͬH"Oh�1��оe����"2)��ʲ"O2����#u��%�(�l��""OPq)�/��zD�k��W�$x�"O$Y�`��3��2��\�p�x�"OZ8����8T�$+Da�/��Ѹt"O���\li��d k�j�["O�HK��B5�����ݲlkB�Y�"O�Xz$�ޱB�=+���06g�DI�"O�,J��	Q{b|��%eLJ��2"O�=a�U�V�P����Z kI`TQ�"O�!�t�M=h��48��'7��Pe"OF�h���&LdF�B�G+.H�W"O ���[/�����y���1"O�-[T�J�-ku`���-��2T"O��+q�I&t��Tk��O:(��� "O�ٲ�?k��L��i��p�0�b�"OH!�bǡy(��I�߶G�^���"O��avH�8d4˵FH-{cޤ�"O����M�Q�H��Rd��	V"O||0&,oc.���=[�
"O8���-F�X�ڕ� �Є@4" y�"O:�S��!J~�aw	�J��9j!"O�j&�
��Pq�ш��=7"OvyBՎ#V�6���
Yu�!K�"O@����ժ2<>��Ǚ:N3�"O���n�"���GF��?<�$ӷ"O�|z$	�3<֘]{�d�8n�`�"OL5ƀ�8�"�a� �N)�"OR|��+Z��ĄO��"""O�P8w��u�:������L��iU"O|��`ߙ�ıaǂ�/	��r�"O@�k�ى9��0 �%G�@	Q"OX�����UkdsV�Q�c8,8�"ObT�H'`\,�P�̾�	c"O����*-����]���0"Op��6$	��̃��  �`	"O��񰩜�2|:�)C��7Bօ�U"O��@�>$�}�����h�^��6"O6@"I-=�,��`�3Q��\:�"O
`�!�F8�d��	69��AG"O$���%kg���A�֑R-z5�1"O
%��o���X���!5p���"O�58W*Y�5�xȖHH�eH �v"O� �A�1a���H��bi�3�E�G"O�3��R�6i�3�&N�`�#@"O�y��>���ڏ"j�`�V"Oh���#ƺ]���c��U!p����"O�@4n��2�� �5k�+�"O��T��D"��Q��Ӕ"Om)%��.��'��0lnx�"O���,�!�.HR��Ę�`r"O��STo�6l<XSG�J��Q*�"O��� ��]���fT6U��y�"O�}��H��qz��˕�Q!U��"O
D�Ңd�����@�t&�bG"Oδ�V)tu���&���5D*��u"Oj��A������d4@�A�"OX�b�m�"K.�0p�@�2q��0A"O����	;rkFDhC f^"3"O�tӶa��"���Ф��f1.�x�"O��
P�0cx�x�B�l�I�"O8�R�Q-e= �
d�X�'�Y�&"O�4[��X|G�� �`��{�H��"Oؑ[    ��   �  Z  �  O  �*  �2  �:  �@  CG  �M  �S  Z  O`  �f  �l  s  gy  �  �  D�  ��  ̘  �  R�  ë  �  ��  1�  s�  ��  ��  =�  ��  ��  �  R�   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6�F{��'O��V���&�;�+0:��x	�'%��"J�[�]�R�K2r��"
�'Oe#W烹�R}aC��z��
�'��;��7�������L	�'�:<*b&K"4����M����9	�'نx!c̓>�D �,ݻ2zX�R�'��@ �F�9<�m�7I�"+�a�'ր����>��Y�
�%&���'��0��3L�r5��M/� HJ�'U����J08fx����I$p:<���'6�D�)n�N]	0��K'~8K�㊵�yŬJ�Da3gǋD|H����פ�y"*@-0NPI�-@�=�D@f���y2-ݘ;������H����u�O���ޗd���)�S0L!��҇���Y�� 9b����2?qEԁ#�]1Ѕ�'?/�tzV��J̓��=iWɋ'Z��(���Z�:H�p��P�'a��G�ԧ��/:9��ƌM.��s�B<tK&C�I�:��%�
T�6P�� L-4\.C�I�p�̫���? t�t�c�ǩE^�B�*<I�u�Մ<���y��U�B�	�x��9��d�to�H���"O.k)�g��
�K�ws0a��"Ot��A��z���� �L0!\ ���"O�=V C�j�Ԙ+ף�%y$�(��"O��6J��r3lL�T�;( ��C"O� ι�s(�I� ��%7]r�X�"Od���#d�P�0eղ&����"O*�0�=K�����?
�K4"O����i�&'$fx��/|���"O�xJ��P)�|��@4$�Z�A�"O2	����6�~��󨓖�	"�i�����}P2lq���-��թ��D�a{���X;0���!Q�ANkJ��6ʆ�:�!�$�0A��<����0S�"O=��*�O�5��+P���b�)C�:\M�Q"OX�����
����7��� �tų"O*-�t����u(�&��M�r��`�F����	W4E��ɂx�Q�r��;.�!���0%>t{��E=V���_AS!�H�x������#v��A���&=r!�$�,L��Pr�����ǲg�!�J$�}��関�\<1�Y�\��{�8O���T�v�l�l9(dBQ=D�X�ȓ7��XN�Z�Y� !�!&`��~������*��z$@�ú���'�� ХK�)H`���
�}�Ts㓱�}T	��͏�ufd1jK��t�ȓ5�Uc��t�LD�B��5/T�ȓ
Ԍ�UmǁCN�I4F��z�Tć�2���cvF��Jx�PP�Z&L�\���t�N�³!�7(�0H�eȞ ����ȓ �|�H�E�?/ƚ� �*�P��5T�S ��j�@	[�bR�d4�ȓC�&$�GG<Tę��+A�
�hT��k�t�V�,�����E)J��'O�}b�C%'!�0ɥO`��� ۢ�y���Ct�CӬd����6L/�O���7.` �`#,b�=KԢ�(4Q�E{*����ȁ,n�ae�8k"4��"O��5�!��:�c��^'��%�'�qOtҧ�& T�q ���2`���"O���q쓟+�y�pA����D"O,!��f[={z�e
�<Ş��g"O���D��W���"��L@��"O�y��M��,Zt���o
б"O\m��였�H��X"&��R�"ON���)�'܈�q$�؆/�p<KG"OpW��g̜]ȶ�N���#�"O�LQ`F�2~9z�0w��'r�>Dp#"O�`�FҐD�شS�a]�Qj�)�"O��x��(�zk��11��i�r"OM����W��C���
AP)��"O�@���)*� ��`F�8D耳C"O"��P䜆L*fA��c30��"O kJL�Y	>��3��%��"O8a�f�Ԑq���Yk��+�"Ob��EւY!�tb�&� &i�X�q"O*���Z�I�|�YU2.�"O\QȢ)Y�HaB
T2�|7"O�2�J�yH�d� ��;tP0Q�"O�����t�Z�Pq��&fX�L�"OݨD�6,��a���ܭ�8U2w"O.�#��M�Y4�����i��0B"O���c,V����"���*��H�"Oh��GAߥ<�X]�vA��AJ\`�V"O*u1)\W��BV�9kH^�+ "OD����{?fa��
+X3^��W"O̳
�:r^9��`ߝj��x�"O��z��F��٨g@F;%�f��v"O� �]g��,$	�n�4)t�"OL=r��o�9��L�t�)�"O"��#	��(��K�u���C�"O�5AKE�@Iq��Ө���"O��w��3,�r�qt%ݹzr����"OH�RNZu�t�k��rZ I˵"O���f�N�W��%;7�C�s�2���"OP�e�(,9.�B�M.u�Ģ�"O��2u��-@�910Mۤ|����"Oh�dhE1qB��ӰKp
��"O~0�7#\+d�hՐ�+�)m� �!"O ])��T&,�y�!��Jk�8�"O�t"���܌�p2��R���9�"O8AJ�"��G�|`�m	�fK��"O�)�ğ8f�E�"Ӣ3d��"O�0����S��ݣGjl.�{Q"O2�іJ_+^"d�U*:Qi�8 6"O�@Ã��7n��]�@Y�9ɴ�3d"O��Zv��d�ة��*Q�Zt�F"OxP����U7��e�]���00"O��I�I�QI�e�#�Q��X��"O.tpw,Ƕ��l��L;g7P��E"O�E[����-�f}"�lR,4rM�'"O����#>/�� :�I2�	&"OP�F�P\��p�O����"O6}C��WPA�tL�'	���"O�$j3ꑙt�h��!'� b�"O��U��1e����o܂3�����"Ob�� ,CIJT�C�*�l�I6"O.mH� 1n���,�ļ)�"O.07�./�ڑA"+�Y��!�G"Ot<�sh�������KԹ~����D"OJ��Äc��I�� /��)�"O"i���X<� ��-',A� "O�d����5*�p�NR�$@�:�"O�P��id��]��cї&�!�"OP�p��@$�	�!�I��L�"O>B�m��P��=gcD,y��E"O�P�/	�Xj���$'[��@�"O�=���uی ����l	�z�"Or�u� P�Z�!u��^�X��2"O�0���k��J�GVO>��J�"O5�e�,X�I��H�9{9R���"O����Ι�*�fIg!-=�iZ�"O�`I��^�@���	f$%���&"O2Y�Ј� ��Rc��3cT���A"O�\)��|�
��dݝ>E � w"O���� �wdƤ35c��T7bm�"O\%P��P&���!�ȟ�k5����"Ob��tԓ*����f� F�h5b"O�@�4)Fj9���[�G�.��"OP:������j���7�m�G"OF�`� �d�6�sg�)ǘ��"O&zf���J�J)ÈR.fަU��"O���hфN^I*��[�1ͮ�h�"O
�2DZ�2^4y��̫-�&��"O"	�VA�~(¤Q7������p"O �o�K9x���댧{���8E"Ot����Ʌ;S�����d�|��"Ou;@ǌ�r���`��Ii<��"O\`�
^v��A`�VQ���"OV�R�ǊTT~�I�N�L�i�"OB���	v���CHM����"OʠP.̯V �w R>6�R�"O� N�s��+>�؄9��KX��0Sr"Ot���99�0�!^*$�X�Zs"O��a�&�� _���i�\��"O���w/?Rf���V���Py1C"O�P�qIX�`zXb�O�2l�H@��'�������柴�IП��	џ���(&.fH��+ղ3��Ͳv��;�jA�	����I�T�����	��l��ԟ`���P�1Q��B����ce�? ��M��ӟd������	ٟt�	�P����d�	L��  d�8X�A�è'ps4E��ǟ���ҟd��՟h�	�����l�I�w�nEC� �RH��0E�*����������<�Iퟬ��ß\�	П��	�L��ֆŅ�Ե�WהF�%��۟(��ݟX��㟬�I����I֟�	���@
e΁y�|�[�n��~������I����	П��I̟P�	��4�I(Ezx�A+!���	�JX�`e�	�	ǟ���ݟ�I�d������ ��� ���㕀Z�Ap��5)�`�H\������I��4�	ğ���P��Пt�	+�ֽ�5�
�X��J��NY��'��'���'�R�'+��'�b�'�@0$F�?-�`ia$J��2%Q��']��'�B�'���'�B�'�b�'S��E�U���Җ&�b�P8se�'���'r��'1��'���'���'�,:�	�4��Q��n������'�2�'�'���' ,u�j�D�O��A0�+2�����H�\ P4�%�_y��'�)�3?�r�i ��+��V����V���٨��Ě�]�	L�i>�	��M��B�$�zlBt�P DTDx0� �{k���'U ��������ΠN��=z�O����
-;���`A�pX�{�͟�~r�c� ��cy���%熹p �T�6VP�e@�n���4.��<����d��E"Q���2թ�c�F���-����!n��MC�'��)�S5C��Q�Cd�h���#����7 �8yӰ%�%&o�9�$�|	 ��'R�����'"� ��;�E�4��9Ӹ C�'�P�	�M˶�
f�6!��� T�����	H|��h�b��>��i��7�e���'T�����;@X�a��%6ѩ�O"��g���]�0*���Xg�(����O@d�c%I*�ⱠR�Ѱ|J�,�U"�<�/O���s�$HC䂳.��%!$����n�KJ}��ڴ<�
��'��6�=�i>�PgO�=�@Y;t�7HD�qB�Fn�0��4����'���!d�=��$$r�����Sb�L0`�<�f��r؇�L|�p%,�$�<ͧ�?����?A���?�2G�/�V4�5LX�u�� b	����D����'�i����ԟ���z��'𠂴.K�]�,����$��!*�>y�܏(�, ��'c�O����Oq
 jVe΅ �	�q�ǭ�Bd A���)Zx���'a~��a(D�n�f�YAB΅O&"�Oru�/O��y1�Z-%˼�"�M�D9� ��O��d�O����O�	�<1c�iTn�z�'�JchR��}�4#ʞH��(�'>7-�Od�OM�'�27����K�48����Q&,>~�w��ZH�{A�ݖ&}]�aDi���M��y	"kB&�?9�'xH
���2�s�	>v\���ɀ�4.ak5O���On�$�OP��O>�?=#��)��*�M.B�T8�t�k���	�p�ܴ�b@�'x6m�O|ʓyE�K��ļS�6t	3�="���pg�'��I��M��i���ҷI�rm��'�v��᪈+ o��;b�N;'>vXp�'F2lQ�i�bЍt�q2�'Y�	��D�O��d�OB�dL�/�p��) �򅓽�����Oj�_雖�_>�yB�'��Y>�C���p6�؀r� ��YU�6?�T���ߴߛ�o�O����i��H�"4��,T�!u��}�j����2Nܚ�i�<y��t���y�&��+`āvⅫ�}aQ@Ԃ4�p=����?a��?��Ş��$ͦ�R���"��`��/�>�\S���ʠ�Qe����_}�j��(Æ�-����"�v�3��)S5��m��M;䪚��5��?�T�1�Z��%�̀��y��P�C;yD8,u�� �$�<����?I���?)���?�*�DpAB�O>'�֕b'$�'B�2�z��Ц1���t����ş�$?��+�M�;BT:��kĎpd�d�KD�<�#b�i�7�ٟTק���O���CD�4xy��'&(q!��$N/ze��̯v���'Sp�Hf�֙U�̐h�|B\���	��r'�G�@��}�GX!��[���Iɟ���y�sӪL��<O����O����#=�^���K#_�$0c�8�	4��$Yۦ���4(C2Q�l`n��o�u���۴�lzW`c���-KxQ�D.t�*�'���'��0����'d��V�Ym@YX�jF�(Z��iW�'���'���'+�>M�����s��Q�}�
������ɷ�M+�o	B~��y���]6�P��P	�x�/�<(���I��M׵i\Z6�؛d��\�f:O���F�.2dAE��&(Jpxc�%O�x11LʟE\B�1 '��<���?���?����?��n��0�Y�w]��,�R�����d榭"@�h����۟�'?�I%S��(唛\_.!����،�O\io2�M�B�'�O6���O�Fp�bJ�a� d�3��:F��5��,��2�=k�Y�(�"L�1��V�&��'#剿L��y��C���<R@��J}�Iџ������i>��'�j7�?��Z?e�6��5�ʺg��e�$V��dTʦu�?� S��ڴ5ě��ӄD��e\'/!�"g$_)?0ze��!ʓX�p��:O���Z&MRa0�ܦb!>��"��� ��$cW#'+��YɵyD̡�?Ot�D�O����O`���O��?� � Q�`N ���E>fOP��Cn��I�@�޴'�.��'16m;���4t�4����G)'�:�&��	XgD�	j}�ebӚ�m��?ѐ+RN��	ٟܘ^j�j��ş0��CK��e!�]�kģipT��w2�D�<����?����?q$G1��ܺoƬ���Q���?	������}�C�l���I�OW��H"j�<etV�c�
ؚ����O���'�l6�Ʀ����ħ�R�$��]<�PlK�����ꏹTJ�-X6��J�2+O*�iǃ���/�?]S�ys`9O<���-K$�#b��Z%R�p�"O|}Q0H�1K����`�
���%�	�)�**��B]~\X�B��WM2\:1�@�-k�ѱ
D6�Xd�0���pDx�E�4spG�o�{��E�3��3O,9��Ċ���1׀�al�hs2us %@qޠp��
(�n�+w�U,'+� �Tf�� �!D)���e�p0Y�(��`��%������	.dP��3g	�kQrP$����ʟ��I_��ʟ$r��'q����-��U���&ʛ���	ş<�	��`������Oh�$��mc>�@��3+�����R  �jU�)�>a���?Q����?YS��a��ȔV�r{u�	�Kʘ��� I��d�O����O��/�	�E���U��	`���8����FE�{��6��O��1���Oę�`�O��D�O�,������F�c�b��oi#֦}��ßH�	ݟp��kB��ħ�?��J�lz�i\&`���p�!Y�:Z���x��'t�៳p�'F�~�BI��c|�p1�@�r�������צm��ϟ�J�H$�M�U?��I�?���O� ���d�d<��a�1�l��S� �	�4"���?��g�I�/:X�$R����g�
=O6M��^� )o������ӟX����'W:y�/I�
�ܠ��Щ\(t\�#�~Ӿ�`B�)�'�?��G�B�rE:@�
%io2��`H;֛��'2�'n�G�:�4����OT�;�@�)9��;�ə`;<L�o�c�M�<����?���f�aÇG�9g���ȁ|q��
׹i�+G��O��$�Oh�Ok��iC��y�헥H[R���D
	q���'�"�S��'~B�'�r�'�����6��uh��v��-�X�+�	+ؔ�AO<���?���䓣?Y�f��:P�����FW��r$�GV��<a��?y����DM�*2���'C��ȉ�e�4���x�K
:L����'R�'P"U�8�	���lZߟ4�c#Y" ��(PN�"� l�F��+��d�O��d�<A��a��+�j�$�-�ޑ �K+�>p����)|n�k���?9��e90�H>yE�R)=�p��Rl�w�8����ae���'t�����?U{�S�����?�ذ0 ��rI�2,{b	��`��MݒO���O8��W%&��!�DQ�+\�1 0��H��B���M(O؀������`������L��'K� Xd���"m�1;1��q��D�ٴ�?���LX>����3�O��TS>7��'� ����E�S� Ac��g2��J�>PF�6m�O��d�O�ɕS�i>1iG!N}f�I�2+
�g^QQ���M@ǹ�?����?�����(���O����t"j��,�	S+�æ��Iҟ���	btEbH<ͧ�?���P��I���}�ǦB;��i�"�'���;���<���?���oZ���"�8U�JxJ`��)Ռ�j�i;�`ǓH�O���OēOp��@�X
*Ȟ�P!N��|����ׇHz}�A�3w�2��PqA,P�Q&n�k�� ��3)�6,��'���a�K#a�j���X5lS�l!���G��%"v��+Jw�a��e�{�����S��l�gO�OƤ�ǣ*@p���T��-n�lP[t�O�u ��D� �PC�J	�{k�D�4|$ P���=A�Q��'dܐ`���۱+��q2��
��)↌
�q7�M�U1P�59���?U�X���Ŗ���L ���0�1��N���k�9*<�XQ��'��'�8�ᄅ�,�����@�H}*�(�Ҁ��8<B��׊"�����剟\�8ӱ#rBD����"B�p��(��%0�E*đ�(O@9��'�B�'"Z>qD
��EQ��j�_Ğ�Y$�ӟ�?E��'�nIi���8Y��Q(�\F�M����'��5 ���0��H�Uʗ�U�̓J���Rq�i�2�'Q哄5,��	����IE?����.Ƚh\Zt���=�l�A���7C���#~~*��c>��6F �C�@�.iM�fԼ��`B2"� +�Y��=?E��c��;2��/Z�@�6#Uh�!2�=�?!B�i(r��?}E���*�d-"��X�DTL�õ�ыy����?��Cz�)�#�H8����(�xDx��(ғ����Y!�:�B�,Æc&d�i�O��dT/׾9�s��OX���Of�d�F��'�d�ɖ@	�8��9���=bLl��'�uR�`�)y�u�D7O`�bB
v@Hٔ��&p������O�ԡ �ƦL��U��}8����lָ��d�2u:�T��C�¶aM˟���ϟ��<����D��{,IXd.�=z�٣� �.)c!�ЀWY�D�^b2�
��Ͱ%�^�;��?��z���Ӽ�G�h2���4,���XA.C�I7Ut����f� 5.T"�'Y><�VC�)� z�Iu`қe�ޘ
��O���h�"O,��G�-�(�3π�
��I��"O��x��}s�-R'��)���1"O�@9���(3�*�`P��s""O�p� �uZZ�P��V�-��"O���䭏�>py�.V�
�Zta�"OX[�%=$�s%g�%H{D"Of�2�Q�~�`(�&�0)�V���"O2�)P��	,�`��M��"O�ppأH�M�43�"��"O�<��1nm"h���U�&&�m�e"O:�ӱ�1f]1��,Ǡ}����"Or<�r�բi�"���a�%9�p��w"O%�Q�M#4�2q�C�?Ό3"O�Xj�0h��1�9d/�͉%"O�����~�蓲
3��%��"O��*5'ԳU�d�giZ�vζm@a"O:X Z����'-x!�S"O&}p�!�'�
�PF�Q-T!�"O�9�l)M��d��Q+|ó"O|D��/�ZL��nHp����a"O����F�hh���n�?Y"���&"OB�%LC�L߈�zVn�+%���r"Oz�1TAאW�0�LMl��&"O��E�P?h�R��q�R��ര"Oj�n�-MbBicf@�;�E!�"O��Pv-B�cԢm2⌜�	�N�"O��m��q����l��]�R��"O^�s`@Ʊl,�y a�Iq�n�q�"O|�s�J_�E��ClS�\�~5��"O�lh�)D�%g4eła�� C"O�3�@��L������]8�"O ��1�]����S��2Gt�l�1"O�k3�P9eؖdj�)
$]���q�O�(��,#�)ڧjEf	��ưw��z7hݔb`*��ȓ #�!�M�Ѧ���dԓOEܕ�'~�Lу��H���A�l,���q-O%Y"T���%�O*|Z�*�HJ
��	R�5͠�H�Ņ�yd*(R#"O,�I��B=�*�{`��/�mq`�|	rQ���
L��Xp�G�X&.\Ѕ*_"d B�	�qHp�e�X:Mc�4h�\�J�!G�f����d���$�<)P���;z{�EX�@օls��5炏}"��:��D��՗ �*�*G�֎LȄ��Qy�)�� ��_"}�yh�-Б�(O:��f,� d岝)�'�NN��"�'y!)��\���qpFN�0]�m1�f��ni3!.��n��]�d��2_���ri�Sb���#P��!������1J�����V�4��k�Q�h��r:����S)G�F,�5
õtY�% };.B�I<��YR�g2'���K(R�!�c�u� pT��?��CB�R�)hZh�8��F�!�츢7�F�K�2C�		(�hȪ�Ř._�N�k �v�y��!?�A%�j��8���#u���.� |�I���X��E9ң��%�Ɲ��,e�� �&ڱ^U�,�2�0^4$�3�O� f p�D,G�"�a'�x�	b
G D�|�\ <���ڶ�\�Kb�a�0�߾��d[�8Ľ��i��=?���냊����DO�(� �f�*����'���y�N�[n4s�o�˒��r[h�|��
Y'8��=�OK���v爎�y'�A�������1��x"�Q�E��`R�Vў�:������BךtK7#,z�����Ӱ7��<P
ID�x��T�s����DQr��J&"ջ\'z�i��%@J�	�e�H�vo&Iu³-��D�S�Ը!wV`���'7��Q�0b���
�9�D��Oʰ���S��\�N����W�@��|"�&��*�F���@�xE�e�3ANd�<��o��W�ӥ��W
$�W_}����-zty���>YN?��T(�`8�睋;�ڭ�/�uɶq떭½M#�C���{ ��w%W�@\rS!�%�p��(Ppg0Pp��W�R�Z�S��g��� pB�l��C�H���=�a�2�	�	F� �O�L�/h�@�c�7��l�� Ӎ<�3�J�>)plEn�퉯(����mW:�����V��fi��A<�)� �"&+|�"D� t� ���e�`�d�R<�Py�+ޭ~�� ��M�N^,J2ߙ�ē*���Z�l�s�zĹ��Ž��S����#�R<����18)�	S�k����?1t��J�P��ѢE�ά˂l�*5:R�!�U�q�,X��ܚ��S��Mk c��P#�ܲ@�U�w���X&aZ}�'�&�U�e��*u�MR�C��`Pa�_�&�$x�'����*C|�z2♀*Vt�ԯ���8	�ME�����>e��{ʟ��Ӣ�ÓQO}��J��:ӎ�!��Ve҅%_o�<	TŴ*�|��䭝�A�Qb%�M�I��)���'ꡚR�'�D�+���@�	=t��$n%q��A�0��"ٰ?Y ��<i�V�Qk�e��$juMT�� H���O�-�a.AK�dE�P5��?牰3�2�kf�R	@wP��9r�#?ɒ�MKJ��� ��S(<���/i�>�O� l�Q�^ h�R�Ñ�p=�碂�I't]#�V	}q���X_}��
�`4J�G�SM�T?�	7#�个�$F=QM�ca�O5q��C�:�!�D����q3�	c�A#3�I'8���'F�ŁBn��<��?�����#B�����V�Υ9�K�'rG����<$QҀzI���5v�F���JV?ѷ@Rw��51 ����'󞙩 �ә��E�͘%Y������0�2٨)(�ӱ/]�0B$G�j�N�ȃ`�\���	y
�Q�rjW~؞d(V.��!K�СJ��I-?A�Ɓ���'D%Mڠ.�Oڥ)�)�"u&%KG�� {����3"O� ���p"1�@!��Q�&q��A����)�O�qO�S41#�L��Oo�xŎNI4&��,�5o���0��?� z���}��\����$ ��S�䀭qz"�'���+���!c�E ��E���Ց���լ0��� N�c�������0<!�@�$0R,ѓ��=>H����bF�PyS�L�m� p��B�uiH�������7��=I��g�ԡ�$��D�|�C�Zg~BmY'	��
��L�i`��������!IN�YTz}��3'�9pUd�<�n�(/Ha«����-�`kW�!k�����a<�I�=�O� �Y��Ǝ�y��Ҳndf@�AgH�f(��E_2�x��.J��@�d�o���(��k��yk���t̆(�b�D6���J��{��3�.]	P@���r"(O�@y��<��<e2͘��Ҟ;����BhC/�h�����j(�$��.��{��� ����w�DU�7�K�0����N�'��D��tHdqQ%j�)JH4�U�,
}hq�ȓG� ��!G	�v.
q�A���"E��P�TE���Bx�f��g>?T���o08��C-V�L�u�ZP���=�2� 2�M?(Z�y*E`����[���M���ۀAIG�2��ȓ\0&�k��u<�+%gO��e�ȓl��<oK�I���5�2^�n!�ȓC��I[�E�q$�jҠ��C�b܆��fp�� K�b���$��Ć�Wm�]�ChHb�� ���/ZxD��hcb��3@�QC�d�u,�/��؆���ՙ&��~��tSB�� )��܇�`p25�pc�-&^�;��#5DՇȓ_�`�P��x��5��!J�rm4ćȓtn}�1-?YG�͢��_%W����D$�+E�.U葊��Ȣ����Ya��;�Ct��5B��	�&��؆ȓ@�T�Q�-̆�a�_���9�ȓ=��L	���v�l�j$��*�XԆȓ(�n,z��f�]s����u�>��ȓ:�4QH��}��SfJ��T�����^*�$ؑ@B�X�&���N�?3�za�ȓP���Y��,V;D(ǋC��݇�R8v�蠪8԰m릏I3?����S�? �`hp.Y�9�|�pU�.M���k"O
b�6P��Uj�"�R}
"O
�!��N�a,�L $�R�vP �"O�[�=��psaO�mw�D�q"O����M�܂f���&`���@"Ol���I4,dx��a�YX���"O2|a�ŉ�]A�i��K*�J1"O4UXƣ\�PS22��G�uS�@�"O����� �0,�t;%��?5yAG"O���T��6T�8Ԇ�I#��7"O�	�&C�k����U�V�iZ5ؗ"OPt�q��;�|1�@�2���2"O�����Z�#��+`���4ە"O6��c&Q�_k�8�6�B�n�l��*O�Dy��ʍ+0��gJ��� �A	�'��"�Ƒ�p�>��NP3��8	�'[J@C�K=�
��Tl�.ǐ�p�'���D@W,��`����!%�� 	�'0x4j�ς����3���ܩ{�'�6̲u�T�Ztx|MǕ|�z���'����eϋz"Х��`_�m���'�6�z�5C3�����تv�L���'m�`�c:+���I�W�n~�i��'��U�	�"U{�,��s�� 	�'Hj��u�>a,��A!��wH�R
�'���*M�)��Y� ze�T�'{<0�Y��@QEC�f5��'
��X�̈32�\����	���'�&d;�!�-\�������3�'@� 0��(�h���-��5��B�'�N� �Ep�ٳ�	�	Md�p�'�p�#��[��P�h�)_	TX�'���C�=��dp�L�T�4{�'�PL: ��)�*C��M
h��'7�P+w�F�O�B�Z#c�T�$� �'�z�B��n*��2���d��:�'@����Z�9���F�by��'@�� ��02.A;���U���p�'1��ۥ��K��4Ip��-Na��c�'�ą�A��)s����	�E��Ps�'ȴ�Kǯ�4@����I�FA>�0�'P�]
6	8^�6|zlP$B7,�B�'<�yW^p�&4@��0i$\s
�'a�y��
6R�c0nŵ&�j���'���yT�d@�(��\�^5�'T�r���0.I��G��Z��'�±�Ge�'_�����EY�~?ܕ+�'r�+s%�)V�	��@N&CK��9�'���2W�r��;���4���'����u
�=%�9q��AYlYq�'nƜ��7z!��ѣ���9�'X�c�ŏ��l�p��r����'ʞy��&�J�����<h	�mB�'Jhx�C,
�3�(�Ъ�Y�x��'5����lșmH�� /��TWJ�B	�'�$��I_�s���<T�ν�'��⠪�'(Pi%� }��r�'��p�`�#qU���������'�yAe�KH��1��R�L�Τ3�'<���@��,G�t����?G�}��'¼���0,�jU8�ƚ28}����'�X�3rb����!��A*/m܂	�'�B�s���#^S&4z�!��\gl�(�'&H �󅀯,� �`@ �%�r���� l�	��T���\��g"Ov諷E�f�lq:� V�DP���"O�ř�Gߌ^��3!S9Z9�R�"O�X�ʍ<!��@J��<?�\��"O6�dGJ� �ヂ�M
t9E"O����޾�"`)��G�_��"OBA�/��a�j�c@���ʬ+"O�j�.�B�
x���R(05�"O�!���qt��q�M
Q�,��"O:A��j¯T�x���J�
|��<q&"Ozh3P͋�ު�qL	{��{"Ov)���(k@𼉵�^�5��E�"Op� �O�_*8��r�C�A�J-�1"O�P�A$G++��%��#/`��g"Opy�T���W9���� ���G"O�p�Ҫ�UR���`�����"O�p ��� ���R�B�P��0xQ"O���D�M�~���g/ �jbl��"O�E�*��I/u�$eZt"O�@���C&�� ��ߓ`~�ś�"O�\���ݎi$j����T�U8�"O�DÇ���T<�P���yQ��"O�h�KߤIBj������k���z"O��b�/�#dB���1�ܭ`"O,@�����>u(���Nx�W"O�I�.�d�<���([@$�k�"Oa�3�ׁO'���.�n��Ԛ�"Oؓ�MQ/l� �ݔf��)��"O����NX�Q�\\c�N�42��yh�"O�	�D�l��,�q� �1"O�aq(�xA�bǋV;��`e"OL�35��y���ٸa���1D��뢉�w~P���j�X�>Ȓ '/D�賳iܷQ�d$*2�X�\�A��,D���2"8D��C�O��Q�J��u++D��PS!��IWh�A�,v��W.'D��8�%K�����8x��	(D�`:ׯ2}꒵3�i�,t�y���'D� �ccQ�FX�W���3�II�9D��Y�@F�(|���+
8�Ե��a9��7�O8Ez ��k&�m9tjA�_�؜A�"O�m�u`�v7n�B�]�*){#"OtM�"�z��x��X"Yv�1�"OZ�(�M�G�N��+A.O���{�"O��ᖡD�C9�dȉf��tJ�"O�UKTFO�t $H"C'I"��a"O���רMq�k5F��^h��3"O�0sd�͕6�F� ��L|^L$��"Ovs�`[�?f�MZq*�@ �p#"O�#d�wB�𐡆J-�P����IF�O�&�Ifhu[X<c�k2e��	�'�$Q���:�z� r˖�b?�U��'���zԀ����{�yD+	{�<��`~��I�_�V�0I�v�<�K��>��-�C�sq6q�v�<!�E�(e�2�1�A֘6�1���u�<��Η&m�������K�����]G��hO�Ot�T���ys�X�tᙑ2�f���'l�Q�\v�T��*���'��}��O�g|H0�Qlc��
�'�Yө_���hX�(��v �'�:�z��B�$���`"�'U �Ś�'��P�ł�T��	j��E�F�U�
�'-!-	I��
�V6��-��'�Z�<� �̠R�Z�g��� ̟,�I�"O T��,�+B����̃|Z8�!@"O�9[ҮA�R�@��kՊ����'FެC0)�-t:�*UlR�潛�'��E S)s�Qx���3|���	�'괥`�G�/@�J`�B�_>_�X�+
�'�j����x&&��Ά�QG���
�'��X"��ޘ\�l���i�	3��u�	�'H�]6-�81�Dl�P�A,-J�9p�'�)����vղ�S��A/2�0tp�'����d�4j4���ʏu �T�'�!�m��ND	�@-�Z+�'ߔ��� ��5�؃p�ػPEp�P�'9���#��U�"��LZ�3���'�*�F�f�R�:vNJ4��'Y�}24�J4VU�tj�a�{��J�'1�0�"�  	8����m�xJ�'8�d�vGΰ;����l�Py �c�'�p�4���qq<D�Q���FPD��'��teΞN�� h��DO�`�'�$!�(b5ڗ�V;t%��'nP�@���E����ǀ5����'v��st��/!� (1d�#0<�}9�'^.�wE�	D�h����չ=b0pq�'/�Ը�@]!�֬Ӧ�6��
�'<�k�a�8?��0��Έ�hh�h�'��8$����a�8p�'�8��!_ܜ�xP�X�G�M��' B�K�ʦ�-sc��s ʔ��'�A�1�ҳ�����+�>j�<�'Op�6K�	�A9�J&f? ���'=�x(�⌥Y-��'��W�l��'Z����͙�/��zR��z0 ���'��g��M���k�j=�UY�'"����jŸ�Qh� Uf�p�'d��i�@�	J��� �S�u�
�'�8ř���&�
isg�! t��	�'�y���<XTp![��~{��[
�'�BmBA-*���ȷ�z��
�'T0��Sd �p�g)B�f$!�'�����խOČ:��T����'܈�[��R&~h@���E8r��'�6`��$l�K�@Mm�1
�'��}�`CܬOwn0���P�upA	�'?����s���%�0x-i(	�'3~X�#Y!$pM2E�Ct��0�' 4 \%Gn�AX$�DdѴ� �'���*�fǫy/��P��G$Y���1�'ZD�@0�ц�-�qr�Cs�u@	�'��N�$V�:)�M=(����'���'��Vb�h��ح5b8�)�'�I1���1b�9��dI� 1�'&�I&A�	|cu�Y�Y+�ř
�'X��Y��]k"�y���P�.0p	�'}����D*:�XQ���3>�Z��	�'����#��2dd}ib��:{0A��'tp�	F]���-��O��d�c�'x$-�oD�A�|���E?n���r�'�4�Rda��Q�L��8\�	�'34�r�խX�P��@��a	�'b�X�/�
/ UBs�X�9$���' ��1#�LЂ�T(7��'6��n�#*�P�͋:/(dH�
�'�4H�heC>�($��$QD$�	��� ��H�F"�*L��`�' @�qF"O�	��I2���� �V(@�v"O,��K�$9f�xU�!_���S"O� 6�#C�.Qib�T(p�X�"O,��e	3��#poC�KKV$!S"O
H�ѢӋ��X1��>v<���"O��Y�ԅV��=j1���!�� �F"O�����`��B���4�|�U"O�D�1@͉m6Q�M��@����N�<Qg얓z{ ���V�]��<:�L�<r�MG5�́C�y��T�a�A�<�T�p�zI�R�_.A� ;�,�i�<��a�� ��ѭAF��
�c�<�pC��ChH�(f��)bOl�[ ��T�<Y�mƎl���hbI�G��X����L�<�靜��t`w͏��F��F�J�<y�i�
�ȝBv���4�yKKo�<92nD�q�(ya�Ν��6�IQ��q�<�u!��[+���AD�:S�n�P��q�<!h_��XaE�ί?Q�L󡃐k�<��CL�N�\� $M-�I�E�h�<�g8v�T �d���{���D�Y�<Y!c��OH�U��n��D���zg�`�<9b��6{nhyC��I��Hz�j�w�<�d�W���oބ9�E�qcIp�<�Dn�2�|�0d�s�lթG�h�<�$�Yc�`r��=a. KT*o�<y�)��q��ܲq�L�H'��� j�<Y5	�9��e��8)u��p
�h�<A�cH�Pn����0h�`h8g&�c�<Iuf͙���rL�1zH(XG�_�<1*�=^� �S�B+6$�sp�Q�<���xU��;4W�6&�#��^X�<ѷłP�ts�J��fSШ+��
p�<a ��X;�P!�B9K���#^j�<�Ѕ��+��1�3@G X���xa��d�<��-�.�>� �F�ZT�0��_�<�īP����MQ��%��b�<I3�Ul{`|�u��<(U̽�gNY�<1�(z<��Tؼ ~�A�EC`�<9K�1�D���V�dZ�P��m�\�<�f	��|��p$LY�Z$ �z�&U[�<�W,S�%�|%@"����ҬJLl�<��d�<n�b����A},� S�Lh�<�$LЍ�٫��	s��<k��\_�<�$�@�Y�ܙC��Cq�teY�([�<QQ�~	4Q���S `�<��V&_�<�w͘7t��K��> �>��U�P�<Y����() D�����BQ�<�G�3�&Y�!-��v�V� ���M�<�bW�6�B��4EӚ��%0Ƅ�T�<���h���@�B�얽S�MGl�<�3�3��l�d�ÌE�Lc�%T�<��H_mV�p�$W�<K�(ål�<��M	1"��(U"�X�) c�Xh�<���[˸��NG�t)P5��b�<i��M��.�ȂE��A��e�2�g�<Q�((��d��+�⌁!`�y�<�"�$��\r�	X66�n5�2�P�<q�s��ј4�/$� 	I�<q�-.��* +ޕ.�Ƚ%@�[�<��-Y)7̐Z0Oѕo��Ae� T�<��F -h��������cM�]a$�E�<cj_/A�xH���e����H�C�<� h�9G �K�t���;Tviu"O"䃑)�	�l��B��Ra���b"OF�x��H*&�����	ESh�""O¸�'�S]��A�/�7H6]*�"O�,��	x�i[��K)0�Q�"Ob|0��b����`�7H�"O�B��H��4���� >Z(��"O@��4�@�9}l�����	���"O6Ԛa�1��DõCwZy1"Op�J��Ϟ����mC�X�8̉&"O���ڤ ����+�4۪�
"O&��O����Y/ː��5"O��V�z	ss�ڣP�LX��"O�
�$��	D0��6ɂ+?t�"O t�jE/7�5QS��\7�%j�"O>�k4�@�q}Z��V�Hβ���"ON�j �[17vĐ�fjڛb�L�C"O�!`���YX�ݨ�	
i�d%�"O���"`��X��W9n~��(�"O��8��B��D���&"���P"O��[�Er^�KEH�|�h���"OD�1 O�5W��%Y� H
�`a
0"Op�(�Q��`�pA�H,z0"O���B�ū30��v#H�x}*�W"Od�BÚ0��u[���r��Y;"OY�ï�(so��1g ��tx:�"O�]���хc�~m�6�P
�1��"O
��g+h�&d�f`%Ȇ�R`"O�];!Zd�%���V�=�
Ѐd"OƝB��[8>�e3$�խ*���0f"O�ܳB��v��Q2�mD��8C"Oj@�0��"��Z�,�"O�p�W`K�q�>(z����x�+�"OB͋�j�O6:��o.i̴�*O���0`G�m�a�Gk4���2�',�������zѱ�k��]�`��
�'᐀#E�P�r� ���h	�S>0��'fH���\�?�� �E!S(t���p�'P�jǟHg4�&��&f=���
�'}0�C�Ò�)���`�V�Gl���
�'�*�p�"�&�T�E��'c-	
�'B��1*�+y+8��ɛ�s�D���'��%���I	>�* *���e��|�
�'�%��d��y�´��m�./�h(�	�';�:��=�j�B�\�s<���'�2e$�R�#� �p5Z�dEl��'��$�ȫ#��m�5���W��Q�'����I)��ڴa��]0�'�b�;�(L˖���)��x ��'�Bq�!gϥ@�JT��5�2M��'�^ٙ�ВCO.�ym̈�\` 
�'���x�c2���H�0z��	�'&�9���W>n�S�A�w���b	�'���;�J�u�H�jf���l��)
�'c|��@H.P| v�@;iY���	�'�-P�l���<(�Ř�hC
�	�'�dH�#iף4�:�+��s�pM9	�',>���@s���C#�[�H���'��xa��1u�|�C�ɝVU^���'��83�%w�8��2�0H�D���'�@0nF�9����G^?B��l��'���q��oC�؂t���i8��'2:���"Һk����s�^;cDl�'�^-)��L�:��в䇐r�i��� (8�aOw�^�����$����"O��A�ψ�]l^����
��HT"OTH��� ��M�d��]$ ��"OtE���*pM����P#xaؓ"O^h�� �\�" �6G<T��T��"O�l �-�8x;h���%� `	� "O�ّG�H:/_�9��D
)-��t"O���R���骁f�@�$��e"Oʨ�2KP0K�Рg �%�ĭ�y����b���C&�Q�ׇ��y���
�Pl{�J�|6�b��4�y�*�9J��#��X�)qf̏�y� ?��Q[��X���R`��y�)ۨ8��T@v$q����ybb����]�$�[�8~��sg׀�y��pj��ɳ˃�;�RC��y��N�6�IQ�{��2�R��y�*J� P ū�S ~D(���	�y2����B8R�CH&��q�1�Տ�yr�E=kh�1��$r��q��yB��4X��;�j9�tT�GiS8�y�lB�]�bY����u��5��,��y�F�;���A�dWoj\(��G]��y��B�nTc�I�b1�Xf ���y.׮6��	�i˜j��H9�Ƅ�yb�W0O��dp���w�0!�ea�yb_�N�48)2A��gO�5:�JP��yƸr�zek�EӔY�^��͕�yr�67xR8��L�#U� Q ����yR��7���[�ɂ�IpxH���y2�B�?�Q[�^�<h���Ç�y��_�V���i��
*�b����y�$Z1p)�p v`�j���s��$�y2 ��f|�|�k�Φi�dOI�"!��\�k�0遁e�C<����Nܹ|!��U�4K"����F���*֎���!���8׺�a���#�SmW&�!�d_�^�����.�����Էw�!򄅯pR�<z���@(���O�;:!���6Z^n4�5�ڵ'��S
�!1�!�$Mo� �*�=��I3���Tk!��>R�J!{1�˱�H ��HD�!�DM(eN�����:'�4 0EЀ`P!�$Z���vΖA����d�K!�«v(�(j���[�Vdc��$p2!�R,PA�hP��߿U�~ͱJי$!�gD�b�/T�?����_�e!�d	2~��w㜯)K>� j/S!�$�#s�шC�#25���HݑfV!�Čn�F0B*�2)���C⊨�!��N���U ډk,x���� �!�D�Vn�9F�O�\*M��^�Y�!�d`�hb�h�9}W�d���!]!�$I�	\ d�B�^Rp캖��"T!�DUd�x�rF�R�UP4$W#.!�d'@��۔�>M�|ssC�1N�!��5#�\Q��]G���A��0�!�dEG�B=���k00P��C��!�$�=M�r\���	 �= #(��0L!�DN/�� q�[36i�I[$\c!�D��1bB�h��<"���
5R!�Dݮ8s��J_�"�3�IQ25!��W�S�����9Z�,)��\�r�!��2D�.a�V�����*3̂#�!�� �%3ԏD;5�V��s�$NM�yӆ"O^�t��:����V�Ŋb7���"O��aE�
�Aq���F->�"O����h�G��1�[�]�ؠ�"OPy+������T�&f��q1"ON�0�i_���B��S�?_���"OHU-ee1Y`�ϭ���qҮ��y��I�)���6H6�tJ£��y��²W	���V!'r��+­��y�� ��Ƙ�#Ěi�Y���=�y���J�HHH��e� &��;�y2�A*��ZD��a)l����Y��yR�ϵp��`���S�pЖA 1�yRO �j~�����ڞz�f8���^�yb,d
���a��@���d̎��yrIO�{�
�xA�!�XĐ1扏�y"	֋I2A�ᦃ6/O�{!M�-�y���E32�X�-ҡ+/`ݣ���-�y�`��`6�ls��Az� 0�
�y�i�DXBF=}Όa����y�I"��|xU�匀�m>�y�홥#q��a� �6$B��y�M�qsX��,5ڀez�mY#�ybE���EQ��J1.7��3�nI��y�f�ehSA+*�^H��y�͔%ꔑ�J�!�FA4F��y�%����_�C��xI�ȓO�&�(A@Y	E�$���J?h{,��k���W����h-��j;=#�4��D� ����JfBYÅ��\���ss�8��Fːz' (��
|��t��&Yl��H"��Y!��[�D��4|]C���ib�x٦���M$�X�ȓh�f9�u�
1g���B �����ȓ'�h���O�8���Jf�أ[q��^���Rg��2ˁ�ʠ7N8��m��Mr3�7l� 8@r%�l��ȓy�piZ���~�jm�юC�	���ȓ,]�ZE�
1�P�$ LmR-��Dn�� pS<#� ��j�6���4ɶ8����d�R��BcO�r�H)��QE����J�l�N�#��:g1�M�ȓ&&��2N�8j4S��V�.'���1_������<�BĲ�AZ���ȓL�5���L$c|����O*��1��O �����V�`��%����X��@�#�L�b�3�� bd��B����r���A&G�k��<��h�0��RS%-�����i x2ԅ�Z�z��x/�3�S~��C�&Ex@��nO#A�Px(���C��;4�I�#g��^�t<�p�̹wʔC��m���q�W=kDN�3AK�`c<C�I
udV���쓇��h�N8TC�ɛNÐ)���
&%�T3�N�)C��(!0���V�}U���K�U��B䉜S���B� �~���nI�55TB�	���ys��HQ�81��`�C�ɕ7�h�Xl���Ҋ<�C�I�%�mZ�V)r�J�(��݀pC�I-]�z��5�	�p$���(PC�I+�p�S�<�t���Eu5�C�	]R")h%�	�+��%*��%�C䉤?ۚ��%�1�U�3+�E>�C�)� @)�����.]��EQ�l��"O��Í�_0@��$Q�X�:�zE"O(I�椄�i:tT��c�N�2�h"O��r��s�l=ȗc�;�B�y"O搠b�\�k�B�{Qc�(Z�����"O2ئF�
<:BH�$��1"O�y���P2l�f	�wp��t"O�����h�P�It��3�v��"OF@R���t���yD)H��$ ��"O\T��5�5p�bP?���2w"O
5���L�x��hwk�gZ�᪐"O�R0�[��R�^;<��B�"Ob�x�G�\���ע�3j�i�"O���A�M�udI���_��Q�"OP��q��{r�i�`�z�ʼy�"O q �[(�I���>n+�	�'"OԌ �G�|��u���]2
0��Q"O�����UU�)���N�
�"O$ "�X�Й���7|�XU1�"O�T��E�zTL��i)�PC�"Oƀh���&��Ԃ̾U�*蘓"O�I�Bǻk8���� ��^����"O(d�{���x� �n�0���"O*�(u�,�l���P�t����"O5��d�BV!3�E����yCb"O�y���҉3���C!�	�Y��4��"O��q��-fkQx�������"�"O��J�l��E�l��h�*����9D�����M$)�$*Ø�^�a3&"D�����7#����fnn��A$D�l �Ȥ���kRyvp(��#D�t�G$54Y:"M?	L�P�"D��E���R��(��Tt�
?D�����C��D�pe���Z�;D��x�R�(�q� Q�Н�GG.D��Z���J�Z-S�/jwx B�-D����-Qp�x��߀8st�R�a&D�Ta1��-<�����a]�f�X����&D����$�T9�䅚�]�$E�#7D��eS�>	��8��Z�5D�x�E�K`p�]��i�\��؉0+4D���eoT7{S���	*7t��D�4D�P�E�H�g'�"��G�J{>��g	3D�d��H�	D ��`��}RU�/D�lx�پ%�򉸢m��f��! �k)D�tɆ�@�p�&ջ�Ǜ$	(�52%�:D��A0�Z	���k�37�b�G�$D���E�s��=���i]49�w�$D�l���E>#�bIq@�܄n� �Y�$D���l�P󾸈q�Ml<�9Q�?D�R!�#c��Pw�̎6�q���'D�� f�&* �4x�/��Pxl��� D�(��,
Hipc�'m�p:� D��%��Jj�8�FǍ2p*i(C?D�P�a�W�&!�4�*L����Pb;D�����Ӗ{�*����,ꦙ �l;D����2����N�^ph�$&D�P�cƁG7��c)N>R^�'%D������a
H	Rݜ̺BF(D��v�,�ԡ
��؛=Nr3��*D���g��(��@eNJ�B
8D ��6D��; �)D
��I�	� �F���3D��˗C�J�]P�)K%$�D�H�h0D�x���PU�b�÷�I�E�>����,D�� B��B�.	0w�,���"O�.��ڱ�4��m��]�"O��kp���%���b+ϼd<d��"O<|�QĜ<�^���el�"Oz�#5H�_g����&�*���
"O<��T���?��
V �''�ԭ��"O�&
�U�|\;Ei�?�Ґȇ"O&<�֨X��\�`@)�)B�I�"O��sdT��ƴBc�6e�z�iv"OڄI�_��.�A��ɯ��!X"O��Z�f�.d�vԻ東X�<���"O�t�'�K6O3K�""�> ����y�D 0�=��bL"p�,��cS��y�i�f�z�����b4�p�e��yB�2�p8{� �Uc��S��yZY����*L�# =1��VC�
�vt�4V�G������#�C��&$���#�Sp�\�@�Q&1�C�I7l6B��$P�e�D O�$+�B�	�=�M��β%���At�M�Y�B�I,4��#a�° r�5�f�
���B�	>O �2�1Yj(Q'
:+�B�/~��棓b����4@��B�I�,�8(�I;p�!ǎ��I�B��1[J�8�WO�7~#�����,��B�ɣ[B�{P�OAB�a #�A�
H�B䉉H���ȁO�\�Хp�s]�B��JYޝ��q���tD¥��B䉷Ry����K>\���Ƀ�/tC䉅�vx ���s
��R�����C�I`���֧�RŐ#�|�jC�	5t4�Z��ȃ�&� �0MjC�I#C�X	6Ne	F���]	ZzB�I�e�vy��!�?@g	��j[�xB�I�q��q�a���IÉ�	i�C��"K����NΈk��r�F��T�B�	2!>�cC��6��hN��E[bC�I4�$�t	H�wx���u���X��B�	�آ	ڙg� % ��<8P`B�0@���A� q&�bƃ�L@B�I-x0�|�eHB�Q�����"!B�),q��XlD[�|B�� �@��C�	��*uj;4�v@ �E/@C�I<W������_8I"E��i�B䉴_��0BQ̋�"�m�ƛd�B�ɬ/ڤ��U�_*Gl��jg0W�rB�ɒ@���P )>u��(���e��C�	�s��`a��ן$�l��3�H�n�.B�I�0�X�anV�2��[ *�LC�I�Ȁ�2S�
*��y���V(xB�I,x"��) ��m�6�Ê �>B�I�*%����o F�7���R��B��4dw�0��F�	���(�nJ.@r�B�	lO`��������rb	�C+RB�ɣz�kA��5f,�}c���s�@B�I*�Μ��K�A
2�2�mç4dC�Iz*I0�g��8�R+A�zb�C�p �\����-��%���K�
C�I�\ �U4	�$��N�<�B䉞	�TDq"��P�$Y�4Z�WC�I).�)Y2�Z�>� �� ٷ0��B�I1Z�
�@R�G��蠤���B�I3b�~���΋�(�<Qs��Ld�B��'RP`5Y��#��i���+�`B�)� $��p��b:Uz��
?����B"OpȘD.^1&��13a��,��s�"O�pg��10
��&�H�±"O��f`Q�gC��s�O�oT~|1Q�E{��	�6=M@x��ٿ;�veȀa��[U!�$O�^��-�q�4<�pZF��!�d�a0ƴ�uF�?S�a9E��[�!�ӳ/F$�&��I�,��s�J49!�d��&�|�IǏ	�Z�$r����)!�ݝo�<A`�^U:���i(��r?Od�1�M�i9��J�Ċ�6���r"O�4����
��d�ߴ m�T"O����A٤�H�Æ�G���I�"O�E86�<D�r��`�1zQt�"O�T�É[�tS�h��Ef.椳5"O��3�����'L�GK�|1�"O��r�lZ����&<*�y"O�БF�0�XI1U��"�8�"Op!����E���5��i����"O���i[��� �%Z*m�\@y�"Oh��̖�k��D�ڷd{N QG"OdC�&��a,�4�!d���q�"OxбCV��n�S�I	7c�z�"OX"�`��)�F���A I��U"O���7&H�dw���j�D��A"O�`8fh�FIÂ;�)�u"ONR�☢�$=!Rb_	/�^�1�"O��JriV�b�]:�!F~9Z"On(pW�I(:���n��d�.�ZW"OⰈ�)lue��rƸ�B"O�2҈���n����NY�ڃ"O4�+���8�Țs��(X)��q�<b�-�W��0��@�)V�^u���,D�r�oR�e5&�"�߁?1N!�SH,D� ����X�@ؒ'H�*|��`��?D�����a�1R�.rꄝ��3D��0uON�G��"e�D)EG���&D��H1�DnD��Wo�DwrѨ �$D�`��O��I�J§�bipp�#D�h�&N�~ݣ�2�<�eD5D�8h a�.wb (��^>|9jX�t"?D�H�G�W6$��#։�� ���Ӳ�<D���u�Q+^c�܈!,��,���H.D�8��lV0Q��+�ON!X��)�L(D�TC�
�;(���	H*Q�t9<D��s���59I.pǌ=V})�/D�����Ae�=��l��dH��"D���V�V!HJ�x����3zE$!z� D��p�D�$nT��
��מrN �K34D��B�֍3�Y�e&B�m�
�	bd0D��K�	<x�V��C�v9%�DG-D�8��G�&fg�h��¥O�Ԥu�)D�2�I�@6Q���
tj�ȥD'D�t�1�ʸG�2���Á�v!T��qO#D�؂dc�7\��1���p�v܉�"D� @�DY�4)�Ts4$T�gF>�yDl;D�l��#V�H~ ���D��.�R�r��$D���'+�AF�L����8�l��k=D���aE�HXB�K$��1a�;D�XY�V+�h��(JL��I
�5D�,�V�ڶ<4"��MG
�����2D����/��iƺ15��7Ϯ$T&D�X·�Ωp�@5�H! }L��3%D����<�Zu�8Kb�W0D�� n�qUH��TS��B1��Q4��b"O��Q�΄L�n��4`؝(�� �A"OT�2g��'A6��v@^w��$"OXdQ��X�!R�g�db�"O��im���x�UlR�a��9�"O&0�GG�53��a+%��1Ff(���"O��2��K�.�8"-l�CD"O�|�IB4g�Ф�� J�Gt�ڣ"O&�R��u�IЕa>m��Xv"Op��T���U(n��d@+a��a"O4�ɖ 5g�����n��R��
�"O|����}(6�{W��%ӌ�H"Oby%�
<ygB��A��� ����7"O��2���*�f�̛Yμ�@p"O"��G��<p��� V��pa"O�YWj]�n9�ƶ�5C�-i!�d��f�jݨ�fU9&�xy�7�V]!�DJ|� �QEH7.�z- %C�<y!�$80��x(gc�	B��Y�U�Z�;?!�䒶I����v�
�	3'�?�!����HL�RIR?n�mS!�$�!�$�|�룂�_c�X�C~�!�$ҾT��Z�iԅsW��!�D-% ���"f�@Q���#G��$ U.ڸ|���OD�$�O���Ę�U{��k_=nO<�ؑDAAE!�	Y� �Bu e���E_��l`	�'�R|��g�|��!i�iт�8�	�'���*ɏl��1��b����]!�'��̙��*gp����ޡ� �
�'Z�݃灀(J�BAE��Q	�!z�'�ȼ���ɑ!X�]8"�[� ��h��'Q�	����8~^���E�D�}���z�n^#q^fC䉗��*L����i��%ܷ�B�I9h��J�z��u�ƥD�6��C䉫^@�q�Y�x�z�cC
{��C�	;F��Q�h[�5�$�	�:i�PB�	�F;Dqpek��&򴝢���9S��C���I3w�:���ҎY�*�nC�I�x:��dj9[,�# 싒-��C�� ?��[��X>=+�%O�ErhC�	�&��u�(Т:��#-L�J+�B�I%cs�Y��P�f�x��́)8C�	
nC|kd�r"�`C���9#��C�I�������J����.P���C�I�!�
Ԁb,|9�|�B�,ϬC�	�D6P��� X帴�FK՝GR`C�	�5��iSde�+w�@e0q�]bW.C�	�gh�`�л*��J�I"]�B�I�o��0rp�T�
�a��2ԠB�I�yu&�K҂R7?�(p�$X}�B�ɷVr��#r�Y3|�PqDKF�l�C��.JČ��d÷U�عQ!D8\��C䉺0������+9W�D���K��C�	�|pt��DKY����cw�f�|C��8!���0G��)0�y��1��B�	.�~0:B�Z=+�,=p5�ـJC䉻B*�)�gCi�(��q��"B��_�\�`I��4C`��b�[��B��.�i+E�E�6-��
Ħh�
B�	.5yD�0���Y��в�-�C�ɲ�\a� /��?�9�3 ވ�jB��"���+K��	X �37@+$B��6u-�l�a��Pg҅pÁ�C� �f��ǐ,=�eHRc��<C�)� h��N�:!H�j��ܘ�>t�"O*D{���?�0A�����N��	h"O�8)׃��� �LY 
� �"O*qiCB�+R���p�K_�e�,�"O@�����;+�=)+;}��02"O�9�̄F��� �M7��e"O�B�F2(��C� %tM�b"O>L@�f[q�T�c�L�jH��"O����_)7��Iq)�1�n�h�"O(�;6 � z$b�i���#ʘ �"O��K�H�`#gbԼl��jb"Ope����~�^H�!��Q^\,c�"O��@��̈́3��b��b(���"O̊���&��u���@?<�yq"O� a$\���\�B���x�Ȥ"O��)��"g@@�ׅ�%i~�H#�"O$���1k��pWeS-L��
�"Oȱ�C�--��%���>�\�+B"O`�"e�	���l��i� �"O�aQ��؈g�UzeAF8-̺ �"Oؘ�s(.ML ���<�<��F"O�9�e�ǩq����*�$-�j�c4"O6l���G��#�L��px�ES�"O~��v�=2)�fJ��t��|��"O(@qw�7u(��9G��
DDq�b"OT�	��Y,}fh`y��M�*�ͺT"OvT*�⎝p�H��a�^v���"O:��w-��J��4@&�^!�	r�"O�kV̞R����H��s�B,��"O�=`�V�A9��߭z��Bc"O�Iâ��"W?tk��E\` ��s"O8!8��Ogl�	�gO�MN8��"O�����J��S	��0/���"OF%`�N�]=B ��ۗY .�u"Ol��daB��H�2>e�$��"OTmB�ʛ>�PtRa�4q<��pr"O�킵�O%Jab��cB� C8�Y$"O��� ���R"�	I?�]A�"O���1����Aᒐ)��@�S"O�9jC�'�T�`�%]�}9"O�`Ӳ�W2��E���2aSTyh"O���&�ʛ2,  �,�L��"O�dt�Zv���0����6��"O�� ���>/J���F!>�Q"O&��b��CJ�	U�
�'-�"O�	�K��O��MYG��)�Up"O��0 �(Mb�۶ �@���ɷ"OԈ�o��7BP�U�<X���S"O��� �	�(	C��Nk���e"Ob��j��S080�dd�E;���"O
]c��S>iȩ���x�v��Q"On�9��W�\��,*S)ҏ5���S�"O�0R�$�J+򹪐��5Ɩ��"O� �*�ئ�Z�g6ݸ�G"O6}E-��T��}	�H��ea�"O
���j����� �h�R"O���@�γ	�8��K�� �v���"O�tx�' {�ЌV�M�v�Py�g"O�B�"�;5:�{� <x����"Obi�˔�.�@xcqE�j86m�"O�Q!��5/2髱aגa8\\��"O� �i����L�q�@�RT��"O�䪗Mqδ���>��1A"O�� ��d�<����� �Ps"O� �ٻ��ؿD��Ť����(�"O� Cʅ^ˬ4 �d]�6��"O�����[6B�k��З�ޭ�"O�E�b��'.Ϊkc  #�`�iv"O���k�c}AR��'c��1p@"O>�:��E�b��X�&n�*~�:A:4"O�U��g�q(�U�ܢag��"O�h���2$�"$� JX��"Oh!����X�T8����wF���"O��ӂË�h�;a�ɼf?0M$"O>pÔj�	^ɫ@�2f.����"O���EN;Q�!i!/��0r݀�"O@%����\Q�Ih�N'v��ن"O�pp&�)%5*�@��>%��jD"OD�BB΁[���T�G:�e�"O���C�.�A	v��̅r�"O\@qr��D	(�"DkX8�� �"OԸ���0D2�fJ�$3�J5�"O@�8#�9�F�x�c�b���6"O�\�E�е���7IM��Ç"O�x#B�`6��ÌD�14��pP"O��]%0}Q�B�[w�0�R"Ol`��LO�)���ꃃRw ٲ�'���H���WgT����4�d��'�R��FA�h��+���6�(��'�v���m�3!�j nNZ1 I�'��2�������h�J��LI
�'j�2�ڏl�f�;�eA����'���ů&@�X;&��_�,	I�'�8P��L���y2L�Z��
�'',��7 �R����d�J����'@�d ��[�q�A�_<F�i��'�4�{�Jѥgծ)��>����'�^ A��	J��-i�A2A��	�'<x1��Ch�T����}D��k	�'""����ɗV���R1!�x~���',��i�+Ҏw�$��EvFf	��':�����!>�0�zG#6g��l��'��i�����	~"�@rl�e�V�k�'��D���:"�p}���u�8�p
�'+�@�h�c�f}��M
i� T�	�'��a3GU=Nk���%��H	�'�<�JQ�֖~#���-P6ڍ`�'����W��D�,r�'ɱ@Z�
�'�^ã��~�x�
&�N�w׊�*	�'����5�@�N4�LӒ���s2���	�'��8	�(ܕZ��i��"��Db	�'�|R��<��1��Υ���	�'�؋�!E��̉�M�{�
��	�'\VɳV#�#^)�횵�SnI���
�'�
�[G��.[c�<�d��l���2�'�!х�8�X 2%�][<�d1�'�|�)�&��k^q�D���d�D��'��|b$�N�F�����>c�2�Z
�'�Xx�A�R�v<���Ci �\�����'�6b3��T�<yò��UŚ,��'�8t9�ǟ�bK
1�f-�)I����'�*$�riL�?��cӧ�++�����'���D��h�R0�w++�(���'�puCqm /��8�J�&rD0�'��`�����!��"��D��'":L�5a׀GJ���^���i��'i�Dn�"K����gޒ��L
�'ra�bމu����&�̡RܤX��� �u���N><-�\B0�=*I��j""O.�!��ř)EΡ��,�'@e�"OP`1$ C1z^r�h+��_�VY�u"O=6�qY�t��%"�T�Z�"O���r� ���bH��<��v"OЩY"W���\
���C"Ot���B�o������p "O*��ej��R-�C��i��g"O:�x0�ʝLCt)!N�D�M�"OLP"W)�4t� ��OU	jHZU"O�����R�9����"�*M����"ODD��AĴ(;�H�3�	�[��#�"O�9�i�2\4�PBg�m-�P��"O�=Ye��
 �He�7F
 ��""O ��#lH2�\]��e�9KwV`��"On��l�e��[#�m��C�"O�9��S�<�Y�����bh��P5"O6T[�	R3R$="���1uM�P`"O�ʕb�4\�fȐ�nN�yB�Hs "O�=���Ԓ#�⍹`�<?˔��5"OzQ��hа$Ad)Z�����g"Oq�c�G?yk�m�4�Җ&�8x�%"O&���B�b�<�"s@	5D����"O����E�H@����4;�b��F"O68It�(p�ؽ��M@�Z϶`q"OD�UƔ9uH���LH�.�̹B�"O���t���-+0 p��P�Cَ��A"O�XH#ǝ"mF��������q#"OV��g!�<>t�S%I�=q�ə�"O4"`NF�!cB��c�hC�Ф"O�aa�	$����]0�)�"O���w�pz���J)D�~l�G"O�1D��m)ā8cD�6e�ڌ؃"Oj��vJE�/:�z��Vzm��"O8��T�S�J�dSw�� ���"O1ógV R�Ű@OUcb�s3"O�y�b,�>NP$Eفnw�~Ar�"O��ڒ+�&��(A�_2E�@飳"Ot�Z��:_���"@"�,G�"O~�8A���i��]`V��A��"O�q��'J���,؂&)"�
�#u"O"�P'�U%'h�EC��żC�X@��"O r,�3|Y���e�t�b��"O� ��n��-��F� H�&"O�IsC.��%�l���+^�rhD"Ob1Ps�Q�����P��q�"O4M�WlK���)3h�%~���"O>���ͽXB�u͐�x�PR"Oly`n�,�X���^1s�*a�5"O��;�H�la޵r7,�J�J	@"OPP23#�*2�� aT��|h8PQ#"O�h��U�w���1J�9[}p�"O��E���*#�GH3:�"O,sGM�NW��EΟ�P�t��'"Oh�9f̂�U8��:�)pgz�R"O|;lڙ9�J�Cd($y\�dC�"O�Y��DI�/J���RM;g����"O�]B7�ǝe�N2!�K62�(�P"O��@�C"	̔����?��e��"O��Y�
ĩg,���e�;#����"Ob�P�'m��1b������;�"O���Ư^&|l�2��\G��P�5"O�(Y#M�cZ���Ђ�y�tP	�"O~��CcZ�&�:T�#S�\y&�c�"O� z,q$��#u��ڡ`�v����"Or0Љܾ2��*W&�=�tp�"O���v�݁c�h�ܻ1r��"O�h�G�DOd|�pƊB�䥢�"O����~����+�����"O��Xp�ؔ3P�h�G�TQ���"OVAXd!	�7����O�4�w"Oʑ(���{8��Eh�f�Ԁ�"O��C��9~(
 ��g�D�
V"O$�ZW�ۧw�*x3��'_嬙�"O���ѣ\����2N��A�1w"O(���ǋm�yGC�>1L!a "O�8s�W�\|f9��"��dF��"O~����_u��k𯋂VY�I"O(�Ԫ��P+Ch�"sN^T �"O��V�	�Z�[#�X:�	c�"Oj\B��֣L3��F� 4S���"O�RfE�a�Xk�HLp�W"Oʽ�fj� 1Ԗ4�2k�7ML��2"OZ�j���{��`j�a��"O���FJ8%;Ļ`����tå"OJH;6٩~���Z$�E/�,y8�"O�z��	x3v��V��o�\	��"O��� 
�H>�(��̏Z�T�y�"O| �c�+w���@Þ���S�"OnY�D�"ض��cS:��H�A"O�����B�LX��܀Ump1""O���f��}�u�L��4�\��r"O�y;u�Q5oRL��5k�=ˬ���"O>��������]�û`�88p`"O,h���Šs��3��&I��u��"O�]e
'm�eç�0$�r���"O�\����(T-�	�*�P��'"O���n����H�(9�P	!"On9ّ�/�jlr0%��\g���4"O�`5^��C���68�Pi�Q"O�`��i��gNy�Fbڊr�&8��"O����i��G��#�&�.��<�b"O�8!��;!9��cl���"Oe��)�2�E1�IH	�Tģ"O��ҰG�[y��Wc�"�PԂ%"O�d�$��e�:���g�i��$�D"O�p���S�l���O*	}$D;�"O��	`j3tB����.Fo�c�"O�������iy�؍7U���$"OnX %�7¸���%<�,�"O��rᙞ?1�4I�*.�уD"O�����a�d�QW.[%(R(�s"Od-��h�xj��ю\ ���"OjM��������Ӈ-�J���"O(�j֢����aLٌKC�JU"O̠�#�knN���	Ųs<�zQ"O��`  �- R\ɃI�)%�;P"O�r���N�����(���I�7"O�r��=x�~a@e'ťv#�Q��"O$T��O_�(����@�P�L
L���"O�1K����T�U�V���fՠw"O����ݫs��1�'aY�Uມ9"O��#�S%%>�P�U��=ds=�E"OeˁC;[��B�4	0�qB"O��2I<����S�f���"O��rc���Y�j%�$g��{e��B�"O� 6>h�h�da�ha�"O���b�ԓ
���;Ƌ�&P8��"O� X}�n0�8��C�Rd\��"O�0��-cE��ze���Q�����"OF�[�O�(@�������L�BU�"O���B�V��ztp�t�X !"O�E1.�0m��z�@�	!����'�b�@7�]8@n@;�J�-d2La�
�'q��r$��Q��ڧ�҇\>|�+
�'#ȍJ� ��w�2���@[�O��y)	�'�~���Q�V?8�j�(�Bn"T��'R�+��)~�\�4��7p��i�'�� ����g���U�ϒ�^���'�2�[�MF�XD�t"-K&Y��
�'�Nd�Y�s�>�	��ߩz�	�'��H"$&D �ڹB���pZ�<r�'��s�k,8s�i3Ĉ�m8�H��'�8�#g��Z��`I�oV�:���K�'����2D� 	Ka^ [��j�'�ڠr��Jr��#����'۴$s�(�+YJ:СD�%�tE!�'�(ء��[q��𤒴/"���''R0��a��g�@ r&� $th�'霹;ǧ��]�qZSe�O��Qx�'�֥a���?8H�!��囅��P�'�:V)�)k�Bi��T+=�$��'Ӻl��iÿ����%I��.�b@��'KB@J+(f����J�"�Π#�'��� �W�l ԨƉ��.Q��'9��F�I�k礪)f���
�'S�53���[t��R׃6U-��a
�'htpτ'v��ś�m�
��!
�'�F������5Kg�>$�2	�'��[`��/�0�I�@����'Vx�'�([n8sw�@�@ؘ:�'�h�q-� -Ӵ)�R*�L��'�P�r��*��|�6M
�#8�ĩ�'�Ь����-�$�ɔe�>�����'H��*���%���a7G%G >�+�'�t<�"�:S(��AA�49�	�'�])�a`S���@4"]4"O�	�a&H�B ,%k�F�E��X"O����$N-(BB�#��S����5"O�	C8:���jë˹?�܃"O����N4hN�RDKO@�dq:7"O`@P��(r* P%�S
���E"OzuHw�&(4 �C�)O�|؀"OF��`�E�L��R3"5tl@��"Oh�r���3�r���"Y8)M��J�"O��+b���X��!
���o7�2"OJ��ϛZ�ț�`�(9'����"Ot呥,J�d��%�6Ζ�xd|h"O��v����D��0��2'aR��"O�����g&lĢP���%lj]�A"O���ˈ*�q�)�	aeL�;�"O���a����y���)9R��"O:�x�.U-;}&�����oD��H�"O��1��]^��Jt��}`>|�'"Ot�C1��o➅H�@�D4���"O 4�&&MA�֨ u��_=���V"O  �s � %�@��/!��(v"Oxe:k�4UwD�
��P�_.�|�3"Oz�"��N&Z��I�BA�0kLp�"O&3���%g#�QKso�	2"O�A�1E�����G Z���7"O0KR�\�"V�9�F��1j\�:"O� >$b�?<�|�0�QN�,��"Ot4��1t�D���f?&M04"O��E'�7P�tm�H^'':�"O2!YG��V*�=5-R�aw�
�"O�-��HM _��t��፞Ah1��"O�!`gE��6� ��H,���"O�В��^\Ҭ`�o�O���˔"O�a;�
W�h72�:�)	��D,��"ORM�Q�5��1d�|�"OZl �$ݮ8�b@��� g��L�"O�PpDE�hRv=�U�������"O�!h�eD4�q*V:R��y�"O\��l� <�����^#e&`"O� �2ƍ�|���0aL�(* ���"O\��dGI)C"���]�l���"OX�.Wt��9dKV���[,�yB߰T��q��T(�j�BV��y�¼C��0(`��I�����Z��y�IL#ySڱ`!g��6΄a�4D���y���\�����+-q8�#��Ѣ�y�&��G�r!C"��L~��eeѤ�y�Uy�z���!Ƚ�Rx���Z��y2)�>yg�� R�k�)Y�y��ܑBDb��#��ޡ+�����y�`N5R{l�"�E5Ů�I�)� �y�ӯSSҔD �xR$˞1�y2"A<����F��yDT�� +J*�yA$r� 7�dh0�
Sm�(�y���s^��jҪ,+�2��E��y�JN�J����Q���(ɀ��6L���ybC�`�H%��S�T9��ȓ�yRLȐ=_�-�d�ϭ`I�A�����y��J4�&�����2p�xxh����y�JM����Ó��q�DA;�y�ج��	����x�qv�߲�yr�s�%1��]+oD�h*��y��7L�*T�B��1sbNi��Z��y"!
	����CnLZ@ AF3�y҆�b0�ٗƆC>�Heό��y�_�Z|��B�
��Iy��>�y�K�:ی��"o��rh���#��yr�˲t�y{4�^(}嬵�b���y�K�s{$��'�� 
ʈ�`E��yr���:)��f6ƔjaO^��y2MD��RƐ"�r�2AM��yҭȤJ�*���_!y��-A�J��y2��-
(D�a��'bq���P�]��y� րw{�]�aǋi]�ؑ0��y"���$��D�Pd	M$�y�tdK�y�L�f,���B0Dqp�0����y¦�Hˌ�����3�U��-��y�����D ���Vk��7Έ��y�b.Z������+K�z=ʗk��yb@^!A�n���@6�[`�ֱ�y�IK����#�<@�F`h炗��yr�L$k���� ;7�~1��[��y2��}ܴQ�c�Z�:�z��r�T�y.�0�3��5/�����y���g3��k��əCV�x��:�y"a�	�^HY�$�1=��H㓮L�y&ߨ�����73���뎑�y���Jt���NW�|V��u����yB�|��0�AG�$e��[��I��yr��[B�����i`"�q�(�y
� �s*0\|ؠ���GdTtj�"O�,a�t�9��ʄ )Nhb�"O��s�	�c��4
7L۽Ţ���"O���A��*S���Љӆ~a�s�'p�d�A8!i�m�����$F�!�d ;Ѩ�1f�΄ɳ���V{!�� ���S��+#��Qd�\�l!���!^ uK��&p����g�cY!�$��V3Rdf�)�x�s��*O�!�Dٳu�z�L��2�	t���0O��癸2���MV��2d"O�Չ�m� 0EQ3Q��ږ"OzTӐH�x�a�v	�:�"�"O�mcA�܍U~�D��g�,�H1�q"O�trV�L�d��v'De
�b "O6x�%��3Bw��'����"O��wO��AD���t��逥pR"O���Pn�d�,�2�](H����"O�՘���a7vx����2�X� "Oa���Nu��A��(�>�$"O|��ȝcv��ptL�~�:��w"OP�� iў$���I�kY%$���Z��G{��iY�5h�(Q�Q ���9���C�!�ҝ�f��#�K�_�x�u��,0�!�$- j��'���g�\�$�.0�!��"}�&�h�jY�8nt`�L�Ti!�D˜��}� �>z��,�&7�!�dԓ
n���'��+�h<Rc應N!��'n^�|S�FS$H�XՊ�JH�\�1O��Ob�=YCb�/HS� ��[�N�����Wb�<�� ы[�ȶP�i4�,�7$�v�<�H_-&�2D�L�8^^@ c�*�v�<	�g�h���)6wp��B`t�<��fS�sTZ�
ٵ$�l��0H�Y�<��"܄A�8TK�[�$��q�<AG`��n܉�Ũ�@�U
U�3�"�֢<�IU%�E�f�9�h�uօ�y�̏ *#�٤�[8]>��t���M��'��Pf�<��9��@	�F�DI�	���$���y��!�-�7=���3)F��~��'<�1�&��� �#D�2����瓬�)�ܙc��v�jE�c�Po�t�ȓ��!c��n��Չ�����$	�8au
��&v�DP���M`t�ȓ5���j#י]�b�)�lT�"j؄ȓk:J���A�����.O=x>�t�ȓAlE����;,�	��KS�/N:����N�17B�A4\�oV�M�ՄȓuWBE��Ğ.�|s�F x���ȓ@Ԗ�Q�`��:%k�`ѾbI8!�ȓ �N�sφ%�j��n����.N�}�Re!K�(�P=p�����ͱ�&�J��-�w��_�ȇȓq�`�R�')�֘
E�Xa~x��.��K R��ʴ�ۃlq(Ԅȓ+�6)+r��&,`؀*�"f�,��D��E��
$�\����R7$�ȓ1��h�&���,�+��\&p�ȓi<��H�)�����l�n��9�f�1Ѩ�=b��18�HF*j(���@`jY�C<j���Ț�)��';�8�p%�3�.��`bڍz���?1�m@��B'����'I5����ȓ(  ,����HV�X��LӅ2\r��S�? 
u�%��4Q����MVfi��"OB�yՆ�3\��̢�K�	w��2"O`�A�5@�X���ؾ6���H�"O�� �H�g�ؘ+˙>&�2t��"O�]�Se��'2���r�^�b�UA�"Ov�32(I�5������T-S�Q��"Oĸ�r��v��k`F_K\�ؑ"O¸	w��{�>���@��"O��T��:����%C"f' ]�2"Oܐ"C,�F	>�)S�9�Ȱ�"O*I��3;8@�Bcc54� d��"OB�r)W�X�`,�� �6F�\�Ӵ"O2���A�X�l"�������(�"O��si�6l�v=��f֛��U��"O���Ƌ:bj
�)�/ތ�B��"O�lYq ��M�pS@�M�>�,<9�"O��b��!�:��",��p�"O������nL�H˼Kʒa�"OVe@c�7؈=!�B-��m1�"Od��˜>  ;�D�[�fH�"O�Y�s�0�r����(�N}�"O���,b�T�	U�		��k�"O�(��CS���iӰm�p��1"Of=i�j3s�&(Stb�9u�`"O�!bs��
1(D� �/6���"O6p*�ˑ���ի{���6"O�9�$�0�se�3}�h�"O��p� /K�P�n��|�	Q�"O6��bA2$ĥJ lW6b@T!�"O2��$�� �������
ܮ@a�"OD���F˖2D剰� 0kpT��"O\�B$'T#c���7*�3FL&�B"O�`�fҡTN�A* j��^��1�"O��BN4oI��	0OA#�Ԥ�2"O�8%hK���TG��)��q"O��9�F߮�� ͝n�����"O��뤈K�#������Eɖ)�"OJLc�&ϜyI�vf3!�2��"O��!D	5A�Qc��`�~�W"Od��wE�8����Q��6N��5@$"O��{v�$H)�-��!>@��̓"Oz٣!Òy�=���7j��u"O�P��[
��Y�ï�!)Tr$�b"O�Ec��<J	 �ZuH�g6,q��"O��V� ��ꦡژZ�]�"O����*3mT5k!Ts���XD"Of��C�??�.pJ�OCa����"O�ԏ<l��ԍD�վ�"O|�X��E�G�-H��M�r]c�"O�p��G0a\d!���G���B"O�D8��F�v�j��Q"Iĸ	�B"O�d)ԉ�	�r���8�ı��"O$����H+�f ��)�u"O��
5��\�J8x��@�mO0D�v"O������_߸���]<|N�ڒ"OȕҶ�ؘT�
jA[�X��}xb"OP����3�j���d���ѵ"O�p���R3A�\�hBl�2"OV�����[~�S2���h[bh�"O�qCq*�5(� ���&7L(i	�"OpH�K�#v9��X" ��L��"O,U#�K����{�o�mt�SW"O�)+"��
e|�cOA�a]�Ii�"OP�[���'Z�jXK��0PP�i�"O� b|8�Mʝ�6drsG��[11�b"Oa8��X�"@0�	�%�x�R�#�"Op��u��Q6�$I$ƭ^���"O��qI_�,� �2�ۯm�.�Q"OB�q�l��h(�j�>%�!��	"�,8Z���#j�ȃG���!�Ĕ�(G�Q��[�+d����s�!��֑{����W<%�h�t�\�Q�!� 39.t#p+����!o�9'�!�d�#t����J8���@���!��XO�:q���T`1B�>�!���9��-���� x.`[VA��!�DI&.�aW�)¨hs���!���`K�A�&�5������=�!���#~4n�:#c�>��*dʀ&!�d��'�6x{�ؓu��]��q�!�
=d���w���T�ڝ�nF.3�!��b�z�+�83��5�A�60s!��F!^Ot�8T�%v.d(s��1\!�D�7T9@��G&�	Re�$h ���m�!�d���e���ƻC�Y鶫޷$�!�D߽y�d��!&͠j7�@>h�!�$Y�/n�y��i�4O���d��3,�!�Ĝ ?��u�4�X�@�� �'��v!�Z�j۠��ӂ�#7XMs!�~a!�d_4V��P��JT�A�,̸#�� "a~h�������-?Ѥ�J&��9Y���aa۳�y����bŨ��P�\�b48$���y����4h eX��T�
8�y�Tb0��E��v���K��6�y�l��tmA�
��j�5�4dݙ�y"��衊�/n���P�GD3�yB��4k������!6�h��
 ��y"LK�t��@`j/%�e�+T��y¯�����I�k	�V
�2��%�yr�G4Kf�H�(<�N��T	Æ�y�aT+-�����K606
�:��1�y2i,g���2�&*R4(q����y2�Ӭ	{�l��N 8-����U�y2�ʹ[Uh=�4'2>k�=�#���y�"Ɨ����aC�53�5�r�ؗ�y"B�9	�(�!A��'�
-�cJ��y����vrv���KT+!�� �"���y�(B�A�%Ͷ��S�
�y���(N��� 0J
����(��y���P�|QC��?�^�
TN��y�+�%|�f�e��$N��Q���y�$�mAj}k��G)r� �*�yB�?&����/0̀u����y��K�H�7aׄ7��k�䆻�yr�.M�zq �R�f j���!�y��<'@����@�U�`PP� �yk�7|�f�R+O�vpCĪO�y" �:�l��Js8�!#	��y2�Y%*�Ց�F��u�m�2���y�#��6�ҥk4��$je )y�M �y2�Q��Qc���*n�(a���y��^5'��ƭ���y�`;n�Z ���Y�`�qcO���=i!+��0h��d�w�d1a����'���iwKQ�W�
#V��Px�V���,�@�8%���`�N�Ǹ'�zt�U��"U�Bl��8��-�|z.�/�-��hR���۷ [E�<�A�/A�&�����.R ��gT� ��:��R�v1�`� Z|B	D�T[�X�`/CX�Ĕ��ۙH(����$4�`#�D�~9"i3�׳j}	"*�1�N��ǃҗ2�p%����!�$�	�)� �l1�̅f�2� ��
t�P�#�'��m@A�E�T�����.@�\B���6ɶ}k��T��@6��$&mN%q��'UD,+5�����B4��`� M��K��s(�ٸqJJ	f�h����W�@� ǒ?}�`BԈ\9 �k6��:j�@I`)5D��+�F	�3A\�ɤF�n���G9!k�`{��Ԃ5F�TRD��ɉ��(-]����Mp��NX)2I�eqq&�"Ԍ���Mt��QB�  &��%B�b�bQQ��S#�0�a�]+�(i�,�fn6��I��hO@9��KTu����WcD�p.|Msb�'�&���D�=+��#A+����E�[��%J���5��|�P�U�:��}I�鞢��}bH��`�����#YT��
�cL7��DY�G��̻e"��k����,�_��[D+J�Y#pʧq�&Ⱥ'�ntp$�Պ)�t ��2lyd�zۘ���%��a9J�h��W�M���͈:W4����	_:0�C�ϼ{�"
�u)nD��ۂ'��H���H<--UJ=��i�~&u�Q�؎�@����#,�0�;Q�S4H��PL�XL$�iCz�'�\<y���,&�j�H5�\�H�'/�8�F�V������`�b��$�H�j=#�'G'�q�C������@2QyzX`��Q'<e^���I�
*j�8E^�����!�7(�z����RW�a� �X�"(�%v�X�E�
���AA7)�|��↉K��W�K Z �2r��>
���`	�'o"e���٦o(�t0�n���Mrdf�]c�Q�f�T�N$PO�Bl$u��f�'o(�`���Q2�w��S*��"0��I�a_�~>�<�����AD�g���i^�r�Ĉsp��'ɠ]�qbڿ1��yC7�ͺo�\ra�7/��+��^7v�Ҹ�F�$Ŷu�)O�1��@�R`И��f�4c��J��I9[��TS2� o�̴�,?cР�U�#���ц!�<�]xf�V��`3(�iᣡ��dp`� e_4���E"���<-�@W,��]���q0���( �Iೢ�u�R���m��Ғ�^9&�hS��D�^���YPA�!,
�y��ӘR�<�e�ݛK޶�"w�ݩ~�:�� e*�O�t��͢m��c��!$�<e��,J%5�����
;��,:���&ͼ�ɵ�H�A��Qf�>}X��Ft�(R&�DT*t�TP~}��J��p*��
.���$��	�B�����@mL�X!*I5`��`�E=x���T���D;� �
�L��`�VDd^����4�~��ǯ�1�$O !�B|R�	��'�m������6�cv��8��2�I�%\$�M��g� I�6%��O&�Ps�̮{��Xv���oUR����	6U����M�d�Q��BRb�$hXp� R��7��`�piͩ&"fa�F���$�<�0É��ސz"�W�k_|�,5��H蠩L�")`��   �nQ��5�:7� 8`w���p� oP�~�م/��Ht��a2�8�δVȚA�2i�C�ЕH�C��T�Lul�)��Pt��d9�,` 5�5f��x(�̀S��wޙ�R�E*T�h��� ;qR�5�U.�HK�RN�)��5CƦ��7$�c^uQ�N�f0�eS�,jӈ��4,�*���!2�G0i��Y��Z?qd,����	���G5m$��D�g�(A,�Ha�3�R�҆�
�м��b�R�	�!�ϭT��������%B҃�����B�}����սBCntC�SZ�Q��g$�Z�lDZ�G�%{\��UDQ{@�蕫�&psFyZ�gE�[G��'��X�bXb�U�}R���dP|L�8��B��"� s��^&$�fJ�/^����'���%T�@�������T�����A�[\D�"$�Z�I�Du�I�N
���U�G����d��P����;X�|��D��*��Dc��'@D�Cߓv8&l*d�D>@�l�����s���1ͧlm����E~���@���@����n��-{�'��r
���O&mo��6��>�"iY�T��4��ũF��Z�A_�'�4X£�R3�B�Y���
R���ENB%<]"1��O�zx�1��R�U�3o�!eb��7�GA� �c���;�nJ6�I�o�vq�kX��&MZ��ʣY�n!�Fב5����P��%ج8�U���j�pI����"IJ���"[�d1�&�W�[�z4�5$@�/��@�8i^ա��S��{E���l愐@eD4n�\�z��P�V1�)�FN�[ZH�6��*F�	c#�i䄘�D5l����s��o��ICW�?^.0r��px�4b�l00����$LjN��G�0C�[1�ƗP�H҄�ԫMyv�d�2���O�Xa҃�� �ē?Z�@X�A25�]����^�lYD}�%L� '�T�e�ɬ�q�m*�d x����(�V�[�\������
az�/��Y4����~k��jA�K	��OBp� �ԯ��O�d�i#�ݍY$ոF��n���'��)ڤ��V�X(��G YL���O
��`�?�)§X�v��*�n�����?&0��A&�;D��*�V$ �x�C�I.�)��?D��*�H΄B��u	�(ΞZD�����0D���ƒ�'1r	s���0�`A���.D��2 �	T��򮝠Cx�s.!D��wJ�C$�Pr��BVÇ.?D� 0q� �N�2��d�\�x�b�`%��<���哙p���#`�_�oJp�"gK��\��B�	b�b�iS%,.<����A̒O,���c,P��e��6/�\�w�υF7�b3O� ����)S����C&,�v�0�"O Ș�"ĞZ�|i9��׊k�5"O��cs��#���k�9:]&��"O�0�$jJ�j)b���B�B,�Ȕ"O"D����;.�,e`��(=��lH�"O�5�sHS8)��u�4K^�>�����"O�L��iܠ�aF+��_(&���"O�K��=hPP�[�l�=9��1�"O�X�BZ%ge4!0��R)�lT#"O�1�G��$4� �p�]�X@�QQ"O�ܐ0A�bC��r�3Y����"O�d��Ɏ�[ ���E��vM�`"OZ�3$Le�ڑ�C a*���"ON�����" ,�k�D��N��"O���U��*:Z����S�I�V%J�"OZdz�`Q.y�p�q!]$&	p��"O�Qp�.��%������@��r"O��S���q��)kb�>Qd���"O�;$J+��x*g⃌p�� ��"O��Jcb�Z�n�K$�� �Z�3d"O �e��.-�z���v�Pe�"O��ic�M1OJz��s�;od�� "O0�`�%�5'��l1���>K6"O`�BU��',� I�I�/.u,��"OƱE"��2��ݨ3HEz2�*�"O���Ǭ�%/[���FYl�|��"O�d�Gc�s�	��fhY\��E"O:H��L; �$Q�����[��i�"O�-P���3E5 e���
oi�"O���DNA.d�F�j�-I�S�D��"Od��d��UK��Qq���,K��ybK��R��̻ ?h@|�� ��y�bP�{LU�RbDD�[$�Q*�y���!���A͌/|�re��L�y��Od���`E�?p�X�9�
׳�yR̝��ZP*e޵w�\��a����y�*R�J�F����>2-^ CS5�y�E�'\<�
^�MQc�EXk衇�Q� ��;A���b����[x���I3R}�dF�XF��u(�)h����] ����ШɎ��c�a�e��5'6]�Uƅ�MsC��WSdԇȓ-���H�L�<Ԏ��7�(#�(݇ȓ�q[��ה��Cn�2��P�ȓU&V9�"�S$��a�0`؉:���ȓ&Vd��b�B�d�9@���"'��ȓ+aج�3σ�-Qt�$�݊�����"i
4�gCެ�HG�N��e��S��%��>sBC�Y�8+l��ȓa*�;q��=1b�
l�>4]��#dH���%���9§Oy�����būƅ�&��jc�^l�"O|�'Η�3|�8"�?�&�h!"O\���T�W�̛��B�>�&XQu"O�a�!�Y4v+��{_bqR�"O�"Y�����P�[[^Q�""O~q�t�B0��+�VF�:�"O��R�J�/
V@�媗}66��g"OIJ#靜$͊)ˤhʮN&���4"O~�� &�!'}VbE�@�j�6"O|�a�V5���G��B�ڸ��"O���!�ځ<��1��~�]S"O �©�=LxB�����u"ONyb� '� ��,�3;�  j�"O� �(�.V�T��R��M��a�`"Ojp㖮PIG�QHb
ևbOV�C�"O�tj�B� <Q1���R���U"O�Su�I��#X�Gv�f"OJ���d �BN#��"O�)�q�A;���ތQ�d��2"O�-�A��a�t=���Z1v���v"Oz��#�	?�	pE�{ܪ9�"O�9e�>"� c%B�X�"�`"O�dIuO8'�dQ�E	��1ٓ"O�QS�MI�V� ]�0b��H�r�"OI�i�?f���J�Ӑ��źt"O.�HSb�I��{e��"Ӓ�t"OX]QG���#�L�����o�V�Q"O� �ʒ�[�t:�`0�<��"O
��g�Ǫk&�H`�1*�n�C�"O8|��	*0�be�ͣ�� "O�q���7i�,�R��7&�q�2"O�Ӡ	��3r�h����lR4"ON�b7KL�`� ��U��Q�"O���ˆ>��4����|��j�"O�mri��N!Ҁ�^�8��g"O���@ƗE�>����۳O�fM�f"O��pn^�&���k�-�	vR0�"Oh}:��p{�tyk��Ѣ�""O,}�'A�3c�,9��%�"Q��-@�"O��Q���a��HУ�x�B�5"O�@x�@��7�X�:u���h�!f"OҐB%@Zq���S�@3B{��"O,��^�r�@EZ��7+h��"O��P�KQ�[`0�����)mm��"O$�Zf��}
�E��QF��s"O����h��R�D�e�	�NF�R"O$�٠��(9��Ԡ熖�>�(-�"Od��,w�P�ғE�m)�!��"O��K6i�����Sϡ@�V��"O���,K�&*�q@ ٘B��7"O<p�3ᛃ	5�����N�|T�"O���=J�ޭ�F��2�r:�"O��x`��e�4z#���iAMc�"OR㡢Ȥ7v��үH�@0E��"O��@��rظ���܋eRZU��"O���EJ��fE�u��uB�X""O�ј��=,�ҷv2�$�1"O��"��I53fȵ��
�fU���"Ov�[0j�"������^#4�hxe"OR�#d���/
b�j���%"��[	�'�8�4͛O�̙�D����[
�'vx+$$W�G� 
a��"�"��	�'�l@�o�.Z�ܝ���Ϻ�p	�''����$�h����
�z�&���'��i�q��0��q	��o|��;�'D|��#
�49����L&_��A2�'�T�2A֏*'@��P�x���#�'S��{���,�@����%K�nI��'���
�B�9�>|;@����(K�'t���OҀs�p%���X�F- ���'�Αkf��8;$=�en^�%�V���'f��QG��,���*�O��ji��'b>�Ҕ�N�1㨈��ʙ(U<���']�H����k��Q0K��y��'��Є(�,
��`ec�`Q�l��'����A��Xb�JD��f����'gp �"��(�X`FL�D�r�c
��� ��Ak�6F;� �DF�P�* � "O�AX��a@�܊"V��v�"O*�(F˜,Ղx	��*�"O,؁��-�d�B��ݲW��!7"O�U�i_�pD1���o\��h`"Oh1so��L/�(��#U�u9rE(�"O|�D��Q�!$ �'�*E��"O����<\Tl$�r�I�|Z,%�"O�uY���G� ,���L|���"O@��p����p
\�l�M:�"O��4��9�Fx��H�f���"O��"�8����Ђ�`IIA"O0���>kH`�I�!�P���zA"Oj`lL=���'�ϯju6!�S"O���cHY=������`���3"O"d�l:a� �;�*� ��9�"O��hjް|�ztC���.J�\a��"Op�!.� �����.���"Oh�FD�3�@�Qۨ%Z��"O80����>P�H���%�Ȁy�"O���5E,r3�%
�̵���[�"O-
�)Uu��̐�Ϭ|�*(p"O����h�6H����G��&Z�j P%"O�mJJ6#��%��{�f	 "O����Y�O$8n_#o�`���"O Ui�Ə�(ز� �Э3���q�"O��J�'v�>E�*F�?�Ah�"O�*��2{T~�ɧ�3l����g"O~��Ξ6}�p�����Lt�d"OD<�⮜�\�@�XS��+B���"O�qid!J�T9"8k���U�J���"O���-�<ΰ���xe�"O��Ч\D&,K�Y*y����"O>ja��|8����+9���"O�i`S��()gjPE�L�4�:<��"O��IwB�2��IrU��-|�Z���"O�����g�VxÖ*X�-�$S�"Oح�׍A>{�l��U��s~��B"O~����/m"�<�c��#e�T��"O4�:��	-,��	��*��x�<���"O�,b"A>y�f��dcc���P"O� H⎃�^D��P Q�,؈���"O���3��{����$��*/��1�E"O ���'$"��⦭�%�p�"O��ӕOTn,)a�
9�8 �"O@MG�ȘO��AQ �="�\EaG"Ov8����3&j6d��!@����""O(���Á�<�iH� �,���["O�!��)��!"t�ʨw��y"O ��P)��8��	�Rjʥs�p�� "O�p�U[�(s�$�
�#��ɷ"O�,�b�J�jO��	�1/�>�0"O�%hT���C�����M�&"O��K%���E���cU���j�
�b�"O��ҡ�!HK�X�gφ]\F�%"O(و�ǌ7�ʰ���+&�	�"O8�ae؟3��X#QI=Eql""O�[a	ƣ8��)�痂
�xx�"O@��I�+��E�g�*C�z�c"O0�"��*�Ȩ�FƐ'jI2t"ON��GTv"��Qp%�3�n���"Of��S��A�x�yc�$ޢ�7"Orp��P:l��7�e��\�"O�u�bH#�Q��U.zTb�"O� ���ç�?���Յ-@]�"O�97�@�xM�A�����!��"O��3D)_�'WF������)@"O��X�C�"!R�M�fd��8�@h��"O���%�ZI�QF�V��~�:�"O.AB`A)�������Q1"OLQ*���7QE�y"����>Q�R"O~8bu��$?Bz�X"ϕ9Ĳ�aR"O�ɸ �^�6k��DQv 3�"O�h��ұd�1��Ά4wO^�S�"O��c�H[nPօ��H¯FY���'"O�Ỡ�@!\zl8'�� vP��@�"O ��J�c�Y҂ �nWT8�6"O���s
�56
��4��9A����"OUp��[�1]�1pEn�2u.��S�"O�ՠ)�l�������&���"O����J����N�/:�����"O���OC?pŴ��p��k��Q"O��[F��j� d_i�.ݓ6Bd�<��\�ZMȁB2ˑ�I��L�U��d�<���ҁ /�Q��]+0��)Îm�<�ա+ ��'�۪j�^A�&.�R�<Y�� jn�L	�*4���5�Z�<�״
�ؒ�JʭGX�#&cW�<�u�S�wl�)ɑ
P/+�-cĪ�H�<���A�(�I�씨cjQ�W"�_�<����/(ve:���+0q���X�<�`EV1?b��b
\$.�~	�"�C`�<�c��=Pr���L�#��`9��c�<&"_w�@[���&A4l�]�<�e�26g*��ϏH����Q�<ٔ�,<q9��L�Ϻ�����t�<Y	�t�D�"`Q82�T���u�<b�C�4��4*f�0z��~�<�m�|�(��Ҳdw�:�i\�<	�d�%h���C�A�-#GF�zT.b�<i�d �1x�y���=���bD�f�<q�kĔ|1i KG���p:���I�<�e���@0����1h��q;V���<��f˫Q�b���(���3&�`�<�&|�`X9`@D�{+�4��c!��-V(i�@�ݫd�-��_<8!�$�V��8��ͺC��)s����7!��<:�!�����ф�G�!�� _j�0��Ǖ�]� ��4��v!�$_:%"%3b��kQʌ��iC&#s!�G���%A�Hf̘��F�?�!�F�hb͒7��0PL1P C��r�!��%d���J�̬�K��!�ď$hU�#�+�+66����Vy�!�d�G �!��fL7>4��Fߡ�!�D���H�ȭR�p���(�/b~!��4~QBD+s�K,d��h���<
�!�D�k6̲���vk<��d��!��&��(1�B�%B=2qt�>�!���<a�D�O�
�bS�
!��0CZ	�Ҋ,_Z�����N�!�	�HW�QägǦ$5�aD ҧQ�!򄙖>Lh@�'̻9�)xCAާy�!�R�rYr�Zd���G~	��b,�!�ğ�T^̙	a�V�xr�SoBxg!�D�[A�hA0$��H�J��g,�3{�!�D�B@N���ˍyK�����x�!�D��mx 7�QQ?R�32/�7�!�� H�8�S�}K����ύ���6"O�h�3*�x�j�r��ږR�$[�"O����"F8���'E,�|��"OX�J�m҅%ì��r!�>Y~�9s"OP��'܁�Q�����=cHh�S"O2�0�́"�P� �?N��"O�A�PJ}~!�/���|�2"O���=2�
�§MOw��b"O��`��ڠ&7��ЀM�3f��@�"O��%��'2����.N�A�k"O&92#�D!A.(���D*%"O��:��&X�0�	�$A�\ V"O�U�$�~�l ���i�j��"O^\u�	%�R�ckH33�f@z�"Of\�#h�X��ī�+ʣ�1�"O舩�L��J���IX�pb�<i�"ORQ���KV!�4� �e��(�"Op;�#�D���K�MN/F�*�X�"O�YӲH
�ʈ���P���8$"O�� i^hܼ�v��d��("O���E,�
wf�$ F��4��Y!�"O��z .��l���ĄM�g��P�"OL��J׋n2Rta�ƍ�A���"O�pb��_�[D����l��'"O~UZ��A�#p��`�DZ��r���"O����B̷x4��$�Z�J�XA��"Oi �S5}0	I�����S�"O~%xB!͢'�>�p���E�F"O��cD�>�(�7�Q�D�,�Cs"O���@��q����㭉*8- �"Oh �n&IϜ9����->��"O�})�+Җ�^-(,
�^�-@�"O.)����%np��*C�,���ru"O&��痫V(:�)�h�}�y���'�"��&8����djɅ5�:�Y2�

o{�<�����*/$#~�&R�]�0���ID~��1�V��10��J��ccR��*$jg����D��cHZ��F�uF59e�O�0��E�h�HYG@�0|��،4�687��3�44C1�l��@�H�q�=o�B���D%$!�A#I�D���P��+$JPJ���4ÒpA$��؟��R�O�to	0g*����I�\���� nW�a�{���O�p���0|*2Ϝ�T(@$�H�Br�@��J-"��A�"��&,)4�J�/h���}n�?7��A��D�h��	��IˊL/f��Q�P�H��ƈ;}2�9��B�
f����H\�S;HM�V�ѫ4���h�OP��QJ�7�0|��L5-��B%��zO�A0�A�O1��^��s�-� Qx���0}y�IL�Y�x�{����dZ8`����#��g2�P�"�><��So̧����䉀X(�Ĳ�M�+twn�q�] HH�6-EXײ�p�Ύ-�0|�p��L���� /~@��b�:�6��A��x��O�^�I�'L{,9�1i�)���qp��4����ғ���i ����*_�4!�U(��rĖ��"K�6B䉏9Rzyg���v��a�cK9�0B�	�H ��;�FK+Ja���!đtM�B�|q8��2ł:(5V����ñ�~C�	���K�!Q� X2��b��0=�B�I�a���v��"p� �A�C#��C�I�֜���F����ӑ��5]1�C��a*4�QJ��911��%Os�C�	�+����+�jm�&Řp�C��-S���s�:�^m���C,)��B�I�(�u8��<IWL���@�U��B�+ԼE)�$#$�&���_�QΠB�x� ��7-ًQ�$E(�ެghB䉨Z�x!�˖*ZD�"T��
�fB䉝m2}�F�'E8|i���'q�*B�	�T!I�n ט�i��E��C�)� � �F�P%���)ƹF�� 8g"O4���ɝ�R����gй�)��"ON)��D.&�]ؠ�C�a�
)��"O��GW�6�0h��ԃ	ǂ<��"O\����q���Q�hF
]�N���"O�]6�ͅ�R�F�0��y�s"O>t��h�:�@,�K�d�� z�"OLh��R=�J �f�D��a��yB[�V~�]�w D�� �8 �͂�y�-Ԁ[R��P��rR�d��y2��6;��h�dDMz��w���y�BU�5�ش�u�����0K��P�yb��I֩{��J :��c^�y�B�9f\H���5��c�'�yrÍ#|8ݪc`L�m|*`�@]�y�n��]|b����Z�ff����.�y"���R�bz�`QE� �1�yBG�	]�jlr5

o�^��W���y�����z�a�I�;⺝{���y�ҝ2�R�SP��*t|�S�����y�Θ�~i�F#"3���QF"��y��ʹ��l�d�1�lbp�ֈ�yRH�-F�H|"�
�X�X`ò��y�M�K��ܑ�����倢��y��ѯV�<�gW9���9�+���yr��,��	����ʵ����y,1ZM���[�h�B#�,�yrMJ1]�f1�E�/�!R'���yI,i��쑓��s����L�yҩ�L�@}�G�
����!c�y��э,^D͡��"���&I��y�%�"�b�s�[� Hhh��&�y��-	$Pc��,��Dp����y"�J%Q�b����}��H���<�y��Y������Ï+�����I�-�y�
P�-F�E���&���ӂ���yoM���������Z�CR����y�Oy����R"�Z�6�*����yXp��F��(&e��r�C��yR�O/M�$���*�%�4{DG��y�DD$:�}���T*BnѪ�R��y��m%E�'ȃ�"�1@MJ��y"J��3Pk�)vp�L���y����%$"�a((;W�h��&��yr���n�b8�7'S52����#�Մ�y�.SP�2%��_�$�\ �Ҩ]&�yB��m!글���.g��H�1*�yBƁSW�౐J܀4��S!�4�y�`��v��!�<U�����"�y2@V+V����@߂j:�Xфމ��OZ�~���/yfx{Q��A�f�p�<�W�M�50�	����29x0HC��j�<IE���9�c�ڢJ.�yڂ	�z�<q�@[de< 0w$Vw�*}�E�y�<�t*
>i2���P�� �FUv�<a2�P�+g42�R�]�	���G�<���Z��܄�d�[�}f����l�<q0j+s�H ����_	�<{h�j�<A�J�GFtu�W��l|�$�Q]�<�ׄНN��QCP�ê��qR��Y�<97����c&�G/,�U�E�Y�<iAJ��T0�hi�@��f-����U�<B���c�H��.�۠E�[�<�5e�c����ѯ�d;�9p��X�<� vX0B�۹X��"1�� 4UB}Q�"O�5ãEP?� ��\�5��	�"O��U��_�sK*W���$"O& @W�C�^��je̪O��1�"O��*CǇ�6�Y��M�~$h��"O�E�Ë,]F�X[�͕�Gp|��p"O`E�K(P\$�9��"O�Pp�i��{��ʂ��\����"D�h �6�RT�Ae��T�����M%D�P�2)�>E^����&���s��!D�4��\��H���C
V�j���e D�8�4�3SӼa�Ç:32li�>D��
5`�.}[@����id��#R�<D�$z�,�(s�n�pG�]�y�y8E'9D���Ƅ�cZ6��6H��
�A���5D��!3j�\���2����]h�lz�2D�8�En�6r���#�.ytpu��(2D�� �%�$�x���A�9@l�,9,!�	d���m>z(BJ �@r!��w^���B/T+3�mh�i�8;!�>
�X�x�F�,����H�"0!�!o����a��s��y�'(\�U�!�-^I�b��/e��A�D0"d!�$��|K���dA])����sǕYF!�ȏ�J-Q�I�`H (r���1�!��ӅT�2�H�QT(�a3Kz!�DD'<l~�r`�̲$���C�E9/C!��7xR��(��ש��q���.�!�P_^�ۃ�
FVPRꉴ�!�$�����¥�ép',��hԘ:�!�DM�l|���;�n�!v'ʞB5!�D�
�0�C6��OYJ�z��\�`!��:X�9ɴl�_ussB\.�!���G�R�׹$l���Y<dv!�DO��ó@�U���Ǝ>n!�Y�Yp5��B/a��YE�ԞP!���/�1� �'O��a2ǔ��!��T�e:�Z�HW0Y<�T
����j�!���Wڈ��4F�(9� �E�#5�!�܈uzJ�
�fE�m؆dSG#��v�!��2�^��m�Cо	��ǲ8�!��qEҼ���-$��Y�a�?�!򄉟Q�d3��%:)�QxWaN�3!򄂁�n9��ǧx��;B�>0ԇ�cb�´g@�3�ȶoY���YV�����&>�2-;�k�>W��]�ȓd�D<[�IU���|��. Kx]�ȓ~R�S�K	�:�̭��CL�L$1��Sޥ
C-��?B����P�F]ɇȓgQ.EcH� �X\�M3��u�ȓ,�>[���X�Ș�F��B8�@�ʓh�谄��E�2�b!�;z?BB�ɲE$n�)��Dm(�:$K� B�k���⟻O,c��T�^B䉩D��,��D�@��p�6)�:_ώB�	�S�H�n$Bw��r��\�%��B�	"g<^eð��(rʺu��Z�{s"B��3��Ar��	upժ�
��C�	w	�0p�Êfю��B�T)��C䉟R2!���5����'U��RC䉧>-�� �B�{�r�sl�5�`B�I9q��`����I�OwLB�	?*�|�z J_� 5~��2��
�vB�	=�����2$zD@����	jB�)� �,��NN��a:���eR~��r"O�AI4�;RpU)GbQ���,0�"O��*�_�g������z�ܜ
�"O������>���ФL���΄�"O�$����k�`�:4��
�L�{e"O6ar��F�H�s��T,{���q%"O8�����	>�T��5�C 5��dq "O�	[�%5�q2U�#m�1Iv"O���G+cw�P�g�K�H݋w"O�m�v/�6�Q�[�0�x1�"OR� �@�,+��!)��E��QB"OT�V�Z� $^tsfK�C�d@9V"O�,V)�Ģ0HS��'i@(�"O�u및�'y�ʨI�I�|
�Z"O 8�C��^F�,Z�� h}��"O
�9�h�:>.4}��-P�+�"O�A�� EQ����ȟ50<��"O��+���2K�T��ß�k���u"ON-� ���x�~��Է]���(�"Ol(�'ȜM�V��6Aםjq����"O�����ޑ�" о>R4��"O����fڊg��}cwG�/�!a�"Of��"�9)�2����1����"OPś��7mRl`��>,���"O�ЛV�\!��9� B�����"O$��(�Y�B�x���qq>��2"O`��@Ɵ~�
��ҜJ$��"O��)�'U�`��KĒ,F\�HA"O��V�J�<T{�)[$Ȓ���"OT����!@6�0���W�"��"OJ-� խ���0��;S��� "O>�0�'ڬ�2�.CD$8�a"Oz�ôώ�z��a�1�".���"O(L2�E727� N�	/��bD"O���T��*���9�l�*v#.,B�"O��Qf��m<�!��#HU`#"O�@�B�_d�AN6� !��"O6=���ŭ-���@�dT�e��"OR���jʒ6�$+v�U�x4J-�f"O&����Y*e��`��A�	)���"O, �fK6{��8tA��\�Z5�S"OL�䍉]�&��p!�9ghx�Z�"O�u2 N��l=�*a[�FL�ak�"O�d8!��#I�ؘB֯Z�,D�H�E"O:��%+E���F����Q"Of��m�M@4�̈5
Z��p"OPBa%Q}}��쑐\#���r"O��xPo�G��;�+&G!dH�"O&�p4�O�]�ǏB�,�;�"O�I�$i��\x�H"A�R�t!I�"OvH!W�%0ؤ3wό�ָ�yq"Ol��5� -���a��z�v��w"O���D�<T�h����Ϭ4�
C�"O����e�l{��c�
z�\ȋ%"O��C��>A~�M(oX79� �"O"P1��ۑ>?ZЈ`$ŻU���W"O.�bf ��L
�ŔQ~v5 "O�u
�-�-[�,��d�`=��"O�[�*h����_�I����]Y�<y�,ɲ~U�%��!��	#�C_n�<��@DF]�%��	,��" 	Mk�<��Y.?��LWA� m�tB]Q�<1E��,^�d!{�kC�$t�q�KK�<�f*W: 8  ���]G¥�@�d��yG�g�Eln-iWf��G����m�>x��w�Ӫ~��Xb�d�9#3~��CK���uj���OĀl��6~fR'�ЧW��#<�Df#j"���f' ,Hr�� !|y�#�f����{�<���hZ�;:���f˒1:T̓;�~3u��3�z�fD�[!�pC�O��Q��5���ZX���ȧY����.ӈG�9����),�\ص�N�X�6�0���!X R���L�X����E�S�A�	�;R��8�G�͑9t�����?[�X��S���s
[
�ʝ`�Ҳh5�8��>���( ��s�>�����m澼��J��޵(��Sp�s����a�6\钨ߙX�q���at6��A��� �:X���Q䄹
����b�	?R���
��ҮM^���iL�.���+�\R59�`U�vO�)���ӓjx��O�(sv�U�"�>�8���( j�:@��0`{FiRBO�P�<> ����u�}Pv��r�<Ɇ��: �$-شE��C^����(��je��c"˓JV܀jT�I��B	ᶦ(�i���Rͻ �ļy�)ƿp
B�Yb�4y����0l���V�1�^X2�,��2n�1BL2m�v�b���F�H�b��כe,��F�,�(O"�# �	}j}�J��<��4�'�0��v�n���_v4�P�E�.:�@ADy#�<[9��ܻE +������g�Ƚr&��G�n�sǊۜ8��'���b��T�<{u�fL��R���
$(�q�Ve�3ן�����;�T$����>s�Ȕ�S�D߹ff��!�)!��hp�ۑev�� foO�pD�q���I���=�'�e���r��۔+"�����"'�(#����EB�}'�H�0*܅s`�F�Z�	Z"��g�'h�H$>$ʾ���R9@�"Q����
CO��;bLʃ.s&�;�*S�/�~�p�$� ®(�b�R�B��	�y�&�
��@+	��B�ܢM���A	˓W8�%�:B���󂛥Ufn��2#��4O����X�FclD9���.;Rk��X]z�EfdH)��O��Y2�(�Ӽu+N��W�1O���!e�Г+�OFQ3�I#"Z��n�0�� ���0��jbU?���hP8��@ j��f����!E�����P�x)���	$.�g�<r`]#�,���S���kz�=���7gI�u��\�~�ٹ�����O��L�m�=���J�啖=n�T�!Eɇ]^�-�c_�PNu�U8�D)��6u�m��d�cx\쪖�Z�>�)��]�jG�,ƇE�kZv<���1t�m�K�etT��'�:�!�
'(����V�-XX����<�p<Y&��1�nq ��Z�c�Tͣ�)�\8����-䬌�ʖ[��Х�	�	�fр�nk��2��1��DD�OM�T���
;�Đ�EƤ�x�_�0�2#���C �%Pl����S j.��%M�N���#��i�%��9[�`A�4)K85N��8P�?�=� J�*��˥{b�S��MT͐�0��-��L�� �K�x`����Q��Mc���?�k���!��d�YVP�sc��=_�t3Q�I3=hy��%%\ON�P��O�"ªe3�T:&�u�aH��l�RL�7 iJ5�S"܇��L{��|B�>.�Y��J4��I� J��d� 1O� !�MޟxQ���d�MA0�T�#M���'R K�)XƁ�x8@pP�ߪ<��{pf��fؑ���䅂���g�#}*�w���#�`SwOt5�� Q��0���'2IP����9ݘ�R���W��O�9����F'@^|2�*�Qk,8@�N_�H+jt"�e����9P5ƃ ���;��4��������EC��HH��hőoc~@��
�8BX8t
���/�@ʧo�u��d>%��:p�xQ,۬M�4���^���W�ƶɆ牆_��s�֍�(��VaM��(�bʀ('Ӕ�P��)i����O��/��BbM��*��;5�t�{b�˨ ��D�O��a�B?[�.�{�홁@@>�{��$^�ސH��^�V��	�F�A�$���X��M���봡��-�����z�,�-ϳHD�� _.9n�ٹ�- ���֝ܲ���N}t�}�'8A��H
X�u����82� ޴(vJ	�� �(�"����$�d0��G����2�S-8vhZ!l�)v�-��@ۂv����hB#F��Q�Ջ[�J�1(�#O�0"TH�\�ax"˖8~Y����5P�2�&�
R�z��'���nvjP8c�Ītf`�`uk�9|\����gǇ1F���G
Q�~�ӷd��|�ڦc��,;��N�gN x�Otx3L�2��'Ć�c懘��X�x�K�%9t|AP��z/��F��s�2l��'�@Ɍ4�7���b��H׋B%8zba(�,�'��v�[p�:��A�O�X�6��(�v��u+��``t�=��ꖱ:,H��2fP���\.]�r-�p��<m��B��O��k��]������\pY��I�5�I/LB��Q�.V)**�Xb �<a�'́b��]*�/��W�dT³M&��6M>Ic��F�U�Or�!�DW�ξ���ޝ�%�$8ҐI�����g��CUOH%,��qwH�L�p� $�9P�@ʢ���M����/���I�-��i!��N�v�(�������ی˦!x"�0Q���´[)J3��0�[�w-�)ke,�-MH���$�	º 碝�U���d��)H9�q1dlB��dR�L��z�έ
���~Ð#eT�[�n�1L��<I���O٨8r�ƅ7]��f��.b�(U�&0tl(c�o���
&�
�P��|
�cƄ5X���檞,f��09Ej�rh#ɂ��p���I�b�,1�1��E�>���W���E�8��pk�+?���V)!;��b�I������A��a<�jF�۶�vh������
ic�F®c8�Q��-�����Q��4e2�z��ڵ�?��gLD�K�� �Ľ�I�)w��'��(�o���*'K�.mX`�`럁!�©�	�z����f��MC0n�qo���Pgݍ:2��*��߶�XPWf�x���S#έ�?y`ID�O��Z `B�5t��A��{��!��!� >�	�AV���`��m�(��2� ��3`���z��-��1�V�c�236�U�r�H6�\t���- 3Bc4)��T�`nDl��3��=��(g��'Zz��uJ�8���e�[��%�֒.9���O\�_��:��Z9�~�b#,U�С���دP߸��aHV�h*u���P�y�IB��eX���f��6:�
#>�O7MH�h�q��4�&xB�&��z��,��lM�].j	�'+��wl�y��II��@�E��"��Jǆ�}��4ɴ�6[!|-��!ui�ixm�S;
���[�5+� `�d\�	�4(� `T��4p���,~��q�MGN�)�m�Aޖ�f�A IX�P��,�)����n����P ���ޟ�)!K\%?�@�γ	0�P@��Ō|���A���0�����M �R��
ə7��1���O18�LpĎx���i�)��p��DA�@R����(Gڑ)�H���	� �XyR�M	G>�g�~����I�^e �㤁ΖHG~�0�
��,����O�pzBk�3P��l�T�ǭ7��U�0�K�"�fc�K�R��o��a�zEdQ� �f�t�L��D{�X�]�P9DI#����MC�X��#&	d��ʔ���]h礐���<J`�z�Z�cq�ZsC�p��ˣ'|����>Zc*rpp�#"�^E`��9}45X��x�_:<z�D`����ZY�	����sG�������H��	4qA���Ѧ�n�pD9�+�
#3�@W�Kn����_�R�q��9!X�O�ʼɁb +�*��p���D�6+�%�5�R��
�%
a�:n�ڔ��OBqP7�Ћ&��q�u�wl�����7����Q�G�.��()�&��(0��T�N6rU1�I`����F>/	L�`�@�',r|�f�\:����B`�%�I7e������L �bR�3.\Iir�MY`J�:h^��%�ۊ?>A�f��iֈ��eQ�hOvE���΍D[��S���1�M����:M�`uC���)ᩘ
uv��a϶U<d}������Y��W8E�Tu׆���Yy`�+��[�
U	GL���eGTi�I�M14ŋ�Ι�W/�Ա�#.醔�t��<.嘥Γ+u�S`�W	hC�����'%{��{%G9�h��&D��>AQn��=�M3`�,ےG	#NI�ԩ�'�����v�҉�3��j&r �3H��0W�\�?�0�f�ǀ;���	�u�¡���ӣm/j��\���9���Gz�P"��k��Ŋ���M�`�gO n��V*].;��E|B�^���S�]?Z�Q3d�K����e�
�6���@e_�@ƶ ��
����)��%r6E�Ey\К�j�&9����q�zUj��/J�@�fC�'�<5:���S����r�O�۳
��¯̶=D{5͋�(d㰪��.��|˓1Wר�� b��4��̷;HSE�xD(��GSA�p-ǜ2�Ĕ�%�P��<�=����(Cn ڒh�m4��V��jt� "+��P���^�PQ�аw�����3ti�M���K���z����(�<F��M�d�<V\��������s�Od��A$S���ɑ�P8�7�F�C<�� )�#��0� ��{�|�����舁1��BD�|�p���d��5x�T���H�R��-j��ŕ-V��㷝h�d��ݠ�J@�"%�N�'Cz��7%hՈ�/�-r��c$W.{/�Y�N���"�)@�pKtݢ�bZ�l���/v��kWD�|]|y�vi�V�N�"4ˈ�j�2���e�6n�t���T ZLDd+5�ݝ)��Q۵'A���yE&�O��+&I�Zu
x�j�RnB����]1b��}��ǁ����iu��M��	F��^}X(ͅL�LA��@�&��M	Ǫ�R�dC�5O��b�T""i�� �\�"-<�I�+�RzrF� T
�`J�Sa��AFY��"E��x��P��$\z��!�P�-WmZ�=�����6?��1jV�s0��43Xy�X����0	fN�#@A��66PaА
ï:X�	���U�jeXsU�>�SZ�	f@� �����KE�	@H�Z���[�Ѻ�����'�&��u�~�'J�-zǡ�/Qd�J��Ӳ���W�
�ϐ$�"%�-#! ��i��M17#�ӦM�ki�!�!K
ߦE)C�&Z���'`�,*�Y2�F1���PD�O�'�-���[�0f�8#�C���w�����8#K�-!v`��w�ћ]�`����1�x�����?�U-V
���SK�/%~p����_�d����*�R�	�M�81��܉���Wh����n�̑Q��O�XՈ�b�/w����I��B}�X�E-	)1�Ht
N"I"Jf��y.��ZG��-H�)�� d�N郧��)vvz���D� J&���>[�T�֧Ñco��ے$Y?M< �e��ny0i&板,I����c½^�@8�F�B`o�՛d�=I68��E�3B5r�Y#B�3}���3ԒG��c�#�6$�5��%�@�cV膎?\�l����hF��*�+y0���%�+R����H�r�L��#O�9V�@���lO��"��� }9�6�)s�m;r�ڌ�xl*�Q�,}����$�=o@�}�A�\H�="��ϼ������L2&�
�i��Y#q�=ѵ�]�S��;��@��R�Z�^*ܭQe��1�?	t%|�	���Q���)N}2�Epe
�#h�`qar��D��U��QP�`�	��	wi��5�m���%x�8��[t�����Æ�_�h��'IL�O�,Z&��0Wjj���h�?�t��a9u�G+]�l�3��1{E�X�T9vd�m�!�۲f5�<� �N�+�F�'�9KF�̲~N�0QM�;td�E��a���⍰xM�����K)���2�+Z@��f�^r��"�;-�x�K�"�h�I,\�u��5;��S؈���eΆ�ęC�ʟ�g�.و�m�	R�D �L]�p��sV*R�zێ��`e�ğ�w�( cdE���3�P/���O�#U��.,��TB�F�mZ���TJ������-� �0���\�:��%�]�����Ӣ H=�	R�g_���)�05���1X�4�8��������!�)�w���aX��O�[�b��=�G�$z�aqGKW[�tX&� }9LL��a�s�b��R��>̤yX�}�bA��!ߓ*I�E��l�O�M��&<��de��}¢�2k��(K=ӂ̠c\�'(�#�Ɛ ,���sm�;��Y{��81l �hK=׈Ԙ��4$/7���>?T���.՝R�3�䚆�\�sCT)�TՅ鉍b���q�ֹ0)^�%�y`\�c�+G�Kqf�3�"�Y��A�U��x@�$'�82(\�E+��{e^�S������cd�5�
m(�ƦcH08R�^z�'��2��� �*��ty�@��\:�d����9#��c�A��[ș�#j����F�Ŀx+0��B�<������R?9˓�Ϋ3�v`�dO�hMȩ��c8}2�I�sӘ��O��ʡ���d�G0f{P�9�G\"x�$e)����i�dŲ'@,r{�!�O���U/� ٸ��e
�U
��!j��u��R/xR��J�^��o԰K��8��N�F&,KE�U�.�D��$����a�{���sF��sz!�DĜU �T���M���co	�q�!����Y���ƙ��(�!q!�X�& ��xg(ˌ)̈IXG�(h!�$QC�5�!��2�`t�p��	&^!�DA%�^�bf�>A����E�0d<!��	�R<XQJ�1�x�;���2.!�$��M^ꈸ�D�*��]��hW?/�!���dD� d��o{�Ĺ�'�q�!�D��}�I��g��2<ʷGC�V�!��Y��AH�#��?zV�K �:j�!�$�30V܀�G\ ^h^�3�"ƍ!�dпY/2��	��rT�MXQG�!���$eZ���B�=[�!�EF>	!�Đp����}Al��G�a�!���e�����n�<97M!��/X�!�t�L$�rlD�_,�T
�i��?�!��A46&� 3% i��	e&ڥ0�!�D
2��d�%!	-[�@aa%�9b-!�d:����p�Xi��5C��l!��E$-���0�
���qD8[!�d��Hd�S3�)s%R���ܒV�!�dG�h�2:
�/�>�0s �gd!�[�*�
��*n��D�%�=�!��\&Z�<@QRI)��@Pa�s�!��E}��1oي.���tK��!�$ �'�*h��
K�1��Y
R���PyB莞I���+W��Bz���稔��y��hgL89�d�#@�����yr�ETT��ⲁ�yЃ���?�y���K <Ձ����@Yt�"�A*�yb��$"����S�75ΐ��DL��y��Q�|8���� �,��`��K׳�y��C2?�@��i"#@ T�2���y��	� ��!� )ΖH�qz�k΂�y
� ��`�BTr��𳯟.T���(�"O���� �nH�A�� P=�X�E"O���1(�I�!���	���XU"Of���h�!(��h�e��2g�|8#"O��ò`�P�"��IE�yk�Y��"O^)��#�G�t$j��Φ2K(�I�"O��w�\oz���i�@"�ň�"O<	��HP��hW��*i~Rq��"O�ax�X�G�j�0&��; ��I"O4��b�?=)ʶ� V Hb�OÙ"�)�����O�	�G�'>��pt�Ë#W�9!�"Oʝ;��P<ƚ��UJߔ{G�tB�'=]�S̙�\��I���cF�x8�͛{�I��@ɽ)����dY��<�g�30Ď�ل@\�����T�E	�PT��W�<�vMX�Q�pa��	�/x4�ï�v�>���7��7hĠ�J�+3�'xn���Z�M�x�sCÇ��	��	9M�|�{S�x���FS��I%�ߞiH:$�� �uO�!����W��陖��O&m{/�P��':�	����C�R���j�1*K��'����!bV�T�}�*�+H��+�)��V�yKc)�3v�(���
*��}xX�0�V3׈�9�䔅��Yٔ&F����
,N�f-1��Uy҇+J�6���� �gS>����� =u����KҸ_F�K����V A'���Z����D�
�/a"��.,x�:��Ã$�$y��j��@�1���.2�>4P�̒�J�b�!Tᚁi�n�Zc/B�u��~z�+~vp����H�õM�h�@Ҏ��V
}�| ��ִΪ!����H���'��-(�UG�8ʷM�2 &Y�0�N�ADjA#~<�Ԃ�&��h��4��͕�\@���Q!
�pF�&	��	� �P1?� U ���@�4������a�/v]@��֮�:�Є%�($�����Ĕ�f�`�����KSV�z�(	x�����[G3�ѯr�r`q�-ϭ;U`�e�'���iƕ!��ܪ���_O̜:S)�,u�vxq�mO-<Xjp�2�Ǒ>W���#��^
��&�Pg���9�Iʢ.z���o[f��%�2�� G�X��V�	���0V�ۀ,)$ D�M�m/t�� �Z�d��-�OԢ��U.Á:�h0uD�N*�lʄ9/�#?q��C�'Ph@*��$g�u��OiƉIC�70����N�+,���01�<�}k�k�&� ��r�	�uF�z������)��4 �*	�A���AE�)�a�8X�s/jr,гn>���� ��鈳G�(���'Cl
pe�(�l:�� #�/h�v�9f�
?&�ll����1E@�6/WZ��x��O��0��c�U�t%
Xѕ��x�� 3�LC�>�Z�{��A�[��Q����3�(����?t(d�Z'}���R�dO�(����F�%E��b�'�O��@��ɜ}��qF͂;�H��kL�n&�A�gn؟vb��Nʖ.�����Zy���1����9�D��̭o'�I�7���&�RL�VhiK6>�F�*Q�3�BA��$��/�*�[��YXE�%w� =�b�&N1>��@�	�]Q~7m�%^<ЃD)8�%9��.J�"QJ��Ɂ;�L�A�o���`�m�0�%9Jx"� �"4���@�u��s�c��F:B�{����x`�֏��;�0(�� D(�YYp�Gv��1�%L���2(�\g��V�
q�t��)g��0ᡢ�u9	EQ$N���"&H/�lq�cq�� C�<�nb�(����@� f!�D�P���!���q��A�Y�b���^0yy1��<�U٥a��u�D��eaS�Q�C�$ϟX� �r.�� ���p�6(�axA_�pn�%�@m^~��iV��.t� ���f���+'���8�K�"sn��ω�s`hU��	��D(g��( sܬرU3��'A�qu�2f�|h;2 ׋躰S�$QH��J�?��+�00| a�V�"�z���8D��wƌ�@R6���g�Z~$ai��W�vh�HY�Œ�|rR	�Gӕ�f�g���'R�j�]�)�B�Iۤ:�p4ru.D-O@��ēf"h��#i���#��K��YP̌*D�8B���9ؾ��d ��,�B�!X�<)��D�	�Ţ��
d�hQ�G�HX���E�2�������i���f�!~p�� l�q�N;Z�y"�A�l�	��I�B��MY'��$h�ą,O��OfA8�d��]�B��׈��,���J2��G����)�?q�PME�((�ĳ�΀��R�ȕ�(F�^�BU�'���P���~W|���E(J)P ��
ق�l����:�#����H:�f���@4�
F C0������%��)c�S,ZCH���0?��K/3ޚ�.�0 A��ގ2��JM�-���I���[y��x� ��7֊�B���6U�-O�PK�S�K24ȣU<	:`�0�BX�lp���}H�R!E}l�h�я��)�3��#z`έ���"�H z(�9�!�w\�#h6�#�'�����ĻF�H��NJ�E��39�'���ʍ?kh�(7 H�h�j��0�ܡ@�����ⱒcoް~��*�m��lL��s���8����m�2D#�����3�I=N3V��S>��B�ǟ+$0���T>��E�C �6�t���b}�'X?�LAAA%���fC"6���[��e*� M�l�0]B3�O��k�j��9>��F�g�@�7 @U���1��k�uP�NԀz A�*=:>��v
a�N���T���� �=*��ڽ!�.�*�j Lej5�'�(��j\yZue]�B�ԝۗ�	� ���I穖�s�r�e]�|�� �Hq�p=a���UY�7m��(��A-3�����9�-��$^��'�!���ڥ]��x# C�o�Ol��a��('C
��Q,6���8u'�ޅb�P
s�
�
�ȏ����D�[�@�@� �/��� ��%�Ր��D�%P˓;v ��|ʢ#9s
�Ч�W�>�v�:ujĵ�nU���A���1��V�W�LP[ۓ&q~��u��d�<�cpG�Y 0\k�D�++�	XV�ÿt�� �5O���a^f�(�#�g\	>Hs�T>�� �ՓS�Z��T)��|�$,z�	)�"^1!�ͅ>O�`���"6���� �U_��@Ӏl֦!EjqC�D��?(d�Х6	�vMZ��5AC���BH�O0�.9&��\*��@��$C��;L�H%S���($KK�5�N���R�$��L2%�:���w�p�Y�	�Y�J��M�vj��Y�
�� x�u�U�jw��+'&hݩҍ�D��[�J���IN�N��� 1E�śEnl���ti�}
.1cT>%h�'�%{��DMd�~�sV�J R��k��^%'h2 ��ӈdR�b��yx�(ӤE�`Z�0�v+H�B(U�#�X-��qX���j���@`D��<��b��چO:y��K	�L4U��aY���a@�T?�:c��넄��W ĨF&>ғ2�
�<�T`Y�'�Ԩ:�f27�n=��ޑƆY�CI�@`��$F+/��	��왖?�xIHd�O�-@d��"/^�uw�%X��c���I(B����.Ó��a�t�ݎGA6M1y��A(B�=I�~��(��U�n1�W�%,p�Ӥ�;��u17�m9B�K3%48��D�ʛb���Q#y��C�X�tAr�0Y�����/hŒ��1��8��%��n��~'
���LX��B��q�ځZ�v��W���j����Q����	��N֚|+��6L��q��PS�P�N���Y"� O%��O����N� ��O�́a�ҋ1���vO��]�Ԁ��
�B[hu{�@l�x�ɕ��Z� �qDW6GNM�v֘[�ʼ�5ʒDQxiS� To�r��U��Di��@A�v�1ǬM?_Vt�r�{��߮(2h���R��46kL�``���"#WBt�3PHS�!Q���3��>6͖�gڲ�?a��<9���[��	Cu�#��']�ċ+Oݡvn؏����`�4%�V�#W郵�M�!�C>}� �d��}� ��P1���|�X{�o�>w�*|��.Y�����`��02�Ś"1��!�0m$�� �mm�ĹP#F��~Rb�b��R�#3맑-, �*���ܰ!��	�m;aЀf�Dx�@�����@_�8	pV�ħ��б�	�m3q�P�\F�U���d]���L\�p�E ��` f+B�ZO�@��Dn�,O�L�¤��t�kBa�"9�89� � 7Ԏ�e�? 4�kBN!X ����*V��K��=!=�y2 Ģ4҄���!:� ��W|�	�W�C���b�x����*?��'�t8�FbF�<��mq�k WƐi��"h"T�#E�[KO�D��	 �v��qC����Q����H'~���+�5pV�;��[�HN�X��I�p��E�P�YYpa«O�$$���$�����?O$��T��J�*�ji
���q����M� (���.!����1��|�xc�Z�UC5�U�)��Q�g��3S��r����^����ҏ[~�E������ye���i��p0�b�,y��ѢL�Sl�x���p)T���A(�ν�&L6l��XpG�-y����}�!vG�*���x�a�l	FN�O��H�A��upVͧ|�<�Q�X9s ��P�0p��J��=]�yKag�	�2A ����Y�E\6s��Ќ҇6}��aaZ=\�u#�
�xm��O�<����`�%���H��V	�~�ۋ�d;z: �cĔ#(��Ɵ�� ��h��>�<�V�8Rn�iP+J3\� �0CM�l �e!����hC�;� ���'d�A�ϧB��e�$A]Z����!�\��'����!N�Y��HrDꚧL��@_�h��5���F��P@��@�\�Q����4)MG�$0n@�.1�����O���C�P�Ґ���O+���Ye-�%&��|�B����2P�ܝP߂DJ�/̧(�2t�Q��)����	$"��\�o��?% (�G�	4@�b���
 G��C�'L�.�L�gā���d�
� �T'�oʤ�ȱ�N�a��L��A�3KwT�3z�!35%˅H�}�3�5`[X�p3g�0WY�T���Y�j�pb,N(�B��5{�(AP.F &ў� �����������;"BkLF�-������sk�t���������ə+O���s�O��N���J�,�����mO�ue�L��OP��1q)�%��	5<"p!A����%�4��:H����Aݬ,���.�&�Y�cT[?�(�1G ���	B���3��U��(��Mn�X� �/
1��d٠k�h3��a��2* :��W#G ��4`�K�д��Br��	 �Hy���Ie�pQY�4�Ī��re4]*C���r�H0�٪
��R�K����E�O?)W'�]"�� ������d<|OX �p� �0�� B'�<���$D���<t.9�g�E�'!�UX�����` ��Ӂy�^���4H�P�+@�oA���h^>d0#	T�ў�@([.���j�e��H�剛,Pl$�%�Ӹ1����M��4Q�������[�(�S�
���d	�剘)X| ��S87����	1]��ђ��l�A��E�(.�����!ŷ�ēQ^����ji�xS�"��t9�%ؼ<<2���'��RdhT�X�b���4-�����#A�v�ie�� (�،��̎_n����6���z�eڙtj\����O½�ղt��Y��d-F��&݉|Y@�M��tj {�b�h̡̓p��yA�!�1b#T5����
zTDŒG��0F>�a���1(��D��yfs���zuUc� C�*MNՊ���
�Z�C���x|�)څ-V�`�8���"��� _���IUˇ���)?9�
ݺ���(X?F��W� V��������D4
�	Q)� �J
��Oډ���"2�n�@U@�T�(Ys���5�� ��U�ގq�@jR4R�i��J�{@}��m��6a%�Z�� � P�նۀQ��ʓ�T�-[@A����'�1NфSU�䘧i���%mX�wz,���Ξ>m��,��WҜ!����9��Y֫�J��%�6̓F]�q �d�ވ��	!l�$@��^�4��v�
N���B?1��F�j����UB��/�����m��Q�`���I�?Z)���J�J��)Ql�i�����b*����4M^V�v����n�Hu�ƛEl�p!�i&��F+4PCb�DF��&,�F��IN4Rtƀ$�T�ıp
���R"Dg8��∶g,HS���JD(!z&�$�h[f�E�q��$��Ut=1֍�8$0�X3��@%H�Rpq�P��0<�1$�j
2ij��)<�� �Ǫʯ �E�����	Ba�3v���bPa�1b1Ja"�;�J
� �I�������1�a�1r�<�C�M�4�ƥZ�ϑ+vtyt�>A�⃞"U �2�u϶�����V(B%�,��p��6s����^���I��>�0C�[�R�ND�@�K!����q��	7S��;�4h�q1$ޞ03,�w�:c��	���G_?g4�K��M�x������������sfS9Glެ�i�|O4d��ϟ�<a8�cf9x���(P1O}����DO���W�A����7O�X��L��O<p�� ~J(�	D�G��B}�Si��dO�����@+d�pLt�&1�,I:�M��Ǒɺ����M�L��|��D���� ?H�X;�*��7�~����OJ��4 �,PQc,Wx��� T�<���H\��A��@�╢
9=��[n�ʟ�y�N.��˳�=D�J�X��S�ˤ�J9�?q�-Ŗ/�V�qӥ�G�fX��'�n?q��-�`J�#4?�|-���K�U�������t:8p��n��i!������df=x�7'��sT�Tz^�AFVf}ZhKB���D�B툧��Q��ӣ��n�' �~�L�ʔ�?��8y AN}��׈1�J�����~��ǀ�z�X4KJ�?��xb �V9�,��T����cƀ�%h|���J�̰<Q�,�&O���CK\JGԑCfd6;7�����(>�Ƶ�Ą�bN\��#^:hR����K�LDн�� �;6潫�o�~�s��A�X����DE����ީՈO���B��)q|��0!��Vp����[�)�n��ŀ<��k��gɻ�W�
�����L	1	���a&?M�~)��Ȟ�@ˀ.mՓ�K���Tc6$�4ؐ<�$װAa�4��9O@k�H�7Cl9{���H��XKF$A6Վ{C$V2Dl� �4i	6`I.|����z2�놢Uvy��2���4Jj���o+P� 7'	�U">`�Ԇ�?c�|��b.B��ch�0?ǜ�kCg͕Z,��:����>��s,I�4u�L�%�[�D��c� 2�%��>b��
�-�&� ]ˑ�ۄ���r��UW�B�S�ްAH	Ǔj	^Ei�$�'k)8 ��^=-.:�O|ت����� L����r�c�j�7�K>m"((�m?(q>!"��xк��B.;�@���x�լ/���G|�%�! �Rc��+�������q[f(z�I?_a�	��n\�4��df�={�гe�زk��AQ��/Kk�����H��(�Vn�1�����<z�4�R�=���Pi�,ۋ�"�(���m:"L"3�4}�	(t�� K&�0��C�5c�t�7�� Cz-�Ԃ�*t����V?^�x<����$	X��'�)+lB�ǂ\Y�L2�+w�g�}��v�ڍ
�@�� ���]�g@�a6����@�`�)ݥ ̔)C���H���N���A��i��$�]�tbd�G��nx6|9��K0)4��j6LO�.MĮ��4��=o,mk�NF �!��f�O����f�7��QD�Z�Ii���d(_>=j&uSaA�F!�=��'��� ��1F^\q�DL��r�٧�ɘ[�ui�)0`�dY�(9�G	�s
R�Yǂn���Y{�x0�`٦�hp��b��RyR&фD�Y��~C��=���d E~n��S)�f��X6���hM���"g�l��*Lȃ����*AzHm��!�{�Lt��C�E���L���B��/�q��'�)A�]���"�>@�P�'$�<�J^�/���C�#�($��q��
I������D͒�:%G�<:�x8��Iə;*PB�	�/�L�H��@k
\�aHG�X�\B䉖3j�X&BQ��X�%ٺ6~C�ɦC�~��2D͓'U�`f�pbNC�q�6�HW��	J�\�t��\C䉐Ƙ����Ffd� ǤibtB�I(Hx�%�a-ҏn/:5 �-ؗ6�6C䉐1�4x�ȷ}+��
��د}\B�	�f^\
�c/l��y#o�'���Dl�x�7�R�N�|�
��?- ����V� ��n��b'd$�2��w�M��'��	�#
%P���ґL�ִ���rL
'���S)P>D�ȓj�t@QIˤ4��m�&�J��F �ȓTyxG�T#QP��[#'�T�%�ȓIp�x�E�)��t�$7�P`�ȓژbQ	�hG�c��ٷ�����	?�yU(�)o������,~��L�ȓI �0�&���>���6�O��!�䞙 S��R�&�����
%�!�Ē�o=��[���w�����Ǖ�!�6p,��si��l��,`�m�	u!�P0��d�g��*dB��@
�5xY��91K���ެqT@������(�x���A&T�$j���.4D�ԩsL_�1���;A�<��i��n:��aK>��N3��i(OJGziz�O�~�t��+�F�~�v���O&�<��R�E$EiM�m8M�@�˪Ә�'��OL�H�h�2RJr����αB7��;G	���B��4_u��aΟ�J�� �O���Y�)>5��A��V�c�t\�C��� ��@c��4j0���[�]N�tP"uc�z�,՛���>�؁��kG�R6�5�	=	Za�td˕Ry�|hE��~�>��`O�"F�X!�g�V�^��S<Q�P"J|�ҏ3�� l}�a��2
��ʥ�ԡszJL�w�'��4 � �(\[N��R�ل�$�����	�a4���#g����$I)Nk���Vc�,<s���G�(��[$��P���bվ~]X�i0/�D�>~\Z�a �O�:�E�Z�|���L�7�v�PO����#\Vn"�O��)�	]�B=�9Kg�?S�@qkP��~���#�O4���I<��o�L08g��S�0�AG�{?�p�������&�x��Ɂ1i���g���g3T�c�����֌_�p'X-rN<E�䪊'�Fac�	~�T-���$�<Q�o�P�T"�h�	�^����Rp�\��J�u�4�3�i�&�z�"�>yw���S�H��H!7Ě%V"4��'n�V��yZ��|2N�O�}R��OyƔ�,,�d�NÔA=�X,O����R�OQ>A��/���T���L��i�,�O��	u�S�?�`�(/�]#!Z,S��k�'������Ӭw�m�7�3aД1c��P�*⟐����~�'FPs�\��ᘊW��˷&XE��
W��Ï}��� ��'6���gϧ@�p�Ja�
Ut�E�@�L~�x�O���"�O�q�d�y'�hA�$�	�'�x���,E�jtzᨑ+%�f5�	�'�eP���1^,�0(�C�>"=��z�'.D@�bԴ!U�d�S΃0����'P��@��w���'���",��
�'F8}� )��gO -H�Ξ�΂��	�'7T3�^4^S��B7�0	 ��	�'Ϣ<D=���W��38�	��'q>�����2���Fe�(+d0��'�p�R������(M��� �'c�h��;a����U,D:�
�'���
�M0�
2)�>Cv��'���R�n\N-�� q-L`�e(�'�L���S¤ ;#n��lx���
�'��s5h�Jd��'!"M�.}��'�`��c��&�LYd�F�?��K�'� pt
��/���;�D��'% }��b|مMJ4�l���'\�0ꆩ�3,���!�>'$r��'Y����&��peE�#%����'H�ԓb������b��Y���в�'$�"goėA��z�Cb��J�'�؀�7�[t��Ņ�\n�]C�'�n���'�56�$��e��2b*D1��' DY5� R�d���l��r�'��l�֪R7{�l���/i}�a�'_���o��~4�� �#U�b �
�'���	�����L1��Ă�@9����'P8x{�GM�]�����9{�%	�'Բ`����6Y��ⓉJ�_�J��'�J��u��	X�6 ��j�!(��[�'_pEx��
DK�-�OD0�Z�J�'�oQ�Hu�Q�$ˍ�N�:�'��ڧ�]�):�(س����%
�'CP��ʈ$J��i��������'0�`zG��ߤ�K�M�,2�P�'h��t�I@H�4
�54��k�'�-J'�Y!FL�I�KW�==:�'w6A�����^l��K16���
�'>�) ��� )�=�2l�1+̖��'A�,�l5|i-���E\����'�%��oЕ`4���"-�,f"�Lq�'a h�Wʱ��yXbbӔ\��)h�'��iq���2Q��M��٭V<�	�'Ȥ���/��|?ؐ
�9;�(�	�'a�l��#�K�za���	8�D���'�����ʍ�ծY�f��&8����'mΘ�"��"F+6��N��(���� �$�a�'0] %-C�m���w"O��z�/ogB$x��;<�6�U"O|�`P*F%%8,\�UKR�Dj"O�����
y@�a*P�<uI0"OμRa�Cav@{�J%�PHk�"O���ׅ��7R�"��H3rs�Q2�"OP��k�0M��8#"_zBa��"O��B��=���(u4��"O ��b�)S��y�RaԹ]px�"O<}(rU��������N8�ȩ "O�9�b�ۃtp}(��_�<�8aU"O��b)Ϛ_���͕SҺ�"O�@ P�o|ΐ*�̒��"OعR6#
F�d萠л1f��'"O���E=kόA��ކ46��bU"O���N&^bEh�>��Q""OD��J�0�p�eN�3|L|��"OHq`�o_�:
�r��@-5i���"OڜjuMG�^Pf����	R\1"O&=ĥY�@Ȉ��]�Z��"�"O�#a��<?�9��˲E�H���"Ox�+���zv�pC��� y��x�"O�]T�Y�1��A���J��#"O�1�c�3���V-�򒁐�"O����T$Iޚ�Cm���E�0"Od��!B^	\f=�D!�8ߤ5Q#"O��U��8wnMʓ�E&;<r���"O.���.B/MŊ��I��q"�,��"Od1�4�U:�h�Bg��Y�"O@�XF���t�E�e�w6�Xx7"O(�6揟f#Lt�tj&@00+�"O����
V���c�*�/-��"O��J������zri�#f���"O���!�"JT��aЙp�IP�"O��c ڻ'��Mʁ"�$"O�\C!l����.����T#�"O���;QL͘s �!u����"O�� E�<����Z���y0�"OF���웶a ��T�O���"O���HG�9�Q��-۲}7D��Q"O�y�����c�m�5D5J��#"O�H8!YE4��!
�5}.�u��"Ou�$DK� FN�A�F)�D�t"O����I��<�v�Ŋ=�e�"O���I]ɾ)������H�����W�@6i�]�R����Dd���ȓG8�x6L#}�:Ĩđ&"R���98���ˇ1���0Qr��ȓJR\�r�G�&JJ��'�Τk>v��ȓ9��б%���{:���!������]߲1���˟�|��q��'D��ȓhL�*���0Oz��)_y��(��"lPi��'XZ��y��!���n�D���σ3ꂈ2Rcƾ.O�Ԅ���ၲ'0}���Q�$X���&��j�A�0Q����,�r9Xq�ȓ{��*��Q�"$�3�]���ȓ�~I;$��D2�В2�U�s�����*���D�w#r��	8yŤ��A��۳Oն���J���2B�j�ȓ5,X��V͈�i��H���R+#K��ȓ�j��lE�xn��K��}��4��3�( ����p�Z�Qb@��M�`<PlQ��4[0J�$�)��S�? �A����(\Pe�ʢf�0
"O^��q�7x#��i$��Ge8�ː"O��S*�(g��}"���&S�٪�"O�l�7T�o��`�4)F�$���'�X��m�0��H*��G�x�N���'�TdR�f	�#�i�MH�wb6���'���cd͑v<��G�y����'��h���$Z�����[T�K�'���y�g���^��WƂ$Z� �'��|��)+D4�A��M��͒�'��Ւ��	+<�HD��+��n����]�.����=.��钂�0:HH�� �,I�����$M95^�R�4��ȓ
�b���P�C�r ���?�6 �ȓ%<W]�z?A�^ZH����"O�}H�k5^���Y%"J�� 81"Ot�'�Y�6�� ��uTlq"O�UZ��Q�!��/��"&��"O����fGv"��3SmS�ZդHxG"O������U��iLN9K�"Ѐ�"Otlb'(�-p���+]3��4�"OX�Yu�Y0V�j(�R�/RӶ�BR"O<�:�Hԯ@=,�z7�Z�r�%"O�ѓ���Z��d�v�<�n!�%"O���e-�A���6#� ���"OȐ��hV�#�8`*�Aˎ.]s�"O�Ր4#��Nx���W���f�hs"O<���U�m����Q��"o����"O��K �!`H��q��D�@�f*O���܎M�hp�S�֙M��Q	�'��!�f�#&pz�ؕ��8A�t��'�"��q�H;�r��P�C����'-jV�G��_�2j��ö�yB�����Y�/�$2J�*��O��yR�גf@P���
��e��D!�yr�ȯt�XC�ဟ`Z (�r�V�y�b�8�$P��T��<��ǵ�y���0
>�q����J'FH�!���yb�6^�v�{��K�������&�y���4R��9to�3A<~$���I�y����J�(�9TA�D@�<�y��k�D�3�ں[�쬉��N��y�.�"��I��1�n@k"�Պ�yb�G?D~�B�CN	�@ڴ��y��r�f�;�e�9���!Ň>�y2F�=Ba�4�RM��~�f	�����y��� -ʉB�o����Fl��y����ZH�*���0k^��F����y��	��т)��c%R-вH��y�-'uh/ h�J`��$@ �ȓ>1>BA*�2���J�g�[���l�� cBlؙ?�l2�c��{��u��w�a:�
�<dKƸ§�;D��}�ȓo�vH�caFo�tn�!%��h�ȓC�L�4�W�?`��Z��L 'Dة����`���_8��H� v�V܇ȓw:��UB�M�9��dΦ't�e�ʓ<��o]�8����`Pj5�C�	&Q���j6&L�4�H;f��O�C�ɲ(�Ը�+�� r�O�|8�C�	��5Bpo�g,l,�Bc���vC�ɴm�A�#�R}P�d	�b�0C��:8�ċ���0���I��MN:B�I%.Z��rO[��z�Ç9�ZC�)� ��������eN+`'�Ui�"O�=��DW�.	�5��  $�"OZm��D�ie��L�%fģ6"O�(��`�9m�a��k�(l���b"OE�#m�h��lB�jj�X�"O,�94EQ�����Q��%*�)�"O �`qBT�j	�shKl%`lr�"On�#K3��iq'�U��=��"Ol�!%�N��&��c A�2i��"O��QHG�kF�ʗaC�ٔ���"O\Ě#G�P
ތ���1}�ĵ c*O\�LφjϦȶeP5E�Fxa�'�.qP�,�_A>�q�MC�1��'%�5�G_`�Jq[���Je� ��'}�4�e�I��������fpX�'n0;B-�#�X�yÌ� �����'������SGPIa"hB-`k�'���c���.+8����A�]'bAz�'�@�R��*_����j��k�'��E�2G�g�K\����N�c�<�D�@� J�ԩ��v���!�UJ�<��,�    ��     �  `  �  �+  �6  �>  �K  �T  �Z  'a  lg  �m  �s  4z  u�  ��  ��  ?�  ��  ş  �  J�  ��  Ҹ  @�  ��  -�  �  �  ]�  ��  z�  � �  a �  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P���G{��O�^����0k��	S���$5&bP��'��Ma��/l��ث���*%�u��'��T9@*�'��'/R�!�BI��'u~,3��E�*V����o�&.�PS�'w܌3n��l��2�,��HLj
�'e�踵D��o��aQQ�n�`
�'�:����F�P�z��Xk�Lix��$@�O�lm�d��PF�$���Re�nh��'��	D!^6d`^A��$�)Z�d���'P9k�س����źV�����'�h�ڷ��|ƺ�UMH�N沙��'���sb���8�Dm��m��Ds�T�����L�@�Q�bn�T2B��>�qO,��d�*f/04��BGj+ri���  ѡ�iӺ��F�¨C�@jRˉ^�]�s"O@�Ȅ��� `H��ԫ'M��3��'�,�<	R���X!�hq$��;A�,�ځ��R�<�G�[��8ף״o�|�I��V�ɗi�����>r�a0�C!ߦɚ�@J�
�lC�	֦-��8�4̻O��X���aP�6D�t��X��d��2�@�.$����I5|ON�'V�� pY`�� / Hu��D�U?�ȠE"O6�zS�S M��E�7�:h�X����%�S�ə2��=� Lؖ5�`%� L&o!��[2 zʡð��6:�<`��Ͷe���>�	�=k,�f��D9|-�G�
���H�'�A�U.C�sW��X��ާh"H�{2�'����b�Q� њ�鐠���i�J>���?�Ži��\�wB?� Ia����5d ��'w,�*4a@�^$Z��2L���-�L>�2 �Sܧ9���7a]RE^��o�9j��-���MC�MY"E���Fb�R�f�1���]y"�a��(��������j����F,{�HM��y2,+���c�#a�\��2.��y⠜�}� h�M�Z���r�۰��<���I�qԠ(��N�i����>o+!��ΛR3�u�c��[���̈́�$m�'�1O�}��qp��&��p�,�@�*�W�<�0�/�� b�2T�䘚ËQO��0=�mG����
��.5�|��gTd�'XQ?A]x ��5�Z���Eh<9��
,n@*���g�����#Nv}R�)�ߦ�z�ȍ�ua�W��2U;�A3D���˒]�0MQ��צ#�00�/D�((E��+�B��E��V��#t".D�L�CC��5�&�`��U/(B!�'SM*= P�m�,!�SC/4�!��# J��aTgI�~��0"� U����)�'%�R$Z� ��P��M�<���'YЅa�Y�|��\�ua��K@&E�H�L���7]ҜP�%~Y��Ր7 F����@?q�`K `؄\��L� kt�	�Bf�h�<�G�#Q�Tx�N��% :��H~�<Y�G[2.�:<�dAs�ܱ�]z�<�a�B�K?�U��!M+
(I�g�ty2E���OQ>�W�ɿJ��MQTL��SB��3�F9D���L��$y� )&-J�L�~�+��+��w؞L1�Ě	�D�����H`4s�)�.$uQ���\��k��y��W�V ���G"Ox �u�_���eH���GUVi�Z��lG~R2OHc?�ɡ
��@�bg�#��@�����\����ȓw���
dNT7�*�Q��Hz{X�'��~"'��;/|��[���(F��4�y@#Y+��S�16�(E,Ƒ!>�'�a|B�T!&.E+��I#_?�<���ز��I[�'[񟰉2'n�.�d=�rjN�{�pT��"O�E ��;���(c) *<:L
G�d|�6�=�O�$<k��	s(G��:'p0�'Z�AN2:"R$2�'!���y�'`5�!C�U>��)� N�jEB�!�'0y#�<K.��+ڧi�`���'�a���o|!�U�P�:�>`p�ǔ!�Px�c	>'q�y�UJ�C`�m鑠ַa6�MB�'j�(��Q�1���3�Iǐi=��b	�'
Z��𢈘��M
�.C!g�ܰϓ�O�:](yE�+XQ����L�b��'3��Gy� Gt��`+�)H9ZX;�?^!��U.i�P�Z0-ќuQL�ɓ��1U!�䉊a��5Qv�|"���)2Y!�ę83�RQB�IT�o�!��
'?!��ę+!�Q�d��"����1�B-A1O��=�|�&�N%��Y�S��	 W�M�<�C�G�|�P���P)1#HA�F�<�vGO�Z��-Y5�L�X2rԳc��E�<���Yt����G�~��T��]B�<� �xqe��^K��H�Q 5�^Y�|�0O���=i�y�NK-5��s&�g9yK�nю�yrO������	S4p�xY��Y��M�}��OZ�=I �m���Wo\U� �m��y�C�99��2��]��2�)Z�y�A	�pE��J�T3>/�����$�yҀՔ*�(��o=b�����y��J�G��q�EV%cKu�dj
�y�/<x�txZ ��8kߔ�����yR���t_&��� �P�؍�􂎅�O����wH"c�ݢH�x����&e!�Dװ���E/ħLu���2�V�^b<C�9$/��[u
V�%m��iR���.�C�	�?���)@	�-9��+�K�#�dB䉽n�4BNZO!�Y��ݞX<6M=��h��D%A�b�[�@ N��`Ye�5
d!��ٛa�Č"��O�JC8�#Kay�I�	D-�Bb�:yav�zá7 ���(ʓtI2�%�F��x�&[WG�$��z^�H��"S�2���Ao?dy����-�D&�~h����JQ^��=I�K!LO2U�פ��UŐ
T�(�r�i�ў�S��(O
=�`B�zg��Ya�¶b��
�'�T9������`��\�=����'8�>�	>n�e���p���#R�*C�	.)~Xez�#О>��}@w�S�58�E�հ?��郙S�r�[d��20G��"�b�'�\C�I[S����@(�8$�.HPf0}��'�F@X��G�I�3�U�y���'��(�T�4�\�p��ЋvFR��
�'�J%҂��v����bQ7e���
�'�0h)V(D)"�X�#�Ƌo}~qI	�'����_c3��J���3��c�'Ն3AA�t�l�Ȑ�ϣA⨹�'v�2�Mh��<� ΀�n.��'�z�PGY�u���� �˂H��H��'נ9RbIѫP`�Q@�ׅ6��+�'���0��(8��Q�g�.�عr�'�����\.v�}xRG+!P��'r.��*Ώ&��\�֩�&�X�'���ÒB��h���&�Kݔj�'$��9��܏�(��n�O��X�'2&Y(@�Q;nt"&��Ff"���'�j��b$�W0�L�ū�P���'eȨk�5��j��@��XR�'�n�Á��?&z@�qQ�ج0�6���'�LM� �G,u���!�ܶz�(=�
�'[ډJ�,�&���x�I1	[�08
�'�>ya����_�
�DI/1zHA	�'4�4b��#y�M����$%3�(��'8hHPhT="rMrQ�q�-0�'߆)�o()��ժ�@��b���'�bx ����6�΄�3��V@�	�'Ϊ���h�|O�@1�b�Xn�9:�'<6=)1'��f�Ni�c��U��$1�'zf*��E�� �����#ިy�'�@a��M_�o�i�L�	hR�<)�'��]:�"B
 �d�5��gsNT��'l�����\�Tr8�s��CZ�m�
�' \��&�Ĝ����QvD�j
�'��"Ԅ]�.�$�V�P�Q"���
�'(�x82훷@?T��b��H��}�	�'Y8;p�,4�zlq��TB�h	�'�zY(vD�6~�ə��ǩC������ ���sD�0�@Y���<l\r"O��b���%p�`�2V��QWt��p"O<ɲA T|�����Q/ n���U"Ol�#6��8��{P�:5c:|j�"O>I�g��0=��K�gJ�<U^0�C�',"�'U�'��R>e�Iş0�� X4���Ԃ��IxU���}�IٟX�	ҟ`�	柈�IџX��џh��?z����5e��(� ��p������,��ʟ\��ݟD�����ʟ��I;Mъ�R"�	{n(�p ��p��	�����˟��	П�I̟ �	şX�	����b�
I"k��A�ʞ������@�	ޟ��Iǟ���埰��Пp�ɶ�� �7��<��I� �#����������˟��	͟�������	�x����B�ҡ̐)]7�	�d�-5P�������Iϟ��	̟�����柠�	7_�,�Z3`B
7��G�Ӵe���I�D����l������ş �	���I"Hy�w�2K�� � �ܕ$lb`�I؟����H�������ϟ��IןH�ɛ=Fր)B���De�aeΒt3�U��ߟ��П8������	ҟ<�IП|�IF$�@㟼�(�pBhT�>�1���<�	Ɵ ���<�	�T����	!DT�=#�R< ���'���	�����ٟ,���T������	������;D��F�#1lySb�Ԡ��	���I�������̟�Yڴ�?!�=`8Q�ud�Cؼ{M�f
e�V�h�Iky���O��n�qu���Ƈ�#d  k'ƾwpw�9?�'�i��O��O�7M�NC��1��[�G!�L��a�*���m�����n�)�4�x~�=K�)�>W�OjAH�H8lu��(-�	AaY�y�'@�[�O�t�P��+�<襫��V=j�`��q��2�S=�M�;7�d=1�&Qp��)Cƈ=�l�s��'m�V?O��S�3012��ek|�tR/��l�Vl���µ4!�lIdy���ւ��H�Lk#�V�����'�b��HO�����*��0��'��s�I��M���N����z���<	q�I�k��y+��n�<A��Mۙ'���3<9rerc	F#E��Q���Uj��K��Q�"�ΚP���|@c��R��{���腆K�������
���)OTʓ�?E��'ܖ8If�W��
�0�\'[���1�'�7MP*d��9�Mc��Oҝ �ΫM��$�r�c�(|��'vB�ir�%@KН�O�t!��L�*��@J�vh�\��Δy&(�ꂪ-ex��=ͧ��"���!&e�E�L�8A���R�@�k�	<�MC���M̓��O��}ۑiُB8�p���� fJ֝�,�<����M��'��OZ���'=��3qdա
�q2▗ �J�Y��V-\�2�O��W�+e�f5��	��I(��D�*R
x�D�L��cd �B����<A+OĒO��o.:_��� m��� H���ɚ3d��m+z扇�M������|��?��4�?��F,|���mF�w��ݓ�+K�^N�#e���<����� ��9~���'�Tgy��b�M���ЪrD(��٢�g���ImyBW�"~"�$F`4=ѫ�/G�p�ŗK̓:x���3��$������wy�o&IO�!�ʿ.) ]�GX9��ļ<	ܴl����'��y�)�?�yB�'� ���L�I��9��c�'_2TK'�E�H��L2F+_�>ў�Wy��'_��*��jp@"Ǣ0���8��b��&�@�ش7Ub��<�)�D9sV�رN�J]C�hE�$���)���|�,O���yӢ�f���?�J �_4
�Ҍ#�BP�d�Aႈ[������eB�p����&�c���S�k��.�jt�	$:��� ����8��pB2�>Lm
@��V�O���*����`�F|��޴�~}�t+h8>��d ���O���]�dݸ�-F�]�v9�R	�9`%u҃T�<Ϙ�9Lx�C/ۚ#���I �R�q�,�3�@��6�ݙR��2��DI�'t����)ր�2��i�T��]��������N�% �^a�$I޸|��x��쏅!�(�@kW�x�8KD� �%��ّ�O<4Ɋ}q�+��zI8b`V� \�+&cQ�[\h�I<���?�������O��d��V��p�N�.���Ƅ��T�H�ou�'�R�';2W���mS�M���r�{1���=�� �Ѡ0e�Q�'���'g�\�8��ƟP��&�~jv�)}
�R�ǱpItD���p}��'+b�'��	*l�tP#N|r@�I308��P�0Lhi	B%K����'�'��	C��b?]��拣$2&l���E�cmt�m�z�$�O�ʓp�`�)ĕ���'��\c���%����	�7t.^�i�4���O��d�*>��s�H4*TŌN�`%:@�3=�~u %�i��	-�ݲ�4{b�S�0�ӗ��$�o�J��`FH7A������[a���'�+պ��)b�g�Ij9�r�K��f�q�#�AT�7�� a>|m���	ן����?��	�T�I�G�lk�m�R��1��pf̩�4*�d�����|
O~J�I�r����{�P�0န�0��׽i��'-Rf�'	�7��O���O�$�O�	ŊIi�!īw�u��I"����'/�	�]�h�)���?a���f�@tNOI��@*��(@���i�b-��Oݲ7-�O(�$�On��Yv���Ofؘ��U|����̛�'��uZ�S��#h�4��ʟ(����	S�t%W�|��Hs�kY;IW>������
�T���l�z�$�OD���OR��O^�韘�� ��(��ɞ���cg��5њٳ%��<1��?���?���?y�6����iV{g�,�퉰+�% N�=�4!s�F�d�O����O$���<��uָΧm�̸�FFZ�AD�2���*�^ȂT_���I�H�I�|�ɩn�h9A�4�?���kd�8�FQw�QE*���p�B�i<�'�_���ɍW�x�S��x���O��dk�dɡL����� �"ai�'����I̟,�	�^�p�4�?����?���d-B=YlMV*��ੌ$v�f����i�2U��ϓ}�,�ST��?7[�pt�D��y�>�y���`}���'��n�4Kx7��O����OT�i��
� ��=3t(�Xƺ��Ge��L,�'2#�1Jr�'��i>)��v����՟^XX�YTʌ,"��1�iozр�fkӚ���ON�d�"a�'D剂=P��3,�;�d�s�;N��[�49S��Γ�?y/O��?��	??���4��o[����d��X6tu�ݴ�?��?�'R�r���Byr�'�� YX��ש�?8J:E��Eڑ-��v�'��	)�~�)J��?	��YX�U)��B�x��m��C�CNv�@r�i�R��j
v6��O|���O��D�N��O�l(E�Ÿ��$�qŀU�by8�[���+h���'���'b��'�LҢ�Tu9��L� �{��1��A�P$u�����O(���O���O
����j�@�=)� Lh�i� r�8�d�Řd��Eyr�'[��'��'���Hy��IU��je����&C?h�$��,��A��ڟ�����`��{y��'[ԁ�O�Xha��~؀�	��2cI����Ӟ�$�O��$�O2��O�s��yӐ�$�O���v/©!�H4�D!;^��P�VѦ��	͟���jy�'�����D��_hf!ʧ��=~�x����=4'���'���'<b��4���i�b�'7"�O��l�H��� �o��1c�'e��d�<���/j��'���|n�w����e*��\�}j�/�&HY�7m�ON��"Dho����럄���?�Ik ��Ԁ܍x���C�Ŏ31��Ol����Y>v���O��$��#?�i'���;����C�2Z�����M�7�L:��F�'�r�'����OU��'.bMD�	YD�0g������E��7m�3$����=�4���(l&�ɹa)΋7��[v�ںk)V�m�������DR�Ĵ�M����?y��?�Ӻ#�I��{'J��l�0��0���Fئ���iy2�]2�yʟT�$�O��d�D����V�,�:q����5Yw>qm�����o[��M+���?���?��]?Y��_����!EN�N蚹��]1+$=�'��Y�yr�'���'�2�'Z�ț��Y��
&�ǹ=�x�J5�G>��7��O�D�O��Vs��_���87����P�BP����>T~fq��w�T�IΟ������	E��-M6^4v6��w�j�J���J�.�ʜ�.�N�l�П����������'�b _-����'~��k�+[%NN���._�'��7��O
�$�O����t��	��I�7��O���N>���;E�T�,�b z)�v���n����	̟x�'��BZ��dU��q�l�1)���PKLS������7b38��	蟠��͟+@i���M���?�����&��M�l�0\�$oD
;�\��4�?Q(OP���0��	!�4����6\}&L�C�8a�
�È��M���?�7��`��'���'����O@R��IΝ@3�M�\�j]���ˉ3 ��?��FI;�?1H>�'���2n���*A���4$�&7�6�U-dܨl�Ɵ,��ϟ����?i�I���I": J��#�G�Q~�,�Ճ#�,[�4nt �������	(�i��,ŉ�a
K��Xe��<��Ax���Y����<�	�h�!�ݴ�?a��?I��?��#�]�ք��!ЂnYO�,�nZ��X�'F�`����I�O��d�O�]	��D Y�a
�>ڡ� �����	��RA��4�?1���?)� ��S~?9���8�v�x���B����q)Ss}b��9�y��'��'���'\�S��b��^y�H��ʒ	�00Aύ��M3��?y���?Q�U?m�'l��N�!��K+>:쨐F�8���O~���O����Oʓ:좽��1��H����
s��q�@�(#�ֹ��R�L��ßX%�H��ß�҄�t�PIM�����¦أRQ�mˇ����O`���O����);c���ŷt��Ա�;it���Ǥs�N7��O|�O,���O��� 0O��'�j% ��ȓf�X���'H
�F} �4�?����Ā�
�%>����?e �O�$`��]��"��C�E!���:�ē�?���2P���S�cm)8�&L6b� ����|QUl�dy���O$�6�[E�$�'u���-?y�U� 9��3�!PZj��T�æ��	ӟ���-�S�'(�f�"�탑J��Ĭ�
R`�n�
81�!+ڴ�?a��?��'F�'�rÖ�9Z���vȄ�Gg��&�_>fB7�J���"|��#C.AA#e� ,A��0S��i��'#"��ePOB�d�O�� )L��a�!��)�a�D�[�'��b���F��f��埤����4iB�I'i����aI�1�0"
�M��{jI���Op�Ok,�^�1�G��*���8b嗦a�	�f�6P�IPy��'Cr�'@�I�� ��
;��:��N��� RR�0���?	���䓾?�7e�Dr���a�dijsɑ{#N�b�Ù����?)���?.O�AP��|"լ,\����e�(Xs� ���M}�'�|�'��f^wE��=N�����i�	�n�B��2�p��?��?�-OD�X�M�S��4h�bҲ� %*T�Ȍh�(ٴ�?�N>A��?I�i��<�I�� ��zG��<l���3��3aa��Q��i�2�'�2�'qX��u�pӺ���O������d#��S�� e(���D�G)�u�	֟��	3Ǣl�IY�i>i3�(�;ft�(��K P���@�4��tJAi��p��"N���H|�>����� �+�U"��<Y&��9l!��)R�X(F,T���Ё���&hf���j�d��q�p�=���Ԛ9p�� 'ΐ� ��p�X#�@Y���8�0 ��J �`�H�~�h0�?"3x�`��R����;��݄߀@Cs A,$R����M5H����k
1*�.�˦�O=��\��j^#:�^-YC�M%O��)������?)���?������$�O��k6f�z �5n[x)LIB��P6����ߺk�h=����f���.@���ÙE��Kk�\�T��\�H�� 8W(ġ'���Z&I�?�=�b�@�(�@� h`�x��\?	�G���DJ۴D����G���;_2ڠkc���G��#�@���yr�Z�"D��M}���b�hM��A������<11H�-ԛ�'}1���`��7$L��46�b�'i��'��
��'+�0�4$�!OM� ��Ϝ 216�!��"H��]yV'
�(� ����><OD�襡�8���R�
�
��,97+C�Gf�Е+]�0�b�8C�$<Oh�Ѕ�'�R�g���S1܈8'�c��׳6'��$&��<���ʝS�x�3�)ɭR�(��Da�<!�c�z�X"B�3c����!�[�<��iJ�Y��r�B��D�O��'_F���_
'g��6�9"`�#IΨ�?���?A�曆�BP��S
@kF��	V��t��u J�6q����zQ�x���Z=��!�v �y��ѡ�l�	Ja�����OYX����m�V u��-Q�,���O�n���MK����ja��#���@`�y��ɰ?*��D-�)��<�wo�\%�l�%f��?��m��L�G� �K<-
fIk��a`$��m\C�ɿ�X�r�����n��������'���O�B���A�V, p��vD� �|,S	L�z�EBRA�6X)��T>U�|�	�v`� -?ݼm{%��<m-�!0[H�rc��6�,�r��W��?E��\����0	,T[7�ǊW����EN��?a�����O>��7��yP��΍� b��>?�d�O����W�E0XYRr��>XO2���K�=6-�4@��4�x�$ū?gVx+�ī���S$�OZ�d`�l�Cm�H��O���O����?���>���@V]�:5ˢi�b=Z����Ӱ	F���f����|) �#�AF{B-��cF��^5
�(�"E�B��,25���*՛#�֘4JRa��hOLU[4� �+�vt��#j�;V�O�TI��'�"�|��'�"V�L�d@�'�� ��'�-�"*9D�$[P�Z��
�AgIC(b%�ш����HO��	�Ohʓ �n<㦰i�֨���$,(��#��a�di��'g�',"D��f���' �C�#U)�8j����8��БG�X���`X+c_8���O�w����P�Y=x,��-�N��\���SQc  !0+C'h��hkC��'?����N;��`�M�O���ܸu�����g�8cl�z�kY+`��o�����'���?y�pCZ:>� �K/O�p5j��1D��3�
Wn�"b+=t	2lp�Գ�4OE�W�$S3������O��'�e��*���HI�L�*�1�!#�?I��?I���Zm�}Ö�˳��}r����Ʉ7XQv4�@�%�
	;2��08�Q�@����*H��`B	�����&>A�T@�9�$S�.[�Z��:�u(�A�	�������O;�B�蛮H� �����:�hC�'��O?�	�i�|��!�,��8�t+V�+���$VX��V�t-���#B�᫡(� \���ɇr� ��4�?���)������O��Ǌt]4���EX�Z��L#�_�v�^��$����<��O�ɢ��5���k�$6�r�[<#.2dP�h�o�|����O?��A�8��������A��Ȍ�q��J�#�OL��$?�{��?i�ݽ*����Q *���J��<���>	`��+>��@'Z;R�L �`�m�'��#=�O��Zw�X/k-F����÷^���!�'b�ڣ�м�5�'�r�'���c�!�I���ɁB	k�Ѱ���8G��5b	�?�$�Ԧ�c��L�D����g�'�j��ȁ $Hj2�%�75�&�#��O��!��V: J�z	\������'2�!�Ră|AraBD ����ٔ$B+3lO����ׂY_���_6�.<�d"Ot�GL��Q�y�A$�� ���ை`�����|���Q��6-ܛ8)�Tk�n�7-AB�K�f�6�����O��$�O�z���O"��r>�"�`ݵW��P�Uz�P�QoD�)ڄ�$e�#8 ���D����A�"�3��6�H�^�.i��"W8N����'��qR��?ye@ԻP��)���?z	d������?I������IH�a��8���g�@��2�	�>f!�Ĉ
5Ep�0�RRŮ(���M)pU���p}�|rd8�g�? �`�F���h�h�$�>X<b�"Of= .ہs���@�S�qi�� "O<$0�͚C�  c�8(MJ��T"O�]���Pfz�]jE�� T����"O�d+��K�J�z�C
@},�p"OT�s	�a#(�Ĵ"x�p��"O(�"��W���{S!�"nlRYR"O���&V	�T�G�VR���"O	R얦֦X!�hWzP��i�"O�,K#SG���;7�*G�B(#�"O���� !d��ߑ綄Ӣ"OR � VS�@x�MF�hE8a"O
-�D��	�RI��E�c�Ĥ R"O����	# SX����	!�Th`"OB\�D�ȴH?p���g���{U"O��Z֢V�*֢@�7�V�⁩�"O���^�>º��%;
�ȃ�"Ou�Q�wܽ�p�M4i|P�"O�q�$Bv8Τi�ֺB��4j�"O��0Sc�(c�r���C�����"O<x*�,^be+!e\�mܬ�p"O�0�� ׅNJJ���e���D"ODh1����X�$����V�v��7"O�2��B?T�t)��Y5T�2��"OD,�c���T��e���>{�Bh�"O��@�d�x��`seL�z�Fub�"O��3EN;@��P�9h�X�Z"On{WD@�(�Y�B�w�q�"O�a��lT�5������ۦ��{"O�yB扐z:9 ��� R"=�G"O�`��6S����W?�k`"O��ڥΓ$f�H�ѷ�ObX����'�6m��E��'���т@��F)��E�&�"�s
�')��1d�^���%�r)�5�EN~G��* 2vc*��Ӿq(33��u�<!kPlF�N��B�I'<]fQ�b���F��(����&��u�O<IUhO=m���|�<�T�h��i�.^D������[<�Pt�.J��ԣo�@��C�'b�%I3�R���?���	3><5�s�X�>1p�ruk�N�'L��:���"U�����{�G_4=���L.�Z�bu�˸cv���I#1��C"\�;N�hkdl��D����a���� ]	�'���&�0��,�z)��o��9$���Sf�^�<i���0q�vd:4�0H�F���͘��7��n?��j�?
)�,�Ĉ;�B��e����	�S?6xP���(H��)��;LO<)Q�`�8��$f�)
U�^�9nzmh,�g+j-��~�Ě�OV��e!��%>�vE��2�S�>���P�R��`%����@��a��N�!����'V�v�I��V;bo!)"��ʒ`a�d�`�n�!�r� +$��v�Hݨ�䘚\h�-������ɭ
Ύ�������g���>A�F�l
��!�.(ld�y&�Y]h<Qt��^d�Dm�OcLy�c�7���i��P�>���� �O�M{�k�]��D�����z'`��JDb C��0=��Ib��I�_�
ًA$4�8���!��]��0�^��u8%ҲC͓X���#� �u��Ě-3P�Sᤂ�h�{t�	_�1Oh�yp�-����*g���ش�yÊT�1��J׀DX�o��k�2삖ɑ1S�8Q�pX�u|a|Ҹz�b10�aT1�"�� jV5� ���'�F�'#���dKF�1O�nM<6Q�g�H�)Y4��XzC�'���Yw���K�,����'t5�0 �O�X�1,�W��vB.�s�>����*|̭	bDǒ=P}����7��M�HXo���y����o��I0c��%+�K &@�1�͛�V�N�#�$?a0H�M-ȜlZ:PI����0�O��,�s�tK��V]����|��F(���Ƨ}Ӗ���k��.i�'��-qUG��ܐ��ȟ:ff4��U�3������!����I�.��"���d��#^�j�|r��[G>�l�/Y��Ŋ�Ӽ#��� AE���gD���B.YSH<14��3ʲTȣ��s�I��׹~�ax��R>-��6ϟ�T�|��3��sJ� tmR��\R����ECvF�R��'�R���U?�F�R�I�U>f��W��8�\A��̸��q��X�qe��<	�I�O�Ty3������O̲�4���Q���$)Ę��%��E��u�<��-���t0���>�h�B�J�Y?���M��B�m�(ַ&Pr�qgNJ}Bg 1�d��{�RAp�.�HO�*7`� UD���gL�i/�%�cl��2��VMĘ	��5����5�4%��U��*0e^��6j\fx��U�
�ʨ W�'�Ƶ�Wf�)m<��3b�B�0� Ór+1OT��3���:�d�a�A�%Cd�3�� ,l���剆��c@%A��Uo��wY���Θ�D�Qj#�	�9;��
�O]��>Ov��0mm��I�'�ᛷ#O�َ6MF1r.�����t��c���2g�'i�4x�Y%N �*$N�%�"y�}�MY1�P%C/X�|U��#�9��Đ
Y�x��^�ΠӢ���������F=��"��ÙR��u��8>]�Xb�+�b<�+3O�"?�1\Uj0X��]4CV�驵I�d���Q��U��D1���!E3n��B`�(gV�p�	ǓTM �k�8�
����G����뗳d3ʓ�ɶgH�p���'If9"�/K�-O�	�򠄗:�>Y��f��H�]#�׹d���O<�B���`a�eVF!#۴?8��"�'��<)��N��F0۶���ys�A�~�	{����b��=������(&[v6��'VLL�1���~����P�^��d(�߶B�JDJD�==�T�ԁX�"��l)4�T�t�������e��@"�kX�MT��r�_8#iv,R"C$b8�$��LŘn���sf� !:�a`cI�H�D����~���-��9;����}�9��Y.b- Ӗጓ#�a~rnI�3ل�p��W�=E6���"ڿ	���yM�cjԚ�d��;%��� ����G�|��*ʟI��;��O�E�:�
Q�Q�@y�S蜠6�azbF�! <��I;>�z,��Y)JV�x��� Gʾ-Q�(R<D����ܴgF�SdHص!e�@Ǔ"��un�\&�@��~��nU󇏻M���3�N���'4��7�^䟼S�Aq������x��e���9QKU���!L�����\5pq�-3�P��8��@˹Jy�T�͂q�tS4�Ʌo��4������)�`�\�}��T�W��536����]�OW��+$)O'z�>}s�`B���^�����l�����K�<T|8��j(lPâ�'�<Y)T�G/-���ӇiK3{3�-��̒�F�jԒ�y���#ڠě�����O��x�V�8^V<���3`����!�Ӣ6�����1&@"|	%KVǦE�F��U�2�YUdQz��� ���Y�-�M��/��� �� �</�n݊fr�I���
C41
1�ۧ,����A���K����?)��������R�! �7M��sxRh2ڴP�j( ��D|7�)(5d�,LטȰ�o��-3����ƝVK���.ou�Y�6�K�>�l�k�l�_��t��0d��i�U%ݫ2 ]1�ML�qN~	A�Ŏ��Ҽ(��g�TT[g� R�H��-̉v�7=�����I��8N� �+C7��=����7\�څ�(��>1P�-g�h86�{ ��2� 3�8�3􊇑e~���BY.GX q��|r6d�m��2sE(�@,6�*��"+Cv�r����)-����DF�vl�䪁P��M[�ݓ
���&��y�=5�W�sD\{�X�zk��5�فKl4zAŷ#)��3.��S��I�7�T}9�'�\xb�t&R���=�8bM<)"�:��4r��aӞ��+���M�ぇ=Ō�0`"ѱip���!m[=�BgeČn�؆K-ZF�QK� 4�R�F�-��Ր��$7KԜ�7�ҩY��N&c�p�`H�l�00s�&������J
^��{b�Ƅ7J����\c�DHc�Lz�`Ag_�Ƭ��C�$a�f ʠ�*�Okl�)h�X!�)�I�衈���C,�!� ��҂Q�t��,c�zDb�|"����j�i��`��9zU�vCָ���'�z6햌1��+�A�0B���C[Z� !��^&0� �f�O0�G�*�~� � �vg浙�R,>d� �޴X�A���ܜv�x@P����~^�<�"�D�,Z��Pw��O�mD@�9V���_M����-��E�� ��GM�	�UD̓)t����{���i'�X�A%~�����"��6
��4�СU�U��+@ĉ2i�&����4N�a���p(Q�h&�cƦ��N�pYd�¬$ς�ʴa�:bd��F	�e���Y�\)��\���(؁$$������Ű"ʄ�ub;�O��@7*Z.~��*���)��0qJ P�2��c�Ѫv骨��37������u1-�1bf�)�fr�a��d.E��x�q
U&',����'��:�"�3Vt�ą�B2�T��4�T1��"?o�\�($'F�}2`�qM�J%ѳ�̔�F�ru�#9PW��P* +OL�j��U�B8��7��4��C0�U8$E�'"�A4�Ed�\D* Y��!��-eR jd"SM.��6D��	a���@�.}�ʦ��oKd(ٔ.�J>�0ԯA�,�>��L6ғ��`��OƯ��Y e�@�MkT �~d˓g�-r��X�P����u��4�P�9��r���Z�VKR�j#�^~Gp���G�,&���k�,�v�����ƛH $uSr��,����&N-�j��FZ'�yB��?y����)�Y�xR�]PF�=��K�2���"��K�PX�ד=#��&%V¤�7i�1����^��D�#��	�px���jh� �w�|���*��!�s^y�ΝEw�7�Tsz��B0��l��Dy筂 ?�O�x�$د����'X����Cuyb/�h�Th�n�)2������_����R�4L�30�'Ubm��R�4����Z �dF�r��Y%y�b���	�E2xpBbl@�yB!V/^^����?Y֤��?��O��!Nq�P�f��(5�^1ra��S5�O��V�i�DW���lHM��@�!�\���M�d�Db�7���|֧y��ڐ�J�
�Y�p@���0>y���C�q�S�? 
X��D�!i̸�17�Mmm*�貤�\��bZ�U��'8�f@
n�̌`�Oݖ���3�6����a��=&쟐x��"<GF7�l�'O���O�-!���4��8sf��)|�����W����#�N�1P�6}u���Ee*ғE��a�)O?$�,ٶHC�*�h [�g����'�
T[C(?A�۲-��O��pQfQ=Ŝ}C���
��u��,�W��W��W������tz��1�. ��	�#ΡwW8YK�'?�bW�o�q�{?A��<�s��i�Ҵq��)��	Yl��7O����g�O����h[78��Y>]�"	�@�\8(�H0$jˁ_�����4A��	M	����M��O��v���C4�L�ʞ��׊��9T��(�j�z~2�	)�]�U&�05���J�s�L<i2�^Ҷ�t�_�j1�m�&G}}��x"O�f��%�ɂ�L�3�57��S�ʶh��-��I�x�0XqG�)q�m��}��MK�4���A�'d��!H��e�4�8UIځ9a�zF.�Z؞�<�y%���;y�Ƌn�������'z/D�$�b��:�rd tg>����վ%_6����><��8�C�݋=˾m U�E�L7 ���'�A�Όi��S�hK����O�	`pn\;��I�ɇQ����$t��Lh���M��г���dKd� G�DC�e�R�!�oRD�@�jf$��5��'b�Cej��
�]:�$��K����OK.��'1����*�UFxB���V�wc�
f�j�t��=*T�iuhU�0�֭bҤV���<�K�Tj�iX�Q�$ Vo���%H\�&�$��&JXim�pB0���$pq6L*�'�JYk0�Ή^�ErD���;��˅ď��<���\U��x��?W�&�;�c�Xh:�S�i���R��	�ax�HÁ�L�R�O���*2C�B�<|��B��=��5dM�B�d�)M<i,غ$��W∧/rV	���@Y�Ej�p䯕����Bp�lD�'��h1��:FY��@�4C��0���yDJ|����. ��&��-d�P�C��'/L ����b؞	���f����J��,�h�g�X��en�	(�{Zc`��S掍y�8<�$\���/��<q��)�S�o���Q�ٔ{"�i��ĉ4�T�d�&��<i��ԩtU�`�,A�L{�� O�>��S�P6=�V����IQ�XثQ�-h�})W��;l�x�D�P'o&&��mj�YE�Sn�*��[A�i��'#�l��O8�̓\ļ���ҡ���EK�.IsȘ�'�D��%���3���� ��T8���?%���b��_�5LM���U�~p��I��d�'/�ď2ݛ��O�u���I�<�U�D�5F.���MCl�D|�4�ƞa�L�[g�it�h
�?��,x2n�lXp�ڧ��F#���W�̢gcvp˂�i{4U�شba�>�S!�9�'^4 ����P!eo`u�ȓ?�u�bt�1�^#Q`�4�7���t����iD�ɀ�p<I��'NC�����h�Xء��Gk�<�S"M�*ͮdq�D Q���ٷA�e�<	�h�4K>���AlĔ1R����v�<��σ.N��	��J�s+��0��q�<�筍l�6�x��G�_�H��3!�D�<q�Ď�Zwj�ʷ�V�<�@0�1K�e�<!&	ǍR5J�B`�X�EzRt��`�<I�o�c�V�1����<Z �4g�a�<1�,6�: ѷ�m\����e�Z�<�MU7z�b�Լ\ �-�(KL�<)@����hQ0��9�t�dC�K�<����)�!2�c���	a��D�<�S���d�f�!��V� V��|�<�eI(o��1���tV��(Pgr�<�V�i��"��-z���8�di�<��gL�bb��R-K,=,LP�`��d�<Y.�e���"EJ�8�^��v��g�<y�M�� ��Z��өT�����fFg�<	1�8<�\ ��:Z���bb�<�d@��sߊ�ƀL�#��y��VR�<�f��9��9b�Nդ�X��h�<�rlS�x�P��Ң,K�x��e�<I�d��i<�T��;.����j�a�<y7NF�x��ru*_x��C���]�<YTC�"mj��مh��v+�	�#�Y�<�� �2� I�Z%lX��T�<	cB^�;!�Kp�I)P�
��P�<�d�/0��(�Ґv��\��J�N�<� �m)Qǉ�?�4q�3�V�{���)�"Ot){�ĴM��Q�s�݆x���7"O0҆�\9f~xtp�Ir}�ѧ���<� gR,:�0<�O�W�6��5�KP�<�� g7�1B��r��$�/L�<���*
-�&k�	�U	��ZP�<� 'F=t2`�@a��\A��F�<R�ҚTtfd*�m��05�Ů�k�<�b��-����'�G��H����e�<fl��!��iTC�P���0�Xe�<��.P+8+!��ݽ^%*m���\�<a���Xo�Q�Ӕ2־qSr��n�<Y�)�~|�8�ÚQ^�@;qhg�<�E�ٝ��y��@T�Ԛ�J�<qR�ɄP�t4�է��@w���d�
H�<y�P3'��c��(�:�j�J�y�<�A�=�����. X��x
[<�yr�K�츩��ɚh.�����y2��E������جȶ��-�ybAC�: ��ؠ.{�^Ѻǀ��y�["C��A��a	�H ��kLI�y�dI�L��1	�f�F��uS'�yb�֓7�Y��R�B>(]�	_�y�E��%��%Y�ڞC~Qᖂ@�yBn��`ߨu��3:��ئ`^4�y��Z�[��㎅���LX.۩�yR�_�F-j���S? b
���(п�y�Je��D���L�wV�LI��G�yb��:��=9`��!cu�8g���y�a��0�h�tɔ��%���y"c��>�:t(@���L�R��%(��yR	��^���ÅF��R�X�UBA��yl�& � ��*@��0x���yb	�C�F p0�I#'U�]����yr����	�`��1D�a���R��y���[H�y��*8"U���W��y�̮5�DCcķjZ^x�Ca�)�y�l.h��Ad�3\;ԁ:�C�<�횞H:x�`5�� AD&P��"�B�<�5T�&
��aU"��|�������W�<Q"��4�z�O�Z!�0G]W�<!��\bd᳑�1Ӥ0
F�E^�<���O�	D��! ���Hzv����BS�<�'�Y<�|�K��}�VE`��Q�<q�]�@ l�jQ�Qy2�h���O�<�M-eo��񫔍_2Pa ��Xe�<� �� V�P�n��eZB�:��Nc�<y�E�LAL���m�UZ0C���[�<I�ꗿTp� IL�vu�;��YX�<9b��@"���I [1��]�<)�1&	H}��!np��%��Q�<��-�k��ᢃ��1��i@���O�<�=BĶL��	,97��;��a�<Ag��9�.a�)%Y�����G�'�xBO�U�|)�C&,�F|;��O �y�T0,vL���6tx�6C�:�y"j�F��<���օX�|�Iv�Ø�y�	ٟ+ސH"
��ZVd�tKI�y�C'�p�a�׺S�X]9A�K��y�(�{`��F�=��: �\��y"�ژ	�)�([&/θq���y��W�p8RA�����qB�LU��yR�Ѓ���ئ�L}bQ�͇�y�eN�PS~�2I�; X�t�W����y
� �M"V�^�}�hq��L	�m�����"O�L	Fi�B<*E	�m
]�"O��[��η
��U!�N�q���"O"�X���,�^��d�	
.���"O�l�G�M�f����>D� Y�C"O�)PA� D[�l�!=���d"OH ��)s��`���|�h��g�$0�S��K�kN�$��� ��}p�J6S�!򄎉,���r�I^� |�1�F�6n!�$�7�`���_�wn����<2!�D�9�|2�li�-0��"1�D!�S�Ow��9����Xe���`^�HQ	�'���E(Ҫs�:@�*��^L�'6��a����TH�!�:y�\��'G��Qbe�Kʐd����~�v�I
�'����aT�n��v�-P���	�'�D�'ւ#`~�-q���� ��q�<!�@�	j�i.ރ����\m�<���U�6�E"�������%�r�<��
����g���8���
S�<!G#`�d�梌>em��#Xg�<95;!9�*6K9yB`�T@�z�<��@Ūn\<�5KB6q�t��NUb�'��x���T���ӚeG>�	�Ì��y�S<��������-z�-��y",���z|[�HȞ|�p�����yB�˲Jb��۵ɑ�l&��K�ɛ��y2�ӫz��D#��9!������y��:u8h)�@��f
�#����y"�U�s�$s0$�eZn�Z�ö�yb@ِ)L�a .8`y������yR._8X���93-K"n��[�d��y��S�zV���g͢h�91E�V;�y�-j��	R&�8IY�(䨆>���hOq�α#��I�����!��Vk� i�"O\�x.!M_Z���-�eyBE��'�ў"~
g�
q����bL�`��dI�.�y"B�{�������S:J�c��y2�ʩn�QB֋<9r���r���y2�A-S��9C6��.Q��QNE�ybI��(��Q:c��r�ҍ�$����yҠT{� pi2d֑ihQdQ�x��'�<y�Pn	�GB�)��/p�d(��'5�r�~�����*y�)�5�'����^��)+��	�D����l��,Y!�d�e���[��h�r�8�Z%*U!��Swo��H���g�`%H�i�B>!�d�9`P+ ���p {G(&{M!�D�l��Ȃi4P�̜�e-��qH!�d.�Z��&mT�,��@��&�!���<K�BFBԕO��V֎q!�d݃cr�T:D�V�XlRlaŅ�*nQ!��:S*��b%��a9d�T�!�� Kr��(�J��B)`��`��[y!�$��� �$�ߢD+t�uj-C!��'B��C�K?�U��A�!��"n���D�o�J�$!�%{�!�ʾA��f�����������'��qct�C"}E��"���t�`4(�'$*`)�3^��4ҳ�\�gQY�'�,֛1X�����`l��b�'0d ����I����3|}��'��B&,H�IT�i���RV&�y�̯\���-�x�)��ǓZ���S�? �L#�޶o�D�BwE�5`�U��"OV�o��I��ӂG� ��"ON4��
J���3�Y�4qC"O��3恋"p�p���B��X�k�"O}��䔍`/J��� �Iz�B"O��C���-@,� �[ъ!m�.�!�D�=U�Q��M��|z����Py�ө�� G+�3L�a��V��y�kԷi�� ��F�`�#L��y�B43G��S��A���Kdn�y��ҧ?V`|���Oh�$�8Ԅ�7�y��ǛV��%I�� �x#AN��yBjӤg=0}Ʉa֖87�آ�N��y�D�p����@1�����yB�:5�j<�&Jk_赫�,˨�y�l��f�_����*Ȝ�yR�X1Mr�ID�ۤ*�~��c'��y�� 8��L(�D��#
=1���y���4V���d��k:�a�BD��y�M�j^J�N��q������y�˞
=�ܽ�%%�- �41����<�ybH��J0Pk畧t� ������y�MY"Ƭ�W�˞6s��+��yr	7l�`K42�r���OY��yb��<r��)�S<,:P@P���PyB���H��(ce��U�p���BW�Ij8���u��98�B�hJ<Ъ&�+D�� $c��Pۥ��&��}ꁢ,D�L4��}���B�V�;���14�/D�@3�F�=�^ٳu�߲[�m��?D�����W�7^N�s잁 6����<D����J�W�b��WÇ��t�m>D��bb� 3*T��r
F�QT��ы=D�x�D`�%hQ���D�םQz%�u�7D�pF)v|Q��U� �`���:D�`I�͟�4�^�(7,U�}ex��<D��8� 	&1~�X
��l�f�R7e<D�k�則��50�cԱ+b����'D�d�����CѮ��K�(Jc�ɐb@"D��9�I����ei4�V����M!D�2h��gd��׬�8Q$��E�;D�`��
�Y�t��O9��R��%D�p㣫�YpCY1�t��b "D��{�	V����3&�?^",��O:D�@�ϧG��a��ȫ9v d��7D�$Y�b��v�%�A+Y=*,t8EO+D�+�I�e̢�*eD)QT9��*D�L
p��F�=H��߽!��y�E�'D�������n8^jS��a���:D��Y"�P�� T)��/D�U�`"D�����C�]��M���n8�:�.D��ڂBENK~��#�g�;�B,D��@8yx�͎b�!�)D�ຑ+�%A�l�X��1��(�r�&D����E���AT�V�%J5���7D���Mۚj�X|r��y|	��B:D�(y����R"�3&@%hr��KC=D����ݛ}����7���e�;D�(`(	:-ͬ�h�K�\zrl�dh?D�@�/��/�Ua�K�+D(���=D�dS�?}�(�t��
%��)��&D�PQv(�8kf�b�8���($D���1�r�^��#���PX@�� D�<��'�_�nِ`a���6�"2�=D�� \�M��
�	s놯���(�"O:��tA�"z{�����-�@��"O��z�\6ƭ��K;L�8R�"O��AQl3L$>T�FI��
왃"O�\7�J�������ՙ�"O*I DA�ox�a�!P=Se��k"O>qы�;��y!�\\\|0`"O���abQ���ƶiP����"O�5����}��e��m&G�X�T"O�-��oF6�v�#����K�B�6"O�A�G�	G������אd|�""O�tZ2�3]���с��{m�ei6"Or�(d.
F#p�v-ɦb��&"O���ɲZ� ��k��j5D��"OU����d��q�(��R�o
#�y���)�T��l�7l��"d�Y��y2�M;J*��F�W�- d�C�Z��y���O_��I�jі#�|qbC��y"j�J�<��
"p��"�E��y�$��)	��d�ƈ&xk��y�gJ2}��
gE׃&���;G���y�ʈ�ތ۔�.0C��Z����y��E�^�R ���Ðu2�u�u"ͳ�y�ϖ�:9@I�� ��l9z�E��9�y�#A�i� 0�5'�^^]�s.��y���-ZK�TY�	^���U���
"�y��K0_��=k�$��N!�����y�fę7Z�E8 �!j�2P�IƏ�y�Z3�*���@�/kD������ �yr��cv�!k�&n�Pe��
��y2k��(}���ʌef�I��N;�yr���ܡ��/?a�~	;�E%�y(X
Wİ�,EZF��xu�Q��y-��Όv�ݚI
���D"U8�yr��*'�>�a�Ĉw���q�	^.�y2�M�+pȱ�K��taqC'�y��P!�����ѷ~d2�0�ѭ�y���3#n�+�k�!
6��,���y��]�b"��!H�v�:�I�U��y�	�'l6!*'ID+g�q���x�<�@��TH��+���.�fe�g�|�<Ѡ��2b6�˩w]�Qǃ�w�<q�c��sYz���N�)?�5@�w�<)T��^�
!A��ɩQު�k@�O}�<�L�"5��qB��`�>8���Gz�<��+�"}.P"5��w�rYy@�y�<Y�L�7Mt0� �-#(��Ud{�<!�,���Ě��$��@�C�x�<�霧��x�A�`�u�p'�t�<�4��x�-ac�?A}��k��|�<��FK�`�=HO�8.&x�Qly�<�DJ�% tt�sϷ84�;�#_p�<IT(�+���s����+eX�S#�m�<���p��s���,0l	3���f�<�!"�$F��r��zW��Ce �`�<��׮�؈jQB�8R��k�Z�<A��� �ܔ��#{4�{h�Q�<�ea��J���#�̰2.(��K�<9����T|���L"�0u1��E�<�� -
��T V�BX������I�<A�M�7Z�H ���!k1�I�ॏB�<���	{@�]rW���-��E���x�<9V-�9A�H�e��D�ࠓt��s�<I� �)`1&zۖ(�8c�T�<� ��$(G�����O+>�r@`�"OD$P�'��s�,%����h1��"O�h�5�ޏ7�d x���7I��s�"O����/%V�@�@�7�u��"OX@�!O�*[Qtk��@!�I�"OH�8�$DZm14MW��4p �"O���jA�p���1�擕]��Aҥ*OD)#�@�:i�`�砇5.���'��Y1U 
�7I�-J��:B�l��'Eֽ�7o
$�պ���*�RM��'� 噑R�lM;D�/����'LZ���/��ِ��"�����'��$�C���lB��c���+:��
�'���3�	yn��`����)�'�~�X�J��������9�',,m�&V!uD<Y#t��S$V���'m�H`1-^�; �٣Ё�Q��t��'L�ɓd�ɕ9ppX�
M�
��'����C�&[|d(
6�]�C�����'���8���^����@�QG@�p�'��|��o��=y���$�2I�~-��'��i��-�2����T��]��'b�m9eK�*ex�#�L>�=��'����c�8AJ,�:�D�*=��DQ�'�V��S(�5��� �2���a
�'�lUy��#$�Ҳe���M�	�'�> '&ߣA��H��;Y'4���'q6Q80j\)@fD�hGE'�8�'ݘٸDIV:wWl��D�%Kr�*�'�jP��#H�N��覎�+;�8��'�)�a
��;o��R��W���P�'� K�Ls��a�ѣ xXL:�'è��R	�2g|��va�8��@;�'lZ���d� r�3&4�d
�'�|�p�ڼi�P���-=<L�	�'�v�i��/�D8*����7����''z�)�\�3�V����5(܊�
�'\� ���̞ F�h9AN�8�� �'�� 3�<�j�(P+���'u�U�g�BF,��K��:�'y�|�ÎX�T� *S�D!C����'!`*녞,60��+�V(��'�Pu׉��}�3��O���(�'A��1o�9B)���O�:׶�ʓ����`�ѩ�2�8U���Yl��ȓfrX#�*9��Ɉ�aǑd�>�ȓj�����:!�`��� c��ņ�2H m@2�Ϭ=*ҬA�I��Gra�ȓKo�)A�r��%8�7g����=���D4��# �O�9�� ��T�A��U��L�+�k��	��T�ȓÖ���߶�D+E��qʔI��o�)�S��42_�3��.7L���ȓF�E(@ �e�HiJEA�bv`}�ȓ/*t�p/�� ��L)s=�	��?}&�B �!��P���;k7�	�ȓu�޴U�@�/�,���6In	�ȓxPt�AV�z� ��!@�4l�8���7p�e�'��D˔u#v'�-|��!��I �@B"� ,U�T;q,��\	�ȓF�١u� 8~J�����#�:�ȓ�n�:Rd.Q���
�|L�����D)�����Q�ZJ�C�I?�8�q���(/ �$pA��G�hC�)� �`�V�DT�Zei��K�c�]��"O�Q��8���qf���;�"O�9�d@\�,�������v����$"O����A�b����#��o���"OI��!S<qڗf�%VP�8r"O������F��⒈�>>� I��"OR%ڳk�.H��A�F^e�4��"O
�)��#T���jRF�=�J���"O씺ӈ��b)Z؂`�QOR����"OΤ�dHF�FXj����$aFu""O���tR�]q�1$��$mj^��"OZ�Q�F�=n���	�T����"O�t��[ 9�ֵ�+�i�"O��5cޯ6>��iE�}�h���"O�h��L�d6By)��O�o�	Y�"Oj	����ö��`�� E0\m)"O�lp5�?)�$�k��	@���"Oމ�`n
0+��#�D�s�A "O�	�)�>~���%dQ�.b`H�"O!�J֍i:zi�f��*&�	u"O�����./���Ǟ�~Rq)�"Oʄb`��4\I@�r�h]1j���"Oju	�����F	x�i�.W����"O�]��/��"`���E�V�!R"O��0!��1^]�uqt��D���"O���Ȋ
,�q��J+ax���"O�� ��-wpȒ�F�2V:���"Ox��S�O��j�H�����8c"O�(���	X����޿3u���3"O���H��y��B~r���D"O|5S�a�	Xa86b7�9�"O�e�#2r�H`C�0� �b"O�	b6+ե"$�t�EJ�E6T�"O�)��C%w��U����Z"O�}�"�S?n ����$W콙�"O" �f�(2p�bDS0�DPJ�"OD�0J��H�@8�!ÆiĆ���"O�9��.�
{��;��65��0�"Ola GLCAfd2&��y�P�!�"OtE��MŁ-��	��+w;��qq"O��dς�Oa!;���U9�eQ�"O�A��ɾ:�4��G}%(H�"O8��@��P���*�f�4*��"OHPP��Y%~ޑ���ەe�&�pW"O�e��#a�Hm#n��i��}*"O�|���4��@3ȉ`vx,[S"Ox�D�P�%�����5SR�A�"O���3��� ߲�� @.?Ot��"O�U�0�l08�Ă�k�6xcr"O`l��@R3@I��E�C�A�!"OjDW�ԍl���,z吕B�"Ot�0�/ #z��
��8�"��"O�0A��T l!j�cw�CȊXA�"O�$(�lA<g@�qcB�G<;�B�q"O �z��[�)�B�yB�#�2�r�"O�(���&�:��0E$r�pRU"Or��DeI�X<Kfc��\��U"O���Ǩ��^>�!���U�Q��"O8�"ӎ"}�츖F��8-��	G"O��!Cl�7v@2k5�R�S	�Ř�"OZ��&�Ɍ �
E� #^��&u"OB��eY�K���ە�Ө
œ3"OvT�`@#`�
�taԚ�܁9�"O�{g+��k����`�<��A"O� �]��e��u���`�?l5:�"O���`F
�̅�b@4-&�q��"OjQ�p珈L��181܀;"J�"O��
ģȒh��hANZ�cK�}R&"O�=�%_�5��wm�*��e "O<�ka@��Q�6d�Q�O
_���Cb"Oؠ�K�9t<&a�υy�F�R"O͹uV�d�s��%G�8K"Oh���#��F����� R�B\a�"O9A�#xE��F�V��:�6"O��V�8��tE Iop�D"O�x F��	������AQ�4�T"O<]	�m�E^@�c/P0<� �7"O�E2��H�l�dn�!%��!q"O�<�w/��"�
��K�O��\Q"O�@�T'�}*`-	"m��?�9x�"O����Z�+��$+��~&}�r"O~��C��8� =j#�*QA���"Oά���Aq��䓷�°3OL)p�"O��jqC�="`6��h �*1�y0�"O��Z`O�*X�$�w�!�%+/D���`l׈hf�Ũ�IJ�lM��`&-D���i�^i� �c�.�����)D�p��>pf�)uBӅ�p]H'
'D�t�ohp b��4Il�Ĥ/D��RN�Dpx�'oZ;��s�+D���f�\�V��sKL�"��<�Pb%D��b��@
���D��RDĐ�W"?D�p�ŹlV�	c� ҇MV����J=D�ȣ�lP�`��M�ф!�(B�:D��yv�G�|�$0��E.#��|*��6D��&�LC�`����9�����2D����֩u�9�$H�?����+;D��&��,�nY� ɔ�At���:D�DB�ȧ<� Z䏇8hMH��U�"D�dS�O>�&H#v.��*{jE�Pe<D�$���1$n8:�˓�kL�;A?D�����d��<q���{1&т��?D�|KB�ܡH���22������,s5�C�	�Y���-\�6�!�dO�6�2B�a�pݫgB�4EltJ��@(S�B�	*r�,y�W��7�N���ߊ6�B�	���,;�"ٽ+���I���9x
C䉅n��q[�?` ���*4H C�?H�Y@C�֍n���e�G��C䉔cb����bR4(扁����,A�C䉹n}��hq#�+-ɢ({1�]��rC�ɵ{��`cg���xT���Բ�'@Z8ڂCN�)֨�g���K�'��$C��Ly�us%�f�� �	�'��|��%�18F� DE\�d�i�	�'Ϧ1�� ���-cs�C�_���	�'�6�I#!��4;�@��Q�H��i��'��أB.A8Hf�|��gA�@�@]b�'�`!"��5:v��\��L��'�j�ME����`Իfn\���'˰����0��!`cKڝ^����'
���Cõ��
2��*X�,��'���p�Y����T�ٚ�'x`���3?y����4�)�'�6����ۆ|,�HBF>@��5�
�'tP{�B
02V�y���8�t,�
�'�XlZ���2��$��a5��l��'``�Cgޘ����� )��A��� � (�"?��*q�ɏc�X�C�"OP�E!�. 0�	_��{�"O���HG4;�ؽx��<\N�p��"O�R���	l�dٛs�@?lC����"O"}���˛T���	S��	�ި�v"O�e���V�*\�S�O�w]P��"O�!���W�+1¥���^>3�ȵ!%"Of��g�/ k�� p�;#�ΨIT"O�x*��_�"���d�3{��)t"O�=��f��pg\-�5��49`���"O�x�A�()��g#Y�Ch��'"OB٫��Qj!�Ģ�(g/�r$"O�Y�Pn�N�:m�����$��@�v"Ot���杄z�✢���"��#"ObU���G���ci��h�4��"O@t�tM�km�}{��W�ҭڠ"O�!{ƭ���`X��j٧lg
%�r"O�5y�ˍ:_戕�lA6`. ص"O��� �	�<���KX#~\��j5"OT��B_����"�B��ȸ�"O�b��h�x���c��+y
�P1"O�4����WVt���ǣ~�sr"O�x��n�@d���'h�T\Ca"O�lQ�ʔ�6�1�H�U< p"O��JEd��)�����Ї\G���"OP}���@T������F�* F��r"O��g!��H�4!��؉�h��"O�4�5�I�A�����k��-q�"O �g%א|4h�b	�b�W"OF����l�<ే�0T�6yK�"Oz���� �t�@�F?
7����"O��zD�Xi��x鰏�<-NC"O��a��TWL~Lg�K�TR̺�"OBl�q�H%�L��N���!e"O���lQ�By�� �-��m�F�1U"O
M;�l�KRRܻ�O)p�h���"O�Q+�
#9��Ϋ��L�P"Ol�	C̃;�^]�$���8�� "O(M�NXx;P��)פ}b�[e"O������H	���fgH�W"O�l#N�k�\J2d"CH��R"O��*��#�B�2T��.��}˴"O�M��?PE�� �Xy��+7"OH�J��)$X0�;o�>IftD:t"O0Ռހx7�Ycm,
Z�-��"O�j7L�zv�B�yRHP�"O�T��B8u�ܬ�Ł� r@�!�"Ot��ȕ�;NP*d�Q�'&
�+d"O�YqboD�IgX�9w$� ��v"Oz�x��-y��a��uv��"OVei��Ɗt�����a�X��"O@�pK'E��9u�o�u�G"O6(H$�c�H%��ҷ Ц-��"O�	�I�	:U���7�>�Z5"OX��4%��#����g��Nt��"O�"cǷA��HCGɽn�$��"O����vF��������"O�9Y���+xrihg�:H�@XD"O\�*� P*V��������Q"O~�F�����j�%N�l(���"Op��Q�X�E䈃PDƀK.��"Ot`j�g��q�������b=���"O�)
�j�a  P�1�K.6�yh�"O�h�W.�<��(�ύ��p��"O� ,L�ƯSv޼�ڒn�%{2��A"O"��夕:Wx�;m��mg~��"O$mr`���LtqF��Ie����"O�=;�.K� ��p�G�86GY
t"O<����>C~�	RlB�< |��"O���W�G�2����g�ۭ|�X��"O�0"�NZ(AR�i��[��(��"O�ŲD���dA��	J�D����"O��J�`��n���x��9d
��F"OƩ 4fΫ���*�DX@\ ��@"O"��O��E�v�!���!\:р�"O�g	�)27�ӕ��'���"O0�0v��eC�`�%-�72�"k"O�"$�	cl��TM�?{�[�"OJ8
�n��.���`�̦-����"O�8�S��l��t�U�Q�i�>%[5"OnA7�!=��+7�A/@���ʥ"OH��Kͯr}~H�2�_-j⡐�"O�U�� �2�fUh�	X�QV�p�"Ot4�ŨJ�ن�a�hG�I2�"�"OU:dˠqdx�5p)��1V"O]:�$$Miv��Z@3���"Otă���OWP$+��"5uJı�"O:}jcN
X�A��n�2V$h�P"O�Ez�`�^���M�	yb�찂"O���FhG
RC�l�6kRE`U��"O�}	����l� %j50�-�"O��Q�!7��-H�f^+k���"O25�2E�M�T���+�	)�!򄝿O4�1G��=v�!��&@b�!�$ĝf�n	S/	1b��
aD@<rK!�dI%3;l]�;Ls��{t��! !�D��[�|��h��q<����M��!��:�2Mi6/I4����0r!��;ڠ� g�hN��h�"�+7!�$�,���sL�E�*�k��!�!���z�(����� 8�Uc�.c!�YP�����f� �
��8D!����Jú�4(����]���E?!�D	ȼe0Q� �e���� hM�/>!�*Ċ<xB�N_�Zē�X�"!�d�+ߨ����C�`}���2�!�d�A� �?'O@�����%=�!򤎊���2�G�����ĒX�!��8'M��"�=*�Ru*t�Xq!��}Gx���$�:�4�k_	qa!�$�O�������U\�Mb3�ǨQ�!�֛H��y�1�U�枩Rr#��E!�S\)�$s���1�څ��□3!���!�J��o\��p�lɽ�Py�H	�4���ɖ#�((�5k�-�yB��8�yb��sEf�?�y�n��a|6|�BJT$k�!9�%G�y�f�<���"�l�%9(x����yrF�/�l
G�4z�jtQE��y�˔	zz}0$��]��dq4ȇ��yLI06��,Z��q��k�,�y�g�	0�m�ҍJ�M3n��f�-�yR�]N��,OW3L+�s��Ʌ�y҈I1vdРo�?��x:ҬZ�y�/Ƒ6&�pR�ǍV�(�@�I�:�y�x(Qթ("��3F�K��y�↴��}ٓM9�$��t�*�y2�G*9��ե&��j�.W��y
� ,0���;dt�Q�曼�*�f"OFM��� ����/.�+g"O�lh!��3Z��h�oն�ڽb�"O��ƋJS��� �3~(D��"O A��	%�Ѝ\o�R�"O�h�%mK3b���!�V&l�<�"Oޘ�`ˢ ɂDzAd|f�"O6ًp�߫Y^�����ѓ\J�ˠ"O�9��O\�P�"�D�X'JMd1p�"O� uo�(|ƈ��,�*u׺��"O�ó朌O>X)��
Q�(q�"O^a���;`�1���%~�X9��"O����FRnL4Ka-%(Ѥ�#'"O��a斷 yݢ�Xʹ�"O��
f	%lNR���k�:EB�"O��ք�rE�8��I�V��h��"O����A"
����� �� y��"O ���!�QNEٵ��x�V*0"O�BJ�:*F.����P]eV`�"ORTj0⒴dQX��$%ޯJ~����"O�a�N�+�2A�D��u?�Ă�'�<��%I:'uZ}@�I�0$~ei�'���{��:p\����!z1�=��'�s'��8>h�`KT�{�D!�'��)��H!M �0]�Cf��k
�'`�1��D��@�fHA'ú'@���	�'~���"�B�N(%��C-,3�\��'�� @ �7� ���'+HRD��'�F=�&3K|l���cJ�"E $1�'�y�� ��fP �����!�Ľ�	�'���c���ntz%���Hk
�'�x�`B7�^`�5j��
�']�S$ K:��3'W!,u	�'��|Q��.1{��ps�ǗC�Ƽ8	�'<��4�A�#��Q��:<||+
�'���CB�žW��4�Ql%je�a	�'��A�N�Hh�!��;d�X`k�'�<@�� N�{����&V�U����'� 0XP��G�xp-ǭM��s�'�N��w�Q8J�,�s�gșy� ���'(|�i����BW��S�Aӗj�0(��'eh-�`m�,Ak��x��A;o��|��'p�T��̝�[��!�CkCjl�\��'��)ڦm��D�D0QR�ơl�����'��f'#G���� PS��C�'b�U9R��.0���$�?o��(�'��r�Hևq�`�A��/�k�'����J�źh!��.7�!��'w\uQ`Rc�r g�#�n�!�'�>�#�a�a��(�7�J8��Xz�'��`�D1� �i 䗋TJ�k	�'3p`�.�2N�~	�wm]y3����'�`� ͖�RĀ;0Y�s�$��
�'ւL�P�kcB�)�hݎt6杠�'+TpCE��Ze���/8PƜ��'C���� (�ޱZ�Ɍ�*PpY�''�Mh`&ͅK=��s�(ޕ)�"-!�'���#Q�J��YƬ�$�<�'ܶ\zS���KЬ$��g�6Z���'%�]����|<���@΍�=��'�Za��yz��7��)B�,b�'����Wf$A�q@ʃJ��H��'�����o�3d�M�&�8=��h:�'\\�1���*�� WO�5�<�
��� ��R� 8`���\�M�"O���3�	?d#�Ar�J�j1�9d"O�y�t��	#f�i�)5lIn=cv"Oe+cװn�4�u��Q>z�s�"O�d覯@�*��Ѻ���6s ���"OPE9��ޅb����ф�-p��"O��2#���A��CS "�����"O����'���8��v��~�����"O�@�� �N��b�GLۄ�p�"O�y�g�D�iޖ\�QG�B��X"O�kr��lȜ,�c��`|@�"O:DQ���Ԃ��Z�1��@"Ol�R��D#0���3	e�iz"O�ҍMy���yCGܲd\n 
�"O"�	���]y8@��f�?��$�"O^A)K�<q\���E��V�,�sf"O��VϜ�K��f+����A��"Ot�kC�ļUsĜ�LT�����"O�sI�9�V�AG)G"r`q�e"O4\{R�>N����/(V��˕"O�as���7���A����dT��5"O\=q�
��|��mA$��PA4y"f"O:y��k��/�Ij��
�E>��"O�qb�5!�h8�g6��+�"O�ȳ����+�dE�C�P͈�"O�`�'IĶ?���S� J�P���S"OƜnN5AVT�h��U��pS$-/D�� ����<��C���IG�@#"�!D����oƢ���0�3��uX�>D��cf�|eH���#!o�1�Ο�y�CG�����劖�9~9��# �y��Y73�6D�P���	�,��Ƅ/�y��:t�`�Q�E}��<��m�'�y��W�2�P�C�"@J6UY!�͋�y��Y*q'��Z/M�*����Ȳ�ybnGlS� �'ۦZ�����yR�5������3���L��y����I���6%B(i�E�y@�w��8�sfp�ti�BdC��y��s����p�i@�ѳD��yB.������I	p��xS��>�y"J>x���i�<���1,�y�.��fx�&G�/4ID`	�B��y�# 4T&� ��h��?ȼ(+so�y���;Yv�G�ٚ3{�yRf��y2�K�Y���B��3�����H��y�eH<M���p��תŲq�B��yB��?�R�D��q�j�(Ѧ��y�n�_C�|���=i-� ȵ���y�CM@�6�X��:d�T�AV`�;�yB�� @c��;��A7)j�� f���y��k�x)T卫M��L��M��y�JϫӮu�& �+[����af׋�y���n쐒 5, #!&���y2C_�-�4�#��G+Ev�r��S��y��1Z9&]��7M��	p"��y/ӭi���{7�)�J�� ���y�E��6�K�L��%�r�9QKľ�y�GK~���g#1ڀ�7g��y�B��kj��3,M�E�D���^��yRS�P�F�D!���7'�0�y��ܯO�J�����b���F��yr@D�QXl�ը�|4���Wl���y���Ȕcb
�+I"��g���y
� �)��ڎ&߂�	����Y�}s�"Od�2 ���
���:�kجs�ڙ:e"O��rg���I�da@-L�A(H�'"O��hd�ߛ<�N9p��*/%����"O�����N`�ܚ��V@꼠�"O�`�〭�&B�#���`�a"O\�B�O�_���˵gT uv,��"O��D�ށWƼ`�'�ʩ	ch�H�"O> �OC���Ra��fh��"O@X;�����ܲ�CN�}L��"O(�dAJ��C��\�%G���"O|u��K��O���y���N��ef"O�pI���y1���Cǁ<����"O�eۖֱ��9q@N/H�F���"OP��ccO8�=����:;�<�q�"O�!���6S�-��HQ�]":U�a"OZH��Y�7�И�#'_X� ZD"O�����n*�V旁|T�"O�邴��'4���CМ�À"O��+s�϶|���(�	>Ħ5��"OzE�@�S�,��3�P�+#�P�"O(�r)C�M�شۡ���
��"O|ͺʒ3'rA���J;A���Y�"Oʤ�pm�2J�r� X�Z�^��"O��C3^��qd�f����"O���� Ƥ:z�|�q,^�(�7"OT�2��	-��h[Uk8~#҄	"OR���Eot�q#�J��2"O��w�2/�����'�yΨ��s"O@�旼p�~e�@��' ��"O�4�uf��h{R0����V .��ȓE'h]ڷ�@�c?b4K�	��~���>	d ���ݦV3�m� ,�"Uߘ$�ȓ@r8�A��_ ����̎"s4���~*�Q3���8��1�!��&�Ňȓ1?B`�&e �"�Dl���@"|r����ԉ��d]cx�Ԑ%��]6B�����6F��n�0r��(}K6Ąȓ&�P�!$�S$A!"���@�'��Ą�QzF�6d��� �r����ȓp&tk7��k� �*6�B�ȓY:$�v�T�*�~���[���ȓD�LaS�@V$|5��s�� 3����F��|���K,L���rI�?I�|�ȓll(#a�փ�L����=�le�ȓ�z��c��&�R�a������-��&<(P�2m�}!�Ꮪ"���C���)�,YY&#�<4�D��-w@1�!kZ�����;AVQ��r>&��!�u"N��c�N�aZxD���� k`�K?.8(��2�����,��A�%ǎ�N3�}�d�ŵx����Lx��2�	/[�hK��ܭcU�ȓc ������-Q6F�#1�آ9i�x�ȓ/J�	S��ɂT������!A��ч�|���k��¤J�9vm�����ȓGu�
L�A�L�:Rȕc�f}��f�:��"L*kcX6�]r�܄ȓL��T9qGC	��
l�/c�^фȓ~@+�hLm<��u.������ȓy�4Йj�#��E��kE�#SVd��S@P�0S�ߪC�0-��
J��i�ȓq���17���sҘ�`ƆG�V�<ч�>��٪�	�y��(�J��I��S�? �<�����Fu[aQ=HAr��@"O����^.y.��En�A(� W"O������!� 51LY�H�Ac�"OF!�RCJ�\x)�FKP�
4�HA"Onux��2Lg~A����f�E�U"OiX�T:h�ֈ"�I���A"O�$Z��U�Y���a#�۳,yJ���"O�y;o��e�b9*Qp�ʜx�"O4��G��f�l�X>}S)��yR�WOWx�8BAZ�]�HY�"AF)�yr	�=s>�ЬǮM2T��
��y��
>!$8C�a?�<�bM@��y�eí&_�m3��2=p�A3�׋�yBC�g�Jhz`�
8`��ɖ)�yR�US���z6,�8M����و�y2�^.zc$}P�BSc体��y�Njr<����0��@fF�y�g˾f�n�Ae\�/qՂ��y�È(���Ն4p��a4��'�yB"�7^\�p3�ۜ �|)��FI��y�&�
^��	k���Ķٱ6�W�y"�I4�`}�!!->�4a���+�y����>.�X����&}+a��K��y����*\K'�S�b��L��P�y�аjx��7f=W�L�)�i���y��C�����P�S�	ԉ�.�y�m�54g���`UT���s�iP��yk[�b1������O|�,��hQ��y��Y�}Ȏ����6�L���>�y2�Ț ��Uˏ�-c�<BQ�Ö�y��_3��P�E�	�5r� b����y���5+S�H��I�,�&ٳRC���yB��9_F �W'��q^dR��1�y�(]��i�/P�u�p����yb�ȇn����t�����ܠ�y2�9k�����p�(���U��y�0!.@"�Bџb躍�	�'���jc�/s�m��&$@��	�'`�A;a��><&�����'�	�'��qH$�K6
�Jp�H��^�&��'T ��0o���b�ڦeō@�n��'��5`Db�?/��[.�)*^�IC�'�;GF�Q���rU��$�Q(�'���T�1P�c�����=i
�'=ր`�p-��Qԋ��p9�	�'���R�
Qd��T���(���'m691��WJ,8���{�@�	�'�@y���8j�+�O�������'�)Y� ;�'ԟ�F�k�'�
�#F��e���@0z���'�ɉ�kM9,��iw,ЂB� � �'w"�X����&�:)K ��'ŌM*� �y�$Pb�	ͧ
�="�'�$�u�m�*ܐ��656���'�.$ ��ґ
~�%�à���'���	�hĈ�3	[�6I;�'����D�~�,�&@ǀN b�	�'�t�$aͺu>v��&K�#B�V�;	�'*��J��)���Iŝ�T�I��'�
��!�^���&��{�n��'�<-��%BI)XuvG�#H��S�'Tl!d�ȓ`���C�*��H��'��]Sf��|��aipq�B䉱~����KF�s�N$�a�̪5��B�)� ���m�/pe�Rt!�9'P�!�""O���Ug\�e�0
���Q,�;�"O� ��d(�2%�b/_�8�z!�@"O����fϾ��K|\07"Ob��0���^e4�z'gO�Rl�"O:���$.?�q�P(\$�+�"O:8�UJU$?t8Q(��I]�.1:"Oni¤�J�F��*ׂ[����:g"O��a�L3zg�19� E= ��%��"O�i�����;��4�΀!""OZ�Q��f@j����@~�t�'"O�k�$�0o�6��f�f��]��"O�Ys7̖�sC�����Ps"O&�
@V�<Ԩ��!#S�}�\�(d"O�xB�j@�r�>]�bR����$"O~p)��ʜnɊ�u!��\���"O���D�x�Q�t��=�ڍ��"O��cZg��1�:V�~=;P"O����ǰ�m�t��C�x
�"O<@x�f�=	�E�C��>Ҏ]��"O�0)��֖)1�Đ���l����"OR��(�l����7~|�ei""OR<IC�F]��"Ю!N�l��"O��kϛ�WK�~ܘ�s/ˑ�yR���m���7醕z��SFǡ�y���rQR0�,lTN [��Y*�y_#"t���p/�e<q��g���y��tN���F���� 1u�K��y�e�� {!J��@	Hr�Uk��y�P�x�z �P���,5 =�o���y"�C�YQ��7$X�!�N���>�yңoaUgU�F�
%%z��{�'�~8� ��*}��R�Í0p�ލB�'��Z� �4����c�����'x@T!���; Y�i���C�c3L���'�4T� -ڈj<���f�ʈZRnl��'t�="�3�i��
|�yq�'N��I��9��83����yH�'Y�[$��8Z�0UH]�(5 Q�'�"I��A��{���AgT�PT���'\p��e�A���Fe�0���'˜e)R�΍lR���� *��
�'��Q�� �^�aM��K�z���'��X��⛺\����O��Fg��
�'/:RMw�ji�f�Ҍ75���	�'���*abk��F�1:�nx	�'��Pk"eZ�r�S1B�[r��'v̠J�b��4���U�d��'��0U(0>���YҫPK����'���0��ZAǖ!rDHQ/X�@(K�'&x��u&
i�����(��HfI��'^V�abo�!i�R|��&S2v�+�'��܁V�>F��:���>0xqC
�'�-��,D�j�2�F��3�xHB�'F�%kw�M:,������[+<�R�P�'���P�J߃Ɏ%��5o,�

�'�ܹa�i͟8�Y�G�WA/�YA�'����VB��5�V-�͗3gx�r�'Ѿ�0��ŃS�����/��H�K�'ʲ`rA�!n��#�G��q�py*�'���ȵ��J"��x�cX�dBP��'�0a�Q���;촥���]8����'�(�ӡhԫ w(�������|��'M��5F*J�b��~�8����� ��:�D�9rȜ��cM5B��{�"O�( ��˾o0���آ9���1�"O��7&��G $��d"��[#�bV"OJP�	�f����@��kB��"O ���I����#��"O6 ��@l2�`��]r�DaB"On��a�6Z��y(����^�"q;"O,T�G%��+�����K�3��	�"Op���c�g>�CgX�r,��f"O��ש�!lz�D�S�>�"Q�"O�Py�K��{�.�WeӡZ��ȹ�"O�]q�N�O����P�[�H)[�"OV<[u���f����Pj.@�8�p�"O�A�B%�ؘw�j����"O<�ꕬ:h�� �]�2�#"O>X�0PtsV B��ʒ"Or����4�8�9go��kŮ�04"O��x�P#]��cH_
&[�ݘb"OH<��EK�`VrQ��%�+SO��9�"O��b@�*D�i'�y>j��q"O>-Hd@��-p� r��
sǬ��1"Op�C��!�iX��N�u�J5�w"O�q���k�L91����X�YU"O���(�##������h�B$"&"O�BQ�>g
�����W�`��w"O���+י:����ŗS��s�"OR��`�4����A�ƥ-��e�%"O���f�T>�a�NW%4��p��"O�E!Ӆ>߰��X�l���� "Oj�`�鏻�4+��҄�i	�"O�(��1}N*`Z��� "����"O(��F	
:'x�j�N�m��"OX��/۾=�B+LC�5V�a0"O��#LpA��HS�J�!�Lu��"O"pA���.J�B}�CNKX@Hbf"OX[�5e�8!�cZL<,��"O:�O[�p����[?E2�%�G"O�g�$���#`5*lҨ+D�lc2m�&�f���ŀzxd�z�/(D��ZՂA6mT��Su�<ZBMK�1D�L�S�]�>\�l�NP���.D�4��.�>�r���� S���ch,D� x�-��]z��FWb@ �)D����
�~��AJ�'߿Xw�-1U�%D�4�ďT)�j�aQ�GZ��I:�m&D�г�ֶY.8���#� �����C*D�@{A����
�`�?���q�%D��Cpa�BlvЄI�H���,$D���ϴR�
-���'l���Bl!D�d��͐|�ę��,'|�5��D>D���ťQ&qt]��n]�M�y�Q:D����G�7r>C��:��Q��=D���seO�Jܕa���]t�5�cN)D�4j�A��g$p�-M�,�T�j2J-D��G�S2A~k�mˡ,C�
�)D�X�gAF^����1~3.�G�)D���'����*eg8��L)D�T�fϋt���b鈤\>���Q�*D��z���B�b�G8)-\ݩ�(D�@�@�. ��@b!��*u�b��f�;D�8X� 4�JLSf��,>�遈6D��C5��e��^�B$�2'�.D��B�W2�Q&-q>�9�Qa9D� ���;R�h����Z�f��Y�c5D�� ��`/�nT�2�,�w�,�"O���&@� ���Sۣ7ZY�P"O`$��N :������Y�b�� "O����b�@pק�� ���r�"O C�܆o^$	�l�k�B���"O�z��ۻbO�2�*F%)�:�`"Ox܊�E;r@���kJ 4r ݁"O �+ck�o��5��	ߴsZ`�c"O�QG,�&�je�R�a;�"O��� �.k�^�J�+X7��A6"O p0鑋a�H��E�!,'�0��"O�4���66���k�̣a	΀��"O p��E���Ma���=��0�P"O�E�b�IP6�8�m�,�d-�"OA�$%�<�� ��ʀ*O�M�@"O���r	�K|(9fF΢m�b��w"O�`��r�P��4����"O�H��J�=@^:�	U`M_wX�h"O�	U�ީ[0~Yj���(b�uX"OV K�	���*�IQ�J+EHJm��"O�IC�"
79�\u�oˣ�Re�"O �2��<$�k�k_9/,qSC"O��a�� Xc֐z�jͶT{&�*�"O|�Z$���`4��R#\oU�"O�8� ��Qd�cB�A�N@|�"O��RǑ
-i~H�&c�m8֙ V"O�Yp�Ֆb��rԀ�5_.��q�"O�e��?r�f��G/��_�N�&"O�kAjۥ����Y--�~���"OV�[!�|h�Xv��0���� "O�w��)xD\}:�l��U��y)u"O����R��H�� � (����"O6��ɋ�"H����O9�ݚw"Op�KT�R$5�BPT��I8��%"O���֚#��'˭F���F"O4@���Q������`��T�"Od��q���"U:E�����B�"O��r�\i- oU�-(6��"O�ݛ��<̬4������D��!"Ox�+�d�5\|D⊊ajT���"O�`@4��4jI�9"`+��^&���"Ofhs��@�D�jIS�IYKV40�"Oz`BR����Xt"h9�P;"Ob�
��F�~Z�M��Ց63��8�"OМ���U9��,�*}n�J"O<i+U�S�u"ia��R�fz�I�"O�XI2�6l�Z���/>�r`"Ot��G�R�]E��F�R"/�����"Ol"���:d~�s�,g���ل"O0�[ �/]��Z�aٯzE�H0"O�bU�R>t`0<�!®M����"O1q1c��t��P�a/L�:�,��"O"���"L�8��=� ��?F�$"Oz��1nW�H��&l@�=�g"O�r�CL N�l=.)w�iE��y���jɡ���Rͪ4J*X��yr��2}� vi�4��5BMB4�y"����uR�U�24��UF@��yB ��)���Y�L۹<�j�1eD���yb� i<�4���I<6^����y���1�������~(�M�4��yR#$͢=Ӥ�݉|�p���yb�P���D`QK�E�z(�#�� �yr�Q�S�,�ŕeeDI�R,U��y
� �Q*�(]�)luY6��,g�a"OZ��iUV�>D�f�5w�Ei�"Om�%喺@���P�۔1a,�j�"O����c��;�ʴ�2��2E})5"O���m��9�JpR�N9GD�ģW"OL�� L�+l� �Sb�$4&rlJE"O���&����ڃ!��H#��9�"O\�3C���6�q�JO�}�� ��D �S�:M�DmP�D�)3Zz���.R�?Q,B�I-[ p�cLI�|Z��3�ܤ����ߴ�hO�I*5$X�`m��G�MU��~���D
2fF�=�ǧ�@3|#O@�P���je
O��J�)2�h�8e( 8�����'P�Of��-U���LJ ͇H�
0��"O�u��$��"��٫Il�X�"O0�("f�r�J��B���0u�0"O�d�GӢV�Q�2'^�G���H�"O,�G&,���l�H.5(E"OP�K���^�80J�Mb����"O�1����q���b��+[wbx@"O��y�V���r.A	E]p�"O�Q�2%D�K�\)3��F fhX�r�"O��������5jAȻ*5#�"Oj�C$4p���.sF(�q"Oұ�BE�#J�61��ɇ�<�D���' �'�r(�����&������a�RM��'�ܴ���E�p,Pb�" L�Ѕȓ�\-�@V� S@�����z�bY�ȓ:���	���0�$��e�T���x~rBN������hF�{8pDO��y�^x̨VN�?y��57 ��?����,�¹����/=_D�+6�3e�4��ȓR��9`O�Zj�3�˘�	>6%�ȓq#�ukƠ0b��ٺ%+ǇuWp�ȓJ�,� ΋�Z����՝�~���_ҽ��I. k�c��R0��V=ْ��Kb�I�G��|�H���t�H��Da1\�aĹF4v|�'#ў�|�L�E�(i;p�կѶ�dlJ�<iF+��U��,�E��qZ#�o�<��IV�։8P*�=^p8RW'a�<���3���2��9�����)�^�<9R�]aP�cc/��svЩ��d�<QD͛kb�3p*J��I�/�b�<!�(@�&{j%k�@0t������s�<���Q�d��@�g��r�m�<�@�Sj����^((h�!Q�f�<q&�K�H�D!n�x@CQʀe�<1��� Q2Q#�g�
���_�<���N�'Lx h���\ú�6h^��������4
= �T%���Z��8�� ����)�i�(邷͋����ȓI_���L'>���D�:_(��ȓa�^���A.,�`��CΓQ��!��2@�vъ�X�����%oSR��ȓ-ɂԂ�LӍ3/Ƹ�&/ĝ0�م�.�J�OЀQ��q�a+�m86���Wg�|��eʯ3��< ��<4�t��ȓWJ��w�D�D���#�[IXQ��"��A$Ɉ�e� 8�ƞi��`��r�#&X$��|�2��"��GxB�)b&g��P�U'ȴ!���w�~�<���5:�����#��8���x�<��K]�B, ��i"�@�Ms�<� X���ɒ����#2A�:=sP<�"O���?i��	��2r�i!w"O.��w��l�^�0���ch=8�"O��������t�Ȃ�=g��j0"Oj���5&Hr5HF&C=7Q�Ժ�"O<��q��2��b6�2dޤt�6"O��r�",8�$E����b"O8�s��.?XT��G7Zz��6"O�� ��J�QZ��
�oK��y҄R�e�u`�.� U��9�+���yb�S7�f\��D
�ʵ̋��ya@����KIΪ*��T�����y=�}n�O�n����Q�y2��<.U0EOD"`~Ji�q.L�y2	�}N�4	�%ǃQ��M��,�y���H���:���^$-`�-�6�ў"~ΓZ-v�9n�G2�}�G��	�| �ȓ �ڬJ֋�K�x�	u�J�K����w?�F����ǋ�*��!K�	p�=���<���O\��Q,C"(ؤ�SE̖�e�I��6O���$;f̸E��'���h�쐀Y�Ov�j�O�pHסr����#�uвP
�'�����锹4���Q���\� t	
�'(�]� k:(���ٷ'�P@8!B	�'I���v�/u`��7(Y#M��l�	�'Ѻ�*F'
�@��M�Z,�l�'f�x�AN�j�̐sw#�� ��'Ӑ%�B���6�7��z����'�ў"~�c 
"N����b
A5T�3�Āph<��H��/�ʄ;�N�&>�hhpFi��0<)����7��%)�˟lv�K�'�!�d�)�$E@F�F�8BҁQ�	�&�Py���w���f�6Ly|���G�y�"��A��Y���G�˄σ+�M;���s��ܩV���^X��A�[B�v"O�0�`�}r.� F/�4�"��"O�E��G�"$}\��Ɍ'�p�iv�'��	S�إ���P(/�`p񅕪4	,C䉤3@����R5=~���%ȇ�?�C䉄c��캱�/�|��@�l�����.�	�8�Pd��ꃫx�'J�X��B��y�.��r&x:�� ��#E�B�ɗ^�(����4Ph��B_g�����>�+ƐN^�ѳ�@�XV�{��Ο|��I@�5�R�0W���f+5/zɄ�vJ�R���at��ѳ y	�8�	\���'1����ċ�@bPzR,�&]�h��	p�'��+�AY 5J�K C�h���$5<O��x�[�,I�M�D���T�'�Q�X;S!�l5R�2��h�^IqVE�kh<a�^.HE��V�V�l�RaHj��í]���?�2`�2
l��R���m;��p�j4D�x��O�#b5+���u@��A?���<��� &D�D�d�7,��A���v�<�5��<Y�(H�".+:tx(��B5��x2N��l�Q%K!I���U�p=Y�}R
�N��D��ϩ=)��{b�^*�y2�C�>�i��bս>��"+���y��f\J� pb�ꅲ2	V/�y��#`j�]��O3G���v���y��H8w�$��ٚΪh�����y���yS�Rg��4U��ru���yK�`�Pӫڨ�z��G��y�)@*rѢ�P�핥+3Bqb���y
� �Յ1��h� o�A� "O���R̎L�����M����Zf"O~�rD�U#a= {��5q��Lӱ"O��K�[�\=v�"��`�8b�"O�ᇅN�R@��W��~���k"OB� �V�h>��{d�����-
�"O����
��\	�f�R:{���#"O�;Eᙊ;�l�3)����=�S"O�!�`Ru#���s�'���(#"OvpQ�HG	Rь �oEka,\`�"O��� ��vv���(��G�H�!"O*y����v��g��2D\�a�"O������F�H��^�T̀��s"O>E
���j��Y��k�
� �9�"O�q	ĩ�H	R8@��U�|Kw"O,���Ғ=F�C�C�4N���"O6�H���(8�bX)R�E�W:z��6"O��@�`3Y����śB�Hd2�"OФ�(�`�����8��у""O�IK�i�I����D�J�8 a"Of�Ѓa�W�Є⍰�-c"OJI *�/(�6�rQ��A�xE�"O2��Cc�"R�ÒL̜Ai�"Ox�A�'�;�mڃM�O��Bp"O���)!��1R�,�5��h�	�'T\@jQ	��x,�yp�̯[KP�i�'$*��6d;`d�؈�	��Ot�ɸ
�'В,ʔK�����D�81J���B��\Q�#úEQ���d�ؤAF󄉞.�Z�(��_n�6F��:�!�d�	0j�R6aP�-��Ô�!򄋺^����N
"��%�����!򤖳��q��,A/�E)E[��!�d� �� j�Dgnr�%#��!򄘿\��ĸ��J�]\���8�!��	�B�"ªųPC��r��e�!�$!-ʆ�C�OL�~�vcbQV!�$X�;�6���.V�x>�����*}T!�d�;��XP�!�,X4@y�n�,Uz!�dŏT�1#j� &�X���`�!��_�l��v$Y�x��h��t�!��<��VJ�lP`�e۲gd!�d[[p���*q*(�+`�F�N�!�O�o�pӠ��Q�����4/��C�I/}�Լ��Α�L
�#���3PB�	�e"��(m�2aoR�F��C�	�*��H�*��9o>̀���T6@C�	
:����L����
��p�5f4D�@*�FV�~�1���z��>D��p�JڨF8`8�Ǝ6��Lp��3D�\�DNޘC^p���ŲCBNak0D����%��~AY!�!)�>�S��0D�p�E�I���1���M��=�f�*D��kC��/&Ċ��2I�1�eA�g+D�L9�#/Y?BC$�])uH��"�)D�t;$�K>$m@<k ����&"D�W͜�g%���bв}Z�yZ�k#D�H����3�v�	�D.rŪ �:D��Ӄ)ܟH~���B�M�H�ۡ)"D�B%��!^^�	���b�U
�%#D�`��߷YԶ�0��?+�=��4D�A����2D��фM2�[�/2D��Ps.ʥ!�2I��˘(TNMpCb1D�0�-�p�(�2�е�r��0-D�$#CJqT��HFB��wA0��r�1D�� @��� ��KV����#A�f��p"O� ��=���@7��8+_�[�"OJ���E�X�d� R@V�$q"O��s�TKD��x��ڲ`����"OT�ӡ�	]ʂ�"B&� ?��̻&"O�I�

 T��8��DX"O�)h��Ѭ ��EY4I�+p�H�10"Of�Q�D�r�sr R��r�'3�T���
�Xv��[|��� ��3�:��ad�^��D5L�5i�ߤK�R���Β���@8�I�$i��4�P�r\��K6���b)#D������+�|��ȓ0 b�)E{�z�� �5t����I0�XL�kW,Dsǎ���ȟ�e2(�&6���҉��+q�0ra�5D��Ck��Y`��¡�Gx�d�hи����%M0)��C�g�7S��g�'�0�'��sT�{B���*�2M��ܢ��λm�qY�ٽk����֠H��Y+�
L����_�o�|�g�(��! w���mgPD;Qǆ�(OnT9�gP���x��DhlDd��U��Ƒ36�W(��a��$�B�	�rP��3�!�-�"a��@M����-X��{4����8U��L���	'��ﮥ���.5$���G��A���B"O�Yt<��y
"�̶yA���1�A���#�%%o�P���	����O�؈7�@&y��U�@��J ���p>� ɀ������ѯN�Hp�U?���"��x
���t�ˇ�L�1�#_]����/ԘV�<d1��N5?Q|�Hw�1ʓuC�Ѷ��P�&PYrG�:Zh�p'���?QBv&ō~�B��g�Zd��/D���G"�J�\@�s�p�����L~'8�ԮĖ8��h���]S܀�'��p�ϿqK��P�� q[���7�V�<D�Om?���ԯI0e�o�1����]Lm�W���W�,�)�?��"*3�I',��R#Q5U�L���r����d�(�e��%O&�͈��V�6X�@�g�Ac���"�n�v!3�eK��M#rl��`�VL��X.ed�h��y�͡\�&�cE�.o�k7E�"�hO�pC#��
�JmyD+��D��i)ǈ
77�t}�&G�Y܈�T�0��y
�"iz��@�	N��ӡ/[Qx��kt+��,h>);�֚���X��|��Ҳf��`�r��pK�"�܅+��<��V����h�m��E����.;]U�m��i��LЎ�`�l�-��xBŅ���9����4m��z`.˨MYF�@�i��[T]�IN� ꦬ�4%E��%�ŠU4l��2Ў
+�y�剉��Y�敯4d��"G����?�%I	P&T���O�<*��౦���~q�#�´J��T��Ȉj�}ʧ�V<[<h�T7:&����f'��D83:h@�w �UЉ(�E�(eџ��a�>h9�BA�S�:��t.��v(b4S�@J�}���C4�0�T9_�e �x����A��3�P�ቧ6��%kኘ�)A�y�"BTeP�c6�QVi�	JN�91	�&z�H�j��g���������t��
�H]�= �`�%*,s0B[9�L)��'f�)q���!�ҙ	3��9}$��s�f^� �F)�`J\4����Y?vi��$�	�މ	s,�y/���wH={ՎR-`��Z���r �8S��uB!;Ul�  ,<�����3�I���?B��"���O�u�O�?�&�[�]�%'&��D)��5�}��O�Y9WCƘ����@8Peh�В�	�X8#r�K��Z��բ�nY��@b�ڐ5`��7+�)�|�-u��I���=@��EN�a�����)=O��q���E�Z}@���dq�5�c������Ѩc��3�gO�?�H��@�(��jVL���I���G�ĩ%,}���<)4(9��_�D�����zV��_�Z�b�M������j�? 6��H�q�Ψq)�.o���� � [�T�B�+M� ��Պ�jj�U[��W:$�(U%�H��zٻ!($���u�U>��4т/P��"D2���0O�LM��O(��3Q��Dv�1�4*��:�� �rϑ<�<x�OT�KE+]%|���� �Lz�����'����X�Ku���0��8S�Q
A=n�ҥX��/�ʴ
��&7�v��18���"��kX����)F�)-��P�Ň2Y ��ch/��ņ1^�ۓ�N�+�|��"�2QF@Pc偹>����I��� A�"S�G�����3':���-Ν�C�h�`BG��MR	��?��L�F�A�!{
���E�&܁��H׺ ��>Q)�8����\�+u��À�>�ĭ�6O2(ҡ�X�gf�i�7�]�3�"�oO�b�mHf؄y��S(M+f��8��ƙai�U�Ǳih
�Q���<A׫���P�1��W5̦\quos8��R�GX�]�v�%>
����pb[�w%j�D����A8"픊?���;�B�F�f<��,��MK���5p�T">AB���U�(�*V�	�F��賎�hy��ح'�IZ����l�Ԫ���2IЦ+���P�	�n�ԙ��:g�����4����LZ�t�K�'��p�����c���s��_N1�,�uF�Q���"P��@�E��T��ܺ+��{J4d�a޵�a�V�mb�$ pÆ�q�6\�f�8�O�Kac�l�? j��3.�:Й㷢_�D�a�ʇ�;�\雓!\�y&�A)�@ؤE�f�ңNT<=Υ��4)���t��ȴ�Ȥ�B� ��6��5p�.5����$A��F4�V�9!̙B!	H�~`��N	�<�6�S����M����ǡW)f㊼�3L�;?��8{~�>���;B��Tn�
	�ȻV�⟰�/ѐJ�xp�0@>n����GQ�D�%鄎�6�����#u��sL�|��d���G�4Ac���X�<�O�"G���q��t�a�rf����
dm�-"��
͑7+c�)��o#D����b.w�E��[�t$�a�tmsc,�"q�:I�a�Jx�X��H�BO@h��eL�\�3aR1;� {ceK
_�X�e����:)����20Y�X� �MY�$K��3��$A.^�i��D$c8��W�kJ4�=�@	Q�R}Jy��E�B��% [�
�� ��SM��W��t��HN�|"��D�vx��� G[�� ����{�U�$̦\����L�O,e�Α�L��\��-O�O��=�Dn�$|�i���%[�� �T���H�(�aQO�J�J��c��V�j����<D�hۗ`[��X�CbJ�*�R�
���{����l�;7/���«Ũaz� �35���]f�`��Nü��y������ڌ�p��GkM��Ȼ��<k�Ę`'�E=r#`��Z��0Q�ϝ�w�P�+B�$����a����µ �o��w(
\zQ��D�5�$�*��X�p�N��oE����X�f�]-"=S��W](�`���
2f&�1���y��!$$%Ad��U�Y�U��Q�ΣE~QJ�'��]���/\�a���W��e)�'�z����1���( o�#V�8�f��,�&L
s�K��"%���M��d�?,�r��cb�$,`� �"OD�aJ�:P�p���+�.X��VME+�&�K�+���``�h�J�"Q
s>���M�)H���=���فd�>53��,?�upB�'On�U"O/A-pi�lM�3�Ԉ@�V:&�ΓW�ܸsh���mYՃ®B*~Y��-(��}(edßjv ����rG�$D~���"�@�S���c������P�2|�Ueݲ^��pC�]K�����&XR�1�u��630�ͅH��E+T�a���B��V?	��˓P���#֋;Y�"`:��Ҩ{�F]9�L�?g��U�B�s� ��`kN�0�cɁ/wH�qh�u%pB�/=�bT��4_� ��@F&>��3xy�]˕
		m� ��-9�hX�/�2����	 �yw'��M,H����?(�h���J���x�闹{��Y*Td2s]6�b�-Q�+�f�ۇ��&BD>{GER�R�5т��9{��I$dSp�V?: ��/S/¬D�C�D�G.���	it�(W�ěX�hX�(�k�F��F@�b�~���']��&��h&m�7lO�u��!YPJD�p̘9cb�5����\13��5/
Vh�ꂂ�d��%{�� _���]9A�DA�E����2L�,K,NC��#dr �3�^�PD�#_w\!�gA�`��q��ߩ7]�a'��`u�#I~z�eq�i	���<(�وb�ޑ7`=�W+D�8�%�	/���0���3�~&��BeŗWJle�����>�nM���@)-_B\A��F�Smn�K5 Y�2δ��E�JV���	�1kne!AMR�R����Pc|���^,G�0��a��i�F֜)��9�2$�L؞��AU�crp��.X�+'d��A�9�I����x#l��-��!�Skُp�$uyQ0�L�	υ&dt�a��Ճ,��8�ì�F�!�DS�|H�}2pŎ*&�~areřn�:��W��X�K��"^D��f�S9}Jq��d��w�JX:7�] }X쨄j�T�f���'�>����j��:��G�L�4��M��8�>Y�6-.Dabx���	l�:�ÌE�'���PeY1T�0HR�dT�D��Pr��1Q%��.&��i�B��+���ɗ���X���Sq,��jYN��q~�����L���kO.
M\5���Ћ��8�=q%(��]}��b��Ztle0rJ�%T�Z�'�T��uC�}TF`�w�� ;������򌙢`NW����b��XbN9I@L�/�H	�ꊢ\"4�E&R�O`F�ɧ0W<���oM�R�3� 4vvB䉲��h�vB�x�̰.K!J�0s��Kl-R=��-͈v��I2��2�Q��R�+ɭ/� ��I�7Yn�+�L&\Oqr�������Q�,"�6�����%bf� % &n��!�%+|�P��I*X�j��ԉ;�~]��ۭD�pc�,�6�Q)X'�48�� W,�0�%eR�I��-v����M�\� ɩ߲
r!������6�:��}��ҏM:��k�h����5-�$� ����eN�1������>or(eB �:D���#�2�l��Nʀ;����ƈ�.�MS���nt�U! gܾ]��g�'��ܲըF�Jp�%��Y��U�B`l]�6��3�`}��Y 	����	X�jeV2z������� �x�0�^�RJ�"=AP�rC�a���R 1��!��ȥ)I�A� ˌJ��"g"O���a�dY!Dw�;g�'������J�B�O?u(���%N�x�K�9@�XL���P�<�ǘ
/!d1!w�ƞt��H��Q�<� ʽ#T�=B�����8v�18w"ORU�w��.��05��$Lj�I��"O�$��n�����lv�| �"O�ђ��	JF��s�L��"O�|[��+O �(��
��,O,0Z�"O�3�!ĳ2�d��N�&	*V��4"O(����,��@��I9>�Ԃ�"O�<Qw��%�Y�s��J����"O�q�R��4@��IpPN !���I�"Ori�w�+�}0�-�7)��iHr"O�]xԤ/1��xz�R:Uzܚ0"OH���)�Jf�E&	X]��G"O��hp-� '=�=k&�NB��	�"O�D��`���y�E*D�/���8T"Or�� �P�j�ه'H:u�h"O\�i"�	`;08�ƀ�],��&"O|�H ����X�rƄTr0�1"O�h�PǊ�8Aw�Be�iy�"O|�t��&�����;��'"O�(Ѣ␣zK^�qV��3r%��"O0m[��%(�\;���"��"OҨK����N�	��
Y"�h�U"O����ꊐV�6p��H�/!�=Xt"O��aA腞��Y8��U*$ܹ�"O�yI�d	)p�pQ����ā�&"O����^Q���i2&��=�s"O1��c i�(�
�U�NQL�c"O��0��Y�4]*o�JkƌjB"O����"J!f���"��}J,Ay#"O��Qn��4���ju@�2`4��"O��
�=I���!� ,I8�S@"OrX9"�ƜXb��`0o4-/6a�A"O���b�=a�Y�"Oh|�P܋Q����,��lX-�@"O�St���NrB݃*�:c�����"O�QSW�;
��lhj�l���K�"O�LzD�_�x-i�zO�P7"OAc�fÆh;x}��ٔo��Ts�"O����d?'MJZ��N����PQ"ONA�g�<'�na���	=�ލh�"O�	T�:O�0F��zG�M�"O���%��vf�yH���r8^ � "O ��F~+D�s7�@�|�rܲF"O�0a�������<4d@5��"O"�H-G�?@��%ũ=�4X(�"O�1!�� M�ZE�@�r��9q�"O�d��h�}�\h�#�^��Rv"O~�a�	�	4咡���!w�К�"O:�����8w�$��F

^,*�"OXp�r�� q"œe����r�"O�٣�������J�-�d��w"O�}3%jԛe��a�N�/a�S�"OZe�%d݈��%�7nǯ?���U"O�y9�ESn\�����k��X�Q"O�` qgӤ&xxP��,"�H�� "OZ�G�T��	vfаYX T�"OL=�'J���Qg�u_� �g"O��$�8DR�J���5UF��"O�x m=���)g��7�6i�"O:���≛�^�2ǡW��vջ2"O��S�,�<2���+vϟ !�|QqC"OX9�4.X6B؜AԎz},2��UL�<	V��5I.��9*����aH*D�Ȋ���\�Nm����u�P�y�+D�� V|�s��[xb!�v�k�H��"Od�
�	&P0 8��=kk�p�"O�\Q$G���n��Bc��(2"OTq� ɍ�fɴ��u��'^,��"O>���M�>y���4F�|J`"OД0�$Y:
�1����U0~�a4"O��c�ܼ(' �ʵ&̋`%py	r"O����-+v%�0��t�v*�"O�@(/�|lR�w����A"O��9p�[9S��;�&J$J�B,��"O:4(��Y0���%��Ǫ���"O�(��/����t��
Y.0"0�'�
�҃�ֿ7{�4��'B�6)�(8ӄ�>}��9k�G�#:| ���F��"Pơ��i���@�Z�lK��B�X(�0�Rv�\=�����Y��?F���s�� 	>D��+����a���kkh �Џ�|՜|��������F���d��M	'�ȟ��h#��u�� 4�"D(#�/D�` �,�2�z� ˊ�M�.�9ġȇϺ=9χ�����4@��g�'��mB4A[<L�,�R2*��h�	�dy(����F#j�]���߷/qD!���(Y0���'I��Y�b��<^�|r$F�=4Dj*	 �]�ݐ�(O��$�58?1@�
ۨ+�};��P��l�)��*3��/M8}cc�O�<�1��p�d��5�à��pB�R1�8�,ǫ_^ 8�� �!�<��q�0����WA�51�"i%Z�9hLau�*D��(�+ߕ%w`�I�L_�(D$Y4φ7��Ei�� ��9�p��B�r�S�96��*C�+�����0�B�#�O�lx�+����@���+Vh)�3_6?�l�BH���T�Ȳ�װ;t�u�S�'|�)��DܠyԾ)�'�B3P]+��Dմq{��q�#٤���
;^I3��O���@�p�jh$/�����S�'�ӗV�& �Ǝ~Vm�%/Ȼ^p�8u	Ò5f��80�ԥ[����������0���+�4<�c���<��7"O>@����i�>���%8��q	�Y�L)��k���x��
����	�\��OB�{į¾3ChY��ߺ�E� �'(���Ꭹu��1�˞lYt6�\+Zg�zU�ܘ$I`�{Q��6Fơ��4^�.��d��|-�Q�ᆈ�Ԙ'����,	�Qj�Ny)<����O0y*��2BkÃ~�D���'�`��ע*y�}u�ɝeţ^����w	�&RS���AP�S?+�'ΠD��&�^�\L%	�1v�9r�'iT]��U�%w.ѠBǰX���'�PT#E�0u� !B��
��:H�� ڧq�-�]�&� d��#$�L:7�M�(���#�1t'�� ���'u��(�2�ȑ?�HKwZ5�PG)�+���N�0w ��hCaiޅ��,�%������:Np�c�'�Ox�ȡ-p,%;%gP���#�&"�F��bR�Qv8a�N8cEIjBOş+2S��Q��f0?��c�,�b�
��%@�� B��A�'�p���Kաh��s� �C��`�+:3=�-[��+\�0Y9 (/%v�kc�0@�蜚�nR��<��B�'И-˅!A0Eؠ*���>���0.OeP�ň�zG#Y�`�dE �l�0�P�1 N�v6�uV<2
҉h�H���``�:{j��`=��k`�G�0��m���!^/��F��? �d�pc��_�
!�u?h�x��6��q�E�� ](����ov�����/l����O
< �l2�a7�Ot��Ŋ�_�!�Cʞ%(��%���S60-Z��3�?���݀ls !	��!T�˳*_�/���vG2?���1&�x���X9\����foU\�'�J���h�����h�H���,2e�* V����8�`���[Ǹ)6Lñg��	�`hϰ���[Q��SL#����d�X5w�:����-?��I�0i�U:�K�re�ړ��X��(�6Λ%�M3.�2A4�p���4I�FY�NA�^ɲ�2#���x���2I�P}k��
^6���4 �%����4.ԑ��ژO	�uI"���M�B]Sq"�^6���d��y'��z�4"@5S�>@����xB��gVd\#a
�S�p��ע��gLx�1�����Qz�-Ưy T�6d�dQvpC���$T�n�'�>�A�X�Py8�PքIĊ����.\��y��ْ%r� C�[�p�Q&�D��C�FA�����D�n� �i��2:KpXX ��L���<r88A�P�ڪl�D�S�ܮ���O@�c�$,���[wc�ʰ����E�"F�٢a�=p;>=S�H�#����Ti��F0�]�&�[sh<��EDH�r�btFG�{�̥�b�QZX��Ɇ�Ahj(�)�Z!���qe�K�v��O�t��r6�`RS뒮l�ur���8��%I#On��$��,c�y�&}��C�h"��yA�K�w�l�1g`�C��XR�	��AIY�-�ب�Ps&�3n�n�<���u(�[��i�",��/��ԉ)��ɥ$�y��mD'
�Z!�\%Ѐ`"2�P�k�B��� �D ��2�x�#)�8R���R�|��Q���*򉌇w'J�rs`�4<���[�jϮ!��T��]�16�K�V�hh�ʸ�!�$ˣVIʱ��B�<�,;DI��W�eD݈L!L��W��1E�V�+��
!RNơ�̟,�b��|�E�ag��25���7��B�2�/>4��G͓>�d�2�) ;Є�q`Y�z�,�c��w��T` #����q��;�z�JG�,�	�Q~�\J�b��)*ŉ��V���D�a��B5i[%QإAU�
�&1��q��-r�*�ŭ0�-�j+�̈��ޡ`��z��B�3�L\��kJ|�lC`c����}�`��Pp4�B�j��.����/��; @�!¬3Y0`�J	�� Ik.Y XD��'d� W�^7�`�@\I�T�:V��w��i	#�J���i�`r�87)�U���Q��j�h9��P��N���i�!#�����H�ll�Ɔ�3,�ѐ��N=\�6��dF�-n|,a�؎.��軅��K��ʙMЌ�=���L�p��vz�� �zx��f�G.srd����D�}�v}x�-"w#���B��%H0�p"��;@�|
�ظ.�A�Dc?\OhTk����l��Aj�[�*����9���?X�8Ȓ@c�m"�ɩb�T�O"v��uH-
2�Ɉ���}Qqg+U�N��BW=o C�I�����V)�$X���	zSyZ�I͏l:~|袪C6���藥P&��ؐv�?=!!�
�3t�1�̵"�L�B�n�K��{h<�L��=��<�G�[�h� ��[0h�p��s��~�-����o!�9�&�F�9��ѷ`�R�K��k$�O�0�"w#�O�8���I�N�<�b�C2I�"��$.�:X2p���,#~J<��ew��H��@

FIR���&q�ד R0yKGH�* �,�@Ő3���<�pE���Q�eR5q���Z@�
0_#P!P�n��uS�	Z��e�
�)���[w!�DU�C�J
��S ���6��SX){��"T�*!��N-o�H1��ղA�Nc>�q5�@hÐX�d�*#fE�]�@�(!"O�q��o?�HG���jܚU�\(�L�ئCw��4�`M,Z�-6��DxB��,K�$Q���?@qR̓Vl=��=$��=k���3'	_-H�����`(C�ؘ�3a@<M��Y�i
�$��Ȁ0�'/*��@�m��|�ЍYt�\c��� jhTL:�� �:�vM���Z1�����{�&�	6_�t�#A�g���N�s�<'��(� ��_��|��)q�4���"�� !���uD̽R�(S	)���Nޤ.�r���܈4� qؗL��!�dA8lV@)c�I�I�Ƞ�Q�-t����107K�&Jm���5�����2�ٙEHb���� ыu�Y�F�0Y0�#"*lO��[b�$�Th�W���4�8%��@G�@0���#k'���o�1��(�섢,a{���}�ʒm�42g��cCҸ'�@��Q�A+!Bܳ0�j6��Ac����j´�,$�ËV� yc֧��̆��"OVH�D"�1��`�C�)`���f���I/�,K H�5=?
�zF+�n@l�$�
q�S hs�N�	d'�9G���|�z�����3<|!�d� �@0��#A@��8HpN��y��E�.4ty4+�t��Lxd^�N�� W�~ϒXQvI� _p04����	��]������t�#���P\~P0�-$zS�a�6��heƇ'�R]�wE�x؞����
�C��oH��Z R1�>�ɉn+���o-@ZN ��H{H���������)�31 �S��L�;>��3��]!�DCL�d��1`"�ѡ���D�:0�T!O�F9�!{֢]���RT�C�Mq�X5�w�@�1�,#@uȠI�m��r�'̤E��ڋ~	b�5��1TԔ����J˼��g�G]�La�%H̠U���I�'VK@�E�8�q��#R��9p�O}��R(�,ce1�� (m)��Aæ�?1����a�9�"��"��6h����1�p�-9� ���O6�R �=ɲ�[�D"(p�h�d�f\�q�Y�/|��'s�R4ʔ�� a2�z ��!���(H�q���<<٠1%ޫn����'e�-� R�X��vAx�O����n�2���)/^X :�-�nC�51ch�!�"SQ�~��deͬt��A;#&�v'$�y��IY��蚵1`Q��� �X�g��c��ȿ_��H@�f=\Ox�W.6��1�BdfF��\�E���AW��3�f܉�UBf�݇�I�'��4���*Fn��Y�����c��bå�~�̛c��n��&Ik�I��?ܖ���̌H_��+ ֈc�!����N�	�7J܀1��ϐ7�<{��E��d33�� � qc��9	��`�Lu�Ã��D��,'D�\AS�ZP�[ ��2��U��M�p���y���&&� #��$�g�'��`A�ԇ\�<3�,F�B�B}���;�	�.2^���af�q4�2��l+�@�b�)���(7��y�㉕>n���"b-��'^,#=�R	��x�4�ф�߷Lb1�� X�2B��.Ƙ��%�3W`�"O$��u�9zn=�"�=$#V(��'V#��V�,j�K�O?]�e�B|>��W�Q��qB�z�<�cTrb�z�$Ɔ"�}s��q�<�e���]e(�Z�Y������F�<����� �
��G��;��#` �T�<I��}�t̊��T?�,T��b�~�<��c�"m��|pEI�>�i���G�<i À�B����|����7�y��)�b���uEJPӕᗖ:�����*as��*�;dϐ#�T�ȓBi����"�?=���BĀ�Wvd�ȓZ���F鏣sH�R�N������ȓP�A;�+�/��h6c��W:D��m�9`���A��X�(E/)r,h��V��q��=�F	��n��W�R��02� pi�.|`~1(c&�&J�Ć�S/�	�����|?>3�@��l�Tńȓ(�0��4.)!�\�[V�6�40�ȓ0����	ݨSƒ�: Ő�u�p��E�B(9�MӻO��*`���'lhQ��J�ĥ��ߝ8���Q�o�Q6���;�V�2%W�.��Y��k��*�*)�ȓb���*�� �������L�Ňȓ(*nQhdn�3��YZ��+�^��ȓ9���W�KJj�k�Ν�/u��A.%zg�Q;~��҂�7 A�A�ȓ���T�^|�h�
�|%����k��wF�dPU�J%M:���ȓ>[�!�t@�u��=(7��>H����M��)~����@y'E�ȓH�6��G.��f�n-�e(�	MrH�ȓx�p|��j�Hr�����p��x��i��]R�įC�Z�r1n�X��!���(�&�=^L,���l}{ (m�ȓ;&�T+Z�.@���$��漌F|�g�z�ty �+��XIG#]�y"Ι�?j�L��e�,�����~r�gfc��}�3MD�9Z�*sBĮC��D�v��;�F��5?�R�J���']��m�|�"T�d��a���Z*+�z8)�#՗ +@�I�|h�Ǔr>PyE��25D�����?�l���c��-��,{Acԙ�?�7��;k:��Ӳ�O�� ��B���eXt�L�����L���E��PY��M��u��u��ɡ i���83��i ���Q�� �#��wfP�-&��'�v���'��TC�2���MS
<-)�T���~B��h�P�aQ�|��	��q��	�F�8��pcG�кqk -g� 0i��ϓ�����!��ͨ�W%]����D(6��<����6��"|-����G�-ȕ�m͈<���I˖=���'xJ�k���0|z� ]$@���0��	V��#�E�<	���<�p���b��i>a�B#�T.��(W�#����r���y��r4�$8B�|����Q��M��$_�`�3�O�^���uϚ�(N�Q&�pG��&�X>���9An��#��Im�xH���A�	�[�Q>!�O+�aY�a�+���.� �����[V�ɀ���	L|j#�ڀ����ŨF�RM67	�!��ɯ�M#�D�q���a�~�K?Γ%��	��o����#��,[��mڿa��5j�mQ�~b���U��~�3ʺ��ea��f��F�9⢨�q`q�.��S��%?I�Q?O6��
(���@�a��2i��^%D�t��2-ލ�?a�'�PBdj'
��4G�K��b�� q:`�"f�_��y� ��~#T�;��А�� �\�H�Pj�2�Y�B�26��<�@��pϠ�<�~�sn��2x�CT �
?$�"jV}ң\"8T���y��	�$��;��V�3&j�;w+�_V���B�}ƶ�"f�|J?�������O��́&D�#T�jP��_A���A)��hC<JU�F� K�q�D���^������)��P����:q�C5�!���5��1�%I�1\�=��@�m�!�$ƕ�0H��N7_M`qX1�Y�t�!��ՏOW�P3 ���js�h%!�� d�Cюƽ�yv�	�[4�<��"O�U���7� !���>-
i6"O�\��/�b�aao�|�\��"O
�Hw ���{R���pJ )3"O,N֔pz��*�x9�g"O�����d|h�闭<4之�"O�����J�@}��'�.ƌ���"Ofh�'L�|�QB����س"OH�P�&\PT`CG�ס(�Ī�"O�t� �b勔ϗ�5/z��"O~pBpǔ�3��X���J��A��"O�hz�!Z$� �2J�1��Q9"O0���!��a@Z� c�B
)��#�"O*(� &��D<@��A_����"O
�"R?���J(_P0�*4���y-�u�
��,��Q>���D��y�9!|V%`�bF�H��$�y�f�~RL��C�f�D�g����y��V95K`j�g��.�HT���yB�T	K��)�6�{n�e0��R�y"뎈l�x�AXp�$�`PE�y�υKڤ�Z�z��* �'�y������ a�Z�pҢI��b��y�G9.Z5q�jVi�|
�
η�y,�	�BY2wLV�h��u���ք�yBAWO�v(VP��0y�*���y�H$�J%�֬BL��MP0��	�y2䒬M�<�	�'���b��nҊ�ybF����[`��#��<e!�y��Y�3=�t�Ȳ~�D��L<�yRȒcPh�w�,�h���$�y"���.h�)��¿nf�c��yҪ��W]��䇔+f_xc�.�1�y���d
�,v���d��x3�W��y�� ���q���&/~�("/:�y2	��y�؁�	ަr�29�q�\�yB�ۘw�8��1�ÝY��L��/F��y��^�\舃k�D��8���y��K+,\�����젰P@����y��ȗ+��U���*8���sW��*�y"��	�p8j
Ψ(��1����y2.��ka��Rԅ̀$����"���yB�5�&I�Ef[$� ���y�iI�-u`��Ɯ��<p��N��y�� vR���`Q%c]DE��J��y�`K/y(��iƠX�G����@b@"�y�&O����  ��Er�m	&<�y�)�0W��j�M�1b�M�f �yCH�x�`pA�i��[4d @����y�3�$���VP�#Ɨ�y����_� I�a�T�sN�\�BIA��y�C6^ژhR��/jX& �i�/�y�e���-`Ѓ��Uw�2q햿�y�eП=m�L�Q�ג`��|��@�5�yb��>E�!�3C��Z��-h�m��yGV�3+�	��H�=U�����y��O�bG�� �Q�49���y���l��ʃ����!��y�fܩ8\6����ۀ��x7���yb*�>���k� ��1ˑ�I��y�"��"$| 1Ǩ��(4dA���y�C(uS ]ے��UD<Xr`���y"J��e�iZ����NVF��	��yRa׈y�� ��[Fߚ��� ��y
� �B1�ױ� ؠQ� i��"OB c#F�j�R��܀VMƽ��"O�̉6 �
p��S�$Ïe4��B�"O�З
�#w��(�bÒ.Ph�	�"O&��a��/g>���`'�*F5���"O�Q�A`�\�Z\AǬŁJ0� �&"O�Q��A�8ׄ��M�l2V"O�� �)ڻ�11�P�G�$� �"OR��R	ܼ'�e�p"����7"O@@��kB!"�nly4��rŀMq!"O�:Qo��V��lB�*B�|誁"O�L�v`�0%<����� yT��A"O�m���H����%K�{���"O���AL���´�ӄ_�9W<0��"O��	t$�-.�\9DcC�Xt��8�"O<�r"����ܲ$gf]H"O�����Ձ4J�b �	�NP�(�"O���Ι3B~�JFI��!9�ek�"O��K��ԬtZ&�r	��Ez�y�"O�y`3�B�
 �%%Tv2%��"O,`WA	�;U !�_,y"�� "O�	�rF�2EZј$��(Y��K"O��+AH"\�bl[4hҦ@��̘g"O@�+�-�v
���	��Tf֩��"Ol�kv꛶[���Hӟa(.�B�%��z�Iי�e�% �>��C�GƆѳb�<o�@��`U'�*C�I�v�r�ӳ�6�,	&Jg�B�	�c5R�[s��P�^�Ӏ��CH�B�lZ�h�B��{e.D"�߈T��C�I+ָ@��K#/� �؇ _�xq�C�I/�R�%]�t����	^<�C�	"v_ I���(����4���Ui"C䉫p�h<I��H"�����2e�C�	���Ŏ�6D��@G�a�<��e"O^Yxƭ+���� k��m�!"O�d:iL1O5��ãI Z��"O(���`)JqXE�8󐴲�"O:U�'	Y�h���`�"ۘ�S6"Ov�H��O k�PP���n�D� E"O<TpU	X��HX�dB͓]�Z�"O�be/�	��2��úc�\LK@"O�|�b/Ch�ʔ�ԗKJ&"O����͂a߾��t�N04I,�ks"O������H:<Iz���QZ"A��"O �Z�^'6���`B�˝
1)JC"OH$q�E,}c��Y"l�:G:5�E"O�``Si��=`��"�Q7=�D;#"O�\9��/I|$��q�Q�@� 	�"O�R�aK6�	!e�c�v=��"O��Re#%e�%0A�U�.(�ڐ"O��H7�SE���#a�N) �*]�"O�h�R#�u'�� &��²��"O��bBI�mS� �0�	�"Ox�P#��T<�oO�n�P
G"O>��5EZ�_�l�;q �7'Z��р"O�}P��݊p�<<h3
�#oS��V"OZ���D�L�U�D	�j����"OZ�j��ǎ��!��1{���2"O��{��yjT��גSZ�b"O`���[[�H����p�f"O��*����^����1��9�"O�=��N]�����	��bx��kr"OH�,�Q�s�C�i�,e��_ b
!�� @ ���5z��6HA'{n���"On-�o�b�Z�؆�˶Na��`W"O,t�R�\�tMKd�T(cK,��e"O����p��Z&g�/K렩'"OB��",vİ F��S�r&"O�q	@�=���c1�ϫ�	!�"O���!���j$�*9�@�"OF@�u�V�v��{e�V�D4��r"OR,1rd��܀G  �F� ���"O~$[�$��o�D��MA(�f(��"O��ubǦL���S�`�f�3a"O�Y���7��q����]B"O�����0m�4	z4Ŕ����`"O����)w���Vdɴ!�jCc"O���E ����<h��H�F�Q$"O�Q�QcZ��u�0�9��$"O@�!�8P�
X3���R�.��"O���7��e���c�D�$�\�j�"O@��N��23�z��	lkR�!3"OP����*)P�Lܴ%3�Y˕"O�q`�Q0^8�2��&$��9�"O<,3��@�HȺJ��� z-i�"O0�8�F��O|0P�D�4iq�"OL}�󎖭����c�<e���"OHx�U�=i�H��!S0@7̹ �"O�%.΅�pI�>l���p-�>!�$��J�G�����
~�b-�ȓ�D=Pa%�W| �RR�1E����(�:e8@@L�2?�\J6-��%��هȓ1�0���[�0	����T�u�v��ȓZ�9
cm�R��i�"�2l�ȓWX��`���d�l��Q�w%���ȓQ����1�p8�T���!Vz�<��lw�J�ٲfճb}h̻�H�^�<�ǩ�0>�L�׬ӭq�* �e��V�<��LٳgH�Y�RP"z��iBS��S�<9�Ά�&��97j�*D�	e��I�<!6�H"@�hTzŇG�JN�Cf��C�<��o��l�|	�����]9�L�0��<�Dg�T�LQ��Q==O���j�y�<� Q�V�P�	�!^.&c�Ī���w�<��A�^�f�2B�[�h
��Xw�<A����q��%�.M��X��cK�<�h�Z����΅&E/X�5�_�<��") �&�F��"~�] 
FE�<�o���2�+X��J�C m�G�<q%���V���{���
R�ce`��<�ָ4��H� ��$g|5) iy�<ia4"@)���,����'�}�<yC�U�L�:����<(aIy�<Y�`�$��y�A�
!Q�$�BO�x�<auAƁF�X�K6�OB��s�EXI�<1�-�V(���^�d�ȉc�f�C�<��bH0<r\x�ϥ0	
���JB�<��o�%Y��)�Nއ"�x�p�Qr�<��Ød�2�����+�t]y��h�<��i�*�~a��/F9+�.y��h�<)s��/��l�䩉1P��Y��^�<!�e�>r�#,M$.�qɵ�o�<�FAO1h�X8+Tƍ'-ET��T	�k�<��C�t�*y��O�7I���d�f�<qĦ1v�^0�P�β/�tP�C_�<���*�8=/�&rw�l0kLY�<�6�!� �i���/$�;W��S�<� ��(WN�d�ƥJ�I���CE"OJq�d
 
  ��   ;  M    �   O,  �7  )C  -N  W  @c  !m  ms  �y  0�  q�  ��  ��  7�  y�  ��  ��  =�  ��  ľ  �  L�  ��  6�  (�  ��  K�  ��  ��  O � � 5 w$ �* �+  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡*������X�o��!�'w�v�'�fT��
/��Q�)N��Ì�D���S��!��ZW�\�l���畬h!�)4�vܩ�N.^W|06矊PK�'~�	r?1����R)�4���ްD��1!ԹyJ!��[��)�-S7*A6���o
[+R�J�B?�~�'j�˥��GV\S�_����'��s����
����U�_/"��A��<��)��(D2��'�V���%A H����6���a�ʴ!�߶�Q
��ʰ�ri!����O$$��%�|�:��э3R���I@���)�3p根��ɻy��4;��& �!�À"��m��ʿm��֣�c-Q���>IH>��\����u�^�w�X����G�<i3@�j5��*r��m����Cy�<�7��|3F�ے�O@Ӧ��Df�Mx���'{&-6�^��8�qǕ� IHUq�'�h]��f�
�lEqP�CFk H��'E��[�n˨OS�x�O
�@��z�'F6UH��3 otU���52%�'
�'6,b�D�|�ʘ�d+��1� ���'2��g��*>Ri3����@��8`�'�z���Z3M���P�JqU�5D�`�W��\�p�b��1wh��) D�{1%�cҬ�P�/���0�L:� o?:��"�ǰ,�(��k��:`rC��0D%Hբ��ҝ8S��u�R�!Kb��$�<i�4R>��h��jTn�C�e�:�.��^��<��a��n��@��蓠	N�J��@G{J~���ʊ��5ZgK?<���f�z�'3Q?Y����;��6��H_`x�%7D��
��X[��3m$A����O@��hO?�� ���d�BQ�xn	��^��E�O\���8R�����0r+�ds��	�}��TS�D�!���nǋok�U�F9�O4O�|[q"Ԡx�Z����	`��"g�=�Ş8d^庂�%h�8$yq�����D~��3}B��tf�a�&J�!��A�Ar�'�
�yB#��r�D���LN�ӱD]���'9ў��YA�4��gV5�*�"O���..kp8�f�5X����"O�l�2�O�p�V0YsC^.6��mr�"O� @�oע<�u��'ޢ�H"O�p DfQ����S���. ��+D"OF��	Җw�̼aD!(X;@����(�O \��������tɚ�_>Hu���'�H��'�0AQdԷYX<ȶ�[�s � �'��d��ɮu)l���e�7R�t\��O�����w���;�"��u���p��>�!�d�s�p9"�h[�y�!�GOުK���hO����V!G#���0�IO��q�"O�	�r��i��9y��W�=h}��O8��1�O0��$i5v�`qG� %��D"O!���'��@��v"��
�"O"81mɈ_>�pA��M��Yi�"O��t�/	{�H��#]�
:pXr"O��#��S��fБ�@��s[�̖'�B��>Qu!�i'!q铼F� X�G�v��Ȗ'���*�&��6�����X�C��y@�''���	��~>E@ԧL848n�{b�Oh�'z�g?y��Bc�Y�p �)��ѫ�.PT�<��̏��*�W;�,��
@���N>��Oq����,6�`�!�y�b��$<jC�ɴ)b��3�^T�|�[#F�"�r��y2�O���$���1��xlՁEE*]�x�y�'�Or7��<�F�ߍ|����m* �Y���M�<�c�M+��T"��E�}v|�	Kyr�I%�OJ�`�eM5rI"�ڀj k7�Ib"O����bB�%8���ƛXz9&�O��� �O��YnɖT@��k�F
��Cc�'����O�uH���= -�,*e-F��m�0�>i����Mcd����cB � � ���u�!�D d@R�	��I����2Y�qO>�	I�����D�]	\�8�.xyR�[W���'�S�O�6�J;F�Tha"
YP�5���E)�HO���^�z[�M�f	��w��� ���D�!�Ď�Ynu��[�n�ʐ2!F%��b?Op,�WGӠ+�%�!g�6'Q[���TD{2�=��"쒍J��	�8Up��f�)R�P��-ʓ?4�MP'CL�s���S�C<j�y��)�釋UtLr0M?�*�j�l�<y��'2ў�>1{ ,�*)<���$ �X� p�&�	��y�'��(�-�����7}Tix��5�Sb�����*�C�3v��QQ��|�1O�����L�n���P3�d��Ì�;X���hE�DU(^�h�B!*ބN. 䱄L��0<�����-K'�&A׍�qH�G��?"!�K�1�>|B�]�x~D(�e�I=&�yb[�H���O��w��L�y�5IҗtR�yW�@�<a¥�(7%Py���hf�LQE�9&���~T� '��'��౎J
aDPEX �����Ɠ<�L"�/DZ&I񗆛4�ኍ�$&��<!c�I8;�+GM�?x�pQ�ȓ&-��kpA��10(8s��6
�"����������Op�A�C��k�k�� �{'"O��T�ټ)�ȹ�7��*c.�\��"O� ���a��!�$,� k�  R`�2
O
7͐,r�ȁą�|�����!�DD�z+y3���U�B�7iF�.��|��x�����P4n�z��0�F��y2��C�X	��K/I�ऑC�.�yIV5C�r���m�����r�e���'푞ԧ�j�rn��%ǌ��6��G�p�"ON��&e��v��*kC��nM����8�=)q+����T�C�L>�@'�]\5zu!��S��M��/�O6� g��#� !��)��6�Z=:D�ig�?�	x�'ذ�:d� lol�Г�Ȣ`E����'��2�H%[nv�	�c�/P�,a�O$�Z���D�<E����
�j��AԐ'%p�	�
��$>�S�O���oN�6n6H����y�l���0O���M�a�<���D��"@l���%�2'>�騥��|��fl���4��'�2d�΃3�f��cS�~V0L
��yb��"Bt���V�\��kP�
'�hO�㟼�'a�L�f��w�D`IeLX��OP�S�@��	4�
�O=x�.ȣT�	L���)
�G�}�HU�y��E��+�i��6Ob���O��[ � �Z��A�[`Q8ٰ"O@�#BM��D�#�:,��,cA�|�)k_�t+t(L�nL䊲���F�ꓒp?�cћW>��+� ��B���NAܓoc��$��Q_�\an
�_G`q�p���&�!��)��E`��̭f&Fѷ$�*b!�D���x��$auE��!�D��"�PZdJ�,�ĐƤ�x�!��2+^�0����X	a2⛐H�!�D]�t~Tȇ�<{�p�Pv�	G�!�d�W�d��fO�Sh��5I/�!�P��P�p�� 1Z�D�6i�*)�!��,Zji�X�yEP�XqG�>Z!��۪\H��(�*t'�t��e�f@!�D�H-��)�� <��l�Pp!��!x�d��g�>.�!���S_!���tbn���#B���X��!�d�,�`j'�Ym��d
�N�!�d�&Wz��B�_�
mJc��f�!�$ɁSR�BC��R��)�D�ۺM]!�G�?�������w��l	�gC��!���,-��Y瓑T�T���!u�!�dB�Oi��y�
�>�H�aֆTF!��P#�V�@�*��]#����f+!�;&8d�s�]�E��8�F
�!!��3��´�N0��p���!�h��r�a�(q��$W�!������c$�Kf�:�;�i�[�!�$7'���CY,i�xFO8u�!��Q��h�5��j�r�S�O��!��Ǉ[�01h�>i��p`�^o!�Dܳ4V��#$i?1���2� ^]j!�d���,�ɔ�@&_z���̞�\!���s~�@T�	)r�9S6��#HK!��V /H��5��_i6�q����3�!�$S�plڰ�O�nCT0���e!��>:K��b"׿j$ƅ��	�ud!�Dp��0¤		�C U�g)V+3]!�^�vI�Ak�;0��]�E�S�GH!�䂓�"@)���
~b�iv*e5!��)
~x%b�,��~��P�Wg�3�!�d��~�rweΩ,�ҁÕ��!�!�dՆu?"��@��^gZaI	�!�ܶ����@%'��Ȃ���#f�!�� ���͂�7����i�$b��6"O
u�,�F{��r�(�#JX53C"ON ��ΛiI����*J�a"O~�Jw���p�ɖBkJy "Ox\ B��0	6J`[�́4]�8�'�'�R�'P�'CB�'��' �q��M�ِ�X ���|>�,w�'R�'���'&��'R�'���'*E���ƌ^�D��k50I ��'d2�'�b�'�"�'`��'Nb�'�z�9��J�����咠w�:��'���'"�'�2�'�r�'�b�'��Tp�B�o,��5C��\�DQu�'W��'|b�'���'
R�'+�'h�-�CGCxp�����+o�!�'�R�'b�'�B�'R�'��'�jY�CW �p`W!�#{놨�d�'!��'h�'�r�''B�'%��'����V@<���6�K/
����'���'5�'���'m�'���'U&�@���H)�hIR�V�J�T�',��'���'���'��'ab�'	 ���l���1V�_�$L�����'���'
b�'���'4b�'�b�'\Z(ˢ�ǩo#��j�O!���G�'E��'�R�'��'��'���'K���G������P�]�R�'or�'���'���'��'W��'a�/�n� L��� ��#c�b�'��':��'���'4�7��O���J�SL�B#O��V�>�yƫ��%���'��W�b>�T����C�������\
���CACx�8,*�Ob�oZE��|Γ,�6��(l��eB�!M��-�O�s��7��O��@�z�F�S�r���K���O�p]�ģ��j3�Hy�	,#���ێy��'��IO�OH��p���5d�H�yW�טcWd��!}�P�h��$)����M�;9BIyu���h�b�P%Js��`��ioL6Mc�|ק�O��D��ie�S6yɈl�ӥV�I��1R�Ӓn7��͖mR��˴I��8�=�'�?�$�X�mb��6;J�������<�.O*�O9mں9��c�iejc���y��!4D�p�&�P��>��	��M��i��>Au���M�� +E��d��I#ˆq~���y:��̘֙O}�Q���2�ΓL�"�j2Kƕ Y��s�P�h�'V�IƟ"~�wg��%����kaĪH%tΓw�6!�����צ��?�'^e^�y"��DHD�� "c�@ΓG#��$i����5}��7-'?-w�����1��p��`ԱZ�.�:r�߿����NPG�I~y�O�r�'�2�'3�!J;� ��÷pj
4���X� ��4B��i��?����
�����򄂀�M������7�[�!}�i�'z6�j��|J���?Q��	�j�B��@ �ZC���F8"L��Gpv=#@�#&eji�s̏�p�6h��6hLH��G�5U�d({vgI� �S6 �7Y$<�3�̄�mc�� ��:o:��D�#y���:�aD;����'�)e\��Zf�Ϯ�h�Ҵ��-
Fkٛ����?A"�y{zшԣѕ �-���=&��qw&�B�P�(#ネN�$�I�s�<;ċЄ8&���ѧ[E�$Z4�̨y���iX���ۧoݶ6�}:5��;j��d`6�]�|�ZE�S�M#4��Ы%�H1p?�uh�(W#6��d��.&lL4Ԋ�DQL��ի0A� �J�2�d�Of���nSm�脁ac�4Bںp����Φy�	ܟH�I_�IܟL�	(��4��Q^Yj ���s�1� ��$�´�'V2�'nV�HۓKCv�D�'�,�:cK&`���0�K��,{��b�N�(���OL�$�8�O�pah�hGpP�˒0=� ��i��'��	/'0��O���'��$�,}DaH�U$x���8�9P��O��$�O��TB/��~�'l̔���k�&�� 4+�릉�'��HH��'�b�'��O��i��H�N� (6�a� �ܞHwB���s�����O���Q��O@�O���͋�ǥ����H��b�9�iU���'�'e�O��	��	8(�Nh��@D�Iz���Ԣ����ش0>()ɋ���O����W:XXd��O�?�LQUMF¦��	ʟ��	1��E�'-��'��O6�va7Uo��� �p}���S��ۓ�1O����O���څ �d�!P �I6�0bQE��Y���n�͟�LFSy��'3B�'mɧ5��D	\�.`KTm�<,�� ��$�c�v�O*�d�O�D�<��[&E ���o�@_\�C4nӽ;�uJ-O
���O��$1���O���� [u�,��T�(�ԳB�C/el����O"���ON�T ���O���1�^bހ�� B;�4�?I���?I>A��?TI'�~���,@�`Ӓ$�RUS�k-��?)���?y,Ouq�	�|Z��?�8 ��M��Z���f�(��i���|B�'�"��-iqOf���f�Ea~�����OF�;C�iwb�'r�ɸb�v�Ov��'����ͯ.3`���,B9䥙�.�e^�Op���OVA���&��~:2�9�� ���3���� �ʦ��'2�X]ƛ�M�~����#�� 8QB�2H�)��h#�q֏n�H�$�OF���O���OK�H��4��L�U��>2?J=��
\�d7�@lE���ߴ�?	��?���o����gZ#G$`f�]>/�|�%%�S[:6��O��D�O��$�<9*��D�OH@!g_w�H����E
H�¬������i�Iɟ��IY4�H<�'�?i��m-��"#�P� )��ώ�����iO��'���%��9O����Ob���D�? �ꐁq�T�CE(C�4���i�RŏH��O��O>��<	jמC�=Aq�L+EF����-�/�fX���Idy�O�s���ɚk�p[���CÌLX@)Y�dT89fcHwy��'���D�O���&�X��,�� ����ܬZj7M��4�1OJ�D�<	��i��ł�O+�X�v���>v�z�F$@*��b�4�?�����'_�4�Bu��d�(�q"��v	C��:��s�x�'����<��dNw���'� Ɋ��^�`��[�#O%h�m�$'}�R���	jyB̐���=����+�-*?N�ab��o��8o�柄�'bH۝��S�|���?טȘ2����-���&�9 ��OX���<��)Kf��u�F0n������%���P��D�O`�P��Ov�D�Oh�����Ӻ�ɳ�K��FB2����˦%�	`yb&¸�O�O�d�j$��7Z�:d���
�bY�dj�4/��,p���?����?�����?�j���96�Z�K��A7bT|V̐����a��b>m��,6���q�O��1��:dc�%K�4�?����?!�G�ʉ��T�'#��Y�*Ŏ���aV]���@i
N7��O0���<9qZ?��ן�Iǟ;I�x���[0ب��0��F��Mk�eR[b�x�O���'$�	�x�4�4c!^z��j��ƥ�ݴ���O��O|���O���V� ȫ$�aC䀷5��(�$�� 	�'h��'�T����w��� �>��p$H�W��k��ߦ)�	my2�'}P� ��r����'�TH��B+��q�D�	/|�m̟P��o���?�-O�1
f�iɤ-����бR� �(b[ZE�I<����D�O�� ®�|Z�	p���t ��^��jFnz�D=+��i��OH�Ļ<����m�	�Xh������[x�1F�R��n6M�O��$�<�B-@r�O����5�K�g���ٷ�S8D�@��@�M#.O��D�O>�$�O�������G��t���
4�H&^h�q�i��	;u:��47���� �������^*��1���J���
Q'$7���''b�'Rġ~*)O@��]C��ԦHt��U�� Br%{��� �Ԧa�I�P���?1�J<��b���e�,�Ⱥb�>�0b�D�=��ߟ���矜�'R�g���>h�p��l-��ŸC���@7��O��D�Op�B�<�Oy�/��s�Ƌ-�)�p��T�!
��ɍ�ħ�?����?	f��w��]�D�Qc��yQ�h����'80\�,�4����O�ʓw�\Y�5���t?�iz��Y8�� ��i��I�|�'��'���'��B��7f8@�fV2j�J$���X�N���f�����Od���O���O��	�����ڞ-��M�\�uv�����;T(�������X�IΟX������$Iլ�Mӳ�57PH��HD�B{�iPcJ��p����'B�'z�'d�I��d��n>���hI�)��&A�G�t�(�M��M3���?����?����?�b�F�x��v�'z���r b��.6
I11�Շ�6�O���OX˓�?�B�|"-O�������
�"�"�`Uř�RZ�I#ش�?���?!��?�L�!�i�"�'���O\� 1�B��3��8����)��Y�}�T�$�<���H�0�'���|nZ�*0:R+��f��1�6��/��7��Oh�dC i��m�䟰�	��?I���
YH	�Ǯ��Nl�C闟5}|=حOv��ܾv�����O���|�K|�B��N��<K ��i9ld���u�ҕ�)Bڦ��I̟T�I�?���ϟ�	��p��kPt���ٶ~�@��0���Mc�bL��<�g~�O�Z�.��EO��C���ʁ�^�)��6m�O����O�8vئI����Iǟ �i��p#��,W(9o�5c��4�c�>�*O4�����S�X�	ӟ�hDL�0x����B`�1�؀�)��MS�F���Q�i7��'���'.J��~r#!mD�ce������aB'���JW;��<����?����?��+.�1�c��M������(�z�(�?;���'H�'��f�~�-O���'(��t���NEI1�*Z�|������	ן��	ݟ��O�h�kӜt���,PT����!�"��sj�����Iȟ�I�����cyr�'��ӝO�4܊�U)
^�B,tV�J`|ӆ���O����O �D�O���q.�Ħ]�	(s��ܻw�� p���w4�d�Ms��?�������O��+t1�x�D���@�`I=c���I0� �sB�y�*���O��d�O$�SÀҦ��I؟ ���?qX�eQ�o��p�U��a�e�<�M������O��Q�>���d�<�禉hd�|I(�
A�D�!.�Ûv�'�B��
��7-�O���O���쟰�$��D�$�u�7t
)p�H�5+��'�"*���By�����X�e��6���2�.	�%Ϥ!� �i���vHq���d�O4�$������Oj�d�O �j@X�M`	�6Vq�۰�A��J��$&��b��͟Q���>I���^y�	b���M[���"�?�ӥt����'��'���u���|@(���*�^�hi@���M{���?��{sPX�S���'���'F�����'X�%��	W:x�����l�L����+]��nZޟ����4�����騟�	�Ɲ��`���OV"e|���@�>9v��<����?����?����i߇6��J�E�'��Ys�Đ��Q��P�M�I㟼�I�@������?1(]7(��jF������C��]g����?	��?Q��?���?I񌌰)d�V "� и��#�."�*�O�;-�2�	�i�B�'D��'@�S��I�g�v��}�e�f�BHQ�v��J��	�ش�?1���?!���?���eu���ѽi��'��˱쓽PܼQ0��%��-� Df�T���O����<Y�7$�,̧�?��o�xMra E��L�2�I�)��㦱i��'��'q։�d�`�H���Ol���|�K�5J(+iȦf�NQ�w"կZc�6�'_�I���㣈{>]��� ��M��"ծ��d��ǤsΙ`�ͦ���ӟl�kA��M����?!���*���?��K�e��L��:k}��:���P��'���IM&�ry�����l`����$&I�<H��i�r4�n���D�O���������O���O(������DV�� ��X$:�h�ΦA��H'���B�ܟ@Rf���ߴ���&Px1�ꁔ�M����?���Zw�-Pſi���'�B�'�ZwJh�ːbUhp5"_���ir�4��o���S���'��'�2����m�>yꗍ��H-H2aoӢ�D��a�B<�>������ʪ:g2hI�+g����	t}��M)I��'Sr�'��W���&�J.|�@�����p�l�@�ʞ�(����J<����?)O>���?�D�� kM��X������zKؕ������O��d�OʓFq��4�v�� ��Р���H�x��CV��I՟&��	՟�Ն�ߟ�Z�i�)�`(M�F�𴋃,��$�Of�d�Of�X��<B���DA�1���E�և@P0EI�S2F�6m�O��OB�D�O��,�O
�'A.��QާC}���*�#z\պܴ�?����:��$>1�	�?����S7�Xr��V7fA\<�7����?q�0�:\�����S�ToE7 ��ؽV�jY�1l�;�MS(O�@��Ϧ�Ү���D����'a@|�v�_X�TjW�J�����4�?���N���c����S�'tH@tRo�1��!zu�!���lZ$p�M"�4�?9���?)��5ǉ'~B��?E�}�N�$]�c� ~46M�7?!�(�����Q��"�::�x����ѱr>����iqR�'����r�>Oj��O������I�Q���_���C�!��T(�7M;���*�T�'>��	�T�I�vi��"�k9,�pl�bF�e@j���4�?���QY�'��'�ɧ56�ǷQQе�R=1��<�u����$�k��O����OJ�Ĺ<�4냨/�^P���L/c[J����z���:�x�'�r�|�'���ČL��ꂋZ�����)�!p�h����'��	柨�	[�I��5��Ojf����J�\ P	�㉭{#�٬O����OL�O����Of�����O�D g( 5%c��M̌}��`�Fc}B�'."�'7��=^&�)�I|:@M[��\�䢍�D����AG|���'��'���'a6p���'4�o
��ӀI\�m޴�Aߩ�.ioןd��[yB"� ���������#F)�k,�q����w��:���J<y��?)lI7�?iO>�O�0L�p喯zbK2(սW�4���4��,o���n���	�O@�i�k~B��3l/�y1��L�8�����M{��?��̋�����O3�M""��J�\�Sq �*N�V�Rݴ�X�(c�i���'�R�O�*O�zq�A5�ѝi
(��2�&J�e�'�BZ�\ˌ���O�Aѣl×U����b��������)�������F��'���P��rL>���C�lD<z���@�x��4�O|����?���Sސ���b��<,�,��MS,N�ڀ�Yo0���U�6hoZ���I�������Y�(����HZ�H��p)N�BO.�d9���O��D�OP���O� �H^�B�ȉ���6�f]bĉ��.����?����?�O>���~b*ӰW��=ra!͗1D<������M���K~��'��'���'�dH�ҟ L����7h���BT�W$FPbƷi���'��|��'��ɌA��7�X�<? Yp�N/9$a�"b��y�IԟD��ݟ��'�����i"�iϏd�f�Y���r��4P�E�G��n��� ��Y�B�R��~b��%6�X��1`�%�b���JצQ��⟨�	��#C�̟���[y��O .�8�{W U�¦D�U�>%�i'��O��Iwv%DxZw�a���*��d�6��PөO2��\�E,���O��D�O �I�O>��h
X"׆�r��x�G�OEh6-�O�ʓb�,�ExJ|�^�$���`ܯ>�,�D��ͦaRE�ܼ�MC���?���Z���_�i�p\��ꃞ��W'O�Pp2H��	ɟ��FO��fi�tDܻ^0�XC���M����?I��\�r0��x��'���O��3Ъۈܶ豓�W�M8L[2�DZ�{�1O����O��@�劑�� Ш�(I���L?K(l��tX"�����?�����k�߱B���`�����b�U@}r-)��'�2�'R�'�B �G?�x�c�V4X����u꼔P��'�"�'_��'=�'^��O�:�əw�ĩ E������ۗ�i���h�O\���Of��<)d�	Z�J��-"���	���&d8F��ٟ������?�W�U�TMD2`�)aàuԖ�r�٫��d�O����O\��Ol-�L�Oj�d�O����O�;r�󑠌�}�b�.�u�IJ�	�p�'��YL<ɇ��*��)r�h��[6�@�dm�ۦ9�I�H�'��b�!(��O��ɜP�? ��Qq.T�GsR]yG!�?*�A���x��'U�@��O��&��(s0IV�W� x��+K��b6͹<	�n�3Z�)�~����򔕟T!h�9���E̕4�8$K��h����O�
��)���m��](�.�=!X�{�ND�6�%h(o۟�����������?��2k��m���]#FFY��\:R��԰�O>��� l�"H	A
D�GJ%�b�4b�p���4�?����?q2��?	�����Ox��G���X��ʒ.�Y�ϫ:}J!���D�V�Ο��I���f, �R2�rF�S���b0O���M��b�`�V�x�OTB�'��.�B�Y�L6~%p�҇kT5NB\�'�(��y�'���'��'ݒ\d�A3'��\ZT��+@��FE�B��I����I��P&���	@?�窘�0��f�މV[<�An����hG�9?�j	9�us�)ԭ�f���$Z
:���'Ejd2!�vkv	`c#��
�!�ȓ�pLi�n]����#qfd�=��Q86� #�)s�`V��O2�S�bj%�l JV2u(P0�Ư��k�F�+�+�J�Lu�G�$d�r�م��H�*A�L[(A@��#E���W̶1jD-�~ݜ�i'JJ5U�ZX�U*�,��t ʑz�� ��*�^���'OwyL�h4F gזp�1 ���aϟ�I&(�C����`ޮ �t!���ܟ���8lq#h_�}~]@��p�LT�0F�3Ϩ%�O�zE��Nמ�!��aE�PP�jO�<K#���"��4U
�^tu��%�93�K��g�=#�L{��V��V�U�s6���L=}��!�?��i��7��O��?A�Ce
�|ؐQ��r��L��0�I����ɥ%�l�0ʁ^~�0�	�&O��DF{�O��#=��bS�>nP�s�rb,[�m��6+���':��'԰t[�FY=bq�'�B�'l�Ƌ�Gv!)�eu|�@gM�op�B�F��P3��mZ;*��(�o-�3���5��|�CM���b�ԡ$C�TTD	1~�Z��`���g⅍����2��
��b`u��4Q�D�e�i7X˓.$���i>]��A��%��Q�n�O��@���1Tn�$�ȓ2�Q`�Z.D�,��`�,U80�'w�"=AY�0�'4@˃$�$Y�։Rዎ�y{���ph ?M`����'�"�'��$nݹ���HͧU�t9b�B@~I ��� B4]"P�	� ״H0F�E>`�!��]�0k^�@��&�<׀81�L�(Dк��&��s�,yB���h5��)�)o8�j�v>�H2J[3w� !�M>qJ[�V.��a�:)P�h8�g�	%.�I����|G{���;W���Y׭ݳ;`�mӲA�
C�a|�|Bm�!I6j #N4Q��i݉ޘ'��6��OZʓ!�jԀE�i��'b�2b�ωTF%Xt�ceց@u�'���C���''���-�fI����9��Ц�H0@h���c�t* 9b���?f�U ���e�'���Sd��G
����:�M�[�
u���J��l|�e�7v� �	���b# ;�DU�	�B{�N���O��
ڂ!�)2W��'e��'��O��d�O����O���֒ON���c��2�&вE�y| ����E����y�}
��.#h4�����* t�m���O�˓R	��ȧ�����'��,,}��
��!㔈�/�u�ŀ�KS���	� x F>L��7��&��5��Sc�i�|.g�v�K��[4-d�6/�of��'8�SS�S��e�@�Z�vi:��Cq��ݩR�R�0��m��jէGO��V�>�V������O�"�n���jA&�`����� T%�y�푮`�ԋQ��ZL�Qz�EP��0<���I)V6�z�f/|I"�+�nޱJ����ݴ����OH�e%Q.d��O8�d�O��&A�,�K�԰ (X�d�i)��j�2>�Zg(L�l��d�0��B1{��p��6O�m[B�%�3��ճ0��-�F��,6��K"�[�r���ˠ�V#k
q�e��\.�y"�Y���tHf푕:�q�t��%�rDmӨ���.����Y���IIvb]���0=��sΏ�Ԗą�0mlܳ�_("����n�M����?y��i��7m�<�O5�TV�����8v�`�U�R5��`�!7������䟐��ٟP����u��')b0�ZP����c�vl�tꉠ	DL*W�vl�K�˞k�F�;��H�޸mb\w�Σ<��R}�X�Ae�9 ���ا'+d��4�A/tz� �L+b�SQdj����ğ1di�$À��L�8�V=:�dы�?������?щ��'��ZUbҨ%>n�� Fө@g�3
�'?ybb�ÍLT��W	G�l�j0��y��x�Z��<�''4���ڟ�z���\�$J��U.@�+0j��,�I)}B�)������'}��8�֢�*tF�c��FP �a��7j�p��h�.���ߌHȬ���*ʓ�rh��I��E�ӄ9'�I�ܻx�I�AL�0pQD|��[�m�6ʓO{n)�Ɋ�M�3T�쯈x� �p�݈h�컇�L
�'�b�'�0Y�Q`� }a� 
�A�q����'b�6-���|u�l#�H��m�4?��d�<�Ӊ�9u���'�rX>�iA��h8c����J����>˪9���ş��ɎU�u��j׺x�J��Ş�<�O��S;iF^�ԁ\5k�A��b\����'����s�I�*|���U*E��M�D�Tr�'�8�!��:�$E�D�E�|l �O�M�`�'�6 �1�IY�g�? �p�Jڧuk
Hx�o@7Fl�����O���DN.�>��E�31@J]h���Sax�#�r�B��Fc�?"R�ܘ��y��;��i��'\�AQS��<	�'22�'R�w�mZ��G��m�C��F�p�ӵ�ݮ/:h��WNѫ>M����G8z�1�u�W��#�y��`G�x7��_5�iġǝ>@ �$�̒O,���5�OpЙ����Ŀ9Q6t�z"���2�K�ix�5c4��y�84a��i��z����i>-�q�UQ>��hZ�"�.x1�G42�l���;���)B�Pt.�+ǧ�1rQ�'^#=	U�i��P�@�r�ȧe24���[Aʈ)�tA z��2u��П0����0��'�u��'�9�p�AQ"Ų@��Idg@0w��%�P��yBp'_sa|Rd�#'X��X"� ����S��]��I��C���+E�	G�����I*� e!كM�z-;e�1x�����F�O2 lZ�M����D�O���F�&1�p�yeO���V�Pp�-D�x�*�� RX9`��,�>��a�+�	�q�>���CyKO�ם�����.GA�X���$+��k#L}��(�����ږ�Z��`����\p׀ݴ[Y,B ��N�D(c�B�s�h�Aa$_ ���#n\�%�V�0��� ).�<E^�*���k0���V<Q�-#S��L;���H�H�*ݴ�|�g��S��Fy �,�?Y��j؛v�'��!�(���S��I�%��u8�Q�d��D�S�OTz��T$�4%[�c0�ޫ"�.iCf�)�U �F@P5���<v�
\��m��X��W��JtB�6�MS��?I)���A�+�O�1z�(��.[l���-A�?٬0��)�O����������V�r��D�[�`�����ʧ&���Q�M��a����� p�ɦO���`G�<`H��C
GlA3'
N�ffܒ� �m#��ݭ"��4JɡQ�� 0��Y<�'� ��2�V� �1��M*V��Ie��1.@�Tcv�
�k�1O���/<O�H:@m�8��l�3�L�� �t�.��|b3鉄kar+��
���Z�x�Lش�?	���?!���G�
 b��?)��?�;n�������1 �n�SF�8ir��h�?/��rS�ƌ[��@ǻ�O7�l��J�<��&�O�ܹr�D	5T�e��cR�0��`�'A�@�e��Q���V���+�e�O��H�*�yI�64`�5C�:Ӱ �53���k���Oq���'��阄w*�1j�,��H"Q-B����C�+�����FR��4�l����O�Gz�OJ�T�Ȱ��H�la�];¤�� �x2��z:������������+�u�'h":�l�i�GK�	���qY!	��}i4K�F!�$�1�@l��BT<rf6�[q�X
@ch�XOFd�#cJ�>i��)fC̺
��$��L��m�2�'<�'�B�'0�O�a!�hH�S���Վ]unH!X4"O���%I�aJ2��ME�YJ��J��|}"^�j�ѵ�M[���?95�
>o~���vb^9,
�ٸ�8�?q�+:����?ќO- 1!Q��.eDI�q�� M��&�
�t�tqUgWJ�8�e�p<�Q#؁k,�����J*BIٴc�U lZ����B^'`�h��	0ie����Ol���O� ��? �4�H&jS��l,�G"�<��������!FH��ʴ���iH�`�iO,�nZ�C���[qJ��R~.�*�)WCJ��`y����au7��O��D�|��D�?�?j���h�')E�\��A���?������#�spi�O�T��E�r�"�҂�ͭzJ�1i����I�o�p b�� O�a��;+�r�p#�	�[f*d�%��'���L�D�O��$�O�?��&K��l����?1���E'��ʟ���Ɋ;b��o��4�h��W�[����d
@�'�N`S���nʮ��$�-��u�w�d�(���OL����5aGש�?���?q�˿C0��w@A	���+�0hC�-0j0`c�Y�'���1�C�)x0�J��d*��\�<C2!2p���Ef�� Q�@4U����"�1v�,+�)qp˕�T*<7�CW>]p�0e���ї
��1
)m�S%�6T�pm ��*!%����?Y�<���(�n̪\�rݛG�ϣ.�aR
�'np����A:w�K�*-Fh�0��'��H%��R����9]zf��Ņ�?B��(M�\��Q!��)kQ"�d�O\�d�ObѮ��?������H���B���UQ�B8� ux��K�>b�
���<R.�1���=�b�Ey��m��z7Z�zF@D�E���C��Q �*Ѯgﶕ��ĉ�\�=�G�X��U{���L/�'��U��J�� �6��O��`��0��֕�?I��i�7m"����O
>��!��<]���`h��l�	�����$��'P��(�(�0�6y�<с�i9V��Joǎ�M���?�W��%9�]P����<����?�S4��+��?�OJ<�mZ�jk ����Z<.�T�gs)�&�C O��lK"�&{�jH�p�0Q��Ey�.�¦%�g�H�g�"m��<[��h��E72�:�"��_�E���'遶/|��R�*]�fd2�O��R��'�07���Y�I�|�BYql;[2j���ώ|m��'�2��3� �x ��S�Pꎬq��6b�r����o����)|Ӻ�pE�,c�R�)��1q�@��ă�O�n��$��iT��'�哞`�b@��g��r�.G�p^����&R�*T�����1#C�Zb�	���X~*�xʧQ� �٦���@=:�X���&��O��2N�7(���e��5(��!�K�9�*8�KF�fb�'p,U���~қv�&�i'��א_{ ��@2ce������6H1O��$7LON]���	5*���9"�N�	�a�Ó ���|Tb��l1��
�<X7��sy��'��(:cH�,[�A�$ĒI�x]��'�r�&,��*5���ӹDj�T��'���B?���9�!Ǣ9m<M��'�<�Ӄ\�6n,D+���6%�@�'��3V��Yk<i��'��mj
�'���#�L�)R����a� mL9�	�'�X�견F0=� �y�O������'F��W`;a���0�v\��'YS�ʒq���1� щ|�^|��'-�ī�!�-�����)�t,@�'�N�J����RQ����y����'�(t�t��}{�<�B�	�qՎ���'aF�C��]6����n^h�X��'�4ܣ�l�9A	��/̰5�	�'5����㒪c�rp� �� 7 �a
�'CDJ��*
<� +��0��x
�'�4�	�kF]ì8aC؋%�y��'`�d:@��?AWD�!%M3&<c�'�r��Ο7M�"(6�]*;T	Z�'R2p�� .!�V� ��Q7� PX�'�4�+`�V�,���aӷ'�D��'�NM��GE# hȢ�E1!���1�'�hș7iD/�����ܤB����'��DIS+D���!r&�$Alp�J�'z@�8��C�D���TO�7^�}{�'5Ɯ��g���� �B��_j���'<��C�O�k*��#*�z�(a�'�j���ãf�t<P kI�H&!h��d�vBj� ��Ӄ&t=PcY���O��(Bt�h�yʰ�G*�����{«5'�ay�JO�:eB�燂���S��+���.�5�8��"O!��1�52O>�+U/@�8G�L	B��^��!�,��BT��'��;��U0A�!�M
,m4�5���r� HY���V�Q��t*��$� �Ԉ��I�G��9�$��D�d��"�$�O�x���6}�z�
f�� �����Ӑc�.��T#X  ��)2eƁ�	,-y���'�=��A'�IZ%U����bC��$�3w!^R��i�K����I)�IԤv�hh��S�<�\w/^�;7&�'dJd��]�D ����%���	 5��� 9uŒ����J�X�
p@���2��$؉OF�5��%pRj�)��q���"��/�(��eˋC�0�ɣ�Z��R�p�BH��~"��66( ��k��Nf����E�J�!*��'9&��ஈ�Y��j�O�8 �k��Jn��O�uЅ��9j9U)�,b�6�0�'��M��&�N:E�0��~|�e�7'�$�����U�MSx0���OҜpz�lp�;���jۤ2"P��G�#"*�6ƅ4�0<��Z/~S5H�q����7-�tYz���
8��ku��06x�&@'?)��^!�<m�|�<�`��O����s$�[ݢ 卅}~��X 7�D!�+;�LYE��J+�}�G�yL%P��_�~Ψ�s��Χ9�����'�|!(��P�T��؂h�Xp�b��R@l��?EE�ÊS�|�I�2*��gy�*�"X0�@#�j��ADSb(<Y���#�Qc�_!=xE�2	ة�4�8u�t�ɣD ,q������DT(��OQ��D��"q��@�`Nv���{"�g;�	
�x8@ O`?��'���a2�ζv�P�gߟV�� �?fs�m�e���D_g�'3x���FX�\P!���L#~�P��[�,�be�7$�%U��䗢]�d��?e�3,�O9:f�&u#T�c�e#rrb�b��O�iP3J�V�v0 #/�`v�88b�I�G��$L-Z�UX�G�4�c�TZ�O�t���x�)�O�ՠQf!��!:(��V�Z���g �d�B���/E�D��P0�ا�ɰ�杁K�숨E�� z5�(H�)_C0���d����$�3 3���^S�`��$Y3L�-��M
	W�b�,��E)Bu3Q��(Ȓ4���<�g�? BT��ڮYd�Q�Y,+�lԪf'T%Iˠ츔M�=e��O��IkAlըb?ﮔ�` C=l��p�_�B+���Q�Z�J�0��B�Q-7P��)�Z��>��~>��B?�y��
�@(`�+���*B @*d�[�4P�g)��NqO\����#�\����"f*�ys7^��9�z)`�/nƸ*'1���pG�\�u*�	PR�튀y�,7��d[�*� e����'`���w.x���∨c��(ӣ
�,`$��)+���8�C�}*`� B�����(���zU��v�ڀ;\�B�E�H���<�F�U�����SmH�!G�������O^��!p�vj�`B���'v�5��M_?B���syRǓ�^���P�#���3{\��;*K��*�#�0�x�!�-q!d����,)B@8C�'����If�g~�Ox�L
#�t����&�t̢ٴi���a�rӬl*���]3h��6! (��]�U�є3�JI�Uś1�*��aݿ�2��4ռ�����l��S�O�@��`_5.fa����)\tj�A
N�pT@�n6/ܜ��{2��W���S��(���7@ F<^������VH��`P�H�  D�Dɟ��g��t�0@"�N����$�y6�S�!2���_ l��ia!�X����S��\̓X����W�ϜK���2%�V��ʵ�Hm����dx�i��-��D)ia�\Gk�XC�'��iY2����VvH�q���%8ri�Ol���0��)yT&��@u�q��.E�"�H�R�E��e�Po�+�RekV��+1�1�RE+��O�RΜ,aE�(���9.�P ����?�L�T`��)��L���!��6��!%?��,`R��S�R�f�3�4�.�؁�S?!�֠��Yd��H�'3�.�O:4�i���@�W��XJ��7H������*�T���*�y��P�Ԁ ��Dl�'n�`��H|�9�U뒛L��a4J��]Kt��O��=>���yZwn��d�Oƨp0g��gVx�0vkJ7�,�q��xΤA�G�E+�qO��!�*��8Ӻ��`a�37��q"�|��8\-*U?v��<b2�4N?r���ł2@P�aC�fC`H��/�*p�-+�>��Q?�իL���ܹ=SX3��7,����Q.В�Μ�7-�q��4��O�i�-'$h C�1[?��栌7IH���N�4T<�K�, ��s���F!׉7�(`�/و\�\1Z�/�Or��t�;�)J2*�	*��6�Qp�ǂpXX(� �2DjL���'7�-K��o"� �=�@F�Q�!Pgܸ'��)r�R^8}PS�3`�b]u�@ty�I]�'Lr�CQ܀ ��5J���	Уx��2�l���:���(����AJ4h9��DZ2t�i;��ٌC�� u��N�1O>��D�X2�4@e�ά/�����C|����!MP.���?@h���@���5Ba�ތo�� �O}�c�DW�Tt̊�#C#��I�o�v�tt{EM׌8�2�2ӓz�(ay��
*\9(͘�lO�|�pl5L�xYB�'�Y��̫��CuFP���'�r�Ӈ. z-� ��Y
8�1ߓL�
쒡�c�R�r��4��H��	�{��F,�>V�pMQ��0Nq�Ѣ"��.�ZU
��H�=,
���|V �J�%�����cmF ���
���30y1O,�	���Py�Aq@D)|��1k�@��P��p��)Xk̓*�q��!H�P�D��c'�&��9�<)P�I�|���0�B=ʎ((�G��B%��c�DM�r
�QlנA���SrLQ|��i�5���YGK4�r��䇗�L�qXw'ν54�@!E#W��az�@�`��8��_�d.J���S'�?	b'�ho��K��8�<tp�HP��}Bg
tT��JcŅ�Ti�Q�F�	��=I���^�$�90�+$́�̜#� �����	��B���	�����3Y'��ϻQ�x��򣉲r�&���%n�|`�?��e�/,#��}��3���jK-C�R	�ŀvb�b��͐:6�	9�&N�v1��0�$5� ڀ�z$�R�onp@��L�UP�牎�HOt=Q��w�!�c��
hU<�$��
-��A���5��m�*dĂI�h�� \�ɵ@H^azR��#V���j(�,�!Gҵ����X�K��+/j]g�ڼ}T⟈�6@D�fS��h�Iھ 0<'�5�OĈ��i�.$C�� �6�:6-(Hܔ�R�Rthp��bC�#S�O�S���+�w��̙�T���F
�ԑڏ��޼�`�|���31�*�Q��/>��ag�[��'�` c�K�+:<0ǧ>�@���y2�Ų|�1*.���f����<�5",n����n��m�X-��Ez�����U0b��A����.1^�� N�^!����0=���9��#�	�!m�0GR�,A�l�4O	2X��𘇤B��|�Nބ5�p�8V�mf$�3`(D��#3��8��i���b�uh�jr�hi�g��P^!*�T>��(�ȼCB�7�`B�i�>>�S� U|y���Mz�{̝?elE	�?=����V	vi1O���F)6����W�F�`<��w����'|����K��+��8��&b%ƽCϓkr�9
��"�ƼA�OJ8�NYa������W�;E���t�5Fq�x��.1�>�Q�����OR8�bW$KZ�fִfd2�HL>Y�nƔ&�2�J�)�3i�vD��&ZJ�#o�DP�㚖*�X�+g�íq*�3��^$��h��{���i�*-�1�S)?T��F�G�^-q���_S8��G-�/��q�=�O0�X�2�zMx��0b�z���E�g��x�W�l�A��7��=�H��z`��:�ĭX�N�*2�ٸ��'LN�(6�ɘ:
��n،c�J݈�S�z��)��M9v:��c��W�X���	�2lt���ŏF����C���� ne����,��$�V�1VFy��F�n�m���Bh�g�'���ԟ ��ϐ��0Yj��A�#�qj��.>p�����%:v��� �?0K�}���p�N}��ʂ����S��m�S�Ox����;��APcH��0'�5h�e��axr�:�D�;5�Q��y��>�����Ȏ9h��
 ��c�6��S.�,t�@DL4�Y�ʍ�(�ވpe.@K��DQ��!�ۢ)h���"��D�N�3��Y��<1C��4	ޔS�$D�V���SA��\̓G���9e�H����*f���$�*B&��	 ��"#$:Lc�`��"O�9d� r�B��0�>l�p~�E�|ar��'{� {���q���#��Ű9�(�11g	�s8� #�N]^��>W��!y��$��k�|�����Dr����
qظ�Z��"�I�(X-[��
�$�4�������5�ay�Y2)�4����G�&I{�j|k`�H K��W"h��n��7/F ó�D0$�:M?� o.pirqB�Z���U'ИL$a֌��ku�I��ɢ<�����dL�02s�^i�b�I�RB���T7*Y��=���Ӈ�'�
�����y�O?y"�o�!~u�� �녎L�k�Q*$W�{)׵'�%!�&רu���I�'r\�u�M2r�r�X3N
d���3�ؕ��b�J?�1��0��9S�*�6@���e%͒ی-����1a-Ric��+���5��?w�8Q��GB�*H�c��?4l:�b�N��$5�f����8qS@��T�~�W�]�}3�3��h1$*��;��D����{k*a˒�I)]g���C.҃q�Bݘ��)s�Fq���!jT�X�/ՏM`1O��O�ȭ�v�
Gܸ9�fNhN<�K��P�F̎��]!5**=E|ř�>I^�рɑC?ܵ)�NU��yBHM^��,�V	=U��+���3�?��*� k� �m�}mb�3f����um������oN�\m�8!�.�+q�IYc���l�;WÐ1/6�̓u�\b4�F�3��dC�k�H'�a�Z��!�#G��き�I4H	X@n�"K�<p�]}��)�@���Al�	� )�!c����}�i6c��9(<,� �S��+�MÊ�Ă���O�a��e�3t�����õK��\�r�|�fs�ۏZ� |GxR��/�����=Hx�����+dZ޹�w�ƅz\$)B �Oj�@�"i�qq�ȏ�2�R��Q��&�N=[����'�>UB��Q4勖��'�L��m�zul�	2n̿��'��\k���;'u����ہg�y��'��8�7�&E^dx3��-N����O��tn���7���X�xaM��Y�9�1h֨XJ����E�WV�	��!�'���O�]D��;n�q�P��9w�p�2��7D\����).}b�L�+ �y�􄗪W�R��#O�}`��7O� [J���d�e<Tb?��O���#H� ;�0�u��m�8*��'
d�I4�a�'7n]��]>��Da�OQ�}�� ��Q-
��4H[�"[�5�'�F�*��� -�m�=�wa��r��I1	Qr�2�&.����� ��& ~� ��Я"���Ha�]d��O�����1dD�-95�Ln<��B�#Ϫ�Px�İ@�	��뚢u�l5	ͅĈO��R
Xav\Q��T$Ų7"�C#
�h�9K *ҕ�y2�^:]�{A�2R�=�G�͉�y�mP�G���"'-�s��-D޽sW�I�j+�����V�B䉥&�j1)���+9@�Q����(o���Y�r��+P����\LQ��x�d 8v�L�;�J�1.a~��8We�a�F+�'>1�� 2M�
yr����)]�4b}�3!2i����,Qbn�s՟�G|r.TM���!B�m�'W0�J���p�}sG�ôb'Xɇ�4b&�h��ǧO��)��ݬb��q�n�>|h��_���S�O{0��"KN,5I��-\�?��|��'�XA�L���z�lڏF�!k�'����^m�3��A����'gNȰ��OG{fɠ�"_�x���'�2�� I�
NP���~���'�%I�D�W�����I^ ���'�H#�lL�q�=S!��* � �'-��Rq�2lP�����e��'��A�ꗭ3J�Q���l��'x�E؆��3�UY�MR	�L��''�41k�*�b��g�'U�E��'� ��ð3g���])I�L@:�'�t!��a��Q�`�1Xp�֙��'��6�T�;/�ݨP�ȕb�xē�'��a;� ��p$-�'m�!V@���'��0�d�~裇/��S.ha��'^~�Z!刄=g�D�t��I�� �	�'*�y�`M���z�Ȳ*��BF|	�'��ȋ�b�TΤ�R2D�&5NL����� ~|8�H	����Ǣ��XP��pW"O����ӆ/�f)릢&I�E(�"O�$��R5����6c�B@^|�E"O�\�Dd�ZV,�w�
�v��"O^�5��&_0���7$�(L[�"O��S���ay$V�2��4��"O�lJ�Mϛ�D�Ԅ�9�l��"O&���
�JB!��cB�\���p"Od����.�a�!�9kn�`"O���bټ�ph�c�1�:�"O�$�0⎏?k��s�b��t�"OD8��L�?)NA��@*P�x�$"O�	1G.��k���ÍB9�z"O44q���Aw$X���[7C*&e;�"O@-C��J�0��Į$`���p"O�9��PT.�K/��:њ�"O��ӆ� ^��B�LL u��"O<���AS׈�2���4#�6���"O�4p�K܉ �x��B*�@��Y�"O�l�Ǫ�\�,����D�0���G"O�EQr �Z��<g�.Yh�"O�嚲N�:jV=  D3f) �&"OF�����%WS��d�Q�����"O�����K�
̎`���ɻg�x���"OdH�c�y?^<���žd�ʼ�"Ob|�hפ^����O:�A��"O���E�n�Ji�%�
�P�D�+�"O@E����uHH�UK��/���"V"O(a�X(E*wE�D����W� a�!�8y���c%��=D���Z��Ҕ*�!��d\)4�Ыxҽ`wKګW�!�ى@ ���&GI�����j4?r!�ԍA��*��E
�a)P+�^4!�F$q��x����C�Ո�˃y#!��+NN2���&��nFac2/E�:!�dJ�X\p6�m���ht�5R_!��p3�FM��q��H�=T4!�$�:>�,�;�a�^`��g��<�!��7�6i�-�����&�2�!򤖳��IkX���:C!��
C����!��%W��)���c'!�DǤ~vP�TcV�@R%u��D!�6fǸ�f�<t!xm���Ěql!�D�Y�29��(�P B�K�h��Ű>���@�y�f��E,>8�$��w�<9`h�W�`�b@���ep>�S�_u}2�'w@Q�4�عE(�Mx��X�T!�	�'Nr��i@�f|��:t˞��J ��'�����,�+7��P4-O�LWp�<���ǹc��0��J�d���!��G�<�!��dl�����g�*��MC�<1Æ?_lx� �[
eAq��@�<	d��!s��mh #Rwj�8�lOz�<	��P�k��"k~�ZP(��[^�<��ĉ8�r�a��[�9���[gu�<	��Ǐ7�@�B���B�P�'�p�<	@�Ya���˙�X�<���G�<QCJ:" ^�1���k��)`�d��<�,�/$p�iu�O&N����D�z�<�%�/m�����* <k��Mw�<�!�R>Ąa`��[��ґ[���y�<�'����}h���H,İZ��]�<���܉ ��A&b1J�( BwlRR�<��ձ?j�ё��O$_���F��L�'��y
� İ����ug���`ǐ�rw��[1"O����DI&WJ$@,��9Ԅ("O�BU�٤~���q�D�,Q|��"O$`P��Ͳ!��y���W;RCZ�c "Oސ��JH0t���w���"�"O��A��آf���Q�C)Q�"���"O�l��옲!K
�2�F�72�3�"O ��h��cƈ�	�.-j2t�{�"O.��Db�!l0��w��6|K��J�"O6�(�'ܷZT�4��*��N`F! "Op2GႮ+Y�(�d
&'������d���i�:E�*����ìm��!�F�TN!���N�� ��<Z*�aw�I�G!�Ðz�u��.Y�R���,=!��N�v��˥M6~�H:��F�*a}>aE�.H@��5��9qP͞�<1��V't8;6�U|��I�3i������8n�)�@E8����'�5�ȓd�@)�'N�dĮ���ad��M��g$��wH�3,�SU&@�l(��p��)��0���dn�<����%96�%D�0�!jo�p��E!�K��ɸ��5D�X�v��q���Ϯ`�&u�� !D�`���/B.� ��ˬA�5j�L D�,J6��WF���ȳ8����*D� �dM֣z�,p�Aſ6�dJg-D�X��1S�l����nx4r�f'�O��E|,]{���;Өe�uC�S�����
,h��O�Qm����C�,���)�Ĕ0�-^�VG��V����܅�LM��@S�	4qw�R�2�����;���� ��. Ol��a�7�Ȅ�h%z�J&A+7B�]6��5azT��;w�dZ���aS�l�E�C�| �<���|R,R"D@��*� ?�	�ȓ[�U�4ǝ�fl�qc�A�xYX��ȓe8&A�旋|��Z"ΚY�j���Z��
F�"E��"�I�@�
� ��3��C�9p1�l�#�')ʕK�oߪgrC�ɲ2#�Ur&�:zP(YR�])>~ B�I�&�M �i��A��@�g[
%:C��'En�Y`Η��� ����"C�ɏ�0� �g��b6D�3)C%R&�B�I\ꪕ��&U�R0&,��/�*�B�	�a�$�7��&�^��B�MB��${ld�eWw�Fi둀=d�"?���i�9G��,���G	$fLq2+(s�!�DB�F�x�ƉJ7*�̑�&�!�q�<% ��n����Rt!�d^�`��q"F��Gr���g�,	!��X.#���A�Uk`%��A��}�!�ɱQ�`L�Í�?R�������>�!� ��ȴ�2$&4���XV�!�� �i��������%x��v��Od���'HT�WG�?�b���B�=��y��	&����ᦋ/	���ddD%|��C�		D8�m�eI�j�ȸ c�*1�C�I-�=�U�ͥ�� 7��"+��B� K�2&�W�v�sT���l��d(���y���P:]�L��C+�!��C䉸d��
���7��l�M��ٸB䉾��T�7M�(χT?�B�	�"�2emQ�H����.�)o\C�	�&Ԃ`��=�H��nJ�3C�)� ��QQ�cG�,x���SJ����"OF�"mP�M=�L�BdX�GndJ�"O��J���/��H�')^�'1(y�6"O��ѣ37�~��G\.$�A��"Oڽ3��Y�g����&Ɗ1��"O�<�aBA3&��d d�����#�"O\q ���.5j��C�
N�1SG"O��4*|�8 `��7 ����V"O -�a2C�:��Ί�)u��b"O�� #$��e�D�Z�� `O�V"OB	�c#t�I���<撝C�"O��9�d͔���1��u�а��"O�$sS�U6�~	s���>2��UP�"O�1�D�r�n�rW@�7��Ж"O\�v E*e�j7j��/�5;�"Oz�b'����,K0��%^�ɘe"OF8	�2��͘���=��)�"OJ�b�&yI�aJZ�<����_��D{���Ђ���!��F��)�Q�&!�䆒^	���E�A,E��e@!��r���	�*&}�9�Z:���D{B�O�Tè?>���!�Cc�5�0"Op� ���8" �%A�+0���'Z�<1�ӳtt0�Q  A?'_���3�4D�$Y�e�d�t�����B]��n-D�<�.�&n�X��1@��E�`��*��n�_��u!�sz��S��8&���L��`G�Ћ���ʀCE�=��yS��)D�i�d�M���amՔ��Y21i-D���O��w���BD��!F��´�>�L؞�J4�W? �$����E�G�����:D�8I��[�&�晈��B�B&y'�;��hO�."�l�f�D?'wJ)D���iO�C�� uj�+��ʑo΀���)��C䉟��3�� ��c��9*jC�	�B2� ��_<M�	�
ukB�	�Wz��CA��]��[6�C�	�Ez`�₉���`��Ղ�2_�C�I:��5C��Y�a�my�٤L��C�Ɇx_�����d%t�����Eh�B�I�`D�	s#G׋8Fy�-�+q��B�=�2�ӧa��jSn!:�
��B�	�o#���L/|q0�i".֗`xB�I�,Z�%+TI�3$�=���Ӛ%�<B�	<\��!�JD�A+�8��^�UB��,���1��^�J1��.��C䉋s��r� G�z�=x���,I^B�I#!���'N��1��L#�_�C�	�-X�9RS#Z4\'�<8��-QB�ɓ,�\@f�2�Vy��آz�\B�	,!/|�K���v�������>cl�C�I�:�Bi#�o@ $��ݫ�o�;v��C䉰3��PZ�F�7(��)0!�V>ijC�	>#�d\�a�0<m��#���^@C�ɤ+��i��X�J��ĭ��\�:C�3�<I��C�j���6�̃V9:C�I� T�0�)�S�b�	cb��R�C�ɄW�\Zt��&�`c�i�B�ɤF����զ*��q���.B�C䉖Z;^P8#�����w\� ��C�	�[�*��!I�N�L�k�T�~�8B�I� �)R����y]b5�Æ8�,B䉯i#V��W�H�'���7f'c�C�	�xt����+�z�#G%��W�B�)� f�!g�Q�K�$�� ʁ'X`)f"O���pꇻ���XG�1B��a��"Oڨ��.�<z�q����5N�Q�"O���JQ*"���y�
�S�8��"O�3��i?�@3q*0Z�f�ۢ"O4�rLM�=����/ )���"O(2v���|LJM���э`F�M"O m!%G�y��LQGע =��F"O�R��K?��0Ss蝍Kr�8�"O���� �j�%������$"O��3#7��9�Q�8F���"O̸�5�^ZcVX+���(K��"O��(�C&"V(� D��Za��[�"O�b��'9*�{5��49*�Lɰ"OHHa�h�;;Hx)��:2!Ya"Oz����#����t��\����"O��fF�4��s�G,آ���"O���s�,)s����@�/j�"O�PB���R�,p�b�4`G��G"O�A�FI�}�t0�� �=>A��"O6�{�ǡO4���I&$7���Q"O�%����]Z0Ѹ����28X��Q"O��;ЇF�KQ�@�ٝg�J���"OLC��Y�n�.d��'=qN�c�"O�L�0U�Ep=R��_�*U�th�"Of5I"c�t}�a���I�ne��$"O� 2ЄœF����ы'XN5�"Op�p�j�;_���Tm�6s=
 ��"O�\���ҝ+�Fp��ڂ;+���'"ORb�e�xY��2��,9TYCG"Of�+$h�,tk�)��O=7� ��"O�-;׌жY�$xJ��U�D��h�"O�]�	�� D,��2CşC�@i�ȓ!�X|�Y�|)��+�@���/��tQe�K�`�B��G���N�ȓ-�a��*TPmN%�q���BΩ���l ��A�nl�((ԇ^"�Մ�B�͠�ڇv�z@�	�.�����g�&���}u���R�͚A��ņȓv!6%��Z�6��6��s���ȓ'@)0�ǚ�_+Jyb�	���ȓ��A�C��6:�-r�L�4m�t���9�Z�r&�i���Ϫ#�z�ȓg}
K�K�F�4�rb#Xx����VO �x7���M�wh�AQ�Ah�'E��t�ͿQ�y��ᔅ9הr�'�qD�[��y0�d��2�L	s�'��MC��L'jqh#�ѐ*W�	�'^��J�m���]ڢ��)-HK�'36qXc�G�7���b��?$s<���'H���p+����Q���!�ޑ�y�ľ]\M�G\ h�^Pfا�y��:ob���Wl�T6����Ȇ�y"KB�B�|�	���-WP���6���yr��<����A? 2D�h �y2m��`NXRe	��vO$�3�# ��y�JNjb(�h�L�?I ��E��y"+H)s�Hb DS3�\2��<�y��/x�6Y�(ˤ-�N�*�,#�y�A��J*���c�Ȓ+��ቆEѿ�y¡09�i˗#�g����,[��y� �a􆈠���(g����Ȃ��y�I�"�]��E��f�:h�%gR�yrÊ,{�:yY�囕'�^ ��cނ�y
� �dJ�����(�I�n�4!�"O^�x�͂w��YbV�ҁqu����"O���cYu�N�Q
Wo�,H�"O����-��E���q�#�(Þ�"Od��&݄yg�t2�"݁K���"Oj|��R;`���l��[4��
T"O�� s"�������@	+L$l[�"O�eR⊗0"���їhI�R���y�"OF8dg[(�";��*{@ �"O19�'��:Xsӄ�jz�P"O����l��m�dP����S�Ie"O�L�Pم)˶��`ٶE8θ �"O�Iw��[����Uϋ�,�tZ�"O����bɻ@s�ђ+г � uy�"O�)����B�(�A*��I�<1T��� �l����y���1�C�<�w�D��(p�D�G�~���M�~�<���ەI�X)�R˄�"�"�`��Nw�<��b�<I2r�)�LV(:JF��Rh�<��'�U�r!�4%�*~����i�<Qc`��@����S��#?�
6�}�<a閼^� @+&����\�Iv�<���Z6`�Nܱ� �x^��aMT{�<�炍+���k���s�h�A��x�<�"�)(�����$@%/�P���w�<�b��9H��!q��8d<�	�nZu�<ِ��Xdn��tj/E/��ağn�<q�?udyr�A��j��#�Nm�<�O
0n^
[R�R{�'Fj�<1�E^�]���YP�QfV!�ǂk�<��k��t�lQ���!m���g�<��&�U�ɂIZg���^f�<1��_MJ���~<�(���VL�<!�'O�����i�)�|$+�GZs�<�F��%ݜ��ϼ\K�1�C�^q�<�g	̙G��J3>����@	��y�G��	��$�5��H����K���y"��"*����Z�@xZ��ШD��y��	��Ԡ�O^>�LY��M��yRf�
�:�)��	`�)�!�y�(3Ĕ��d� ZI�����y҅})iC
�x7�����}�j��ȓI�\�隩 \��{��_)��U�ȓ3� �ЇI�F�LA	U�9q̸��i�H�E���;缬Qt�82Td��ȓ
�`��)I:\� ��AՉM�U�ȓ�Z|�g
^I��`�5 ��a�4 ��Q���t*�x��M1!�@�
_�ȓO%��+�f�%?S�u���!J�؇ȓn�|x���&f� ��#Y�<:}�ȓ3�<�	v#WJ���`a^�-�f(��;��� !��pw��YmU$r5H��ȓ����l�d��x�����X��m��k�$�2a��QYw*��BY��v%Ve�EB)A<z	����L^X!��H�4|�U��9a��M���@#y��D�ȓWJv9�ҥ�_�]������Y�ȓD!"����Xr�9�!�( �ȓ(�b�Y�뒪%��őT�H�aVh�ȓ>v8A{���3<!�!K�l��хȓ7����g��*�E��'��p�ȓt0& ��|����#HV���1���Q���x��M"~bp ��#�nXⵌ܃8N&�	W� ����S�? aa��1R�؉���O�C�"O�<+����yzZ�HmW��)�"O�E��/�� Ҫ�����!�C"O*�Kg�_�~�إ�KΪ��"O�M��D�v�x!�N��9�"O�}PqH	��tĘ���S��<("O�-B� ��q�P�=8|��A"Or�Xq`�.g-�ar�+Ө))9�"O�T"���M�`��jV�S
�L�T"O���a��mW��hA� x`�	�'�j|��ț��� 	G9���`�'����$I2rA<�+�ǚ(dly�'�,YG�X�z��9! 'tZhC�'�䵂!-J9����\E��
�'T�ݙuK��1'�=H "X%[D�D�
�'v^�h3��2m�4URTZLy�
�'�pM+�œ�H�$�lZ�LZ@��Hɂ��`�*��q�FjQ�/j�0�ȓ]�F�G�*� ��t�#\Xlԅ�8U��A�-�X�@���"R�$���i��)��Pn@�h��Í��b��ȓa�XI��^=F�X!��E�F��ȓD��)����Q���`��[-6��YD�����L�~@b4`A�Z=�ȓ0f���I�v`z'��>�R؇�O$5����'3t��4%K�o��ȓV���;�N�(A��1��R�P��ȓ/Nr��ԦхL���WG^�( J���l+Bu��ɮ?�����j���QD(�Go�JJ2P�0Aۋ�v�ȓLA�9!����l�����ă{ANL��9���(܁f�����`�)&�P�ȓ6.2!{�ى!L��Q�G�$�ȓxwb!����6
p�@�(?V}��?�F�x��K��^��c�%k�|�ȓ$%�<��Z"�<�7DV�*d��=MY��X?e����v�����8#p�v�+r�R��͛�������($�&��4muh�q�e��G%D�px�&��H�x�j0���B�Lmi��?D�4h���1c��		��г7�$�§9D�ty�I��XB����&�� �'7D�T�m��L�@�Y��>6�2L�T�)D��1��Q�B��9A�J�
sR�$D����V�N�8R�F�V_�}�v�%D��āN7{�V�
�t��Ίq !�zy��k*N�Hs���5~!�×3S�=�E �4=��TXD���:`!�C�Z�8��!t��,kaA>G!�D�"f����2D��q��Z��W�@!��)w���EBF�"W�1���#9!��N�~���pM�Q��#�Kp�!�dp�fu�p�N�t�4e��!�$��T��ت�bZ�_,�Tk`��Oo!�$�0z�b��B��A/����ĥ>�!�$���٢3�ƵGu����:�!�D_I�8�b�Kt6DSBU<!!�U�H��4����q0��'��!�(�D���)�'V�������!��{��e3��>"k���GK��!��j��sᮛ���q榈��!��?"�� �q�׬R�
Y��.�!��*6��vK�6��� Bkc�!�ķhް��� ]?ܚ�Ij+!�� ~��%B��..��j����(��@"O���[�* �Z�	D���c"O��@�%��c��B�*S"y&�5��"O�@��9X���#ɵ>,��c�"O����\4�P�A���3���"O��Pr�[�J�&IC��:>�p���"O|h{c�\�h��rנ�7+��qkv"OD�#��?e�B<��
Ð[��l�"O��Rg9s5�<�s,� �|���"O�s�	=a�YQ�Sf�$M b"O�䂲Ni,�c��u���"O�)�l4/,˂��?e���%"OZۤC�*��Q2�MOXIW"O��1��C����s�I����&"O����C�r�*�sv(�yڲ1��"O�����Z�#�1�FB#2�^5�"Oց��E�h��T&�)�lQ�w"O�	j��ŷ3X�{�FZ=���U"O(,bo[���N+l[�X�WJ�=}q!�ӥ>	�I<6V������n�!�$ŀ=,4�wE��T�Y�(H.�!�D�3M��HgH�V�0�Y��N6i�!�74�B鉶�\�Py��H�_u�!�@�	l2e�	ג1�ĳ"	�o!�D
��2�C��S5tdp�4'�8?�!��"#����ܮ�\�S��o�!��Ʋ=D�|h��T*=� �(7D�ar!�~�-+t��ق�Jde�+U!�-Nq���ā^7K<�j,J
�'���A"Z���WI�	z�8�y�'b���0w�=�"�F�jnxe��'K&
�&�93Bm*^�8ݪ�'�`�C�P� smB�\˪\��'�p���V�~����]�&s��)�'��+���xՊ�<�8��'4�K��$?C"����Z�\} ���'Q�#����Xb���T��x�
�'.00@d�x�B� �?2��
�'W( �ǩE#'*��kbk�DS2�9�'�;��HL0�Bw���>��y��'��(�͌1]�L(`�C�=�nP��'�q���/��*���d0l �'�� ���8���%.�
Ybt��'j|l��C*<�$�S�J;X�$���'�6�bB�t#��I��8b:J=	�'�  �.%DUD����8*��4k�'����f�u(Q����m9�!��'��[�J�H��i`�A�l�*���'D�!�B �T���	BJ��v�(|��':�ٰ�Ύ�(�Fѵt��Q	�'��a"�(�c� 1J�H� B�~E��'R`�HE�ΑvxP����"��Q�']*%�h�0f�j�J���;~� E3	�'0�,��Ka@:���o�f�!�'����,w�l!+���2v�2\��'[�q�% J�L�jԂ��|����'J���Ԏ�K�f�8��N�m����'���C-�/�c0��^V���'�,���ߊn��Ġ�G�QxF�R�'phA���Bؠ�ŇC>~�!�'��=�4���
�o��;� �"�':vTk5Oz��� F���1���k�'����� Y�VN�y
�;'�ld��'
\`�����$�am���Ո��� PU�%���^ �e#���F$��y2"O����NA"	��1�g�HTZ���"OX�ط�6+����t�Y�[�\��"O�p�Q��B� 
�V
�L#r"O�0�Vp�L�k���
u���q"O�l��	L�}"dp��o�I�^x�g"O����G�6�@�T@��k��3C"O�|a�E��XzNE��.
�bab`"O�eS�ݕr��[�JM�:�����"O��å���'�tU���=b�X0Sp"O2��ݖ)�ĭX +��O�P,r"O�����dZ�Ăwj�<T㰘��"O^Tp)�%4������*��j�"O,x�d��?�<�@3�@�F��IP"O�$�ʃ'_�I���)fy:S"O�Z!��`Ifx ��;k+����"ON{hF�I$�A[�,7�dJa"O�,�W:�\�РƜCK�YBF"Ot����F	�.�2�O-G��!�"OTi��ŅhR@��҂qR�1"Ol`��	i%K�&��W �9C"O�\����A����%�_���A"O�q�D,(8���XqKƇW����"O�%�n�1��C�IS)���P�"O�j�����<kP(ک/�| xc"O��E��|;N-q�N �!@r"O܄��,�����
±x�"O$ٻ��
�)�M� �[vd��"OԸhc�!/�@��� 'e/�]�2"O����ߦ[��'�V�[�"O�3v�&z���7��:�h,�&"O:!���E���N�n�pt/�!�䓇_�L�R��K��7�Ɏf>!�D�HV�Z�H��@��	{�N1!�$O�Sw�}�v)�:UbV9k�-J%�!��ޔY�0��e��d^�U{���;I�!��]~>x����6k���k\�	!�!g:�sԣ��H�L�Rǜ	8!�d�H�� p�N�>��TE�,@q!��¬{���`���3����Y%!��_�W�"$�\���dӗgW!�D�4JrQ��aY�<��i�J7qr!�dW8}�@5i�K�$��:�ȱ�!�$D�Z�򰲡��'80ZdAu�ʋ\6!��v$�1b�gɛ[�X"�
^!��p�@�@�%�+�M���'�!��Y�;Ѡ�P��*6���h�!����E,�	]�(�P'3)!��·7r�D�tH�YA���p��[@!��G� 调c�y6
�BT�X<]*!�p��J�LϲO�A2҉��.�!�Ɩ��ׂX�:ƈ�Ńq!��Re�mr�M��m-�8�mƂA�!�Ā2X�4Ai4(JtQ�0OΏi;!�D�5U������@�D�Y̇1�!�D3L��Y� � �N�DD#�N�$W!�dS�j�`� �I��L����ʏu!�Ğ�n�x�#V@��i�_p���*O���G��5c���V��/E���'��,��cK�$�j�jV�P�<�֝Y�'�`�"FDBG����ɀ ^F:	�'7�1�s`�::@D�\xr:	*�'�̌����!���1Ԁ�y N$p�'ix����� �D@�<��:��� .$+'�tw�e��DvbV���"O� �@(LdBZ�Pc�F�]��"O��A,�-E�\� �� 	BB"O����덁0�8��@NHuV���"O8Ŋ#��P����OA�u�0s"OV�Kc  �R��Q/Dg��4"O��T��`�J���F�K��U"O� �j֘aD$�����U����"ON\�����<(�uAJ�,d�G"O֬{�֗�
��fJ�{f>x��"O��Bt++YbzDTD�
0[�(��"O<��WK��Qzu+��Sm9��'���t�\�^m؄2%�6[Uր��'�NĲ���pt2"�_A�D��';��Q&kZ�7��ˁE�J���'�X�CC7/q����
�p����	�'�$�`R�Q�>��i
3OfY^��'5�5hU	�[´Q�B� 0ZF���'��0c&*Z�P�Va��'��W}"��'Ԁ�r�NI$2��y"�`�D'ƅh�':�����אL�h,��B�<��#�m�<���߷��{�E��P�6�釦h�<a�k� tc8��ua�.- ���@k�<��A�o��X1D�(U����
\h�< ꏔ�J@8��\/��٢Jf�<��3�J�9R���~Y��ȗd�<Q OT���"!�ފG�`�Y�(x�<�W%U�!mJ��O���,�C�\]�<Yf�2z�P��fM��)	|��K�p�<�'/96p6�p��U�Rd{ʒq�<�3�̋?D��l)��aV��l�<�EA�@��l���O�=�J�Z��^�<�$o��Ċ�e��Hr*�2�BW�<��EJ2=��yd�ˊWe,�xŭ�S�<IV�&�Ls��Ձ�ؐ0�
�N�<�V��(}���>hB�pE�CM�<i1
�[@6]Ar�\,��Y��d�<1�+J�:s&����1��1�Wv�<�%'Ht̂"�\.D8�:��o�<��i�)QQ�=B�e�$==xH�a��k�<��@�&Dupq�@K�g�,�%Ug�<�5	�\��ѷ�] n2�b�]a�<�+:^�:!�� �<��L����v�<���	�Z���t���}�p@Z��B�I3P�7i �D�f訤�0�"C�	�Z��(�Ux1($�Tm]W��B�Ɏ,r��h�		x�Ѓ�Z��B�	"��!�f�#<��y��lʹڬB�ɐ5���;WGP���9YA'HcHC�II�� �D	����@Ś&��B��p���K3��C��mPq�BT�B�IL����vK֣�=*W-E�WƘB�ɴn����P�դ�\2�݈d~B��d�t٢f	%9Z��� �BB��M��X�c���,�{�Ż2Z<B�I$4�^���kZ�!�
!2�D�{�4B�	�F}4�84![�ke�RF�GqB�	1Z� ��NV�M�)�r-=�B䉸��#�F;�	��FB+5M�C䉏gl^@�"#�<o`��ih�?�B�I�rF�([@inQ���US��B��^���c��{�~I#Q�*�B�I9`:T�㨍� ٙ��R2t:4B䉞N�, �w�� '^ ��nSB�)� j0�e+��-J!jD�=	���"O��(a�\�$֨��ǜ"&���2�"O�-ىj��5�&
 h_d1�"O���eM�(O����Ɩ,qRp��U"O�P�O�~������:W&l�s�"O�=��.�x��C�cݪX j0P"O"�b
�5����v�B"4̀2"O��yBM�~o.����&�X�U"O�Q�bM�-4�Ri��պ;���"O.93Ê�,T��Hp�)E��[�"O�{։G�n� d�Ȩ%��b�"O°��h�%؊�j��26>ͪ&"O�K���%�f�JR*	�~T��"O~}iV�
~���A��Ը�H��"O2�+떐A���j�6"ֶ�{�"O����F�j'�fjR:�K5"OV=!%�̰-�d�熑�d�\�A"OZ�
�i�r<qG%�6@�T�"O�����=	�1���p"�x�"Ǫ�HߜZ~t�aa������"O�xڲ�ڢ3��W��`���	��ybH	7x"̻��S*��(�t#�-�y�BSLe�;e�ׇ~r*|R����ybg��P�V)���K�T$�X��y�G P8�xɂ�P&-��aBCK���yҤ�l�P�B�S�5��eV��y�τl�
D��
�7K􌤃�U�y�gS��*$AV�H4s��p3kĩ�yb�('I�8O _�6��"\��yB�M'CH��&D�28���Q��yH�z��A�vE�t�`
�nD�yR�T(t�P��E�܉#K�(I1�ǹ�y�b�4o�(��ҥP*2��z���;�y��K�+�b�CD$�?,ܺ�`"����yB�	5�
�cVBߪC�<��OD��yb%��,�4���`���a�C$�yb�áx|T]z!�� Q�|��^��y�#ѲA�$}�1����P`
��<�y#F�YZ(e���G�\�f��%��=�y"�*Kz*���ȁM�A�4�W�y�],\���T�֔@D�4'��yO���,���?g��C�E��yrʖ�YcP�;�ռ
0tI�B�^�y�`��9-��s�FT8	+&9���@�y�+�<z��D�1�2N�.axa�A>�y҂�̪��@�E��y� �N;�y��[�Jo8������<���5�y�/M�꒕��E�Q��MPw���y���o��a���ZC�����T��y�����:U��lҿ:��cჩ�y"�U�6a�rF�A,^��S�Y�<aҁG�x�Ȝ�f֘{�����F�<u�ї^��R^�x���ס�@�<q�$C�j�d)�JZ3��ő�UT�<�s�� 1��$�ь,�81���D�<�U��+ �BE�g�B�.��b� �D�<����g=`(�k�>m�ejF�<�C�*e��`S���*�Z�j�M�<�C��>�E0��\T�
L�G�Au�<q$C�.L�H�Y�#	�.V���
Y�<�`J�*�qc�H#������TJ�<�&e�Bg�@#k�En���$��<I���)#�ڄ�P!�n�ѳ"����m�%�u�Bz
d�z$
��i~����S�? �Lr@�*q�:��"�݇K�(��"O��,=}슥�Ǌ�x�E�"O~����T�~sdA`��L�"���G"O^)Y��,����v�A�I��"P"Oh\�JߖS>,��Չ7��a`"O�H��L�7B`�2T��0� (z"OuI�m<L��a�+�
0�5"O���5�1�r�@�X�����W"O�a(��C7�����+s��)"Oe)߷"�0J��x�� "O�<��>a�쩑�C�p�A"Oĝ&�����(�"ɏ����E"O�1�b�,z����!���}o�i��S�R�s#�FbŞ%��jJ�?����ȓ\�eJ�1k]�t@"!+M��ȓA��4���lO@�!PC��uQ�X�ȓqo&��PM!���c��I�(��b�b5�%�,9�ڽj���_:���F�ZUJ�F�s��2�� N^Fц�P\�Ÿ�OLn�A*�L�J�	��al2MA�ѪJ���E�:`8긄ȓE�
�ig���ZE�'��9>n ��ȓZ)�i;'"�2��Z,қG$�l���%i'�����'A.A�Ve�ȓR�m{%�^K�Y ��+	��H�ȓw���:g���\�Wl_�M5��ȓU�,!��E�4�TH��b�f����ȓO:1�ǐDЍq2.�������{�������J\$�/��K�(U�ȓh����m�%:m�c
Z�]����=h�$��+aЁA��,vL���G�6Ĩ 'T+h.��9���1.�����l�3C��>;��(��k�"o;F<�ȓ0��A�k�}A�y�oD�vպ��ȓaI0(���N���sEL� D�(�ȓU߄P�@AG�m.,u+��?<ո���T��9��΁5����O˹��ȓW��X� ���B�
ֱNgH]��{�0�{�;]L.�A���7r�ń���C�c^L&�H8`��^�(ՆȓQ%�m�P���T�l��@��ȓs%X�@��,wZqQP�����ȓ}�������!���
"��;DNՅȓnN���s�Q�..�d�ܶ3�<��c�I��L�	!j ��'��8�ȓ-�}8��T��N\{��߀S*¹��h�����j�"7�#�M��dm���1� ET�T4�A#߯_QP\�ȓ a-��j�@��S�JP����ȓH�v]K��MBv�-B�
�${�ʓh�2Ǥ�3b��=��*�Hm�B�I9j��)P#J'R�6p�`�D�R2�B�I����e�*]�4�P��ū��B䉧3��Є�3Tf ����B~c�C�I 
��q����	���8�-�w��B�	��@�r.�'�����O�<��B�ɿwu�|:@mM�7����I�I�B�ɭo
�l����+��l���Ê��B�	?��(Å�٫b
��ht(C�3D�B�ɣ����-܅kZ� 6,B�-#�C䉒mA�t���R�#n6�&�2>�C䉪K2�L3�D+P7�91��<<C�I�S�J�9���/9I�9q��
D�C�I�t�v�1��+?B�)�_?_�B�)� ��i6B�aѰx��΄���"O��{� U�w���;ы����"O�d�Q[<I	���7�.yi%"O����G7: B�k���)d�6 �V��5LO���BA(ǔ!�c��"�!N�<FW�S�@�HQ�s���2��K�<1@��_�h �шQ�#�z����]K�<���	g4�P횠Z��e�S�G�<!b䊬j���"#�
�E��Xj�DMX�<A��FFB��m+�,"��	M�<�e^�R��]8VB%/=Rܩ���G�<1���;G�\�%�Z 3��u��
�C�<Y���.~!����#�N�")���C�<�$i�"NF��5)�u�V�B�<��N�h7>A��L������Pw�<��E���@`���75N�)���g�<�u���m3 =�`����ƄS��_�<Q�M� w.QH'�ΚA��sS��Z�<��-N	������9K���@NM_�<�D�:
ǆ����\0ZL��[�<QcE�!�~ᙔ���v*��6�PX�<i�o��O��R^�0�T�����\�<���+QE,���ꙋ\In<2�c�<�1#<�æjB$T�)�gu�<�WC��]wҁ(E���P�"�"ɝJ�<�ai/P�J�áiي_b���G�D�<a!/\&x��RN�Ȟ�P�
D�<��bA!_F3V��=�BЩ�U�<	2�B!żx�@3�n�f+�h�<�%�S�\��ya�T-S킥�
Le�<��	a n9�m�&[�̤�a�_�<�3��$/�|۷�S�o�C�p�<������5��*�^� A�^t�<�4EKIb��(rT�B�\�GB�q�<�V!�8 ]�%:S�B�*�pcg�j�<)�tڀ�R�݇<�D�Rulh�<����@��A7om�ɻF�W��yR��>Ŝ�b4�� GM"�A��O?�yrI^q]L��a�C�;�|�fS$�y����0/ȘiY�ʅ�$,�|LE��k���	2FR� H�@a&��8�� �daA�c 6v��r���4�Ňȓ�	{"EN��Hɟ>�p8��J������Ԍ|G(��%^�qPv���}���f�]-G:q�A:-s�!�� �8�r���4"hpH�f���`'������(�B�	�HigA/qk���ȓ��ȗ��('��Ǖ<�d̈́ȓ14�U�\Ze���V�����,+(����d���@���6�0��ȓ��@S�O�0Ѳ���&B��ȇ�/xD��w�S�b��h�"¤nN���oc,�0˜�iu��'�^EX��Jq|�P�H@�8N�	ԦC;`w��ȓ]$����Ļ9;
����
d��!��3-�P`� 1�h�e$�4L\�ȓu��3a/��$��j#�D!S�@Q�ȓ�L���7'�Ҍ"sQ�	]����?���� �P5@U$E����ȓ.�����Ys8��U䞋YAV(�ȓ^+�!���0UX������	����ȓmtX�s6i�T�8�j��H[Q0���Z6꩛���h�X���B��p��(Ò��Ś�"@����q����S�? �y�G.O�	bP8�4�גb���"O���D�&@� wm�)W�$"OQ;a���~�U��EZ;Exv��"Or�3 �Ty2�dƷLM��b�"Oh�kg��	4�"�
7� ����"O�]���ɺB�6��w �$t�� �yR����Pːe�����)�y2l~Nv�
�LN 1���$�܆�y��D8rh^���n(�vX Dn�<�yR@MP��G錡��m)"hۃ�yҁD 7�&�pdB'�<0
�dS��y⚞D�l�%զ$s�A	��L(�yR�ְ5~jL1ŀ�L��u��� �y���0o�QsG�]�GP|�)(\��y�/6vX �V�P&O����A��y�&��h&�D�!k�5�r���!�yB��Vv�R��A4�@��t���yr�Hu�H(1O�b��;�m���y�X�)ŪA��*ͽ|� �
�HE�yr!�gA��Ee�")I�E�u���y�n�Hxz����%,Kv-��b[*�y�i]����+��ڱj,�.�~9�ȓ&����1؜cĸ�DGY�fg�e��@�D�ʦR�r]���!� x����(_0�+���dN.��eI�_���ȓ���XB�P�Y�x��π�K�����]V�1Q�b1T��A3Ԅ� `E�Y�ȓ5~4�f�BȮ۶	P1;��8�ȓXN�X9a��F֍:b�
,Y󴉄�e����>�᳅	�+���ȓEvm��#ʄc�s��(cD���ȓ/rx@R�a�)$��l��E({-X|���ژ�b�=228�韭G�D���y"��.=��	s��'yȜ̆ȓ���y��]4"E��J�&��ed��ȓzO\���
	j�>eaG.��`o�8��Q�t݉�#f��i��]P�х�#|��d�!~����
�S\�ȓC��2g-��fJ^h�)�\�(ц�2%~���L��`$Z��@��谆�;���.F�0��;CY�#�]�ȓd�H�ö́O����υ�3[J܄ȓ@#���!�F� �g��0�V0�ȓ}�P��KT;!�TP��)2��u��\A���T&k��S�g	+>@�ȓ��`��(\̢��cF�U*B�ȓ����B�&-��# G^�wh��Z��c�@�\�
勂.F�
�fh�ȓAęH��Z9<�|D�6�" ����ȓ.v�a��'�2��"P��s6E�ȓ4P�����=�D�T�RK����� `b�=`���G�dzB剒N�#���d�n:0I�߬C�	~4��Ď�.h]0�i�ㆢe+�C䉌4�ؘ����h(�X�0A�g`C��2ަ �vFW�,ʈI��1g �C�IJ�ĸ���	2��x+�C�7%vB�I9J@ cK�,�Vm8v��&z�fB�ɡX\��"��*Q2���"�bB�	�2x5��-Y{�|��DN?o]|C�	�j�hR_�i[ʌ�$���Q�JC��Z>΀IC�.����N*�C�	}�̬�!(ÃJ��2E�2�B䉕0S�m@��!S=����$pr�B�)� ���@�V�aT�0�΋!E��]�4"O�M! ��i2��sŨ^>���"O(93���a)�a#�hϣ`� ]05"O8Mj���,k���E��X� D"O0�R��#:D�0ud�WD�da�"O&��'�͇%�)H��_()nj�"Ot�@�/�1�N8�!�79��7"O���C揖�,�Q�і	��@�"O�D2e��.f�1��;h��}�"O�X E�P����c���&��D�6"O@I���SK�>x���_=U��9�"O�e�Eh?2�k4����X�"O �����Ke��)be��
�"Ol�P��W�/�tM{�툑1�V��"O(hs��1q�q��kʊ|e"O�qhr�ϒQ�$��KX*�b=�"O�<�֣��$���iPL	�Z	�""O
��r�L���0�i�a
��r"Ol8Yd9J��`H��(��u"O��۔#Y.t�RȢ���-C8<yS"Oa��Y�N@P���"J�.T���"O�]��j��f�@��Sf8���"O���'`�p��q��+*�%"OdM���0/�Z2I�Gʼ��"O����Ȉ6�p,�&ޯ<�Xk�"O���՗;D��@s��9��Y�"O�	�Ȇ�6�`F�b��W"OHY�� �lΚԩ �\.:���H"OY��`ҿE=�-:%��-0�8�#"O2-�P9��MiGaώet���"ON
t��7Ut�"r P�?l���p"Ob�J6�U.d�Аsn�!0n�4"O�`(A�R���!��V�f!"Q�%"O"A˳�Փ�J<��l�'OT�s#"O���w
;"�=c-ɫ�����"O�@�,[| dB�U.P�� �"O]!t��B!�_x`�"j!�䍻#;��iB�/Sr S��.1e!�dT�AG�u`7l��-A�y��D�S!�$8d- `Ad�^�Pf���Ԋ4n!�D��m��b�K܈pS�<����}y!�d̀ ��d� � �S8F��i�&}c!򄚠A����ޞ�҇�!򤐫K�P��P$@�4:�'F�-!�d�Pa�Jc!������K(N�!�DW't���ic��k�9��ƌ�8�!�D��R��fLEX��ˑ�՘$+!���[�Ȥ�$�)�ȑ%�8z!���3�P+�c̸ ���A0���!�B"�Lh��.�;6� ��c�)s!�䟍+А����J�[�-h!�dʉ5����� �>��0�ԫ�9M!�$
�(�����h` �K[w.!��\��h��kɌz~؜�꒣9!!��X?]u`� �v��ДC�q�!�M$k��@��*�
�|)e���!�đ�|�����Z:(ǂ��(Ϯ[!�$:wC���A���T�;R�@L!�Ē�b2����B�4U�A�,�!��5l����w���M������@ws!�$Lz���䠉�_�P�@��eR!�Ĕ 72ne�6`ڏ2WX����)=!򄒗t��J���%7VeSצ�[V!�d֌m�"yv$A���`�RJ!�� �D2u`Z�<`LY���A]���'"O�|�r��*8��� OE-M4�}�V"O����L'�*�S�#�<d��q�"O�+ ��H��4�q�I1��`*E"O�h��ËNg��g�ѐ5��� "O�}��ٙC��)d�Y�]~���"O܀z!�Y.W�J�HvB[�c]��"O����煊'�4]�Ł�&ΘZ�"O��9GAц�b,z�@�!%�X�"O����BQ&&�|�q��fe�	ˀ"Oҕ�@ �T�; ǁrJb���"O��Æ� J؂���΍;�h�f"OU� �Ol�ը2�ށB5���"O���g��Zq�xȄeL.|N��aS"O��#Z^t�ā*_��!�"O��B����D�&�*r�$>rH�"O,-Z ��u�`��aV#x��"OJL�רO
R���B@I�@�\X��"O�H;E����b�Z��l#�"O�IsԀW�hO8SD-���P��"O9K���6Y�Qa!m�w��yX�"OvXZ����Br��;+�hH� "OX 02�N1A��fٖ( �zS"O
�s��C.#�ihu� %P�a�"O^�rGN1���Z���O�r�"O�թ҅R*G��Y#U�E���Ĺ"�!�$F�f���mw���w]�!��<�%ił�69��`ϨS�!�)Ffֽ1 �C�����3Kz!����yQcV��mC ��!�$�(6�>��0*Z�.�:Xb���yk!��(R�e)RN���Ô�� �!�dW1*2\ñ��4 @��w�]�O�!��T�N%���%�C�k���R(�&�!��I��(Pa��9�rYARfύAv!���5x �h��_!>׊�Q���-�!�,Z���M�$hְ|�"o��n�!�DLC��ʵ煠"��l�����!�D�F2T��!f�*ª�Y��җ7�!�$<��H����4�$I��M՘c.!��2�xuJJ9\�x��B�A8!�Z�M��آP@	)zq�@�U�R!�̌<��x���'(��C�ݑ~"!� �F7�"��? ����N!�$O
R�~�ؗ�OI�+v!�d�4-���sM@�DD�
E�M#�!�$�/���0"� <ڐ�pJ�;�!�X�kX�-�'!Z]d���C����!�$	��Y�i,���U��=�!��\�n�F�c�I^�On����h���!�$G����%�IQ�J�(�8�!��6:���7��/*�ł��J�%�!��^����Pb��&m���jZ�!��0{ƺ�@6N�Skt����ߒs�!�$ۆqZt`��a�%q�e��Ė1|!�ͼyZ��f eiD�2���vs!��O�>5��,�wI��""�;l!�D� <P���.��!V ε[�!��=%��e�ȗI��8���G�!�ŀ� �y�Lr��0��N�#Y!��/��,@��S4K���hU�>e=!�d��#��UQ fǎ>+�Z����!��(ȍ�3���S爊�c�!�N:�.�s��
[��`h���^�!�� �XK�Lާ[�,L���R�F�A"O|Y7Ϊuќ �eHZc�Z� 7"O�Y@5�;3�, ���(�Ѳc"Ol�b�Yc)셃s�q�lτq�<ٰ��.X~��y�ǂ�G��l3#��W�<pd˗6�fXU�\���Q�gJV�<��N
i��l:�"ƥ��T�*\O�<I`E�&hi�@��$A�F@���q�TO�<���I�	�e�",�U���Q�<����?�qR���uaAK�<��I�9-���W�� ��gG�<)d>t�ay�EZUph3C�m�<�ց΢ǦM� �*J���BSP�<9W��>8�0�E�����%�WJ�<���Ƽ!� �X�ݷI�`e
�)a�<���2k�傣gK�Nj�Y'At�<�%��62(3aK��$���eXe�<����@?�HR����?�>Љ��a�<��ם~/��r'!@(�%�f��]�<��L������)Q�f�##Vd�<���	��9(P�W�,��P mb�<���B+�Zk��R��"�:Ji�<I�\'�T��v�
l+6\��b�<��[v�	@�u�@m3�TZ�<!WZ6����⛀d��t����W�<����]�j�9���vhA@�l�g�<�����A2��ۣ�R#X� X@�f�<�ѡ�=S��Bg��{=�+UOd�<�`�'M���W+�>4n"Q#S	Pg�<�RN�yw �$
��*��g�H�<��ɬ�L�����0:.�Ae��E�<17�M?Yl��hA�1Qq�����L�<)3Ӑ��9��M��S`"��0��_�<�"�3GU�yG���0T@�,�Z�<��H	�<�")KB���m#��LS�<���);F40v�z���R���Z�<��mA8V����X8HD�IX�<y��'���[��܅*�"����j�<a�O�X�����
�*h���Éd�<�C��Z��t�B�J�T�*y���_�<!c��{�V!0u$ݔ`�����B�[�<��n�=\���/�Ő�a�Y�<�BK�J�&�#���	{nHݚG
V�<���:3'�j����u2U{��M�<qs�T����q��V0f���c�E�<�A��[�2×�ԐZC��r�&�B�<Y��2h�Ĳ�`�TPr0��d�<�#�*[�10Y$t�҅bA� b�<��N�`�u�Ɍ#	ԑ��\c�<1@J�d�20h�m�y�ѫ�g�C�<�h�8��kj�"lGa�$�:D���$��`]� ��	����#D�`�Ŭ:L� |ŭ��ͺ��#D���rDCaC�d�+g.��z#�%D�@rgR,OlrB�Lʬ�Y17D�<p�J�-�̩��T�7�����I3D�lp3��#��q��R9XX�)��E-D���f����uyQnO�ZD��p� !D�4���O3T
�͊ Ŏ$���r��>D�4afӸ9�V�:���1pT�$�>D�H3C���[9gh96T���=D�l*5��7>���j�iI�^�Fp8��8���<�Ol\�q�O8Z�������֥H
�'~# �<&��Z��?�F8���� ($j�׆i����&�G$	)0�"O6u�a/��Rz*08��;��,�P�D&�Ş=
l���4Ri~���Z 4�ȓ7��dqc��<$@@�	���<<�ȓ4�Ja(.gkj	HS�W�n����&�z Y�[�9� ж����9��X����T�/�r���[a��d�������Y�X�t��9�<q���))e�\;n"D�`3�
W2PC6L��I\�P§�%D�P����Z@��M�"����$D����l�?<�B�r�]�g3L�ⅆ?D�l�EQ�*�<2��� ^�=J�i=D�䉀N>=<,��tgW�²�-D��cՋ�-՚u�FD�!�DH���)D���g�_ W�d| �<��`i)D����7I-Z�x&�%Va��f�3D���դJh{����(7���s�3D���Hҙ4�d�lm���3�0D�(�
��pD���I�oK�"�B䉁�V`:���f�v8y�	�;^C�I*k�AVT%�|E���j���d=}b@߯,ZPD���U�I�'�-�y\:
V�h�D�I�2�a/�=�HO�=�O��fE�(|d�1���1�y���XHH`�#��9;��a@����Py��9b�Q�5"#HfA�ׇ�^�<�C΃�|��XG�X�F.\��gOP~��'xPىDkE<..J�	C��n`�	�'��4K�Ҹ{�\۳|���Q#�>���d4�\�
�����M�@(�숹m.�~�Y��C�@2�`A1AK �J��3m8D��C�b�*��\��J�/�L��';D��XpF�R�*�;��G{�J��g�9D�X��J��j�FF�8<Ԩa�6D��2�G�-���Į??*,��'B,�hO?��N�NL�0�C�4$"�x�w`%�!�H�y`<4F!u��8�w%�i��vÉA��<��ꁷ�dIB��9 G
[!�d	5_�n1	5�֗!'��0���L!�$ą0/��U��N~�T��1�!�$�� 6  0��r�]��"I�5�!���'�2��`j�؊�E�h�!�D�RmΙ�+�UB�� �!򄉕p��b�7��2� F?`�!��t�����C�	B�6��5)�.!�O^�=��T���(i�.��O˱b�D,qT"O� �Z�CՌ�Xe�bw��$"O�e���O���ꌥi�����-�y��A�>��mH��#a� T��nZXQ�<���i�I�U�)Vxj�; .�'/\�!�pm2D��M��E���cK��rUISBv�����j7x$S�#�*3�d���m�V�hG{J?���k�R�Z����s=�}�d�s���'?�Or�=��#�.�s�܀J�=��n����q.�A���1��3En_
�%�'�ў"}r��x�J,�&���I4��3f+�m��hO1���	BE�4b��	%e[�t�`uB�"O<���Hv(b3�m�td�Ӟ>Y����%�0H���j�6t�D~2��5e�8��ҌO�(�"iJٌ:uBB�	�'�&t�sB@RF�Z�#?ZlC�I�g������32������NC�ɟ%%�IZ'�/k�Es��͈^@�D/?�M<E�$�^8}֔�1O��v�H�e�}"!��  �ŤP��E[��ȻZ�: ۲^���	R�D�����z)�u�[�&��dE{J?��
�^�Y�.�n�`Z' |ӾB�	�;��Xs�G�j����ׄaC����'=�O�qO 8��\Z�
�R��* MN]Sfc-�S��y���dy��`פ3�B��D���IxX��p�	NR��%�&8H���	�ON��$WB}҄��1s��B�͜�b��/���䓋hOq��,�Æ	0\�:tA��^�[p����IW�O2�l���_%��Lwn�	��)D���m
�X��܃rc�;��!��,�6�S�'9�Ӥ��=2���Ɇ�%|8���
4�X�Ӭ�i>�H˗-À�
y�>!�l���S�W�	:�B$'���'^a��Z�]J4L�V�X�U�3�ԁ�HO��'����䣒^�<��EW�`#n�!�y����:îQ�Q�##�'����<�}���3ZS}kŌU�0��"�AZ�<!$�W� ��2���>!{��V�`�azbܑ ŨH�̘3���C!̍�Px�ik2M��@�$EA�w׊7��)�
�'��1z!��'�V�Y�[�=j�j
�'
$b@�zZ^(��i�
��	�'��.ͮ�L�xq
N�R8Y	�'LX��$&�]���Y�
��9����~��ʔIK֤̑lE��2��%��	xX�H�ud��Dx�Hy`Ø==��E2�?�O:�e�dLR"IS�V蒥�EaS���1�ȓ/�x�@ɕ�X���a����	H�'x� ���C��3�#
_�A��'Tl�� AE�1�S(�5T�<h�'�~�a�� �	=�.E�J�Hd� o�<eH�~����(L�X�Dؑ��L�Qў"~�I�R�l�@�b˫`��А�>I&��$�$�?�u���D1A���<����l�<�2�ןO��@��%Ў [8HSh�5s$�<�O�����I4Y�}ّ��v7UXх��z3
C�INҶ�ӖV#H45��^$9z�����<����N�E��S�,�6Ȅ �0>�f! }��A�7j\
�E�X���ضDRN�zO��S�3�	:Y�2�S�F,,U`p���Wn #>y��i7a2]��l
]��R�ku�!�Đ�*}��+_�(��XRը�# g����	��y�Y�$�Ӻ��"܈v�"ayd�W���A�W�<It��^�PtL	 W�Ti-�m~�r���=���"! u���U
0ې��4�
<��2���H�iC�X'�
z�Z9�=!	ۓ%����g�1�����F�[Q���J�'�H��!�o56���C?���(Oz��DC0m��pC��
�8�6ϟB�V�)�	���I<f�Vx���Q&[�RQ�[sP�����>�Ğ�m���r�L�r�&�"��ZX�<�c�(2�$�)��+]�VX�U��h�<��+��-���$��#t���r0�:T�����	�S<��@�9>���3D���D��-k�9��Ȑ�6�:b>D��q4�ȑwjJ�'ڒV� Y�r�6D��� ����ݠ���(�H x�`4D�P��&!D�ɪuc�1�$t;��0D�챵턬aD���' �vE �;c�/D��j�@��K��}s��T	�Ѣ!�:D�(�������a"-E�
��7=D����΋�Eq*4�U�E�?ߌ��S�9D��Q�m���`�eH*�$1��l8D��  ��� /"�48���ШU�����"O|MnϢV��4+�d��1�:��q"Odl�wMT#�i��9Y�ș�"OZ��O�WJ��E`Kp_Th�V"Ov
��Q�{��d`r�D���d["O�u�T�]�z:M���"C�D�"O� �O�]H�1+a���W��mA�"O�T�T���c�K�*�\9q��y�,�i�BᲦb�"���z���y�D��p��Z6ԯY�����5�y�&�JG�,�A
T�����%�y�R	6S�����K�V��7�R��y��ȵM��=��o�>C)j��q���yl^�O��d�'͆��2@��&��y҇�'�.q�ҫ�/z�*�Y���y�'ӄ��e�#_	����D�y���ֈ��G�'8\p1�o��y$��j�z�[u��+&�r��BE?�y�D�=�x�b�eY��r)�����y�k\�h�4q��H���ѠGd;�y��2vv9a"�";��"�!���yr(�eӎ�z��,2��2����y�y	n���(�(�@u�˗�y�B��0�#%�7M��{D���y��:R8��b <F�*D`s�[��y�Ҡ����֫��C���"�J3�y����e<~�ZG�W�0��`b�P��y�N�w��iu-��>)ִ[���y��� uP��0�R�3�� ��,Λ�ybc�P��&K�$�����ѓ�y�� ȚL�fR�n�&@qڏ�ymA�^h�͓�E�u��y��Й�y�M��q�Ȕ��b:]hְ�`#	��yR���+ج��@�ՙ@5h`��yBA2r���􌛽w͘D�O��yҫH}����q��aA+�Y�����n3L��h'@��0=q�����TȀ3\ldE�dN�l�<�6j �Dz=˕��6R�$��!��k�<��
-]���fN�"��5��B�a�<i�d�L~|�12�S ���C�MG�<�"�H���@Ƃ�K�0!�#@�<�B�قz�!b�K5@|�Q}�<	����t�ҍ�Q�T?��t�T��A�<!���9)]^Xf���FElJ'
�J�<�uN�{@����-�����D�<qӠ�|�K�5����?�B�	�Y� �R��صU�9�L3)�C�I7$D[E��n�Y�κx�xC�Ie	\��iM�#^��t�X B�ɯz�zȣ �É,!R�2�� RN�C�	�%������X�><�5�J�i>@B�ɟn��KP�Ѯr�|xr�BWq&B�=�@���Xi�� �a��!�d�G�x���k��E�O�$�!��� r.l�v�'҈0#dΥ'�!�$W��F�bS�2T�ڨ�����!��	""�l�1�ͰY��P����1PT�z",�51V�y f\�<��],hD�ԃ�e۰E���Y�*D��b��-t/�uS�B�_�fq'e:�I�^�lYwŚ*'�Q?a�F#]�P���Y�Y5|ႰG9D�,#T�^��lƖg�ţE.�A�2��E��<q4/�8����BW���1���Lp���!�uD
C㉲|_���e�
�$���M�9'�h�e	-/Z�����Ro�p����+�	3�ǒ�@$Nt�R�4<O�'G��F(V\��t�� V��`M/�pa��HN����"O�x���=�d�C���O�\k�|b�J�B8�bH�S?�!`O3<Y>����̎ B=���!D���c MNZ��2)K�wEڷ�]�9�x)��<aD�_����	)'3ȸ��%�v.�ps����*�C�k_t����� ,H���QdAt��̒�E�*$��D�H��K��0@�UK�G5y��]��b6<O]cr-��z��E��Bv����\�^����Ũ@�$�$��+D�p7��8�p��f$CV����:�	W��� QA&p�Q?��k/P�� ��0����8D�\[6 Á>��!
���2
�܉��@�d4�K>�� �gy�.H�3�2|i�'p��-+2��:�y/�6�vAY¯I��8C����y���K��(8�k^�V&�3�Z5�yRgÊjFv��Q�	&_f�I�mJ��y2�G*=7D!0b��!*��ʅ�yR���{&��"�+N�!�L��o�&�yb':)�ԥJ��ɍ2���<�y����2�p��E�2�h��gW#�yRe�<>o �0�$��q ԁ�)Ǵ�yc�/ s����j7k=�Uz%Ǖ/�yR����3��l���T�M$�y�Ѕ8ߺy��i�e5�j�#�yB���fP�á�*���@��y���IQ�R��!��5)����y�oԺf?��I�*ٛ!�d�{6����y�J�@���k�g &�$j0���y⡝+!�z�l\�W�4�x0�#�y�#�%{5TL)���,8����)+�y�i[�X>`�1���2j�8T�vǕ3�yҌ��L�� $M�0S8�R��0�y��B�E�Hٗ��
q��1�b+�0�*�PL>�Bk����B����/��,�l�;�F�}a�B�I�B8���m�9p)�� �)�]�y���,�,���''*�Z��!T�Q�G�{	j��	Ǔ`�ZUS4E�`z�-��O��:��A�>�p`
mQ�`�j0:��)ECz����>6,�u4������D-<f��'X�3!/*_r�����ӂ��$��ٰC��m���ci�(�@��{��+T�>E��'?V����Y6��ǀK�w lͻ3�T���/��)��o/�3��K�>�:B��Y�T���WYQr���!Q��ͅ�q�x�3�P�y�o�*JU�U+�O��6�Ma��� ���t�kF�����*i0�h�C�9���`�ÿJ��a-ٳ=ax�&Ɗ}�e"DO�	j���"%J�"Sg��?
��%J�bM6c����@��I�$�h5KL8�񟬙u�Hn����c�)�����>�W;Y>`9q˓4��>Q.@y�+s>i@@@D?Xdb�{�A��-RV�zeEӇV����=4|���WT<�|�'��󁓂+����ѝ�b�Dٽ2:˓Gu@0����e��x��?if�W���R,Ovxi˗�ВrR�U`(� n&���4y�a� �ax"�V�\����V0lP�F�4$M-��K� *��p%��>h�MK�P2^��3¢_W3fL�&�7"B���]L��(!�����ڮ>E����|2�,&ƾ���Q�6�<�*�,8�t�R�Σv`}KCl�6�³쇨���&42�" yP
�r�+��tb�	��H5��-l���L	�x�n�(��'rvE�E���&����1�ݗ�.ɠ�'� ���ܳdDB�c�nPZr*py@���Ea�)Sf�'� ј�������dX"{��
W@Y/U��sa�޺/�ɲ_�r�f�[�pF0+��SU� �%J���'b�x�fo*zs8hb��@1gC�P v.�l�D�����2� k&�'�4ɇ$�"q�P��ԣ.ڀ8��ˑzDj r���|�Xꂭ���Sk�ҝ
4�Z�8\A�ώ��v%�2�]�=�nX+FM\&�輄��48)n`zeGW�r6��H�5]&p���P~`eP7!�,D�@l��ֳv��hEW�v*�R�'��ŀ��F)�uGE�v���O6\�ƙAUAF��O�hB♄8�h�z�敄;�`!1)��v�ta"�	�H%C��-J��(Gk�c'�Б�r?��G�X�:�|�'�8�5ٷ9f���D͐�I��Z-O�Yw�6E 25ã�� �lev-su$A#L|"����t��+�̙V�Ɲ�B��<X���; hʈI,�I�����V�d�}+3�~�V���D�fm!�61�Ĉ�K�*^Eʓ�ʐ�G��*_F�����%�c'J��`q�û.P���D�$��i��_�kE����*P��{CKĚ3W�dL
8��*��=5�B�*�B����π b�hG^�"�й'�-uZ�0��ɜ{�J����_�n��m�7���Y-��aЮ� u0~ŐӢA�an�I�������O�@8�B�5L���	�bd�\�'IN�`!FK$9���OQ>�XuI�2J��Y�ү]		3�M8��2D�0�Q��s:�%�p��i��hP)O���T�dY��_�3�I�.˾����u�sbI�6I���dI�-êٺ��>e��,H�e���f�t��@�?�?��16�v���!�_h��Bl@�'��P�Q"7BLx%>��M��y
����F�,�¥�D*D���"M�x�:Er'�D&-���vh%?��ΚN_�%
M>E��-K1@fh�. &
�z4"���y��1'#\�@��(K��r}�=�2@΋P����$4T��I�dDr� ��L�?j9!�$@��L��oT6-�|�5�τ(!�01��b��}�D��aM�=!��&�b ���Զ��/E�^!�$S�`�
$+�-�b�T�B�٣z�!�$ �C���"��{!T�{r��L�!�Dԁ VL���.ʥ&�������!����l�l���`P/�r��G�Y!��'2���v�;[��0�'��0!�d�U?�,t��?q  I���A�!��IT����+pC�igeF��!�13�\�sC�{�d�0qx!�D1(H�b� x�(�rS��i!�$�&P����T��E3`���!�Ā�wS$4C�ɞC�`�
� $B�!�D�@l��P���3�P	�D��[�!�<D���j�Nӧ+���[&N�S(!�$@6#XnX��i��X�ؠ��� S�ɧP�f�r��'q`�����F�D����7=^�0�{r�.�`����-�n��#�֧�ܵ��*D�F�bT�Y1B���lڻ�V���'꜄IGȪfeR���H-��dR�n	6u���O���]3n�IŬ
w�]k�eѐ�~�� /]�~�:T�БFW~y�f�W1��x�+S<Kj:@q���-}���cL�'"6٣�FB�Qp���ǋ<?�zCB�Hm4\I�V�,|�'z��X��	5'�R�N�q��Y��,%<O br�Ϩt��y��le��BJ���6���I�b�r5�&��(q��p�A��W!�\�nףkz�S�(Or��6�F��~���D<4�6{��|���=1�.!qgƼl!l�'ym\EB�O��U I�}��� %�/=���Ñ�R����@I��p>ac�@��� �3k�%F��1�ő1�;A�O�>��Ir���B01�+�O�(�c���#I��!1��ҼCC��!K� 9��� \搉�o�Hh<�E+���0 �C� �Q�����O� ]��9�̓!;��8����h8�ek�� �(0���R��ᡱ��s�& ks��;GZ�=،L��ȉ�>�R��DZ�>Иd�uH��8�\��FG߽l��b$�Q(3#�aa7�ː_�V�fh@�D2�
C"��t���emT<n��j�I�e-L�Y���	Ԝ1EJT�?j.�O�%��<`698v"� �� �yݕU@�I��0�mу=�ȴ��%�^�H�9
eK��ϸ1*B�J2�'�r�cV� �/��8��*��%�z�aȗ=`y����0���J��4�v�sv�`��J��^*f�����'m�]r�o��X�4]S�σ0zv*S�,D��ŏ03��}�W�15*���mS��L^}��Y��	a}����<�'ƍ�#��|���ιP����   ���ܫ�&�P��d���<Io��R��2�֛1�����`��v���5~x�)+�<����"��бM~�OL�XЊ��C��4��N��R0���I�Ez��`;
�ЅY��=��U�&�ZI&H��UIXГpHC�`$l Q�)ԓb���b��%�O��iE�K+(���T�N,�:��ܜW6���bL������O�S�}@*���kF�.�D!̓8�u˕�gA�jũ r����x�<��䖽,a,�Rf�Ϭ)�����Ct≟YR�ѳ���#n��Ȣ/Ob]��O߬���	2DI��dL	V�[�aڤT���2EK�) �֩B,����[9�pe�&"[ Sp�
�R������iq���D����r�,�g'�e6��Ɠ� U�V��7 uN�X���%��!"��4i� a;0������#_ǐ�pէ	1�T9��Z� �az�Äh�����@?iI�F4����=0%�fO�I�<�/�2l����e�d� �G�n�xP����ȟxDiC��	F��*�bC�ED 	""O� ��`��YDV0�E ��}���ز"O*�"��!Pt����H/��8��"OP�Aȏg�x���螌��"O��`�/X,j��VJѹ���B"O�t3kÓ7�vك�g��Ji�� �*O�}A�#����&"_��k�'Ҙ��mV�jJ�1�/D/�Ԡ��'�1��� C��=	v�y���	�'+^����L&�!��-A
'�:���'�
iB��8��|�C�����
�'LH����G&@�BdN]�4��'	
�D��\_ԩ��(�( r�@��'�Z���ꉼ�h�ZңC1}>��
�'�`��c�S� Ii��U�jl"�	�'u�]!�I�2}v�[Q��Xc��;	�'��p4�3�<𚁩���8���'N�  hά1d)��t�bA��'���b��R�/��q9�
�x7�i��' ���!˜ 7[�(0�J2Vؓ�'v6��.ռbh: !��C�z#|���'dj����6?��=2���O���;�'{F�S�
��Z�8<�q�-���'���FL�E7��ْ�]��t�C�'#��%e�!~lT��"��#{`>Y�'��}J�o�	0�ALނa��A
�'ㆸP�W9%#0�ۑb��^����	�'�bq�"�V
^EF�� ��?H	"���'όe)sK�2 ������@���'�8��ꚥt�����ͧ�4���'�H��0n��<�c��0E�x��'=��2�6 v��R�!8��'���Q�7x�IR��(  Ā��'�h����5g���aM�!sl��'���T�� ~��p��A�z���'|:��E ������:@����'֞��& 6����'���0��'�`��fʸnW��f�V8@���'� ����^.܄u��dC�csZ9�'m"����HA�!�7�ҕY.���'�p���&D�͐���1C�v�)�'���G̟	�ZU�E�?��\@�'�d����E�ܨb@ �:^�
��'^��a��6;Ɓ����c5��c�'����V(P	�¤��(�0B�9��'!a����d���@��FdA�
�' p��OY�;h��c�E�)��Z
�'d�1�s&���~���)C0=�&a��'^�E����Z���b��	??�q�'��A��;��A5A&�4��'�>�ˇ��(����Ć��A�$y��'�V��b�ڈqm+YV����'-�U���e��!�G�R�h%��':�*�\. �d��K�@��'��2$�|(tX����%:Ю���'�B��@��P4(l�V��X8F���' ����\F`L�2K]	D*`"�';D�u��9uP��"R�F�CJ��
�'GL�Y��Z x4u�!�
�4`��'�2B�ڪ9CJu"�˜�VH���'����ak��n��T�ءT@��"�'�J�ᰬ�� ("\�5��J[���UrEy��R����X�t!8u�BŒ+�v����/�!�~��A�@�B|4Y��r�1O~<y�FR�p� 8و�IG�# �0J�B֊�M	���`�!�� �I��Q�<`�o�pkJd�6Ꟙs���Y U��9��i�g��8�D�#U	�i��#ƀ���D݉9��
�L8t`~�4O�;h4�X�ڪu�p�sG�7�O�ѧ�(' l���ݻ�v�`��'%*p�Lܸ�b�H�8O���3A�)(l#��_$V���j1"Or��EAD� �VI���<��PG�|��ޑ9���(�`ƩZ?5ڐ�Վ0�"���� ސM�2'>D�xbE�<$�r6g\�+��1�$P8��{bl�<qևF�����6J"���$�>|9����3Jo"C�ɤ)����Ն�Z���v*O'�����	\g|h��%�_�LY�E��������$+�D-<O�� �(��<�dm�<�!��1ttYz� H�f�pb&D�(V�	�utD=3ҡ�ǪT�BM$�I�à@�Z��	�����J�J���H�&N�D�S0E؇`w!�$_�3����RK�]�쩱��o��(+[H�I�nQ>�f���cшT�:v�m��D��s!
��u��$����
Qj�c�G]�����p�Z [�(Ƙ,������}R,��ȓ,̮�*W�Q�eJ"�/��]��YT�<����4ۜ�����/ <���T�<Ar��9�h���Y�9nT<:SdJ�<��NêQ
��D���9�BEK�<)�ŕ�m��]h���6�
��'�S�<�Vl�(H���ڡ��n�xI�-UK�<�E�Lj� ��C�z�n82�a�A�<��T��|�w
L-M6f(9U�A�<9�$�r�`x��@Ţrhx��"��<�SLޙxf:1��G�E�r���\w�<y��~9(��`� �Y�h��n�<����Q��ds��7W����)Yo�<�U I�zU�Y:@
"�&`P ��C�<��E#^`u�2��'��̫��`�<I���+S󜹡��@s���fA�^�<���ͻI��P��;\�ń�Z�<�Q\ьD!fG�_-8�Z�NT�<A5!	�qYr���E�J��ёsJU�'�ԁS
�W�g�.^`���A�Ԉ9�Ԙb�ʓO!񤗘v��-;�B�X��isP'�8!�Ig��3(���7�~�S�M�;�D��q��(K�<��	)6D�+uB ٦(�'�6x��iE�4��E]�f2���'^8������)��w��XQO� �3*�*䶍��N�G�OK�\S�bӂ�	w��k1�u��'�`�C JMm�����J��	�f}X�W�����(��5�<�3�2GPT��]�^ɀ��)ۡ�D٢+A�����'b�<���#z��`ڵdʼ,!�PAr*�O,$[�L�<�j��`nF�n�ܬ*��'l���ŧ��ɮ�[�Z���g��}����{���W-�:�y�O�|�s3��%P1p����,��	�I�r���]HX�%?�X�XO��D6�0�撼5���xӌ�F!�$�!��0yT��Q����rJ�<f,"0�KSy�K��z����4� ����'���	�wG*�y�Əc�����ܡ��T{�'b��贅қ+��D��`�\V�1B�ˋNX,���K��8�0�E� �#�����%�)��@���d�m��urtF��RC�	�#䏾*�yb�SA��3�����Pv��|J�G��4p���Ί\�qP��M�qph���Ǚ��Dr�W�^�>���
��y�]2�p<��/��*�`D�F�	�p�n@��KW"	c�ԊqbF�r �L��U�9�PF�-��?���� G�V�{ �D)B�Rvb�I~� ���^�J�E���4ID(�(u����h%񩑸%'[��/#��5���8!�d�&����҆�-�8e"[�/�޹1�jJ�*a��J�O�U&�!�"���"N�P!�)�'�F�	7�b �h��U��~�K��E�J�YG�E(.�pL-��J�.ɣ2kN�������B@��B��$�i&�Ⱥ5��m#��sD�K��FK�?,��PvN�?+"�[R�
(�l�8'D�K4����#���aO�vE�e��	0:d"���g�-c���cR<1m�˓��U�c�	�L�Д)WL����	Ћٵ9��� �10H�-A��y��D�-�pq�r"O�8*��=ǔ�R#��O��4*OH�q�>���	-0F�$k���O7H�t+L`}��Q�w�t�OE�X���Iݣ��?i� Q�r�Ȱ��X?"���j�!�S�p���/���3�^,T���, h�џ(@D]9SX�RJA�*yNE�w�$�t�BI	��˫��1�^�AN޿j��` �O�
s�T|�bE�����'mJ��b�7�������0r�DmH+O|�"��ڠU�ơM��|*��۷G��J֮τW �@����T�<�0FU%v�6��BM
�@�J �rja���� �eU���g�VŮ��C�|
�) ���,Zq:����+Tþ��c��:�z��"�M�h|Xr���;�A��'nD�9��pK2}{�H��(����� t:�1�Mٿ�ħ㎅!Wn�1�>l����[����C�*$����9g��#�\:Z��'��+ЯF?�ɧ��i f_�(���a��\%@��� "O�@��E:;�@1�dԬ�
�yQ�DV�@��i:��ч�S:$�H���`�%�4��ȓ�R�I0`�8|#~���̓�h��,���e��7\����X�l�ȓ:~���T ŜZ���`��tG�T��'����q��C�(ڀF�\��|8bdpV�c�܅�P ��P��[���8��P�-��ݰ�@�*Q.�ȓ-�lҧ���D Q��á5�����)&J[� ����dʴ�Vt�ȓ#����g�N�z����[�~�х�/�~�㏟"`����
7�z���P![�
���M3���M\���5��Q�q�U-�
LC$Ň�f��CR�B7w�B���m�:3���0��-��^������� B�ȓm�tH%��  �����<s�"����V�u���B��P�WcZ'O���ȓd���h$�5n���	�z�1�'��|�1n\؞t@`c����)�R��U��݂��9��*W�j����CB̧V�f��,��kd� WbU���qLְi����u�i�N䒃J�Vx�D��#�O5T��fO�o��@$�L8()�D�>9�AH�K�tXB��ƪ3��Y���Ԁ"�p�;.^����E'C�T�Y�C�U����Q*���W����V��u-�Qc�%R �iehH9jT�`���6��M�"�T����N?i�$*�;@���*�7�R�HgB*Mk�y��L6�F��B�+Oi��/���n�*�2�BED���UL(�ح�r���$SN�`��_b��ɖg,^��W@�1l��&���xB�O�+�"��~NEA���H�� ���ɋ��]�w��5d������=%'<���oږ}kz@+a�'*�����L., 2-�c�#�W�Y� ���"bS09C��Q�@8��^ZDpb���N��)�?�"����P� ��B�%�1|���O��9��_")���sI� 9+�]���Ja��5��I�>�l��BاHd��)vI^!%����ơ;.�Mꄶ�U���H���E�A.�(qx�)��<	'A+�<Y���W�"m����h�����/~н"#LH�Je����-֫9��ẁ�]�2��,�����j�FyBĐ'9���G̟���r���������GKQ�3��<_t��iYw��Li��B��0Q+ט1�-�4.{�-���S��~�!���L��|��ևa�b��Ԉ�9J��k��<�dUx��+N�0����w�����V�`�`�#��3r��U��o�� A*��e� )PL������1D�H�bǝ) �p+�H-Q{f��れ�(tة����h�Z%W�;,�P�b��<����_b�0�O���J�@׊IXP�T��R����H����!�z���* /��#���[�"��Qa�����z�(�x2-~M�J܀���È��g���n�3�� w
M�3�?����G�ڂ~92�0�N P꒟:�@�$��x��Ј�	��59���"[�Azy�7�������40=�eY�˗3{����D�!�:H�ؖ��`��N�\��T?�낥͝?�hS���<����K>~��c�Ӯ���Q�k�<!sh�S� �pLإa�n��`3�Ę0K���E��%Nc��'�&K$�&��DƏc�yx@��wMhX��兴��?dNF�bh;C^�nƴ�Ƌ�a�����6,�u�.OR���΀����I(z���q`_Wl�B֣�j<�B�	�>��rF\�eV�se�L�=����(S�-`ʹk6Eq�� H�#OL(�q�b���?�N���'��Y�l#�}��p�|�c�iσgZ41��&Ch����G��(���R42tM��c5#���=�˚�Er1z��IEA8N�:�ᕡV=�p�	�P�!�C5��I �B�s��0��2�!�;B Ƹ	�� �?Ш��}q�'�HJ֏�e7j�s�lB4s����'f�|��!�Q��1A�a�u�
	�'��y�b,�h�M� |��r	�'� ���s����g��&����'Z`Rv P�[����S@��0�	�'��H���8�����^,E�l���'�(�+W x��#K�8V�x	�'>��Re ΰ �Ȉ�$3 8��'?��(��*x�HU����8��<��'�4!�!�/U'�%P`KnTI�'^J�"��=e��WԎ3|
D/D���Uh��B����Y66x䩐Ǧ-D�,���S�VЁ��f��e���C6D���LT�dh��G�M��	�a4D����P�%;5!f���m,�Ჳ�)D�X`RG�),��[�ĕ�v��M���'D���e�֏NKV���l] <܍�$-9D���v�ԯI�<�A��JLX�ro6D�$�D*�E�R�y�]����i4D�j���H��T�_��H����4D�����
j4��j"�N6m�>���5D�`4��wvrx C
$֥��7D���AE�
P$\� HG2}��$��2D�L�w��w���p�B"�~ɱ�i3D�,IA؏$�&��Pl�2*ULi�W/D�P�#�RF6(fa�'
(� ��*D�ĺVIZE8�ǉ
[Τia�(D�D2f�L�V�0`��I�����'D��P��a�� C��ؘ�2$�$D��1���/YP�����5A�HPbK&D�|+R��{,�I8�w�d�pa9D�p8���7;����E���%z@�6D�@����	X�m�p	^�H�d�X�4D��@LG�F\C��?2j(��!3D�8���Q44��X��UOFI�g�0D���c�˟D"�����9.�H�� +D�4ҥF�,��!�GIĐp���55D�d�1!P
4nΐ�e��V��pE΅�0&�
[h����>���ę0hV�JK>�;����,��<�|kF�  Apy��������	�+*έ��SCb��6��*gc����}��X���)!0�禁0��кV�~���"({6�R*i���	�<�wC�
���~�RH�DF0e�z�#�CX@P��f��7}"��P&2��=%>���?�r`+5/É(q�4��,=�DP�a�{���'ɂ��g
� ST�3a�1������'Ȁ#}�͙�)�P0:1BA�%���1�1ݞݑ�
ç p`��`E�(�����V@�y��WC����IH���G��t�R�F�ĭ�'�Z9��T?m%��:�k�d	�s#H�O���o�|�Gz����iH&`*����5z��d�H�RV�'{�	��0|:� �k%���e�W���f��|y��)ʧV'���aA�:D�]y'�ޣh!f��ȓ/>�)�� �I��A�`!��MF,�ȓW������ޝ_��e�W:�6��'ў"|24�Ҹ��A$���X����<I����M����3G���ǭ5}2��Z��OƸ�5*�E*���IV61���e̛^�hY�}���i���A %\����.p���.KN��I���)��0�dZU?>A*W�D<Eb���$"�S�� <įF7��=�7?��QӘ|"�)�X�~���eNĄP�6H��[� ���'#$�&�����i�?i�bn<.��g�I(���jΦȸ'Jmh%�Ok$�2"^�?�`|J���xl�O>A�#F.�z��>����\ `+6��G�؀1&�Q�<!�[�}�ڙ�cgD�Y* ���ʙq�<�4�� "Ȝ`��e����	Mb�<�աB7 ���e�,�t�a�<)�S��VQ�LJ=��t[�'�^�<��l�!�f=���ߵ,x����t�<�dK �S}D�A'���.ڴlP&$t�<��W�4�>�6�
7Y�^|�	F�<)�� 4r�B���mŴ{�����|�<Q �Rv��ԏQ3q�Pi6	��<	&ȭ)>��Z��[�fe����J|�<���	,���iզ%*`�@b��s�<��(��6B����*�z� ,�J�<����E_����F�	^UrԧSE�<a� ��:�d�Z�̎�i���
QX�<�����H8,	�Gr02�� El�<IT$�'UQ�u�A�ڽ��a��g�<�DG�v�2�;%H�iEȽ�W��d�<�s�c�X���ț8F�j�,�T�<y�lz� y��R^��q�f�<!&JT���[�B܄�n�`�<Y�
_-&c���oåq��D`�\�<�vG� U�R�jr ��C:6`�f��b�<)s��\/^����B�J����r�<�B�����WR�ĪD�4T��P��o�*�.��9�`A3D�3�!v���L�C�p%1`,,D��˧c�*(_*ٙr�\7eT2E2�j)D�P��KM; cl�jd�ܘk@��o)D��3R�F3%\��[�!n��&D��s�sv��V`̶}�mr��&D��$cY�h�b���o�2����%D�̉uiÅY!�APt�]�?��ri>D�`�҂�.�M��N@
a�� �t�8D���b�ͫU{Ray@�'_De F@8D���KϦv4>���L�:z�����4D�x`��b��Y�Y�|02�3D�Je��$+��H��V >�rp���1D�����t] ���V�F�xp��$D����NIi.|�H#���ah�� D��T�S4��1�$L�Sw�=D���ǡ_�t1����a�gb���.D��TM��hP� �$���d?D��ण��g��" P�H	�]С0D��zv��j��{ �"O�"D��C.D��Q�*\&;�`��OL�W%<���-D��2�jV5J�<9:��^��4g�,D�8b��*,<�ቧ/�roP�·f)D�4���ͺ"6X!B�L��B����+D������K����c�.+����%D�`{�%4.�X��jS�idP)R�%D�p �N7d�0.�*�~��b0D�ة�Η8�ab5�dV�-��B�ɬDaTY����t+�8�0���}��B�	�t:�I�AS�iQ�,b�HD8_��B�I�U��B��3���a��#tB�	7H��u� �Z�9���@Z'_8�C��,�:!�ɯnS$pR�@C�++�B��-F����JF��i��J�	��C�?f��8@&u��6��Li�B�)� 6љ%*�E�"5�7��\䔝�S"O��Ȗ�]�
P���P�}��բ"O~��Q�D-m���Ɛ��8a�"O$�y's2���aQ9=�Z02$"OZp�#�L'6��jsAN%c4}�"O�!�R�ݤh�Ax�@N�-��@�"O��
�͑�4ج����b��yV"O���NK�.�!� E,���w"O:��w�-���[��	G^5y�"Ox#%U:b��a��4w���"O�l�VȈ�n=����
^0δ��*O:}��@�c&��p�B!|p�b�'�N(�Jγ&����mxp�h�'~F��T���}�ܥ+��D�$\�B��;^�軖F�1`�9��f��0H^B�?.
�{Pb��!3`�[��\vC�0y�h�C�',���, �.B�	�ku�]��L�*)v�;��D	3P�B�	�w���j���S&U��a iԪC�IK�l�	�DI4v�&EJE�Y�c��C�ɢ7�V�!H�\� �3�؂U�C�	�<,�a��kU�,
�dh�'�G�B�	��ܻ1�I�V��j���>�"C�	-�P1P3=uu MI�n���:B�ɳk~������75�2I��RZ:B�	-a
jA;�)A��`�݃l�B��,���f�X}�NMA�� �B�	�8�#܏�
Uz!�ſ%��B�ɦYhY��'��=Zy��eޢ1��C�	�g���0�%|�M"��)e:^C�]䞜�e�3PB(�b#��2@C�/N�����o�֤�UJ�+ �C���mЦ�
�#$�|u���C�ɵW�dH�U�0e*������4��B�en���E�̜"���D�C�	�'�L����X|����8o��B�I3C1a+��:K0����J�$d�B�	'�.9C�	�C�����'\6'��B�ɶ/3�Tx��" �J�c�f��})RB�I&]萴X�f��*37���<D���ă�^��c4/JX�PA0D�4h�)�;�Ժ%.�,!�jS��-D�c���]�~-�E�Y5(� �'D�Dه�H�o����sŇpC\���#D�(�+^�T��|;6A��_;�]�V�6D����K�T��*��%*ֹӡ3D���d@�4W6 �Acém��us�3D�Ⱥ1-91�@�8��4���x��/D��s���:$����T��?��(�
!D�С��M\�� h�/,�q�Eb>D�(�W��'1�*mb�*>!ò�	�=D� �Ϙ�tV�e�v�E�3-���<D����].�0�!�NNru+tk;D���&�!BƞaKUm !&9 7h%D��5-�Z���F�,:���&'D���F�����)% 6��l2e�%D�DX�ԱWpp��7)�2Q��J	#D���W�K:�T����γ|�$��$� D��R�M���[î���W�)D�`�#�L!_\��P�˅v;��)(D�4���8sE�)ؐjD�wL�ya�'D��R-S��Y0��-[A.���N'D��Y%%�#2P��e"G":�D@�f�(D�T�v��>yʥ�ŮϜp��I�G�'D�� * ��H,=mz�(��1+T��C"O���5L��.��aPb��
�M`�"O|��@T�N/ƙ��O�&/˖0��"OB9r�H8�J�SF�;� ��"O��Ht�$~h�g������"O��I#`>Z5�Y���	Y�����"O�,���Q+5��b���$��|��"O���#X�f�H�9�!��b|t2"O�0�� P�.�p��@_� ��S"O�TÁ��(M:�P�	S�M&.\1Q"O��Хa��tD<��Th]3�T�:A"O��B$�Bt�)b�N9V�˴"Op2O�&�`�
g� ��Jb"O,E�4�U����^##�"Yc�"O��p�g3R�i�n�|눁Z�"O4]z�8P�d=�j�}6�l��"O������p�ܵؗ�C�b%`F"O����.0���G�($ !�"O�HqcƳT��<[4l�S&΅��"O��XȞ(yt�#U��/	<K�"O���3ڑbꮸ�1�H�B���r"O�	���	[�x��]f���U"O@�xenmx$�%w��I[�"O ��W��l"��IG��?� �� "O�I���a ����"O���P1<H~��OB%/����"O�d �ȼC&4��C��	���k�"O�qH6�]��S&Ic}.���"ONɺ��Y2Y�9�`ɰTc��Kd"O�xi��ʖi�� �-�i�:}��"O,��w&�/�L��f&�.s��]��"O^D�BfP�vU�52�#LK���q�"OH���m6���Fcۀb���)"O�X3�o�,̔H!��[�x��'�dD� G��]e����κzQt���'�~�2�*$�ʴs�D�m��h��'�=��fZ&dV�b�C֫k�Pܑ�'�a�,�d� ,R��H�qER��'�0�Y�aL�C��m���i&�Љ�'ET��ddצ��r$ȃ=c�xl�
�'��1"G�؉+��Hd�]-]f�1�'�,�(B��e����d!�|t��'n ����_���J�Ad`XY�'�r���@���
�&.��5��'�qР��*=B�s��4(�8�1�'k:Y��/<�PÈ��n���'���`�G@�|��Wg�w����'��,���*<L�������}9�� 	�'1������*�z�,�9"�t���'��3���AҦˉ�v-(�'�6,����x�6,�v$2�0�k�'�&U�5�/#�6=C�e,\5��'߄]Iř;&�^E�֧�%$��A	�'��q;�Ɍ&�
vn�5
¡��'v��Ӏ��?����oZqE��'���C�ϟ?	/L噖i�
���'��)��Ӓih՚��3M4��R�'0m�蘱ASh���,9�u�
�'��mŊ#ƺ`Y��*-��%P	�'��3FƢ��L�5�C�h�i�'[BL*2@Rj�|�gH^
5�ֱB
�'gFX���S�6�d��%g��3P^��	�'-|����N�t����"�-�d���')�	k�@ 7���,�\�2|���� ��������	��@�&K�Q"O~yBP�j�x��W��$A/6-��"O�񻅭S�4�����J�e^�C "O��h��:�3莢=$r�!"O��ǁ�h9d܁!��;%��S2"O��F�)ǈ��D�ת	���"O.�*n�5�@�Ȓ$E�ݡ"O�$8�E�c2p�c�\'�L�b"O(�s��X ̙�Cf±_�@�"O� `   �d     �  �"  �-  �8  �C  �N  �Y  [d  #o  z  ��  �  I�  ��  ߙ  #�  w�  ��  ��  A�  ��  1�  �   `� u�	����Zv)C�'ll\�0BKz+ �D������b�6�F�y����yb�҅w+~]�SO	"d��G�	�}<��2�"��3��M��1�cX:\'�N��r�ɞ=n���)H ���+ɀ>
�[`e�-��"6�	92��b��=CR�t
�i��d੭� 	��'�?9�g�x����mN+V��ea�.ĮOwRѺ��F����)5����t��6M#)S���O`���O���&c����g�6O��TȅN;B��OF���Ŧ�'��j[�gf*ꓚ?Q��_N0|�V�M ]�8�&���?���c����'���'��C�$�uW��5k�����&Էm�f �5�̩c�8I5dO=-`��F]��Op��&�	7`ڦ$(��

��Ȧ �b�X�yӫ]R}�<O��Of���T"��A/D-�iU�.MrY8��]�s;b�A��?R�"�'���'a2�'��'k���{�@��r(�MB�+�U�=�c����q޴Yڛ�r�^do��h�4)� y2�i�`5��Od^���K�x�q[�A�)>tj(��8�W��XI�+�	�W���a՜@���R�%3f���L�;P�	��J.P�h�'V�]����c�2�o��?=�'YNq��'��b�(ꥢ�7J<BQ�3c�yo�(E�N�r�㈲G�x��o�QDFE����rܴgΛ��{�N�����m3`�ZRj�\̾��B��+��T���(�%`cӎ�l�,�M;B�J�g���Z�a�W,T�P����wj��4�I�<V�Q4��/s�aJ�@�:ӠT��V��G|ӂ,lZi�6��q⏭	n`��S�9XxӇ��Im� ��3M�ar���M0��47b��e�1H��D���?A�"��2x"�� NJ&�,�(���3���D�O0���O*Ql_��`	kK�����	Ą��*ё�?9.O\���O���Z/4��ρpKt&ך%B���	JG �#I�&�<�&6G>8=ٗ�IO@�)k@O���^��dV/rK���1�U�#3ֽc��1?�b(h�*ҶQB��	$]|˓��I�p�pm�G��_�-c5ƣ	�H�D�O�D:���On�Ľ<Y�Lkj�El���<M�!�߉[q�����?9�!�_z`�M>���<ͧ7�I��c�<�{ԈI�[�,�.\�?A.OL2�K����q�'�yG�8w~�٪�oH;W�D�YZ�����y�bP2uM�x �� �q��i�L-i�d-rԦW.Jjq�ŗ7V(�;Pa���d�5X��u"̜TW<$�f.M�t/h@��-Ȍ����\��ikQ���V5��E x��9������M�w���|�6.҈-pR �0M� �K2�x�I⟰�����D�$)��y��G:5~p3t�M&�hO��D����"޴��وX�X@T����8>�\p��,�<h؛��'�	;t`9�Ɵ<�	ǟ��'��	�"E+��5����UF9�7	P2H���ӌ�	#�T�)%@��{����?e{����Qa2��8(@���=BǼ��B�7�rMj�GN�(t\eRwU�+�NTұ-3����R�O����`X*5�Me��:j�����xӴ)�'���1���ȟ�'
@���zFtH�R�@/AKr\��'Uў"~J2�Nl��Q���i6��7�?���b��gӎ�O�)៴�-Pڤ����+.e�<# �\� C���g/�I��`�IfyU>��'j��Ӷ|^J��2P�K�Npˆ�Z�Lz��S�ȀC@-�WK�*^�n��W3ʓXx�]�Q��.<jr)"�@� ]
W0R�"�p$��%�� ǆ��~X u�̖pQ�t� ߜ)\f���H�V�ļh���!��d�����D#�I�>h��+D�]�V�j�I�I��@�	ҟ���l�'�1O��Y�O �V�]�`%�_f,L8��|�Jo��ImAyr���6��O<�I�|��z �C�W^8E��o[�����<���?�O��0��ߏqq�Mj�4FϠL:����*F%O�1�\ �7��.AE�D�SV;.�<	��������`��v#����^X  yr�;
�e`�*.��͉'Φ�ם��&Ϧ���)�M;��iy�BǄH���	�y���$/E[�	æ�s�����?��}�b�Co���3a�C;��*���J����?A)�R�o�!;i�@�K32���Xg��-$��)�4�?i��ivx\�E�0<�t�s]����&�MC�'k�tͱB�_�x�n�C���B�������?'
��&���jo��.ѬM��SD���>ٸ�.��#	����_i�����H~b��#0��0 �$R5ч⍳;qp��k�9�,c�O�X��礗�ըm���_�"w|��O�Y�0�'�6-NR�Q�'J���3F^�e>�U)��A�2̈�&����M�	ɟ��Dy�F� Q���� W�a���A��"?�p�'��6�'�<6m�O@��e�[�k6J���f����'OڦQ����I�FL)c����	���ټ�QƜ�+��@˱TQ�̊��	" �ݱa��6R�R��*<�z�O>�d���"���'��35��Bm4#���.6�,?eB��+b)D����BE��UBFT>�C��%+��݊-�:80�族��{���Z���l���DX�^�"��'���'Gd����_��a�qC�<~h�p�|�).\��$2��
c�ěU����OB�nZ �MI>����+OV�
Th�#I^��Re�=
=9�b��w�^�l�˟�������'#��|�c(@d&p:�ɲ���.�SԘ�I�%B�)U����8i�(4��@4��<	���p��8E�V�W�\�mนj�~X��@/�8H�MõN�I�8pIdC���K�8@��	szL��,W�;��$�&�����+�4D���DFxR��������1���a&�Z��?AI>���?�)OʒOvX�Q���;�q2MO� �| ��C�O��m�؟��ߴ\l��]>m(���M���?I寉4r4��Ҧَ,n�}����?Q��u�ؐ��?��O5�y����ey@e�N�b� �aR��֒\��*F䁱<�Z%i�钽�����Ӓ]g�M+�"�����h�L'/~�qiV�6BW�|Ò���Tq��V1b�R���,uQ"� ��ؔx�V�!oT�	�8��-�!�d-#����
I�>8ʒ��'J���OnU��a̝e$���G>h��%�|.��&�6m�OF�d�|"t�M��?Y@��^E�(G�� 3��T����?���z��{�Go��1)U�ѡY"*�b�'�l1z��r���������x�'����v�G�hq&��1��7q�>� �!�(a�V�E��,��z��+?I�������E��5O��k���60w��9��܊f�4ػt"O,�C���<wjP��/J������h�D��۞;Ѽ�#�(Ļ6�͉7hdӪ�$�<�p!������?Y���$K�<��ف���<$�x� !�C$�mˢ�S �L@P �8;�L(�F�|��'6���1�GA?�ݢ&�Ax�(�9�
���.��;������B�(����L�Pc�P9��)F�s.h
�5�b!A�T�N���x�� !U�C�Jf�HŔ'�	���jɟ�'4!
p��zd� 5"�G1��'�'O�V�,��r����d��Y��EY"d2���:l���')�7����ɷ�M+.��i�|�s,��:����qe�X�uOO�W�8i��i3�?	���?���L;�n�O���>%��
�&>h�Hl�5a'N�^���c�a��$���r�$�Hx���F�	2 ��i���0dN�H���L� Q  D�F��j� �Wx�<I  @�s?^m��B�^��9�uU,����OL�=)���ܝ0\��#��a��|"��,N�!���	1L\c��j.}�6/��'��6M�Oʓhz����V?��	�g�V�P��2t@�Bp�Y�$�xH�	��8K��_�$���|��F�)#A�mss���I"4Wv1�C�u�����,bt�����(��b�4NN���'V`p�r�� Wu汁3	΢$(��3�@�$��П��'Vj���Hk�M2$NA� 0�`N>�F�F|q��R�d�A�
�}ڢ��<I��T>i���R���ِA�XGfȱ��Lvì���[y��& '�7�&�i�|���;��q���-�����I�\-v�8���?���D�(�<d��������B�0HFb+�F�c:K�T��PوJ'́���H�:��&%��{'Q�#L��t�R�h6�2R	��Dp���
�?E�c�M�Q��i��B:[RDx�,#?Y��Ɵ�ش ʑ>�'"��3��r��8��I�;��?����~R�`�
&@Z�*���/��u{�ŐG�'B-k�"8l�@��
0�VjTH!gZ�kcN�(>	�I���������P�LE�I����� �;;=.<
���0+�ѥ#B<7?�܀�A��'��!���G;�C� V�'uU�`
ŭ����a�%�TY����t�����S��ۣ߬%�,q�A�Rx�s�_|���I�5K�w�H�%kB�$�+ �T�Z��������h�"�'�ў�a#GT����q䀿bW��-Q�<�E�H�!����f�G�J�p�k��џ\����HO�	�O�˓I{�A�'�J|j��]U����:w����t��O��d�O����*�$�O��@�ni{w@�:?��E�5Iԭcx�"@�7wIj4��L�?k��7M�njJ���$ʓr�p1C��*N����19����l 08�8d��^�nZ?*H�c�⋜3\�aė|₋	����7�I�		�#��p��?a��D!��8�5���=ժ�3�*	?��Ԇ�I}�%=j��7��W�eز�֍g0�&��#�4�?�-O�=��]i�D�'~�}�@m�{�H0��oL�\>����'�#�8,���'��ỉAY�5��@�uk�U�n�6�Pb%���\b�J6�˩D�U�b�>VFh���򄜒Qo�`K�ǡmmX�[U��&l/�\`���S�8{����OX*��PJGv��Hf(s'T�O�H6�'_����k>�	Sկ:YJ�+�%��#�Oz���� �F�zl�!�)bꦕA���=��|'�'9�iC@(F��#ž7�ʀ����Dш"�����O��D�|dh\+�?�6�Y8J�Z'���'\%��kƠ�?���}B�I1AX��&,3 �O�^_J���?Q�OLެh��Y<���\�t�RA��O����e֢d�d%�У� !�p9+4D�y�'4 2��s �5bv��疶m��e�'��H	��?Y��Is�pzsfڥOb�寧X-:V����y#K̰=!Q��`H�(S�P/��O��D��BD�L��@G�T�`���zӋ�Q*�F�'�B�'YƤ)\�'���' ��,#����� �(�T�:3C�&O�R؁`��X��D��	Z���E��d�*�z�_�=�h��B�M�za耊K�e�>��,�A5�y���L�uA˓ak(� �=�n��̀�^��\��C~R`��?)���hOxD�'c��+��b��S�lI0�"�2D�L�Z3.�;���a�Rqj,�<Ʉ�i>5�IlyBjX\	x�(7\@�8i�R)HF}+vF�,40��'���'�z�]ȟ��	�|�+�8mX\����(1�&P�%ڊT-������;jPKϚ6ZHua6DӖZ6R�<)��KD�? &�z��O��D�����8[��'�ү��L����~A⌛'�M6�A{-C�)���O�M{��A�D�Z
�V$JH"Ѕ	&��'�ўLFx��F�9���Ü ���8�-$��=�yҍԾ%�p�&(Q(	R�x`/�>��W����'�ɤG�Z��ߴ�?a�4���!D�8����W(ÖxW@�����?��͘��?���?��39�hTj�EW����i�z}�W�V�l#�/��t�Zw��?@���Ey���/;x�R�)V���e[7��&P��x��޾MN��5X0Bm-� ��jS�M:(T�F�I)L�.�d�Ѧ��(O䄋U�ϫ0��g�S4Y+Rͫ��|�U��E{�Om���@B�,S�D�wj��(P��?In��Xd�99�B�P�h��D��CN����4��$V$�7-�O���|ru�?QR�ʣfFղ��&�妘"p����Iԟ�1� }ʑ3�0a:^H-ع��i1R`��4F� Xj��9�v���*Sr~��E\�m�0/Q3S}�|4N�{�h���O._]<l5��#J΅Yf��d�"J�O��5ڧ�?�q��5�|�Qkjp ��A��y"nZ�N�j��J�.��A��-�=��OĈE������0q��������4,@�Rm���'���'�:Qz3O�v��']R�'����9��A���9\晨U��%>�`�3��?6�u⠢�
S.�P�1�	T�cZ���'JM�(ާz�L�sÌ��(7�����z�>��d�;��R"���O��0�%�p?1���M��dـF�1!{8�ؤ����'E�p���?y���'Z��2�])%4�i�k�&p���"O�m o��Z�p��V�Z$��Z�����4���<!f�����u��L! Ly�N��L>8�@�ܙ�?����?I�R���O��k>����ـ#�4�A� �@�>�CC�`�\0�4B	a�-"tE��x�I��Q��0B��P��Rc�:$�����i�l���V9%�d-"�L�M����Lأg�Q� bV�Ҟs�������*P�Љ�9F:���O�=)��$��n�\�T·_��Q����!!���a���
�R�	cU� :q�'�6��O��S�f�Z�P?%�	3m�)E	۲5޸ bBP�jC� ����� QI�ϟD�	�|�����%��Da@Z/"����X�a�"
;<�:����8#����	�!%
]��(����I`TtHb�c�.j�~�R@�տg ���g�5Oў 頋�Op��??5 D$M2��5�px�� �V��X����J��8�Kb�ޔV�P�%*�O^a�	�\R�0���oc��3�Ѵc�D�$�<���Qқ6�'��Z>��������$m�WF�݌9;Ө7L<��'��ɘB+�#�����J4 ^�T>1�O��eP�Ѥl|e�1�|���O�Dk���<G4D�A�%8� Z�j3xB���t1�T+^�=i\��v"���������O��d4�'�y���>Bx9CA�Ƀ��5�֠�yR��=kn�8��?��r��Q��OQF�$l/Vvt��'N����&��}Û��' ��'��a��V�X)��'N�'���5&ݜ��ͅO�)q#����6�S�J6>n�Q��ے1�m��iW	v:���'] Ы$�_Uxpi��q.��Ӵ�,p ��A�=��w$ܫ��O�ށ8��Qp?q��K��t8�a�N��F��դɨ���F��	z�g̓7�DM�%��_J��;rC+��̇�lc�9cӭ�c���(���p��'#p"=ͧ��|<(i:D���-������Ɏ���#.�tz�=[���?a���?)P�����O��,���s��t���d���Z~�0�s
@%P�dA��x����I�g����� UU��2��ݡ$0�LeD��]+��QD
35��K�d��h/�}E{�׊s�Z�Z��U��4�c�=4�������?ٌ�3�f��zF�'q4����<IN��ȓt����U��k:��!��wc�e&�@�ߴ�?	,O��b&@�~��'��Y���L��28P��Q��VTğ���+��q��ß��'f�L�atu����$ڇ�?�Q���[�jQ����	��a�@��+���3�>�Q�@3�$I�	�@}q 3�G'_�d���'��/����dØA�'��I�N��(��_�t	��% 8
�O��� !cD]�a����ƣ��b����OL '��?�v8ʆ֭ר}�w�'���&n��|�޴�?�����iN�L�v�䛊%������+=���1B�U<��O
��pG�
.�XY�eߒ��X�l�2
zD��d&�4?rb0a�����ra�Bc~�b;�!ц��t�H��A	䄣!��ZB���)�,<�����|*���'pq��q�ɧ�@d9��F�Z�y׏�9|[�Kc"Opܑ0��w<������S<U���	��h�0��s��+�|]�3��$8�	V,s�l���O���x�V]Ke��O��d�O���h�=S����u|Y�n�@�h�H�F*uԨ������$(E4`�b>!r7����X��8`	� �X�bg�h+@��#I7�� 0"!k*��DD֜+���'yB|��!Ѽ� �񛣢ޅ"�z���+�%#�Q�'���*J�d�OR�=Q+L c5B�R�Q9f���y��k�^a�Ơ>d:���JP!�?����SΟ��'�FD���J�l�S�ѭ~ݬ�jW�G�X�2�1�':��'��O��'��ɍ�btp�%�2 ؐ]J�ƒ�W�F�B��L��C�+�>p �٦�Ij�':����%"i�%B�^�K�r[�%_.���Z��]��0��G*-Q3.#?��ւg�T�
Q���J)�w�(5%�P����D{b��*_g�A�-Y3"��$��y]�C�I�h�LĘHƒ��Q1��ԟt���O,�n�x�'Y@j�Au�P���O
��&��*H�oL�4Ѫf-�O��dL�R���d�O2��Y=�F�C�h�Ѣe�j[DIJ��
ئ��1= y)�T�T��m��剶ȍy�@(-��(6�ِf��1���2$\���.�5�@L��R�*��-;YΔ]H�i3��	���s���'�l � K��C^��	u��݈L>ٍ�d6�/[
�@"J�fit����߼Tw���G{�O,�6��6?��tjN��7EV�C��
`��uoqy�K��X�T6��O���|���8�?�R⎁d�nD ѡ[�v)�A�ӪF��?I�ZdUK�",
�*TDdÛc�n��g�L@��˟���/��%��U �G �1�Z-������ȃ \C�-[�h�>�R��_�=����@�r���A�2�G���q�S�����)d2�.�ᓪP����L�+O(c%/�G�&C�	_��H1�d&��Ju��:��?����_&PD�U�<`�s5(�Oym�Ɵh�����I7���X^�|�I蟌�Iܟ�;ɜ(P#��L�ɲ��\�р��͑�2�	*S� `0�*�3�5Gl�i�[8.�B���k8~�Z�cOT�M����F}�;D�+��A�I)% �I7Hn���Vb��^@��lڸ��$���"��'���'���S���>�PsC��H�`��$"O䠄*)&0��W-ӷ�ԒP�<{��Dퟨ�Ķ<�q��%#�dR��2H���R}2$}cd%�?I���?Q� ��N�OH��}>�97�E�sg�!��P�,R�8s�H܏E04����)q���p=Y&�L���t��d�S����.@Gl� ��C-V�`��E.3��T�����$k$�c�
@D��2�ԒS�'�6��F�ş,��_�
�2�B�$Y���j��!���'�:|�UG�$%
����f�Ҁ�H>!V�i��U����mݦ��	�OB1��cB�RQ����
�+ �MaG,�O�D�{�����O"�S2e%U��S2ML�hD�ϊiI�4��̎�)D���
��E$8�Ҥ���L��ɰ)^Vi����Ui�}
�dF��֨ɕ� oZ�g̊k@tZ�ςk����g �B0%�����O~�D"?I5OQ�HL����2jd�%@LC�Is��J`���A
�eZ&*C"�[��9��E����Oxu��+�X��t�tE�&D]�U���'��I�RRm!ߴ�?y���)�[�����	LX�a-}X��e�{�<���O��D�ZqT ��h??�Oz���K���pdР6�e�U�λK�*�bj��R�މA�Z��ᓼC�(Ie�#2=�!˂>,��D`�8�ɩ��S�OK��I�
���fCC<���'9��ңN�?�B��<m�Ha���PE�O
f\��䑨jE��k ��o��2��i��'8r�a��q�V�'���'�R8�2��� H[^p8��*��@��(l\`a��i�IK����F c>�:�'�'!(�D@8+<��u0���Ҿy ���ΠY��F��9�E��뉝��O[84ʇ�Ҵ�y����P�p�Aa�S������ذ�?��OB))S�'kr�I�&���`�*��`��X���y���h�+նĴ �T�E[]t�Iȟ����4�����<ɂ��
���f��u#�(KK�3����E���?����?q�������?��O�,D�#	���	Z�����!�nQ�M���'��q~��3R�[�ȭE~�*Չ��+SOs:.���]d�bwN9�İ�e��v6(��"�+�p�ȩ�4���[Bn\�ծ�C���Є������y�'��hzC�/J4TJr �?T֪d�H:D�̃e���0j�J�E�p�r%$�������INyrf��N��'�?yg
.5�$�B�ʼ#贴� 'D3�?��;^p����?Q�Oeh��Ê7�����I;1�P��=.�Z�S4�K?�ܤPq!J�WR#?A'��8~0����͗==ZM��S�N����t��TQ�`�-܈V�t�4��O>�q��'�R��X����.�Uh#
Ϝ0O|IpG�3�D/�OX���Ո�����C?]? LB��;��dG�aD��K��dp{EB�?i,O����Uɦ�	��̗O��)S�'�"����W�Ԙ�&◲s�M���'��JG2WK��:�O�<_��In�8	ڸ=@�ˊ�R�&�'*z�x�5�5����.ԇ%O:��'||X��P 8-�@c�ccӸ+UJ	-��z��Gz�f�)fS��*���$�@���x�ɏ,"���O��}򛧀 �lY�)ʤ�m�0* .kؽ�"O�uj'j�S�|�Y�Y좁[��I۟t��D��K��h"�m6J�����Q7U��l�ݟ���Ο����Țu�h���ǟD�I�\ͻ�,�ulF�bJ�1�$c����"�ܑ`���+6c^[jh 0��G�'l�'q^��b�=P6�	aPMX�Q7Cq�X��`�f㗐2���9vc�(��O�ZO
�[%�>[����RM�alHc�I(�?�3扶7w^�r�jE� ����>=��B��8��P
ʎ-�>8�^~@�ʓD����G�Ik��aR��!w� ��<<�l@Zvo�=E���	ğ�	��l��ğ ���|ڄ雼B ,�bG-�Bm��//G��Q��F7E�rx	�Y=X��Uw���Bh���O1A�° 3�	;=�Mh��O�N�J���@:���D���Oy�V��5l�4�dIȠ��cR7k��'wў�Ex2��/3椌�Ѫn/n	��N�y�a�{�H�S2��4#d�,�7k
���\��v�']�I-1�R�Ҭ� ���?Yp�v���t|��u�ܲ6���O��:�O��f>�U˅�uQ\|��Ñ����3����ktD�jE�V��d��իV>�j��ğ3;ت5��%�%z��H@��+:��qrb�F�(�҂���(� |�����cT��=�v��⟰�	p~r�ϛ )Z�r�M�&ri>�CGS����?iӓzz�s�o��p��}��a
:�]�<���T>�Q�|Î�� ���r�X,�rZ����IOyAH�`A2� ��I�|���2��l)�h�YL�Is��"��W�O��dF�$ `��eE�x��� c���"|��⊝N��h�F@�t��"��S~ҩ� R4x�"CD3[����퓥>�EA)C�FE ���Ø�r�7����	˟,D��3O��r6i�'	��I���3B
��"O
�p�d	6~4�I"�� �&Lx��	-�h��xZ�AQ�Phe{W�f�P�P$�'��x�W���Ҋ���8�Sܟ���Yy�� �55�4KÂH6pH'��ui�\�}���M?J;tuQf��I�t�ڒ��%A�p�$M9&���Ѷh4r�$� ,b���	���#��-����1r��TCBI�O`��"ړ
�PE	C��m���gA�w~� ��'����5�-v������v��Tk/OH%Fzʟ��U�,��a��bئ��5��h����޴30�,��[�ˮOҰ�r�͑�?!i��l�]��v�sȕ�o�84z�b�+:�T���FM�I�8�ɼ#ƞ��fP�\���sdD��?�'Znx�2fW͚�ە�زx��G|Bΐ[?l2a�]!J��*e�]����)gxm�@_�k(Z�3�ԥ�O�#��'FR�i̟wd��^�`Ls��˞e��x��L��Ǝ�b�Xxc�S;*16�b��7?��T>�K*O$�����,f̖�'�]c���Q���؈�M���?�,��9Y�l�O2�״h
ĹPTD�)P����h�4�D��r1��[f%���W%z���!��	w�I��t)�2D���
`�ߣK�hP�+�yrB74� ��R�3d�3/�/�" ��/Rxܧw�XF��'�CWǓ�?{��f����I������$����z��Za$ދ5!�H "t^�kp�߸*V�#�l^�ў�؍����z�{deV1Vj '��X�D�d�O��DS+S`��VH�Oj�d�O���F���+r�T��R���B �dǟk�������{���CBb���)��m���PL�l�&遇�xd1���(�����Y���)�M	���8�B*G�YQ��O	Ҹ�p懲��ဘw�p�G��(J��C�������O$4K��'���<���/F4TA���D?.�n��emAyh<��K�>E�l���� عç�?�?���i>q��Dy"/Q�@&��м���0R-�*]4�x���-P��'���'7$�]П����|R�d��~케�h��H �Sc	9bȤ��C��	+�F�RӪ�;5|H
ej�k��<9B�֓�xCR�C�uWY�#/_7X{0и��V*���P��	���V!o2��<�[�(We��\��,�#�֡���#Ο�F{���![����&BZ����
B��.C�	7�S��� y�<�#���d�"�|����'��	��$�鯟���z>���].~�6��<B8�%(���O��SL�O��D�OΘ�VnM&
��M�
V$tQȹ)�,�j�씈���$d��\�Sk�K� �SC?�Q�p� � ?S�8���ϛ}t�����2y�ڃsu��:#Kז{D���'

��I���v�ɋ�����Oc>�01�X<�y���֊/ǎ�"g�<Y�0��0�Ǭ��^y��b	��ł)�5��|B6^�l�"�L�2�|���M�!n$��e�<Y��W�ٛf�'�2T>���ɟ����V{
]� �(M�0I�a�T��q��'�4%�W��g<�I�ʔ<e{�����yt4�|ғ F�J�8��GOs?6D�բ�<)���V�H�a
iAȹ���J��Xe�BIQ���.�Ti�fʚI�����9�.̨06O��$�'y����@�S�? �h)QoˬXA�a��U�D���"O��(�c�A"���B㎏U~n�:V��O�Fz�O;J�CC �G�Y�����)bd�'�'&ґ�!˔�@v��''b�'��t�',����bђ8�T�P��ݯ`�)a��G�-!�铋Oc��z��*7w��> �. ��>��	{HFIA�MԽ61(��m�h1
)����j�[CH�Q�N��.��Ĳ�I����>'�nZ<�Ѩ׊��O� ��`�]j��ɔR�j���OУ=q�'��-+��@�(����gW�`DE��'�j�ç��rj��g�9@�m���'��"=ͧ�?A+Oh��q.F�o鼤��F5!�͹�	��3| U�B��O���O �������?i�O hv-V��D9�A	l	"��uO�~�� I� qVxӓ*�����nT�EӰ��e�1U;Jak�,B"˜��t�ғ0�򶣐&Q�b���փv�O�����'}Ȁ"A�E78]�be�1��1��'pў�E|2����^ت�!��;��S��%�y�@ӧ;L���7E��X�m1��A�������IZy���%�Z�'�?��O���s+�z���L�59��� ���4���?��h�t=���G+.��)�ʞ/>��%1�m��7T&��/_4fp��!��3�.�փ_d�'m&�SF�R� 0�3��ϊ�.i��E�k��] `�5Wp�<���:�ȃtmS^�'�0���?�����V*��+%�߄G�Z	6,_����4�O0�G'��,X�1	
:)�!�r�'�j�gSn�{c��5;��u�uDǌq;n��'�2�'b2Q�p�O2"7O���PH�*b	p�Y�▏JQ	2�U���?�*O%ԧ�O��#��Ԥ<H�`ؓ.L�y�ҳi��'0�%>�"�X�nm�Q��+�9fۼl��*�/�M�i�t%)�'3X����?����?ɚ' P���V��4�2IE�:D���7D�F�'u&��2�'����I-����u"0����ص�'�� lPjЯ�D��r�]�?i����UX�''���O������y�4k@�Q0fHX
"��<���S#		���D�O�����O���0eK��s��n��y,��RJ<�P�X�
��`jS�s5rA�#�?��e�8u WS?5�Iڟ�������PE��+O z)� %H�[rP���a��'���B�'��dީN����uǋ(;�{��U���\ tn��+a�܉�4a���S��?���8��X?��Пp��1G:6���KY=��Ȁ� �Q�|����<��L�4��,�u��'��d� ]��i.|�2��� ��1Z�n��+���Q"�P�#��6-u���@��Ҧ=��4DH����ug�O�T���	o� s�`�MU���b(.�X7-�g=�	�yWD�m���M#�'�?�R�'l^u��4@�L��+�<!�Ƚ�bC;;�z�y �i9~�*G�'W�$~Ӽ����	��'���O~��2����$D�;A��8��.D�` m�|�.4C$Ɏ��YR�	l�(�d�<���C`�S�X�����ɸ-�h�d�ո ]�t�&aP	~�	��OH˓�?q(O~�D�O2�d���Q3Ą��@�Cj� ��VCh��ʓ�?���|J?��Ɵ�]Ba�b"APM�P0���"O*ғc��Qk�m��$� -���B$U�؆�I�z?�91�@�p���R��8��OV��䏺�ęU�W�>2ͩ�&��!�$9������+!VxSD��!��6\F~���LZ|�V��"^:!�ϱG X�' n�bDڔ"]v)!�$�1%�
� �2�`7��/b
!�䆇4�(��2Fߚz3���[�Ș�"O���`F�
Q��X8"E�6P�C��5KT �J�&�/֘8s��eZ����Js
t'iN�3���"�˓���r�A�f���I���(Zd�3K��OL���m�6o8�)�}���n���ŬE��}k������'�9��ۅylH�!���4	����@�-x�Ƥ0#~�&$	2��r�@ϓ:���jrc)k^�PC�,mg,�Ȁ�7
m��k�B(.� p�5G���j\+�e�XRP�b� Lf�Gȅ摑���3~|"$'��D�eI2C��`k�����H�]80[�nH�v2l�޴Y:M@�xtG�
�!Ұ��E�'�"AKr���דza±;"��Bd���ǋ��ӻ76.urw�'A(�j�,E�m<�O�t�FNԑ*��I�A˾^�DIZG�	'a�HٰIC�\��+Ie���e���Pa��µ��X≌ ���d�ͦ�`��Im���S�xQT����߻fr.�Rc�&D��:���4yB4z�a[�e�x��J��hO�ɒa�'�b�� 7B8�����L$��V.���%�������'9HpG�[Ɵx�I��<���l؃X�$�%� a^0�9��BN�!+�)�>z�Z�o�$?-xh�|rCI߹B��d\=+�����9C$I�Q!��\:�i����'[rN�W�� �|���Q=� �-���i��ռ󦢜#����`U42�a�F�
or�7-`y"m��?�'���x�AO8wi�Z!�L�a^6�����y�kG=@�82��>\�.���f��~�'H"=�'�?��O|Q �+�$~4p�JçYk�	�t�W�,ot�AbIFǟ��	����	��u��'�8� ��=i\������m����4�ԥUV0��4cU�I/���єuE��S&"�&�(OB�� ��W�N1v�CwdG"O.����	C<|d$�q�¸q+6l�GՒ������}�4"L>�� ���@j��M)V��Se�>��5���M���h��ТuK�'xm�%��LùH� ��r�	�ӆ�j��&�Q�3��k���b޴�?	+O���Hc���i�$�fgT�kLiB$�I�q�~�����Of�D�6 �����O��S,��r�Mƀa�dI�NĩY���!��ȚL�b�UbI$)�"���Ov�[n�s����p�z]��@S��p��%���
%��`�;L����"j���'w��jش�:S&��Z�Ӗ��h��� ��	�p"^�B�ʙ�(@B���R(RCቇn������R��e`G#G�4��r�����'�6,��i������I�K�7�P~���;�.g^�z7%�= 1��I柠�f0@=�a2�K�F�K��R�Pk��~�v�O['�\�$�ֽq�f�&��J�9L�Dq�$�K���Y�L �6dˌ���YƉFH7v!�@D(��ēm�B��I�8G�D�i�L�K��ދ	Ğ���hX�B9jj�'�l�E��1�X5@�k�4�ʝ`�pcQ���(ϐk�!ۣ'٥oc��[ ��yϛf�'��'��:s�Y<'���'�B������ŏ|  <*-X-�~� "��(��|�U�͸�H}��N�*�������TU��rP`��/�T�GI�
A�eQ��%YpA�`�I%J⎩����O��Aa�f�Ua�㈝f��e�� ]Y����J
=�V��<�]ݟ�w�L<9�D��=D�Zb�=*>~E�m�R�<�%��8eE�;@|t!�EJ�$�u����'�I�.�8=�B�W�k^�zaEH�@�R��|n 9���?���?iB�����O��;e[��cD�f�����TD�1P��>�iǌ6WO�Wr/�d�`�I�>6�5SWg@�^E>(�W�/+bvr5�߲u;؜�4@��I~e�q��9`B�"T�I�C��L`�ŚQ"��b ��,��ɘ�H�O�m���HO�b��Ge��W�6XX�&�Vo���O7D���	�yr�ɲAL�tB��e�*�M������1	�4�.7��.΂�����5V���� 7*9��ܟ�i�'�����|
S�AR�#�E�[j��A���V:Dx@��C�-c���s�H�bw�0CFe��pD�<��� �q�p. �T�xj�#�=B,QBƹ�n�Fv%�Z�,�5�!�S� ���M���O�D�SlP
&�~<`��D�>��M�4��+lO��:s�D;p�tI %�!�Dہ
O�`:Uc_�@jԩw$�R�#·G5���<�b��������O�<���i>�D3UaJ]Ȃ���d�ڹx��Of���g� 0h�WxP�RV#h4 r���S���>��Tǔ�;w�4��]8+	&��wjΡG
���㌹g�Nc$ ��q��rDT>�r j�5��x@#D�L.n!� �.�d��j��DhӬ�F�Ա�r4���ސIf�/`��	$���Zl!�ę n@#�m�u�����HZ�x�b#��,�"���.N���"��B|�(P �bӰ�d�O���3n"��ё��O"�D�O\��w< �;p�P����P˓�{F��IU�\�֙��
��<��Q��D��ZR"�'���
S���	�<���QG�Z/B`(�ԅ_�/FX�K@�Q�G�BQ[���py��Z ���<� Y 4_>}�$�O
�y��g̴�R5��g�|q��!fQ|Hn���M��*]^�@�S�gy��i�嫵!�?*{�L�RHV���=B��O��=E�t*ԇJ�ЈZqaφYaʤ�"L@��~��'�6���!$��ٰ)�?=�'���S槜64b2�ɔD

Z���
[�8��r���O����O��d����ަ�����d�$�.7W~DJ�k�8����io+d|s�˸d�����6�P�E��8]}��Vm�b���R �[!f�6�'��;|��0!7m�u�'��ai@ ��-�v�C%m�����M�wX��d����4�?+O^���<Q�O8[�bU8�B%�ڥ\w��J�"O��K������B1B
0�L[ŏ�I�O�L�!�4��䖁mdx�;�?�4G�n<PwJ�&R�YJPf.N$vEs��'��/	i��'�b��;d��`	C��y^�i�P����:P�PT�ǧH&	� `h�Q�z��IC�vz��X��ޜW��w-)}8$ՙ�X$0z��nT8F�����!��O��D�W?i���=YJ"pzU&�*��(s�a?i��?1���'���'g���Ks/�a��Q�f�:�)��Px"ʉ�7�N��H��r5w'�C��{#�q�l˓=`B��iC��'���D�8mZ.Sz�b��$T�:1� �0,�����?��ɟg�����O;<$�8�0N��l�:��X �ʪ�DU��"�.(`��ī�2o5� AA�x"�ۛR��<9ᄎ=}h��Y�FO�x��uKK $\t,ۇ���^�n(�B��*e:���I1$;NOzH��'�R��ui��I�9Ov�C /�ZF@9��NX��xB�#<L)E,R�l���+��Dģ=ͧl�Q� `�F�~f2 �D @�����6��O���OJLӇ ��Z[����O@���Oǧ_Dz��@
�:t��h�.F(O\&�@�3��Ҕ,G�_�T��$�?�S�_��4���'rHz��ʔKn�TR�O�d@f�c��
�G\t���D�>L�րY��Wer�fM��`�n���=� *;'I��w�D�Gn�=G�tp�ß|�'�4�"��|���'#�a�6'��c�6�觮Xi�Py�'��@�ԠU�^\��G<���'��8��|������,��i3��";�����$38�;'��.	4R�	ǟ|�����c[w��'��V4M<`#��Îr����vEP�YHa�6%��l�뀓yG�L���td��"��$ĵs���ZR��z=�����+^���-�d`C�#7|�fqCV/l��a�F�[���&�|���JY��'�o�>iᖠFz\�$�O�3�	e�'A���@�%u.e (����A≧DK��遄��	b�&͛MMR�L��4�?�,O��S���A�I�kQ��KŎ ����>b��d���ӱ�?9�Fn��{��?i�O�P�B�敵P��,�f`],+|�b��O����#1pr$�����2�"QP��t�':��O��2l�2- ������)�Z�0�ތ�8�*���4]W"�1q(h�xҲf>�P�2<}ZR�Ȓ_'Gry�c(��p{����"ODctP�t�y��,q���v����bν%}��i@�d\���TΏ�:�FdX|��9
�D6��O@�d�|�q哑�M����#]=��*��V�J�����R�X���'���ȇ̚I6�����>f8L\�v�M�h�$'V�h�� Ё%�u*N��F�x��Ft���5G�(�kZ�=Rb�`T(�3O��i� :��b��JL���I�s�'����N�ɧ�O��)jt+� ����8��0��'���At��!Q�MYw�Ƃw8�ǓD�Q�X���'p����­W1��M1C���K����'h2�'���4B_�I���'���+F�^s��]+�ȇ)D>^X0�٩QEH��)ӵݶ0뇤��e�B�ZU�	MU��!+�#B�t��a�y�p*���:W�d� !�C�*n<�B�=h<��Eo��O�	$�i���g��C0���h�+yP�F��:E�'~P��S�g�ɤrn�	�2���4��#�.{�B�ɬV��T�����r ��5M�jͺ��ğ�k��4�hOp�q�c֬	��vA��!z>�h���>���HПD�IßH��.�u��'��6��D��7c/:m����G�̬d�U�`�uCdߎH���x�)A�{�E�B��,�(O�u��fO����9�;�eI���N}$@�c�ύ1�*�0��ъ�T���`ϟ�dQ�H.��� ��M2f+�0k�2P��
x�V4��'>���dQ&�de1.	�A
��h��	.��|R�x�*<���kM��ҭ�4����'�6�8��Q�<TmZ�l:d�P�Z&��-PZЃ��b���K���?1Gb��?y����Th�A$�����U�U�`qg)Z7�>]��`A�%
N�pR��7bPu���	2E^(Xv � >�@�1�JB*s�0�{%�.�6]r�i�w�6��ď-O�`���'3>�'�9�`�#7Q8��Ԁ��o����'\�D`��@Č� 2٠aB�'�� ��.A�{^�I������7(�~��'0Nay�k�����O�ʧ-�;�442�uZ�L�q�yP��Ϫ i�@��'�rHYc��s@P	]`�v�τK���YƎ�h���u��+�Ƀ�	�V`@��]5Np�OR�� �z�,��Ɔ¯G+�yXVfQ�<�-��5H�I��p�F���!��5R�d�x2)C�?�#�|�������
�1w���P�"��<.�Q�'�<���/�&�㐯��}�d�b��Q�`���i�87b4\��PS»(Л��'���'@ވô�T0���'���K�,ǘQ0�l�D��;/sD�'��\0V�ǖ\���E�1P��:���+$T|K�I$���f��
`�B��[�)�X�G���]�|	�K��w�a�"��.��O����Ċz���0�N�)�H���_vĠT��,J`�'èT��S�g�I�-�f�J�	����Po2H|BC�	�3*�4K���<��!��lǂg�b��˟��4�0O�d��(M�<@g��/.N�C2�O����v��ǟ��	�d�ɏ�u��'�:�����V�cjT�ŗ)zD�y�� �%��:�gJ2-�)�� <ILuD~���7"n�11���:�i�1��MШj��~�I��>=���T� �����'i�TzE��+W�
gZ�*��O��8ړ��'�KY�(�f�R�Ҕu(����n�<��_��D-���_�!#*h�&_�nꛆ�'��ɉ-�L0S���7M�j��YWc�)`\�l%��q�Q�	ܟLDm�⟨�	�|ڥ�w��3&��)8E���T�ˤ��V܂q���D�om�5Q��I�:jz�nn��C�Z(Hl	$�S5)��:���1Q��R*Q�z��E~B��!�?I����D_�x�������@ ƚ!�qO,���^y3�9�G,X��,��.��~-��DZ��ݚ���8p^Ɖ���C� ���%��O˓Af�	2�?���j�TN�w����j�vt:����,lʁJ�A�(�d�O�AB��+x|\�,��P�|�3��Ӕ��U?���皣rr���nO�%�����-/�$�&"���iW:�$��h�(U�|Rv�ͥ(݈Hxwk����BS�c�	�^!&���O�}*�t�? 4�iT$^ 	f�R\�s��J *O�Dx�(ƺ7�t�1a�@�Af�$�gQ�p�bG��9�X�JǶ��4B�m�1(w���'���'��P��N �}x�'}R���ӑ£f.p�p��_�5gty��
.���c%$J�TZ0���Nl�����1:���R&4|(�J������h҅[e�f@�"�VP�ËR�du�U'�
e&��a2��|��g[ |E󎈜~`x;�ᒸH�|l����4���I>�Ĩ���>O�q	��>?��\�J60mZ� "O��Qn��GIV�q��?7��w�O��dP\���ԟx�M�i��D�-�Ч���:eY�mPD͢=� �O����O&���޺��?�O^�=K'NN�Ӽ2�̓ lvL��ۨ�xR�C� N��� D.����$�=��%�
�'F���U�z�Ρ0 �<K�hi0.��?���'m� 7B� R����#%��	8Lj�'���`v拁J����ŠA��ي�{2�oӸ�O��IR$ZߦY�Iצ�
�G
]}R!��
ǆ"��%lڬ�?Q�g�|Y@���?�O:��P��3D���6ꗶ�x����&�y�7����Z���#���K�'8�Y�f� �Z�� �,��;���"_�ȡP��G)2	Zb@ڧjJt�S�l���|���?Aӕ>!�K�5`7P��"'�$���Eq�<����{��1�I[.md�j%Jt�'Wў��M~��B�R(>0��P'��hP��5��[� 6�
��ݴ�?���򩒲2�6MS�yd��⇉\!6`(%	*+J4�����T���K�R����F�6I6�ڄ)Ҹ>X��a��Aj�t%즄3P�V�3�Hz�(Aԉ'z����
\���}���Ga�D;���s��=#bO��?�ƱX�ߋqV��[�_a��4Z@I:�D�.�2�0��I �4�$�
8��sEՇ�!�����|Ct�M5��(4-��#{��D{�O �<yu$�Nd:�s�C�08�����	Y�qFp7��O ���O*��j_�L�����O���O�CV6WsҴ�`�Q�VZ!��X���r����� ��t�1�x#�Mj��0@㛫F�� ��]Lu�u�34L�B�����!���TgM5D1�ĎR��X�!�v(�Q����숻M>i��П�>O*i�%)F�.�Tp����&z(:��u"Oڔru���l@̄�G@��V�y��>��i>$�XD��8�vp�'�5s
�!ʄ��k@pt�W��?���?1������?��O�i��\Y;�t@TM^\�ځQ��^��x��k�Up�i7V���������p
�'l�-r+S2�^�[�a��}(wm�2�?a�'�69� �� �|��dPaN���'��ԠU�P�9�rms�@�@�4J�{ү}�ؒOe��������ݦ���K��h���?�*x�`X��?���XY�����?	�OB:y�����*����C�U�ZQH�y�bp~иs�͔^�J���d�A�#?�q@�20jt�Ǆ��H	RhX�i!����X;b(��@�!y����e���^���D�C�i��I����d�@�;���u"O~5��ʢd-�y+B��i՚`��
O䑊C�!D2. �Fm�"dpR$G�,�ȒO��xR�Ϧ��Iʟ|�O��|���i]��@���N�B��W 
��z����?����e �qa�[�SU����5(\�ЖD�����	�����$��A5PL��F�#-��'Ĵ���4p<@H&Q�V�pabnK�s�pz���	aT��(0@�7wj$ꂤķ�M���;��I�o1�'��i dnx��vɉ�#�{"V~a!�$-W����Ǜ/�x�Q2~_B�F{�O{��<�'a��F�Q�B�X�Z�a��j�6-�O��$�OX�2E�ՍX#��d�O����O7G7p{*ux$�G�'r�)g��xSv�
� >?ѡH]�!���|&��ҀY�Q�����$�4!�49aJ�7	aZ�0�O�|CL�~&�P��l'��Y��]�Y*�Մ�x��'-�3�S�g�X�nca�
�9��pu�N'w�C�	�?6��p���՘�a�M�u$�'�T"=ͧ�ē3d�{��g"(%�/~^�48���y�dQ6�'F��'���xݡ�	ӟļ}+��0�e'��uy��*���RUf�w[@i���H,�2+�0U$ 1D�-ʓ`[�Q��-��Q��i���@	&��~_�ɠH�n��b	�`�L��C!ʓI46dc -�3m��)�oe�d������Hr�������!�&��!���t- D�`�%���21��
Nה^��QbJ9��MkO>Q �ޚ!A�v�'���#��(p��&{~|9q'�]>t���O�#e��O�Dk>5	 �;dV��8��\�kWh ���?R,�xP��ݝC�<Y��Vy�hR��ǝRfQ��P�`ѝu6�XA��`>�Sf�ɜ{��3���m6d��B�3OS|T��M_�����B��_�����_[��/T�t�׶4�D=�����!�� �M��CI�T>���u�_�rX��B���j����
���8	)T���p�rw,��<�P�|c�'��6��OP�Ķ|� ��M;��H9B.08U�E�\nV�q@�
�s���'���`EZbP{�D�v �8�F'H+l�8 SS?�R�G�a�8እ^���\�CO;�ϧQRa��A�>{/�D֪'fЬ֝�T�m D�	4=�����K+��33��"~lT��0�x�^5�?���|����ˁe��D�!�2j��k�aˊ�y��(i�L�J�!_d��#���4Tq֣=ͧ\�Q��k1�1,h�b��Ҿj���XF�Φ��&�'P�'yX�鞰dSb�'������3-B#i���pf�Ӥ@+��glȲ/��
t��U������:H����#�I$}rJ[5�b��e�π@�:�`��C�M�j���X�jú ���݆Ac�丏��>�CJ̄��XT���6У<,�OV�����(��)����n#&�AAO�0 �l@��%���� �D�2�q�/W)}���O��Ez�O��'h�E��gY {�ԝ�"A��b�.-s�&��ps�Ѓcn�OZ�D�O�$����?��O=-�f�)���C��ȍZY�uz��ř�x+V�zP�AN�CH�d��*~��
�����n�J�*Q.>B���A�U��x���V��~BL�\��9�$�?5G\LS3����y2��85��̐Ə�,`�<�MT ��'�`7m4�$F�YU*��OޛƄL�w��xA��Har0�Cc�7L��D�O4y���O��$d>98Dc^�;L���"� �l��q��>"�i�*�,�^Y��M��*�Y����(mp��y�L���Fl�D�!��@�!:n��񂍐r@��!��[�'%�i���?��O~����L p��Q���%6� �"��2lO��@�Y�P�bs��/ �
O��u��B�@���˒�Ь��h�rW��Ġ<��n]:�?ͧ�?�(���y�r]r����-�{6HX�%�,DI .��X�I�O�l�"��Ə7��{W�>/-
=R�nT/��@�O�����%�M^�2#�Rn�b�N<���?�
y	3](f�f\�� E7k"�0kY�9���Rf�[4k���Z�!U <Y���H=*-�'��#���?��IzӦ0�,H��R�O8J��)P�"O0Z�i��f��p�B)y�m��ρb����C&��Vx�@�ڝy��e'IA�Nޘ�
��'E��'�B�<ڌX�P�'�"�'4�;6@�)Z�o\�kA���VN�X.D�b��*C�A�f�i�&��Cj�V�b>	�P�Hal�&G�}
��×��#B��9�(��lI���v��L�t7�F).f<1���@�0�ƬH,�r �����O�t��=�Q���3�a0)O�A�����`��O��;�Hv(<R��]8A A8 $�oj��ȓV1�D*�,V*<P2���L����?�V�i>���t}*��G�^����*ot1�f�N	���ˁ,Q�-N���O��d�OZ�;�?)�����J�8�e^0Z��+�O��lP��bH(]7�1��H lO�u*���?�T�I5�+��h���ُ3p�"��rr<��	�/���Xkk5�<�&	W+WI�`9�h�O��.���'�d��!�5o�.�s�bˍ�	�'�x�&�()mf�8ֆ�v(��{��x�t�d�<�M�N��̦���M�,{"�1rÊj��a�Ԝ�?1�I�}����?��O@��S��[�^L�"ٔ0��i2���w}��*�ÛX� D�朻C �t�D�t�'G؈R7E��o�@i�!��kO:�ks�02����Gq�Q�+\$�>���Ra�'�.���?��O�&�/9,�%�f%��K�h�`�d�OH���҂u�.`�&k\"eARL�q��=á��\M��f �&GXZy���R4f"�xԤ�Of�-D�����|B���ߛ@�6m�xu���o֫-���I�l^�G�����؟�Z +R���IGk��Hb4���X2� q�D���,�\�gl��_h���넻��3�8(HMD�lt����X�f��-��wШ���'r!H�M��q�,�I�*�
q����x�$U�?9��h�6-I� ��#�$k2��aID�?[!�$�>C��9y�	ǑQ�}�����sSb�G{�O� �<��%�x���3��?a�v��4�;/R@6��O��D�O�\|�
�$�O����O��S:]��E'
L�E:q`�P N��=�4��F�Z���k,��T�3�Ӂ0
����';Y*�o��zq�"�)c��4ʵ����i��nڮ0Z.:��
9]U�'?�K�lD��y�(��*��l�y�nȀdƊi�B�&�Ԡd�Oq��'r�x�l��H���:@\���%�o�<q�i�:�x�D7Iϼz�$�g��w����x�C5$�Mce�P5_6m8��F=��p` '�,�d�O����O����O��Dw>E�c�I�n��3�@�*SԾ���uä|��#SB�(S�+Va�E)$ʄ�Y�Q���f.�� ��;���V�&�a+W s���2�ƻDn�i
�VՖ�$	Q�4 `l:w`W�55s�q �š.� 8;%G4{l�U�2'�O8�$$���'!2��0C?N�R�[w�X����
���S�? �$C�еv��\�Tn��^��S����Ц��ITyb�4.Ɇ�'�M�ꗑ���wm�.>"��!�#ȍ�R�'c$Ȉ3�'*�>�R�@���(]^��d��+���F�@�E.r�"%f�Q��5�&�/[m֜X��1�(O ��A�v�AtK�2`
�t�P
�Հ�'�G邱q���)q~�����(OPe��'�_��X��cr*[�DF�p9��;�K4��|؞�pjW�),��G+�2�p��ì0��ò��#NaV���܊rL�����%*�(8��My�8��6��O��D�|ZbK��M�B��Nf)��oM�&f�iɣ��(���'�Xx	!���
�X��3)҉�~*���'*hl�[��qv��R��	Z��$����#ԁ~v�*B�ĵDg���
s�'9N>��N@@�V`D���0z�H$���H�O�	%�b?	b�H�� �(��u^n�90�:D��֪�IT��c�'��M�H\AQ�7OجFyҏ�H/��{���∓�J��4l�؟T�I̟�c��,<D��IɟD�I���V�dYp�_<;5�)%�܊�.0Yh5�(}�P�S�CC�� 2.�H�'q-=i��f�`�`�;SFR��(zTF5Bk�u,f(:���|��(�V�U� ��XO~���Y:��.+�4�y7�ґLk~���A�vj"*J>��ٟ�>O,S��N}������b�� F"O8��ɾu/�!aD&@<j�^-��>�5�i>�'��8s�Z8[v��(ň)m�$�j��=0����?���?1�_w��O��dh>)
g#�+Y��Q�0���a��;��Յ�$J�ej T�-C�	���+k3Q���խ�v�LI��$ 6!Җ-�CƁX�laː�K.B�Z��XP���ͷXd���!��lIm!888�e�*4H찑�'I�����D�l9�IJ�0~�p���!���>����ׅ�\)���4%qOP�mZw�7F/Z��۴�?Q�4?��TAp"�(��*u8�h�3�'�r+�3"�'�����b����"QWع�/Aܴ�ʑ愱^=$�YI�2uSa��_ɰtp�j:ʓ�~e�����!���Z�G1l� p�����Z!�T�RK�(5ء�栎�+Rȩ��D&ʓmJdL�	��	�c>m��/A=��yqf �}}�C�y�r�j�W#*���Á�G��C�I�9�:��A�\�G��JU�\0�)`�CY�$$�	hݴ�?�����6|�6�Ӊ
̒�
W�J�6f6t�0�lF:��I�4R��N���e�:�@�2T�>����gBW�� � �L��"��&ΎE�	Ε�ē%"D��$	ׇm��ä�
\N%I3��,|���')����Vn³��8�e�V�]Ѹ9%��Qv�O�<'�b?!�ӅA�{�E�����6���E�(D�<�! M��X���מ¤�0F9O�DyR�ΑU��ԡ��K�$���JעJ2��m�۟�������橜�-���I՟���������c.a�a>a_r������P�4�[�(zBY*��I�A���i�O�~�'s� A��OB���OZ�0���d�);��<x� ���4q��7J,A��K�
��>Ũ�b͛�y�"1J�-S�nҒL�<P襩�0,\'�Lȥi�Oq��'UnUYd+�&\P�r$�ɻY�V\
�'nܴzN_�%��2.�`2x�N�,���4�pO��XciŴq�����~.`%�B&���Ɯ�$� �H�I蟨��6�u��'X<����r%�; %xy�4�Ï| ���@S )G�s�D�m��L����
&{���1#� �(O�����é/��!�e��K�LE8K�Oxꐊ���~x��7+X)Ǝ��ǀò?�p��>����� Ӥk����:h�����{��`�I�p?ib-�2=�H 3�X� �����Ak�<��@I}����hGj�< ���^���|2�ʙL"�7M�Ol6�_�&P�bV�V�33�L���q����'�RkB-"XR�'��i�m�&�Q�˂q��I�%��h�+B0mM:�J��'C�����V���;�ꃧ|��d �C�.U�hcw��%F���i�I bUl�CACEj�'�$1���n��!"-�@��tq��0���
��`Э[)�h��[�`�2\�voW1~�2�h@ň�y�� 	7�Ε��1.�@H'�i�R�'E�S�+�@o�a(�P��i��y��B�i?n�K��?�쌄�n�P��5B}�!Qҥ�Z��|�`���鞦lƶ�3��X��n�Ys�Ƿ�'j6m����SV�f�,_�ִbU�E�,���r�O�|�g�	O�Tk2�.�0�1�IC�I"
\��d_W�)�S�䒭01��%�^�����*�C�I�+m��LB<b���@
t���4��XGyR� 0d��� y�z�#
:3dl�ğH�	ݟ(��
.6�8L����t��֟�.:*�mc��b��p���=o�"ң`�.���m{~���u�Kz̧L~"I�-�O�m+�k�e�������.�F�z���Q�,)���N�Bd����-3�pm�%M���IC�'��ϻ!P΅)��3DV�Q�ͽ{�9��>�dͼ{���L<!��фd��й����t���Fp�<��L6v�@<;P+Cs6��Q�\l?)�%摞��M�)� �1�U:
*`�8�� h��"3��u	ê�͟��	ßh�I��u��'��6�B S��¥cn�̚F��0�*����M�C��PJ`ŤC���BQLO�E��2��¾�(O�P�N��nR�+�4m�̍�0�۰m���!�ĳ;���ҷ+Q402f�EH�����@�%����SX�c)ȁ*�v�����M�v��O�Q��	�F�>UNU6w+`�Ç����c!�O�O�`�:"�v��c*L�4�T9R�D��Q%����ʦ	�O�ԐC��`G���+7A��:���&�'���Q?�T�aqŗ|�"��ȓZ{��`�Kj)�CO�F2��ȓ'3
���v}�5���ם�$�ȓ<U> �D��4�̑sa��6�ȓ���ȍbg0%�e;X�bE��>l��c��D�>	���#���j|��w8����-�c�,s�maR��ȓ"J��P���]�|!Q��!����> F��r�I	�#ؠS`~X�ȓG#͢c��8l��h��p:���@�f����h�j|HR��%96��>�^uYq	�	��9�0m��:���K@H`��/K�0���:^줵��-?��c�d�<0�h���;,�u�ȓ��ݸ2��J���/�4x����t-3GJ�(W˾�Z0��&��ȓ�"U#���~VY�&��'*Ϟ\��Op�h�����H��B�#}�Z��ȓV�XH�GIXl�da�a"2\}��6��=x���t��K�Ȓ`���ȓ ���#��< Lҝ��̚Tf���ȓ���BM=h\h�(�J�R�tɇȓX�@-�uO$I�2��%��.E
��ȓI�H����/@s�]���ˤ_�>���.00�
[QRћr+�"vs��ȓf��Yk@-&�yS�hX�y¤�ȓnt�����Mo���0�S?����ȓ0�>�qA��I�F�T�T��ȓ�z�sc��?+�m��N`�>)��IE
h�GۨFC�Ű�)�>pL�e�ȓ��Y3H�'6Z��� _>�>��ȓ~�b�!W)��I�F��,��:�����B.E�G,�?��Ũ�Ɨ�[����ȓb�v�h��O;8b�VM��TȒ��ȓi�*!��*��4;�*R�\�J��ȓ����e�����j�	K�e�b��ȓO�:��6�N''���B�OY#d�쁆�H>���֮2� U�n�u{d�ȓ���ڔ%��/ ��4�ΗV�5�ȓDʴD�)�ƨ������ȓe�"���E�{J��M��攅�,X�Jq��'|���Y��ӡ�4���1p��e�����'W#h�Z������Ä}�P�m�� �z��j\}C��
0�h�'%����d��3v(�͘�l&t�������V�<i�aK*� ��B>��۠��I�<��f��]x����ѽ�q;թ�m�<�C�P�#��@��W9~�~3�� j�<�Q�[�����������Nn�<��a���p�G��&r0��U!@�<7�,N����2Ժq�`�+�,�D�<�w�T�@�*$J�ϳ �X �%fHA�<�2�ĐO&����Z7c����/��<��J�c,�h�Rׇ4y2����T�<9�S�U�6�!�ʒ�����LR�<A�n�?<��	�5JY�j�E p�IM�<� �!�0�˃X�<����NX�1t"O�H�b��<_��(a�CP� t�ܱV"O�t���R	J��Л�(X4P6I�E"Or CB�-\V
['J�6خ$+R"O�<!�W�q����d�����"O��y��.�� �m �L�8"�"ON��f���}Ȗ��m�K����E"Ol�`5hN� *��l�h�ā�6"On0�b٣/3����>Iw� �"O�ة6�� �^�h�$޴aș�p"O���-vB���ʐ9[D�a�%"Ot���@L�_�L�T�ņ?`��r"O.�8��۟c�.�f�/A�F�� "O�L�l>CJ]��Ɋ3~Vy2"O���%d�!<���e�,?�rm�"Ó��&�3<ifqA�:[XD��"O�!�"�����E�n�C5"OF���,�n�����Y�@��
w"O8\"Ȝ/�8���*ϐ���"O`�i���%OT���ț�{���9�"O��A��U�FQ���[p
L+�"O"�r5U�GctE(����iX�R�"O88pl�#pR�J�LM�'�JQ�"O$��D�Vx
�EW-�b}*"O^Y)&(�/D�`W%ϦM��3�"O2t;3&��X{rd�N�:�:4�A"O��؁��y�I�bM7,�*�� "O����VЬ��]�2�*�"O�e�㣎��f5Crő]q�-�V"O\���Ҿ1������,
I,8��"O�m
��:u*>$�c�
7&.�t;�"O��W�
�W������̧r'���"O
`bt��[����*5��"O& �'�#|a6� �m��E`�"O�hzS*Kߢ���k�x(�"O�e�P��&���IfJ�G.�ʰ"O^E�F�H�~���Xhӛk�t%C"Oe�@CݖH�̫�'Ė*:&؈"OrQ�/U�,�(d�2L	�B�"O|�7P�gy$�f��r^��k"OrXj��
�>h�AA �[�� "OK�.�����M)P\��93`\�y�e�ͳcͨB嶤���;�y�	P"l�5��p
x}����y��� @S���{��E��A��y�Ѧ(���p@]6_ޘ9I�d��yB�J����a Є&�dBf �yb$�vq��p�<\��D�yb G�7#��e^73Rtk�T�y�R�8ҦxK�o�R���jBo��y�Ɗ@�Რf̎M��4E��yrBɼ.I(�"E�-��!lA��y�e�#m�R���ѳF�lΊ�y����F5
�D��F�Z0�F�y�DΖ�QӇ��R��s��;�y(�UY�w�:KѠp��Q��y�I��s@F	{�&B��!�#�y��]�X�0��h׎'��Y�7��:�y 4G���Y��Lmpᷡ���y����F)�e��V5J��)���y�L܏E�A �^�D�u׀>�ybB^*��,Y�ʞ�5%� [n	��y$�.U�ԸK���*0��('��y����G^�� ���p��tr��)�y
� 6M�r�8a���*g�L��hC"O$<�e�.2f� D�^I�6"OzQhQR<C�e*�	�X����"O�3�j¬"�vl�ʁi����"O�| ��[�T��� m-~XI"OB�ra��4A��8��D�:�R���"O�)�T'D�+;������|�UB1"O��c]��B��D�D'Id�!;�"O0A�7dM8r�����cɕ*P|�3�"O�Yj�
�qIN�a��@?0n���"O�M�w阜$���RW�	�2m�A�f"OL)����Fʠ�fľU�)r"O�r��uw����EI�@D��a"O8��+�-��Q�s�K�/��R"O�l��&�Q�`�Z��
2��0 �"O�ՠ�  ��$��舕r��9�"O�<"�ێuC�X0��H3w�x��"Oȱ3U��](���K@ܪ"OrG&G-4�x`#�e�U��\r�"Ot��GGɲFL1�<�<�`"O~A褮�4Z�49k�l�)��шC"O��c��A�,a U�K X�0�w"O�铅C�fl4�5dZ2	Ćp��"OV� �DKY�D��SD�J��A�7"O^u�pn��@��P���R�&��E"O�AmŊH0���s �r�2y9@"O����>4�KBL#b��,�"O���l�?C�� �N��e���"O����	>��)�3.��xM>ɰ�"O�ac�X�O�rГd��oFdp�2"O�-����G��i��E 
ۚ1"O�lZ�^�,,4�ӏ�5��hٓ"O�i�Eʫ�x j����I \@I�"O���a�ԨW�F��$�i�"OL�YRΉ 5��2bX�uy��8�"O�9�fL�7 �j|��͹
�Bv"OU�KwH@��@�	J��� "O܍����&<G��)���~�Z	�%"Oܙ�"ȕ�o�0�iO���85��"OQ�v�\��\L��$A�O݆q��"O�5��E?[@D3u��R��V"O�X���]�����Ċ�>�0��"OH�x���9���@� 
}��]ɓ"O�!C��B<U��d�⯊��P�q"O�с��H���"�9�"(��"O��
6�	{�,�i�L�#���Rq"O��oƅoC�mb�F�f��#�"O�xK�E$
Ȟę"E�"~�!"O@��3�"<�#5�m���"O�h�5�V�P��5HH#l�ʳ"O��J�
ŴPR�'�\�g��s�"OJ��w�Ū7,X=�u�;d��"O��15��J��A�a`P�DT�0��"O�$��,Кs�"������"OH$yס�h�Ȑ��0@��2�"Ozԫ%�!D,�}�l��JϤ"O䝰�\�c8�PbNӭ;%�Q2�"O�]���N��xz��E�%����"O���rHU�p����aӇGPPy@"O����
](�A�u B����"O���e��R�ŃT�L26��r"O| ��cU;HD�:5NP�qf����"O�q��P,v�ԩ��H�T���e"O ��	��=��-kgMD%!�􄙂"O� ���C�ۓ]!ؐ�#��fԞ�0v"O��Q�a����)�� Z>܂�"Or���cԙ;U�x��ɑ�+U�ia�"Ov��u�U�ws �Ւ��@�d"O����	^��;f�4I��U{""O��i������~�T�*�"O�z�]2$i橀�E˪:m���"O��Pk/MV���%�?	 ��"O�S�MM�~�aFg���X�"O�u�0��8���#Rl�*�h�"O�pl˗p�PBv	[84��"O^| �jG9a|e���A��q�'�m�C��`*��ƛ/��-�d"T7$Z�[�A�<3:�8d�#D���'��";¼��h��%d�G D����J��&
b��#�D�Qy(L#�$9D�l*UǞ�A�Tk�朑.J�c�+D��r���Kx�!����4Tʒ���c,D��xԧܸ;v%bve�ax��'=D����������a��1�d�x�7D�� 㨒�O��P����zX�uP.1D��kc�D6=䄵:q=Z�՘f�,D�T#��#~���a��ZgǦ��G�)D��S1AL�G-|ɛ���_&T��b(D�0�˔�8J��[%z�2�`3�9D���a�E�M�"$��Rvp��&D��¢e�d1r6!�~�n���O9D��A��A�2A��6!:XH%D��"Ҁա\��	����6h�d��J!D���C韗�Ta�QC��Pl$[�#D�P�k��cl�9�VB�4OD�(bQ("D�p 0@�� ��ZA�\��YŎ!D������"1� �$�I�-��P��+D�h6��	�!�H�-q���P�)D�!eG�����d�P��sXB�I�)CBP�bmW�\	��� fՠb��C�I7E� ����X3
��V�*<I�C�ImZ�a�Q�2d�ȳ�ߚ�B�I�F� 4j�#>���wl �S��C�IuZ�;P�W���j2��<4��C��4~ �U G
9�47ƚ�;6�ȓB:4x[�O��$���5n�����F�D��6c�#?����$W��*0��O�(��Ƌ/��@R��MBJ���� ����6��Q�J�C��ńȓ[~Nq�G p$�r��ޑ�ȓs)2��p'� `���+�Q�z���ȓ]�~ ��ޠL���sw#ښ_R��ȓ�ԭ�f��d����I�0�ȓA�5��$��صÆ�۷2� ���4$�rv ��������P��XF0i��εH�1�Ć&D�B�/-Q����;k��Q"�ߥUDC�Ɂ�>X1ɜ�GZ�)���\	
ҲB�	�0�4�c���Kچ=`� \�C�B䉳wx�����+}�rx�o_�(��B�I�O�Ȫ�&_f���sW��`�B�ɁFl�"&B��"|²E��WǐB�I�n�h1ڇ���=�L�t�P�~C�I,]���!b�>Ud� 9g��7O��C�ɖ	Fs'�� a�h�4A� df4B��!uB�;�Y
tM<!�D��$2:B�Zer=��
� uj����B䉳H�^�#q�.�a�E-̞u��B䉾0�*���` j��(���էkXC�)� �H�-������S���I�"OؼR�^9�pB�Ch��"OԴ��A@`.=�$k�W�ܘ�p"O�Hp�č��:�y�
?���%"O u��؛y �"J�-S`@��"O&D��j��b���*w��7n��HK"O��j�܁A2Np�1�\��u�"O2�s �-"^�%�H��5��"O,�s�ūs/R5�d+�>-a4p:2"OJ��ń�,=L!�K�Q��$*�"O�hH@�H.t�4=*�鎝-�	�"OjP§)�X3�Hh�'��J]�G"O� ��J� /*�0�S�dr��(F"O��)��D�4�l@hA�˴�a�"O �1�g||4�� ̦[�0���"Oi�R�FF� 5kf@��F��tb�"Od}�w?
��ˣf��F�`"O���F�
g��L�K�T*g"Ox ��@X��U@&CI%8���"O�����y �	��@Ͼ��m"O���B��J�Y���
��"O<�`�A�2P}8�RTņ�9��"O�'I3;Q�0I�D�6��"OvU����9�LY��^29�(�b"OƉz� �Ĉ�a�	����u"O,���:��p��
M�K���!�"O��:��T"Y���ٴ	M��0}HQ"OV�ɗ��Y�l�	�h�+�D"O��@�ڷT�U��%O�QB����"O���'�9]���7B�4 �h�"O�8�F쎷T�p��G�7W~��"O��!�Ά���R@�gb�@��"O��ؓ*��bRЛ�ACU��""O� 8�#�RA��Z�4 �"O$]�Q.�#�Уg#�,l����'"O��7O�+b�M&��$�X�3"O6�+s��\.Q�d�P%Q�ԱX�"O���D�o�R��1)֌�ZYH�"O1;��Ǹ`"�AT���Sքr�"O|�6�8"Qb(`�k����92"O�xZ�(�h����ϋR~~1k�"O<��u��5gA�9�CDLW� u"O��j�T�|}P�

�V��qP�"O^�˶JX�e����F���It�pq�"O���U���_���Ɛgt\@�"O����W<9��
D�\�30��"O0�5 	0��Te4>yz��"O4�A��]�0�����E�to� �"O&��u���	`(pF�Q�T<�%"OT�4G�9/вl�C�B2U����"O*$�c��q�
y·
]���+F"OҸ���7@�.A�FK@�3F���"OP���B\�s��86��A�]A�"O`�Ҁ�R<	"E��n^(:�JL�"O�pR�M���S��RN��Z�"Ox���ؾ	�|- �d��Z����r"OzX���! �����f�xyp�"O i�a��B�Zp�u���ص� "O��G�N�rV|H��%�(?f Q"O^l�Ʃp�&H�ӄ��JB`���"O���>�`��3)�)��Z�"O�X�TiĀ,�V��)����a*�"OrT�R%P?7�H���"m�ptH5"O�mp�&�
L���'�3d��H��"O� ���7� &
�i��C8�,I�"O���v�; Z�a��Gԟ5Hz��"O5��j	<P�9y�h	�"Oܕ��A����u蚩~٨���"O�|�Mf}�Ġ%�Md�V��1"O@XY��XCk��`�T�q朁 "O��`���'_�h����2W�BP��"O&�[7��-A삄Kgؿ_����"O��dL|0�H+f��p��"O��@U�M�c��4��� �585"O>L�th@�s����K�3y��Y�"O���Pnא\ltA �#L^|`��"O)#���J�~t*t�	�T����"O`�����zS��Y� FV���c4"O�PIХ�7ڭ0���X���t"Oȍq�n�~���c�!�����"O��"P@)t�$ɳ�B�-��-�$"O�ld�в|,��Zp�@�B6���"Ol���Qp�6ဃ&�)�"O`�5�_��8��V߂h�W"O�}u�ڌ6�\08 $�0U���3�"O\�z%�(&��습
�6z�V�;"O�iR�j�l!"ѐ�jҗz��Х"O(�7��J6�arHF<M�Liz"O<�#E�D� +��۸@& �ۥ"O>H�"�' "t`K�bFNu�lI "O�s����c d�$��D���yg"O��9�mb��T�_-�
�2A"On��D��@��b��S�R�<���"O�ŧX����G�:Ɔݚ�"O*��]WJ�BW�+'����"O��R�f��sF���J�W��Y�B"O���@K��rl���.dޜC�"O�E�Wh�|��U���C0�Ȃ�"O����#�!T�����)`�*�"OF(�1�R�q� ՠ���P$��"O�k�G��Z}�a�rH�@�"OHP�Wlݮ?�`i�@ì�""ON�S���W� 8)�m�3� �U"O��3� ���!ҌA�^Lx�"O$��W�Z��	 ��M�\=�"OP��vd�V��б�n�u��9�"O�u��b�v<��w���a��X#"O�M��N��^L��TW��v`��"O@�(�8��kC�2�4�3"O��*0���f"�����%�@ZE"O(`��]��1f���1��`�"O�ݰ1*��C������ñ_��t`"O��sA*L�*�6�s,�H���"O=��a�~DV����Ξ>&�P�e"O�TGÛ�f�BR�Z<5��"O�pZ#	�$?L@���%dv���"O�Y���э����!�T�@B"O�hK���3 pu ��IA�μ�"O���	@)Fv�x�˄e�f��7"Ov�rHN:���*�<�M3�"O�aF�PظI���!��$��"O� �'�Y���@c��&vv-��"O�����
ah�$���*f� *�"O"�2��� O��Xa�Ѕ2���"Ox)���$&�����m�zdq`"OR�yE�B����6�
��,q�"O�P����TD�4!I�r9�p�"ON5�w���m�C���c2�q�R"O� 4�b@o�>(İ�a�O�%<0ɩ�"O�xJcA^�z��K�%�>H�l��"O�a�/#�\�3�d8Z�L��@"OP� #��$t��۴��[����"O��+�"�+V+���2�9D� \K�"Of���+�n��D�Aܸ�ΙT"O ����}:*��Ƌײ8��@�4"OJ�p`�S��p�SLMz���7"O�$p��T�d���&�qՈU�w"O(q�Ê"�l�D�+�=�"Ol��0H�<�&����ձlP�)p"O@�M�#"��!T�$)�D���"O�8��oZF��D�'��9�`�"OL���S�Y] �2fý+���"O�� �.B�Js��"��O�JI��"OZ�An�LN[n֫����'�ց���4_�z,j��MpD�[�CW(J�"W̖1ID�4�ȓ|H%�7�Ėo6Y��M�Pxل�.�FY��"��[:�bR��&"�D,��#~���%�4j��� b���j���!�S�N�N���i�A�p�2ل�;�@9��ɹf��0��=���ȓ ,xR�VHZ�QjC�,�̇�M�*m1��B�<BH23k�,����ʓ ��b'#_�sAB�%�*V_�C�I3<䨰2eLD�ʼ���=U�C�I�9�`9�aD?
P�bCZ��C�	60�v5�!�>�`�
A�Y ��C�	���\c7l�0
����b�
rXB�I�Yֽq�KU�b��2b�^B�I,J4��u�G'��(C�R�B�	�6�^P��	WR�tAa�C�B�	N�"�:��L�����ρl B�	�p�#3Ȃ�T�D�ңc%j�C䉌p���4�[�'��(�J����B�	0�0�RVH�-������>	�B�+1,�PA@+�[32��G�{	�C��+�xkd�K>I�B���$]��rC�	a�:캃�߰DD�2��i�\C䉫:�^E�R�ӯAM�|#7�DI,C�ɀ\�A)�ٜvRV8S��X?[nC�ɔx��}2��M�g�-(*̉Y�LB�I1]ņ��'
�d�����VR�B�ɶP������HI�Ӧ�G�OB�I�L��F&�f~訉ՈC1yҔB��.<��RE��A=���2+�-�8B�I$VJ��!���Q	��醵6�NC�	�bx&$�ʖ8�ȠjTǤQ�B�I=iz �u��|��hK�JC�`B�I6y���s�U��
eH���!btTB�IS�ށ��	L[��de�A�RB䉺7��e����j��k�NF;Y�TC�Ij�(���zLL��Q!ʮd�vB䉊w�X�I#�M�%�F�{a�+�JB�	�2G��f&�9
�xe�4��.�*B�	CJ���ٙ:ܰx��-{�B䉖i����P�
Y���r�7;ZB��ipT4��	�+g���� ���L.B��A^�P�@��.�v�x6h� 	[ B�!Z3,�4*�.B�>����
{��C�	�j����'�h#�@U�V��C�	� �|���nשs���Q$/��C䉟4��9�)܍��!����I�C�I#&����H<��)J�����C�)� T�s$-�+�.\h�K�o���"�*OJ)BR���8:���u	�'(HAP�n�溈Iau����'��AC�䈅�,��nJ-��'`!�1��7�� [rH����J D�����зKTV䣖�ڋ{LI��<D�Hh�J�
���#�
W�3t*!�7$/D���s�2��I�J'Pi�����yA]�I�h���%E��Q�t+P��y2l8<�\a��GV�B-�h1���y�k��;C1�`� Ak�$o��yr+L�h��08��:8���TF�yr�ݛG#<tzqB؎Z�*�3 ۋ�y�m�&^ڍ�3a�<D^�T��S0�y��J2x[:���K�Q�6l����y�@@�[�zA0A`ق~r��d�ѫ�y�!X �H*W�B3���;�y�H�Tǐ1
����kr�Q�L��y�iX/e��p!�eR1�r�{�'&�i��<j�RT��N�A����'�`�(�"��N�|�Uiڞ	P�Q�'� �r����A�5C��\�Nx(�'�N-����[Ж�qw�� /v,z�'����?	��q�+� �l�
�'F�48 a�&6�����r�
	�
�'v��Ui˳��)�Ĕ
���r
�'��(��`�n���J�:c{�X
�'5q�S�C�E�	AU�8\�	�'L �eD63f*�#^���@�'(ejr�K�H���c�˭A����'��Xr�-�]��`�BU�w�V��'BD�X2�J����嘨g�����'
�fG�%�QI�W�����'+d�ⓦ��&)��J��<��:�'�hǥѮA8Fŋ� �wa��'1���ǪE�����D*��(�c�',�Q��
Y�Pl`�iٵ.�թ�'&P钵��3F�PK5��LP"�'J��� Ŗ$c�
����ޞh��'�Q�C���i��\�4mч|��d�'.D�@��Ǔ l�	��%ȺmΪq�'�r�á��B�d���.k�
���'R�8�����n[���'~RXx�k�I�҄�L̨M-���'Dv p1�H_^�Y��E�3��4y�'�ȴK�ⅥV����G��#��H)	�'E��pG�G�V�&��ꔺ�D�@�'`�PCgJD"o���f�������'!tp	&C�	X�lPQ���,C���2�'���I���8���2��qL�P
�'ӎ�z�_�+
�X�B/Wno<���'�B5UN�w�}P�5Y����'�)���>���FCگc�9�
�'��E�A&�8���x��Q	YԔ 
�'�C�H�3T�&t�B�Oc���	�'���1!�] z��d�R�}l���'�L��5�� E븍��$w(D���'�"8�'�2;-Z���aH=rKv���'��|�ф,M'f�x�D�h8z���'܂TCt,Kr B֋^"1zT���'S���Qm��ip�x+���+�4��'X���MM�|�; K��[3T�'�0�G
"Ft�!�-#��$	�'k]C��ȅQ � z��5���(��� L��� �utإ!w�O�x���"O0	�.�:b�@Ɇ�M��Z%  "O
��nϿ6f�M(�DE�H�X�"O���-L-Zi�ij`��(x�~$�"O�0�1��$@���V�%��"Ofp�aK�r�^��F�Vl���"O�l2h�L60p
�DI?7L�lhr"O8pzsB	_����U�E�i	u"O�-�����[Z��7dIE>�p��"Ol�Aadި7� �X��>-�$� "OL-j҂��X��$�B�u�A "O|q�7�F
"��رj(Jܐ�"O�3�L!&l�,� ��0"O�qBeGڱ@X���t�� �l\ӥ"O�<�r-�'�:)s�MQ� ň|�d"On���ьպ%kC�U�ڰ��"Oyx��ťo�*,����
jH��7"O<X@���*3|�k�� Dk�u�"O��a+P�8�8{�I�!j�Dx�"OP%�d�P0dd���G� 6dE"O����� ��	��Ξg+�왆"O�� F5<�
$�c��}��"O6�ʔ/4L'hũ�� �;�Z��@"Op���\���a��1i��D�"O���OD9\��ۄ��1!2z<PT"O�ĀP�C�P�Ӊ�]	j�hҘ>	
�u�HM��b��b����Հm+��ȓj=<,Z$��*L����a�#4?�=�ȓ	)�� �!x����1�̥8VR��ȓB� �6�T	.�yBCo�#~	 ���+���ɀ�߾�δcu % iq��A�sB�R�Ny����6����H�(�SP�mJ��Ԃ^8^�PԄ�n��+�F�9�ޑ�3��%�D��ȓ�ąX6�޼@B:�h��i�z!��u)֙�`菸)���B�� i�ք�ȓo�4BR[I+���P��! 7dI�ȓ>P,���� ����� `BЄȓ1^r�rb�3���ƩНT%P�ȓ;윀�&E�2�������:��T�ȓU�>0Y3f�^\L4"�L�P�ȓf�{�Ek��*��HǬ��I��ĨB^ʔ����3�����N�!���G!�|D��7��مȓ/�~D�c@0hY��"����A�D�ȓ\��a��8�\mZ���$y�ȓr � �B@H�$�bL�N܆Ʌȓ#�Ɯ��3t:�Ձ��ށ7�	���xyǐ<wK|a��EI%T5���ȓ&@���&^6�jаV�ܫc72̇�>6x}�֨�5/X��'#�@���X]�w���W����.KFȈ�ʓp�t�v��5 %��fj vvC�Ɉ{Gh�`��X�]��]����BC�	?i����F�o]`�j��L,9h$C�I�vZ�%�fEI�Hɒ0See�wʤC�I�5�~=��$^���`��ה*��C�ɋ(��|�Â�&}b��5�6��C䉶V���0Hۦ||B$;E!X�5jpC�	�d�LX� ��+dH[��
:#�B�	�h���$�эVpХKw��-U B�	�i��@¥��p�}��T�c�C�	�\\t0�#.\(�٢�W��C��#��8S�>�J=�!�W�(�C�)� F`���:pAb���K�v��B"O��cC`
9*"�
��&<���3*OVe*�.�R�"�2W��y�!(�'v��b�f�6�к&�H`��x��'
��рn	�Gmȕ���%fv��'�F(xAiB=hz�ɥ��H.�9
�'��`�5�H�pt\�pŉ�2X�'�I�J	�|�^$R�iɺD
�j�'���3��Y��p��8.�ݰ
�'50��cY<6�<��P��,9��
�'xZ�aro�4J��Tڗ%U�;�X�A	�'�����e�^%���B]Fݱ�'v�%�7,	�zSژ���/�U��'q�0V��u+�mfF-+p~)z�'�h�c�G@�}$H�mUcT��
�'6�4ʦ.��C���ƈH�!x
�'h��q�OċR8����?�f���'�f���� �!z5�u�Q<1�&��'~Zȃ��̈́.�6@i�n��!�0x��'�.� ���wӬ$P�H6�H��'�4�Q��Mo\��'H�@����'��Գ����Tr�����[}F�q�'�ݑa]C�
x)��D)4�
�'��F-kt����"�  @�'�t�4j�>I��5kgE7|�r��'���&<S@H`��ϐxJJ�[�'u���!�Q�5$ٲQfW�jk�;�'�=A�(Q�1��3V7_��<��'�����:7�hp���a4H���'��A�*��:M9U�ٝU!����'���򁞕+��zdeN┠��'��4���$`��,��c��F�x�:�'#֠�mW�]��8у�K�=�(��'mf�� cB�B��$J79,����'�Q:��(	O�� �c�(3�|a
	�'��8��d[~f����.�:\��'kr�У�.��Ei3�K�,����'A �d|�S���66���'6�����F�LMࢌ���,!j�'8 �0ӥ��2Y̒2�J�=M�	��'mV��@�*O��[�e����b�'�h���oD+$�$hRCN�|:�:	�'0�+�f�"Y���A`�]
2���'�`m�d�f�B�%����#�'�vx �cM�E�P�[��}��Er�'�zlb'��|��t @�{�����'�Nu�'��#(�Y�CJ[+m�� �'w� B���F�xcaS*a��|Q�'�И`��JLPB����!`�1�yR͟fR�s����E:T!�!��y҃�$�0xxCa�*�8��5*4�yR���+���*�V�dN	�y����f�VssɆ?(Vȝ8���y2"�0�����Т�ѦE��yRa:"�N�q!�S�/�8����y���?=�yY�H�(`엕�yb�� tmHT$��,�D=�H���y��B"_i�[��B88 9FF�4�yb��4-�4�a%�~xZ�!M��yҠ��n~�	F.
� ���h&���y��Ȑh�FE��K=v��HR��<�y��L�_oDM9��J�m`.�#��%�y� E�nԪ���ϔ�kΖ����yr�Y�
#L0��	�4/@�4�%җ�y
� ���7h�m�0q��M[1ZV��"O�e�MF;g\$Cu,дa�F�C"O������(�V�Aa�C���Q"O.���(U;!"�h ��i�n��!"O&���{�$�)G)[��q"O��xD-G�k�,Uɥ��+P��	�"O,ő&��Ve@�Gѷ��D"Ol�#�G��v0���sI��-�\��"Ode���!{S�!��0��ӕ�y���~��EǬ�*�1�R���yRQ�H��l'c�9��M��y2�ҭm��[
@ O�h"����y2$ʆw�)µf�	���"�B���y⯕�N����'�4��a7�8�y�K	w��bWl	�{7��Qp��ygQ([G,��Ɓt��$��Ǌ�y�MS�m�t�7akn\�j�F�&�y2 Ը]�|Y�e�f�1�`��y��o����dMY>���ɕ��y�K@�&^�t��n�)�݁w��7�y��̺B�|�����1�ݹFa��y�w�t� ��ќ|
x�F���yr�P;��c͘.{�>�H!�B��yr㜧8`��H��{-℡@#S$�y�	�8^[hyB��q>�Yeޕ�yr�NpO�(:3�_%aA`��*�y2eҢ!W6�!#k]�M�>�	C��0�y",D(bX���E��ӏʉ�y���u{���ï>
Ő=�dF�yB�U��LT;��E�	��rtM���y��ɸ�b�2�%� ���G�%�y�D�hi�xcdo�	�$��'���y�m~'����\�gLb����yr�b��$��4t���#���O#~*d��K�v@��]�p	A�c�|�<��脚D"iq!�&W��prACw~¯,�S�O�$@���'�Y3ϋ�$�(��'h�(�퓟%T�����+0�l҉{R�'�����cH-45��y �Ĝ1�\`�'`�z4)��(<��gƘWCʽ{�'	�e0�z��t��ΛHE���'a*<��ː0�
�I׫O>B�R���'k��h�Ĥlrf�z6��9�l�"�'v|���E�o�<��%	%��`c�'�x�1bO7�(�a���$�p�'~�Qa�+�,�d0���f�J�'ph8p�FW� @i`�k�D %)	�'KN���M>$��H��y�����'�@t�ɕ��ś�N�x�X0�'��ܻW��&��=�P5o�h�'U���gB����ȶ�Vfr���'!6�Z��<��Ʀ�u����'�8����{ܺ�[�"W�a�Hu�'�V�Z�-���� ��f�4a�����'#�i�WM�?#Ր���Ǔ�D���'"D10fD�>���R���;H*�*�'�� #d�);��0K�8r��a�'��R�G4b4���j�7��|�<)$'��.-�P���i���ha^v�<閎�$C쀓�mصip<����W�<qs��u&ȼ@��2��$(S�Y�<!�k^'�	��l�
�\!RD�Q�<9�n��K�:�s���N�����L\M�<��M[�
��4�$$EC�����"I�<� �q���
_����U��'B���"OV�CI��ݘI�@��#O-y2�"O:q�"/�"��;`Á�Mν�a�'���H�'�v��nR��0i��l��Rʐ�s�'P�=0���:c)&�� O�"��h��Ą�!�pE�D��G��`�O�
[`e����y"B��]Д4ɒg�=n�Q�J"�~� �� c��}j NQ�Ah�H�"���l��P^�<is�A�*��&�vBV���DFR~�!�+�N<���39���'�\���T�d]l��č1�M;SƓ�/���RC
�0;4���!l��X>B�I�V8 �˄iL��p1c~>L">�s�N�[t]!S�"�S$gkp@ql � B��#oϝPC0B�I�#t�H�F�ڷS#Mj7 б+S�����ۤ\ZɧH��R2�\��:��� �	�qb�"O`S��D�5e���3��4
��c�>b`���	�N�zyc�ل�f�Z$&�	Y�\q���3�y���q���*F'�V� �@�kA1�y�I-X���qAA�+9��ɷ�H<��Ox�V퓱B����隒}ժ��"/����C�I+|�ЀW H��Zi #ݡ6��əRj���?E��A�N��RH�YLi�Oղ�y���]��)��M�e'�|1�N��y� ��k�o��] �$���y�n���DЈs�۳� �7B��yrI�����ח4BɎ��y"NA�Hh�u��q�������yb�H�9�I�Wa
^F�C����y��7Ӱ��R�WX���q�Ͷ�yb#~����� �Tr�H�7�Pyb��-}.Q�Ԣ�YFn��D�{�<	�L�y[�h���&G8�"�Kw�<�����Ybd�ZVh6�z0Þr�<��n�5|��a ±t��4�e�Rc�<���+m܈I��j܇	؜�&�k�<1��P7Q��}�K�T/�`� �P�<�s�؟SL���a��;y�壅
�N�<����:G�Ba�Ï��2��Je(J�<��Ȍv���5$X#�	�SL�L�<�j�An�:`�|�\���c�<��;?��T%�$N~"x����^�<�#�Ĩ�$��cn�T���De�X�<ɤ�$���ڶ˞B�Vd��Q�<���p}�h�aC�"���YVI�<ѷF�*��i�Q�C�Q��)�5D}�<�"�4�H@X&���-r���pe�{�<Q%��6BT6�8�c��a��C���v�<9�
� r��`!&��h�t�W Eo�<�b�ŎV�&dKN̏4%� d�<ٗ	C�k��4��nĴ0��a�<��H�X ��Ґ�C&�����_�<�����%+�iP�����]�<�t�݁�:�{�&y�v����_p�<q&AT�2�b=�!��[��i3"�p�<��ÃLR&����^�����V�<	�IL�
w���G�O��PC�k'D������*W~��vD_�V9^�V�?D����¼X}��Q�Z�%Z��p�(D�,���T
v,�0�,��<˵�'D��	 (^;���&,x�)+3(9D�4��b�4*D��AѢ��|��8��6D�����5_P�z��R5Ҹ�(�&4D����R ����f\�_WlB�&0D����Ŗ�h�|u�#�gF��0D�� ����׈�r��+�HlaS"Oj��6LY�t������b�έ(p"Ov`"d��u���j	�/y�M"O�� "��vJX�2#�e����"Oꑱe���L�0`��ktBZ$"O�`Ґ^6]�j�����,det �"O���W�"O��� ֪�>Q����"O>���_�d��53�2A��%#"O�AA��P�P��@���):r���"O���EI�{n,u��̩b0R�C"O��ɑiDP�^�zV��*#����"O\L�e	�' �(b�
ҿ�<��"OF�)�)g��b�Đ;J�#r"O�,�G�ۃ{�Mҁi�d4}��"OD�c�1m�4��	]�&��E"O>��L�sРr�A@���Xt"O4bB�TР��Lc�J��P"O6xI�D;,�t������t"O��꣯ùl�"��G늬'qN5J�"O�]�EK4>��ن̎Hg�R�"O�<J�9�H�
�7oI@��"O� *H�o�	���DqA̸y�"OB}����'A�$	�J�G��!z"O���A�4{;�L�0jt�
��'f��\�l��!��'P�6��Ze��4A�zT�b"v}
���Ox`�1� �DJ����4�����SSf�r�ƒ�~�A�l�/�) 3嘷0Q�LB��K(�>�Hp@6r�r����U$8��E(��dKD�Jx�(C��(.+�"<	�e�ϟ�Ӗ�*l����%p^�h��'Z3!�p�1ߴ�?,O����<y���ҙ)X�����<��Cl�y����ⱦ]]5Vh7m�7M�U�.�VAwӮ������i���T,�un��w"S���=1��xR�i�џI�z�شJI�%Y�	*<�[S@�&��Pw��$l3ZH�+���(Ot0�cǌ�U$k�=|\��3���'9j�t���	N����ea"2z���M�$Zt|���dM$Z�Ҋh��I&>�m��hP��K�(X'C��a�2������������R. �2����1?��x�]z|�VE���9ٴX�ֻiH���	8 �l� �������dCϦm�����M{����D���0�4�S��F\��s���m��L��fåG|:�(�Z%>���%��'k�ݠ>�S�?��M�/�@L�S�M>k9 $B��5���AQ0�$,U��k�Iޭ:��$��(��z2D�|�1lw��9��?m(�,w��q�Rc`Ӏ�9��'�<6��Ey���������P=�`1`�G ^0�S��x8����O�OJ"?ya��U��d��c���*!�L�'�6�Hͦ	&������;A���S.��5-K�\[���w_�qr�'��| �̰y���'3��'E�����l��/hL�R"� q�<���ށJ���@�ƈ�ؓ'M1 $�	�����b�i�6XM>�&��T�\�ا��?ߪH��R�<��V	Cu���sMCf}:�h���d�0�X�ƃ%<��La'a�Ƽs�ޅH����'e!h�ԘWH�F}��?�?	�i��Or���O�s�� B�*�\���9�o��?ܤO~�=�|��4v�xT;bG�-:n�ٳ�S�p8JI`�-c�|5l�ϟ�ܴ�?���:(�r�ʥ.�j��,j&���}�"�:��L�q���+<O ��x}l����G�v�VM2�GՌp�p(;���:0���$�9ӵF%\�(�����c�W�'|��ө�$Z����C���gܝ�-B&l�@t(3W�� �ǝ����c͌o�'���2�cR��V�ְ,?İ�p+�f.���@|қ��'����<�?�O��L��I4} �$����&34�3��.$�D��cH��q+ǛR�x�hdį�0�e���M�)O:x��#�����?ɬ�΀��b�2=��s���I��cs�9@L������h&0j3%�P�r �G�z�����6/��x�	ݜ3�Đؗ�] 2��)�5 'ʓso�Q��P�#��V�;�Z�ڦ�
ֺ{b/ӓv�(�÷#�6IM�<�v�?��=��`�I1<�D�����~2ݴz���X�����q^�Bd&%��'��O?�$�%;?��V@��,M�U+�	����T�����
�M�"�i���\�HV��B�/d1�G���jf8��O����OF�O�b���ӯ
   ��     y  �  H  *  K3  c:  �@  �F  FM  �S  �Y  `  Sf  �l  �r  y  ^  ��  �  (�  k�  ��  �  ]�  ��  h�  @�  ��  ��  ��  �  ��  @�  ��  ��   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p͓��?����3&��H��� �R�ѧ�
R��%��	����J�7eBr�X�׶�yb���U�Lx[���l��}��ѝ�yś??_N3��F�s���; \��y�@_�-��L
͊q@�_+�`�G{��9O�qYAl_�|Ҁ:%E�g��PE�'��	؟��Ŗ��Pk�3a���ޞR�C�:W�4Zc�ćI:Thw���MQC�I<d�����C����oȔ�C�8�t�a�JU�`��Y`OZ~l�C�IpT>4h���z"����HX�ȴB�ɨ:ghU�k�[^KX�_�:���"O�6c	;���c�K�g��h���`�O��8�Ш% ��p�	���A
�'#�D@'Z��𤁤~l0 �'�`Da$L$RUˢ�̗q��=��'@���fbʁ���%��uJ�$�HO`�=�OO> 8&�ؚif���W�]���	�']d+&�A�x]u*�(P<����xr��"~Γ"�t�K�<D-B)�t�B$B/����IB�g�:�3����!���90h6j��	rv�d#LOD]�3IP�>�%�6�ö"B��Dgӄ}�O�b?� �`!wCU�*�I!c���h(�:"O.���b�L��Η�8!I��x2B@�O駧y�dP%1�jⅨ- �v� �!���y���8*љ�hW�x4��2��P��'��})ƀ�i8�� Tƀ'>`l%R+Ʉ,F�3q/$ғ�hO�ӿ$6l	�R ��y~�#��H�!��S�'��؆��I�0`0���'3�H��ד��'�
u�F�O&���0�)�ހ�`OXd�CЍ1�6��v!�(rlrC�$6�S���'p ���ӭ8�2���Kڹ!���
�'9~���KM>�qT�4���	�'�����Q `f�-��Э?�n���'i<��sJ�5Z�tA�fI[�<Ydޱe^D��/�%��a#2�z�'
�~rÁL������8	㞁:u�����I�o�Ad��7Q�~�R���d8�C䉯�ܼ d�|S8Ă�N�$t�B�ɘHr��C��#ߖLXB9	�	L��8hv�}F�$'ڧR���Q5�>D�(��O�@ D|��i�0'���;D�4�6�Ak� �i���]�~Y���:D��YOH�u.X��UC�5:���S;D�8k�&�&%�x�ɒ�ڪ-��4c��9D�r��:C^�D P��<�p�@�,D��q���"d���*�<K��pb)D�$X�'�|����j�#f,��%'D���b'Ú&.��#�� H#�1��!%D�����*y�7gS)��ٻ�-5D����D�:8$�ڠkQ ��"� 8D����O(H�ʽ���i$�j�)*D��H��1l���EM��i1S�(D��i�C�v����B�Ťgj��sh9D�ԩ�����D@W� �& z+4D��&E�"[�	А�Ի����	2D�p��g�Rt�T*�������Ñ�/D�����1M�
08�P�g,V@k�d/D�̸%��!Z�eYsd�(L�0�c.D�pX���
fp�#S�;+ل-�#)2T�4[0�Y�C��R���b�(�H0"Oh�Ц�V��z��I�" ��`"O�)��C̆K��%2R��:!��	"O6��t��1Y�6��I�t�*��5"O�Փ�-�2%�亥LO�r���"O�+%ِ+;�aF��#_�.h�R"O���ț>f2�aL܉{��ձ�"O���h�&=��JŬyz���"O�|��kK 4j�I0��S�Dx��""O$��@��"6�1���Zp�8;�"O�(+�U�P��	/ �	"O�����K G��]��i]�p�l�)�"O���wh��� ����5�$H"O=�� +�H�O�R̪M�"O�8�(�Θ��!��(��"O�!���E�,����=��$%"O6�q�E3�~ɩ��C/.�D5;�"O~���˻}T�S�-� �;"O�t �)T�f�BJ�g���"O�4ȵ�K��%8Q��f�j��"O�5�G��V5Th����)ή�J�"O@�k�,B=t������B��ؑW"O0�÷A'M�zKã�&F���"O� �$+ްc�: å�[�N9�A2�"O6�7#�"�<�3$�9_�:!�'"Oč�b�/�d��^',q�""O� L �FBS�JF�e�.#j�t+�"O�X�2Tq���*bCہ]���g"O�T@ 1U��D�L?L���"O���ጦE묈�� ؑ!��D��"Od�
��Wp�Fa�Do)
��,�r"O�����&jj�-`-ٜP��-q#"O�ee��[0�(rl�"ϰ9c"On��Ǐ�+o�T��J�	�>DxB"O(��f�1N�~�J�*�D�,�S�"O��*���Ӫ;�|�t"ORy�T��8�i�({��R"O�)��eZ(pNa��)�8Z8*&"O<��F�R�8chS�]��C"O`i�̉��(8Bq���]�Q9�"O��R�M@$lkJa�F���BsIBc"O��wc�3d�ЁBA�4�(�1"O��S�,��f�l����6.���"O �:S�T�&� PZ5�Ё%�ik�"O�'lX/��gH0�]"O�� �O�(�hY�A���x�v"Obu��K�&fb���O��s�Ҽ3w"O��Ac�a����୚�d�!��"Ob���,��z�t0�pX#9�pS�"O� ⃆�~������0E�&d)�"OveȦfY=*�*	b��L�<ʚa2�"ON�J�G\:x��� ��V� �#r"OLmFj�,Oz�<���X�P�zQ��"O�i[�c� &���ӫҩ�x�@�"O�`G�� u�2���>k}�R"O"��$��K�Zi�N��XO<�"O<T��كNed�a����0K�P��"O9Yw���&ա1��NG���"Op��
�/��"�@"A�2��p"OJ�a4eȵ6� �Q�)#���h�"O�� 
�D"���MO` "Oƥ(bgO sk�13�[-JNz-�"O��@��Q����M��J"��S"O6�1����I.�IQLH/ ��P"Or�J	֞@&�����R���"O�ijt�@�lcj�S�*I����1�"O����j�&�y�*��.��}�E"O���/V���Q�Ӳə�"O�|Q`v�y@CgT ���ȣ"O�Ԋ�nQ._��xf�-1���"Ov���!�"
P`�{AK�7 SF��e"O��@��;$hYaQ�W�jD>ic"O�cw��2�J�#	�<b���"O����Eכ	Z�Q�F�L>O49ِ"O�Qq�+�4𒩀�K�1D�0��"OX�%L�<04y���Fs�
m�t"O| 2��/07���i1�|"O�yx2�HN�Vr�J�p��D"O��S��fS"0���ܯF�!"O|4��j6-&�r�
�@`�d�e"O�l�`a�6J���E�ߙqY��pr"O�]n��f���rH� `��}��"Oވ��,�/�,�˲,N���9�"O� ӵʝ�o�� Ц�\1t�u#�"O���	^4������f�Łv"O���J3{��z�뒓/� X�q"O���V�J�H�.��"��"���`"O|%	w'[�?sF�f�+(�"O��z���KZ0��IU�7
ʁ*"OvɲAۊ*P@��3(�/�Ye"O� �X��ΐ���:�G7r�i�"OF��Ĵ,8a3��P�M����"O^�1���l<@�"�!��@�"O0��D�u&�|����!�v���"O�ՑEl��{�b����@.�Q2��'��'<�'
��'�r�'��'�z�`��1:��:u��_f�9��'�B�'8"�'2�'��'5b�'��͉��μ2'�(��c�Uv���'��'?��'22�'8R�'��'זd�g���I%�R%c�Ƣv���?���?����?A���?����?!��?��e��hZ�S᎑2q@x���^*�?���?	��?q��?a��?����?Ʉ�:lrJ�w[Ь)���?���?����?Y��?	��?���?�ŉIo�D��NAz^ {t'���?	���?���?a��?1��?)���?yǇ^�f�`�i� �Zh�UU`��?���?q��?����?����?I��?�6�՟y7ʤ���Ƕh�V�g��?a���?Q��?y���?q���?���?��ݸO�^�%V#�@l�h�!�?���?���?����?���?���?q�/C�Cg:D1��O	}:�,�����?����?	��?A���?���?����?�E��*L�*���� �{XP��)���?9���?a��?���?Q���?����?IT�ɲR�]B�EW7LP囔�L��?����?��?����?����6�'≌V�f)H�gP�PF�T�4%η4���?�*O1�����Mc��ýc�f1 b� ��A��	>����'�86-%�i>�	��M�����	Fp10�R$D�S`E�jz�f�'��p��i�	#�H�)�!Y�'SM���l�8�e�@hJ�"�^��<����;ڧ��܀HZ�!wؽ�BJ���)c�i ���y"�����ݶ�\��_%QGR t`
',V�mP�49B�8O�Ş�8Iڴ�yb,
����� F;6����yb���9vt�m��1B"�=ͧ�?����I��;�J�]�h@r�Q�<�,Ot�O�]o�W�<c�xB�&�8K���zՌ�?�$p��g� ����M#�i+�>!�OOӲ4��l�s���
 d~B�٘i>�8pHU��O*���������3q����%Z8�ɍ"��L�'}���"~Γ-Ϧ��QGЧ�$|��&Г[b��Γ>R�vC���D�����?ͧByD�rўY��[��f����g`�6G`�|��^�{��6�)?��
Z���g�c����d
�!����F�`+�T�����Y:��,%�tE����|�J�)��y��[/\`���mR��y�O��t��Á���aQ*����/��	�P�B�����A�����8�O3��m!�(�̀}!!���+��X9W�2I(��M�6>B��h��E	(�2t�9>��������n8���$]+xmC"O�*2I��^-UY
�Ѥ�	UF��pB�����s7�}0���M���?�����Ƒ���_�L�x�S�gU$5� 0�S j���D�O�hsD��O�O�)2��X}��0٣-Ǆ ��<q� ���M`�@�Hx�v�'NR�'^��f/���O~��Аa��xAs�ѽ,�`)��̄�j2��՟4&�"|��PCԥ�"gK�.����S�
z�49r�iEr�'���:!�(O~��O^�I��`�ڳ��Q�Ƅ �hM�\��?	�ΰ<[/Ot���O,����q !��"+d͸`g��Q8��av�6���R��.������<�̍�+P�ǥO�\��|L����v�w(7?����?���?���X����6bM�I���WS���)��?)���d�O��O^�D�Of!ZcI�_K	�6Eϋ$�=9���i��B��,��ßH�������{�,��'"��y�AN��x�����n���l�ٟ��I��x$���	�����'oպ7���5!X�S��؟t��:��Z����|�	ٟ���ڟ� ��z���'oB�9�lл씤sG �&�F�@2�d�\��?�D�O^�d_7k���!�x�@I.\ ��TE�*b�d��Ms��?�+O���T$�n�S��X�S*\\0y����H?z�p"�B��ذJ<����?m+|�����!M{��<�X�B(��<�&�'�r�[���'G��'c���',Zc$��H��yR�0:-���ش�?��9m���H�j�S�'-R�`ʐ.��zUFxS��\��l6�����ß��	ڟ���ʟ8��y��h�d��G�n�m����c��7��5u�%���䟌��H��E`g'O�b���x�+�M#��?��lw.�1)O ʧ�?��'P���7�S�	�2Q#�M�R=���6�IA��� J|B��?���:�<��D��Y��P�f��&�vq�R�i��
�(�O0���Op�Ok��.z�X�­�
p-p1,���'~���^������@��py��'X@Q �-�d�ab� ɬ���)C&��e��	����	���<�/O��鱏�7a��쒒�ոA�@��Sm�����(�I��T�	XyB�_:m;�S�qj�ԢCDΘ��)���#��ꓣ?a���?)/O����O �S�T?��&m݈�:��3���Æ�RUn�>i4��>��!�+6K����j�Q>�*fB� ~��7�[J�A�s/D��R�f�-'��N^�dR��)�m��̠��X6v���,Nie|����p����NR�'���D��&�t���M���K�>#���9�m�=	Nuғ)K�X�,<����.pPfY<���+H�$�0`xPh�Q�� d�Pe^A^��pfepC@��t�#AJl�W�ג]!�љTc��s�ĳ�
v*$�����O����O�ܳ4LX�.=�|A�b� Y�D�Q�ͮ|�JuR�e�G�	�޴�M� 	�([�dLɋ��;&��X��ApZ=@"`PS��`��˶p�t���7-w�t��几1Sq�G�O%�*qs���"V5�%���V~��P���'��6������r��?)  H�8t���Ϩo���Ђ��<Q���>iƄ���(�h�	��Rd�Ċz�'~#=�Ā:�?���J�T���Jܾ�H�D#��?Y�e΀��%I���?!���?����.�OR�X&E�|���\�:ɪtS���3<$ne�7������Q�F*?g��ӱԟ��D)Q�Ř'w&��l{�	���X�2=`�҆��	�2�1f��!+s�F�N�$��H`�RVY�$\���'p�DsD���w�~ܹ��I;'|124�'�<]yG�'�6M���<����]�]]�m��c�6kЬ{W��gR!�D�O���ж^UD=
$I%b6���s$�O�'x�I�b�',�	�x�@� ^w_p�Y�b�"�H��%.����'2�'yC��TR�'��fԸ$W�\�2�
B�l��i��-�]��_.
Ć���	�')�B�С�Pn�'���	5Ǝ��ɹqlPs���
"���t�&`�,�F�HD.��M����K=Xr�O�}���'DF7-�]RjT���"�ܡq�\k<pn�͟<�I�����ʟ��	A�S$�'��5向�Q�V�26�]��M,�L��8�1өUN4���I��|�(Tmt���4r^�\�hkF����M���?�)�Z���-�>���a DDR�� ,۸+����O��G:8�Z-�q��.-�tD`���b� ��4E8v-�Bʐ>T٪"EŕL��%IT�6�d7����G�.5��B�x�0%1w�؏Axx�Aǐ�9���F!��J��[��'��~d���M3a��4�'�欑p���}��X�F�`?F�j��'��O?�ɘ#��{嫏pO2Q�5@4Q�"<i�Ńj̓u��F�k���Ĕ3K��T��,�#��X��ɲ/�E�۴�?�����`�P���O��� ��й9Ƨ�m6́DZ�iw*���тs=h` B_�xdE�%!��8@%�)����*��h�:��ᄇ/^��pgď22k�=�G���@[�'��C#$�+�gۀ_�q�g�E3� ��U4��R�V�-6Z�0��'�Z7�������I��y�T���@�qM��[��˦d��<Q���>I n�Oq�I���$+Ԙ�[�MR_�'@"=��'�?��V�UH��zףQ�u��K���?a�\�PXɢ �?�?1���?A��t��OV���9?N8I���"���U*߰R�$QR�_*\��8"��J�8��ݟ�P���
�'��,���O!]U���@:F�������/n���[��_�.��Ս�����2@�5&�Y��IV,���F��"Y	A;�~��<5b��ĝʦ���4��'z��'�Hm!w
KN�6��M����'6���j�xB�%��!L�slƃ"#=y��i�"S��&dι�Mc4NF�?���)�F Q����?��?��Ƅx��?�O@�i[�f{�d��v��q��qq�_��!k�Q��lZ/	Ar�����'�(OD���N��;���k2��7�A�0�M)dL��ĭS7]����c�R�8s�8�A���͚v�2�DZ�R��r�����p�3ֈǔ?�(=�}���OP��?�ʟ���w�ʉ��옷hQf���cE�'Pў<JՇ�8���Γp0�
W���pܴ�?�)O��������	؟|�Oz���"�H? �0蘳灷(��p#f�)n��'B�B/[�Z}�pD?��X�P�7�|�*%*�vl	!"a킀j#*�4(Zbb���9_���� "E�@0#�̅�,��kO
�g���X��j��z�򤈪W�b�e��n��\�O��9����s�:EZ��քZ�@�Q%�'��O?�d��i��F])f�JQ&��B�(��dO�I�j4��&�g��Q��]�M����"kir�4�?�����Ů�>���O��d���� �i�
O��� &z0f���9�ů�� !V�1�߉3lv|YQO5���:	hk�s�:������Ҩ�SA�N8���M���|��� qޑA$�ƙD�:p�0l�f��;���0� ��ʈ ��'�iC�O��|3��2�)�矨��[�?�RH{r��D�$wM2D����T�p�t����'3?Z����/��LP��4���W�]l�i�P�P0ɢ4��-j_!�����)R�" S���Ʃ5-(!�ʺQ7��󂀺.�f�A���?G!��
�AH�1<�ڐ�0�"{!�d6��!'��1�n�ׄ"�!�$�8g�yCc%K;m� �(���	0�!�R�~D��Po;fz�u9���\!�
6lQ����GD1cp5 ]S!�߀`���Ia	3ObT* ��m!�:d��
��[}8�q+D��{!�$Þ Kͩr�[�t���E!�$�$.�v�[�J�F�r`´JND!�� �;�DC��f`4@L7n��	��"O�u �+����b���G����"O���S�[)�ȵc���wj���"O �+���I�\��`ҩ!r��"O�yR#�#:���)�,CI��u"O�p2�C?s��0���t9zm�t"O2iX���kމ����6_9�s"OnY� "�9;��țVd� X"��P�"O�A�T�^�N^tT�2$�6ED !�"O��xF+�)A6^Qن(}��<I�"O~�1gǾp�%�Ӈ�7 ̙"O�UW"
5	+ @�l��H+(T9e"Oȥ��fX(Q�����\�h��Tc�"OZ�`p�,_�h9`T�ʔqn`�"O�uAՋG�fx�蔭�	�h	�"O�u�6��^���:��vl@�A�"OJ��p�L%	�y��J
�d���"O���ѣ[�W���`C�y���V"O���1�,\�T �^��|Z��M�<IJ֛/��B'J\�E���h��^E�<�F�� Pa����pU�d����.t�	v	*?��	S�OP�}��]]� ��F��
[f�Aw��#z�.�ȓT��R�f�
��`3v������o<J��D��7,FN����U8��r`�](?�2w�̝W���f�<lO����"�;\,�y���8+�50t��!pEj)���4es�L��j-��I%�/o�@�P��p�e���8�	�.�f|"R.��S>��X�Sy�'Ζ����7�F����3] �0�ȓ3b<qy�K��b�&1+��d9'��~�ѳ����2�d\v����Q���8*�;k���0���Z�!�$R�!9�!BP�
+A�p�RM�,e��6,�
Pc! �ʠh���'�F��RGB�x;�f�?	iL<(�/�m�#)��G��ڳ��[�J��0���,z 8�5�ޛ9t0i�	�'j���ț�D1$��4 �(�ja�}2���©kd�/�Ēp��"S�T���Q)���ɄL�%tX!��&]ìŻDN(;���v�eÌa�1�J�D�����.g�@S2��T�I|��Ù�J �eh�l���9�z��K�u*� �Ҡf٦�	fdR�_	�lyAL�m��c�eZ� �&���޶Wt���$ō8�>���gP
bB$q�&��?
������W�|R&��)�0�S��vӨ5&Ζ<@8�e��.N�h�q�J�Pxj�m�Q+ �pJ��������J!���Q֤H4V�T1��L|��	�TX|������<�<]�bj�1[���3�"E4M�0��%3cFX�uf����Ҍ7��O��ɒ�L!`k��*@*Vg?Y�����H�'#,�bT	B�z���8d��MgF��4=*�2֡)Gj&p�O�R����IF:5!�@݄�����J[?��%̒I��K׋�=�BpQ�[V}fO�����
/X���nل�HO ��_>)��Lѕ'��S�[�H�d6$
�=K󌎢 �IF}"�B f��]��@�4VL�k�"�'�*`���,���>a��4�D��t���']��	��� ZdX2�A�=��=	�=�%jBbZ5s%��ɀ��4j����	Y?��Y��p�/	��2ҥ�:�����Oj��8z���x�'��CD��4u��Q� ��_���޴3@�YT��c��� iG��5�^��b�'Q��ɐ�ihF��oAc��<
�.��]��V���#Ё؝\r٘�Y���]2�)�>��֬'L��䂹���D��_�'��HQSF�9���Ag�W�,��,��u儙�W�.�~�����Xq�IG}�
!#��iFמL㊍��lȮ��05*�f�t��d_w��㦫C</��l��l�,;J���-�z����5|O"�㤯K,F#�] E��$- �d8�Ϟ`�.�D~��
8J\�i �"ˉH>��p��QM.�2A��[��p�Gɒ,:(�� 2*4�t�
d�C���!t�n��hҰ�ra��7��.U��@Q���ҭ�G��]�D���+Ĺ�r'`aP����~�.�W�BqV ϋD�+�a�����B�^E$M�M{Ƒa�J�!�����C�3a�z�kG)[�,ʰ��,}4=�ɀ�wy���S&ْl~����	8t�Ѳ�#�3��c��I�<=^�AS�K�=Qӓ>o@��f ǽmly��k$��Ukل&����@�٦��=i� ϭMTp8��V�=����c�	�3R��{e� :�fΞ<&P�3�X\N|���A��}N���u �++�M��\�'�L�q6��C��Y[�g�0}?�q��t�? �4¢kά!�h�*`Κ?.n�C5�XC��~�MǼ�h�QȌ?��3��O�u��܀\H���d�T,8/
e��V��@F��k&b�{U ˯v:d�Sf0�@br٘ �ҷ%�Z�� �'x��T�'�,sъ��G >���
 q9Q����`�<�r��+W����Y.�ɡU%���Or�sL<I +��<�4� /U��iEh��D�Pѳv >�O��ݿ
�@<�t(��
{���Lؾ���'��DȞT<�O��	�?�
����� �m3 Aξk_*�@�	y؟4#C�
4� Q�b���� �2"$�yQ��P�H2T*b��� �P,!F�w8��Q�N0(�(�i���ܼ��6���@�B	]�f�&�����E7�)n�4j��hT&�gTZ��$J�P�FIa�
O汱B��0�Zb�ňF-�t^��K"��2c�F�2v`�3s�Y�D���>��Q��0z�|@
'��|z� ���6D�P��<��(4�ӈ~DT�c!�ˎ�!5#A��BLŀ~�R��:��K<��έ:�h�S����E�Р�w+Zi�<�ۼEdD��e����N�*��[f�<��[�{���! DC'�p"�	B[�<i��Zj�Z���ۇe��8��o�<A�`�"c ��+ ��)��0�jm�<��̈�%B���K&#�+9�*C�I�]	�L���).T�yӣN�d�B�%C�,B�b[==nfM�P�s�B䉤p�BP�R��p�B	0.\+%:�B�,���CKոz:�m�U�ƈ$HB�I�[��3Ƌ��#(�]0a�U� B�IC�MY�N>5b�U�A�DCWB�ɱp�Fh��m�����<B$B䉀c�R7Nڒk1Di9�h�Gn�ȓ"
��͵IA,�%a�t�ȓ6Ԧ�KEV�I�ɶ݇ȓC�*|���=0���unL�vp��	�J���f�<x�ؑ����.b`P��ȓo��0��kĿsE>��&oхZ#�X�ȓ~�b  Ę��x�u��T��,��q5������x����1�X�YX��!ʩ���ž4B����� p�r��ȓ_�� �4�B*3	
E���9Gx����%p@�� �2?m��C�d��Yv�݆ȓ�>�y��^�LM��C�ϔ^>t��ȓ�f��q.��R�0# 2 ݇ȓ]�ʽ@�G�)rnp��L�y�f�ȓ!%|	{�)�4W�Xc��6���ȓ,�.!Ȕ�3g�!#�L�t�R=��EE1��iT;1n�cU�Q,h��B�?��U�pH�;AhP�k�ɷ{��C�	4��8�+z���@�
�b0xC�	
Ϭ�ௐ�:��h�FgŶ?:C�	|���!!/Z!H��چ�A+i��B��.Sp���`��pl��3��a��B�P�|�ɑ��B�t�˥���c�hC�	&!�x5�G�k�-���VC�ɐ�B�R�Ӻ7i�!�C�b�$C�ɲp��y"���w3���1��)9����1t�R�F�@t贈�(�9L�!�DE�O��b��3%�$YQ�Ŕ(7!�^�c�H��m]�Ad>$���"O�}��'.n@{�C� N�;�"O�<�%k�
�^!�b�3d�4�:�"O��m[��8� � +��"O� s�
����34@� �ޡi�"O��)�j̿,�D삠�O{�v�"�"O���F
�m��؀g�+��Q�"Ofԡ��Ý^�`��f��B�HK�"O�����J���	��O�@$��`"O�����?�>$s��Y�Ya"O� ��X�����,���σ,�Z�٧"O&�;�D�9o�A��i6���1"O��[B�\$$X�	�fP|�&@�5"OР���?S���a4��r}:7"O>�j ��A[r�z�M3W̅�"O@����ԿRg���:a���"O�	
B�� >q�t'Çw`@s"O���� Ű:6(�jv&�9dmp�8e"OZ���䒚��P#EL1M�����"O���ЊgI�'��$&#�Y����yR�P�zW�ĮQ�ڼ��Oȫ�y��R>)�Dl���4R<��hď��y����X7��0a��WvX1���yB�Y�BHbc!� z�$񑰄�y2�T�[(,���#)Z��$ �yR��Y`&A�)#@<�&��y�F9!�2�cɵ*�d��H	�y2���,��1�L�~24���Ȧ�yR��3M&l��#B�|�B�1�J���y2�۳/�����ı@J&��S�D�y�TN��]�7	W7-�
�BcZ��yR��9dPj���E��+.�]�!��y%ˡp�@Y�H*T�P(à7�yrF�(P�Y2�Ο�ww�)A�`�"�yRn^�#T�c"�5u��Re)���y��O�tys��:k��Ҵ����y�e�
zu�B5*ep��ԈI��y��Q
>��;G�����Z��y�.4gޱ0���D��X4���y��)MЊ	���L	5��yҩ;�y��B6O�P-Z�O�9yuΉ{��R��ycP$Z�9"�na�������yҩ�,'JL�p`��.ex%�����y�	�.�����Ɏ/P�p��ݍ�y�@��(�Y#�ן-�@@����y��*.x����&rN����yNE�|� I��_4y�\�DS��yb.�	>�^�i��,�`E�g��y�HVV��b��	�(<)����y2�ѾZ�4$���~�&����[1�y��غ2ôlj��N5AT@�83F�yb��'>��o(��e�ò�yBlI		n �P͖5�`��u�]�yAPJ�Di��/ͥc8�x���y"�܀1��\8���w[8�3�y@X,�$Cs'Q6s�xb���y���/K�T�y���S��c�	�y2�*k�XX��b
}�
8�Rd��yb	��b��`mĹpy���@�,�ylM�[����jpP�3��yrI�x�J@�s�R�d�`����y�͖"dN�@���:Wi ��j^*�ybM��N�@��$V��AQ@�/�y�(F�@w�9`& �=�>�P�#��yB��+'T�ˣa:'�.��,�y�$��x� q9�M'&�eRgo��y�&�(Ad��Q��ì%=�4kv-�9�yb ��:��7�F�[,����uB!��I
&��Xf〢g����G"�l6!�d�Q�R�)�|���R�[.j!�  o,e���=|�k0�B !�D��G;��M�n���B�S�}!򄂴yo��Q�ǎ{Z�4ҥbƗ0a!�S�����M:iBH�5K0S_!�� �hRŃ-J�n���NW�,�"O��3���Q�ȱ��A�yH��p"O����64vmɑ`�$�N��$"ONu��-k���ؑ��3jl��"O����Cˁ{֩�`��x&�L�a"O� AM�e��n	/�Pa�u"O0L�cZ�9���J ����4a��"O�y�1n2�8��Ԙm�F��R"O�q���85�L�+���s6�#*OI�p뛐i�С`�ߑ2� !�	�'^� I�\��mb���<z����'Hze�@�	mq��{�B�.u�ʕ`�'�X�k��Ȕe���"ǌ�k�y��'`2��V�HZ�		F*�f��	
�'r�%��a��\�F��`\�I:�'�pB�c_�Y]<��ă��<Q�'�訡$�J��@#���f��J�'0�é���!���f>��)�'�@U�6jn��i��Բ	������.D�R��.L�pS׀Q��fy���1D�؊���K��y�:j�J��.D���2��*R?��z�Bm�"a�T--D�pXR�]"FOȬ2���1��\#�(D��b艕p5q�G��7�����F'D�Ls�
Ս>���PbX�0t�3 8D�,a6ĕ#j 
�Y�dǬ]�ȝ���(D����"�v|�UEN�Z�-	��>���M�Ӥ�6G0Y����6	("�����?A�D )�И���uPpm���MD�<���ڐwՆ�k�O ĠX�tDj�<i��Ū�����GR	q�I@7'j�<�6�A"i��E��		�48agL}�<��mˊ�ס�����eLW|�<a�ԧn�h{�� '�H���w�<���	a�A��K�;��Pxvću�<ф�J,bW���V�Џc��)�&�w�<1(�(>�1�K����諶��H�<��y��%�@�½K����(-!�ψi�����A-�ёq�^R!�䔂!��Qi��`�Ҙ޸�D"O`��R�K���K� ��"�<��"O��)����]Px-R���6�T	�"O���t�3%���$�0�|��w"O�-3���XE�0�ӡH�iY�"O�F�\�ARS�ȋ*���r "O iB�a�'xӄZ����,�"�*@"Ov z��f��!�!i�=��Ě�"O��"�H�n¸��j�钇셑�yҥ��6$`X3�A˽K�d�
4��y�ϔl����._>|5���y��L�Y� ���ɷ7����m��y"��`��,�#�T�]��\���?�y��.f=�Ib'_�kU�2q�<d%��F{��T�Qr<��4k��{���ă��y�CZ�Ae#�m�:k�gT��y� ͝sT���!K�e����@*B�y���:#�6��AgN�\[�4(�GJ��y��+©s�C�Q��i
�d9�hO��	�6�qc�D�P�1ëU�2l!�DABϞ�@�?�f%飫�!5c�)�g"���-�$sd�IT�Ov����'���	��ēV��u23��3�*u�O~6�R��0>!5 �X��\�D�5d<%a��
m�<1$E�FR�[�k�5䈄��`t�<� ���s�ЕFFn�Y�L�ش��"O���!���qZ��ɨRȪ�2"O R��^.pC �`�#S�KB�'��'2&ͱA�"4�x��H�6&?�90	�'
`�G�o\X\�!���}�D��'u`�q J�$��%r�a�.
���	�'cƨB�b���Z9Q�z���'���d��7Db���ŏ9Pb��'��T�a��,P�0a�+�J~:�i�'� ��P��88Rt�P�C�@%i�'�z	8##�
ML���Dn�C�09[�'8%X%b�0��3���n�8Đ�'�@�C�?<�]�e�D�a��51�'MJ�y�o�]^:=q%ϟ�S�}��'~8}�/ �~�����2Tm��3�'9�,�`�̮Z@a�b�ά[^���'a�Q ��j��=����"f����'�U�����v��U[�f`r��i�'�p@�2-�E�hLp��ڨjF��
�'0����;S�Щ� �'r}��z�'������ u]��r��o�Ĳ�'` ��5`մ	n!9Ri�$2.j�I�'�=�u�.>�$x��W�&�D���'���R����3�Q9/";�'�T)k���ݒ��be��+&6 ��'����[�l�F�X%:�xs	�'����t(��<�L�wfUhw�p��'��mBth߬/��˗�]�im$���'� DR4B�Z`���Zyp����'@����l�a
Z<:0�qkH8��'��X��K�U����-[/v
����'B ��PŞ?o�E ���7YO�t��'ǒ\�_j8��(AL�P�1��'1l 8G5�B���8G���c�'��x�f�̹.��'���9����'�&����Ȣv��Z�I0$@i��'�����ͱQ�@�[��3gn�i�'�`|��jS&L�x�䤚+�����'�^0" �W�6�s$��%��C�'������&6�"�q��� �����'�B�6��H��@qE� �-��'BF!Pg�T�ePtI7L��	7B4�'�L����~�Bu�v��-�T��'뾈�KO�6�A�O�[0�0��'���Rf*���Q:5$^�
*4��'kFhaE��=2����P~�N��'F:��኎=�h�q��	j~�+�'���I���H��0��H�5Z�j���'�R�P�,��;p|M�`��Gq�4��'1���#��w=\�鷏��D�
8Y�'�J�|���+g��h�#��y�h��0���%��cda�cEO��y�ǚ����!�C�n/`�eY
�y�2}�b����&oe:0C���yBI�:T�6����P��܉q/"�y�!��a"���Cv���dT��y�FZ�9�=�A��1!���W"U��y"��$�Z��2�4vwr�� Е�y2I˳F6V%��$o�tÄi��y"�O�S���s	�0]��)!�K���yb�\�h�M	'��
�|Q8����yD�v&jQB�I[m ~eX�I��yr�͑Z�f)h���_���H���y�\�k��}�`�V�K�(a`Oӽ�y
� ���4�ʷh��
�Ȓ6h���"O e�`(��Haf>�,�1�"Oj0"$҆O@��[�e�;7t7"O9���]]}�a���v���"O�hK.X�5����� .Z|�j�"O4�(���<j�Yȃ��b�4���"O��IHN(~��bA��|nf�`U"O�8�V $b��!Ht��dq�b"Ovx����%�
A�5.L%H,R�"Ov��5*^�<��eD-V�W  �b"Oh 4[�+qz��j��]�ȅpD"OtR� ��"vurD�!}���u"O:}���D�O�F��t�C���1��"O��J��v)�F���V��j�"OT�I b�+Y�H:�锽+'(�C�"O
�Y�,�@�d�A���4���"O�[`hB�tq�i�p# p���"O\�sT�B�Wl��K�@�N]�5yS"OԀTCI�i�RH93gB�1���"Ol���dă_�h�� U�g��ɕ"O�A�s+ںS��\[�7wv���"O�����ʩ ؒ���c^?oZHT"O��a&�:do@QXF͓�DA)iQ"O�9���&,�<)чk�����"O"=���W�2������, ꕀ�"OBy�)	�=o��R0O�y"O2����H�8+�KC�]�j("O~�y��ay��@��:��B"O���p��0�lQ�@]=U�F�(u"Ot��G�(#`�����,e���"O.��i5+G�$
gˆ�*�� j@"O��&��P�����I�(�%b�"O���t��;D�H�sOτH���s"Oy��`g^�z�l�-}��LI "O�]ň܋9��T�Q�D+u&p<��"O�(�0!��gT
%yPʇ�?$��	"O���Ug/,��0�")6&��8"O����M�2��}`3��,�=�u"O� !Ga�mw�6�������,D�� ׫5T�������n����j)D�,!��slV��� �� !V�&D���N�A5���b��s�	we(D������j�����"e���3(D��pE�ٿR�H�RQ��4Gz��&D��W��t,\��P�I��@���8D�,K��S�P� ��+�t���7D�dP`╉8�l%#u��y>`¥J5D�p�&'�5\�V�s0(�^d�`�%M(D�L��cX]��B "�"�*0�8D����/���^�����[��(�q7D�H(p�պBAv,R��Y;���ӣ�:D��3��4!L�d�QELQ�hd�%
$D�hp�P�E��q�wgטn�:��M"D�@�ci;� au�3�؄�B�3D���dL��R�N���	�t`���u�&D� �G�J5:_�  �d�7�Z��f/%D��`��}YDI�A�G�#̰6�6D����`ܖ%�sbٖ\����"D���rm��f�hu��i�pb�&-D�<�e���q��q�i�?]w�ab0D���I:-g��[��X���2��3D����l������� �f:���1D�����[�8[���RA��sql�q��+D��B� �%d�,�����s�:𸗀+D�� f��喊z�r�%O�*y���v"O�	�e�,E��DHȣ>r�!Pd"O�Y2T-!g&T۰=!@��E"Oԁ9T�l�����Le�Tm"�"Op�(�/�\v�yWC��;�����"O�I9�Â{Q�]���w�Ȅ�#"ON�g�E��(��S��)U�de�"O<Lk���]v	�Ah�58]
t�"OB��HY3$���IV���I\(�C�"O�X�A�,�q;�&�J�s�"O�=��+J�Ll��C�O#l\��"O@\�B��)˸�z��C+f� T"O�p��cU-X?:IS��J� sA"O�`���������⇃aYju$"Odف��<\��e���B3m!����"O"��Fe�~���𒏆�f�uzf"ORmi�?R�6,%�ֈrY(���"ON)y�g�QR�A�(׫E���J"O����Ø1�.5�G'֘G$���"O��s�Ο�eS�D�NH�*�B�"O�s��Z"c�ʤ��&ٙ]�jȩ�"O�lpЗ6BuxD���\�*��"O��:�N�K��� �(��C+�CU"O���!�
�n�\�A""���"O���!7X��Vo��c��a�"OJ�;B�E�C�n$�t(�:&�m"g"OEqD�z�~`��H���pS"O�<�ҍ�&yyJ����Y���h��"OL<�u��6� ����9:���c"O���f��'��#� ˎ��D"O@�!���Zu��� ��uv�as"O�!��l^�U�FEʃQ^�u��"OD�{�+��b����3@GI:�"O��A#�y�puHe�:$U�l3"OUA��M#l���KS���"O�M�`��4�8���F�)E����"O�hyTG�:b��DR�Q)B9��
w"O|%a�OZ��1�!N���Z�"O
��*�
dؕGF�M�h�"O^!�0g?T�LMpV;`(	w"OJ��A��j#�S�z�>lPP"O:�:T�0�DX�ˑ9��3"O�-��٧ ����끀epxd��"OpĢ'j,#t!��ր}�xy�"OV術���(�����$٤W���+�"O${�	Ց	-�K���v���8"O�����Ŵh��0*D�+3�v1��"O�$�J ul���/��)M`�u"O��e�%-�AC$�3O3�Y��"O؀���_�+Rz�R��[�3d�R"OmztG�%?�t5�'�<���"O6Xhb5��v䀙-�� ڀ"O��r�[�5@���b i�Z��u"O��T�Ŕn�DaP+��m���c4"O��R��G6%@�h H �Z㴩Ȕ"O���4H�$�L�q�إ^��e2�"O� #�g�,��ݩ�![�|��1�"O�5�q�N���
�"�,L+�"O �sA	:נ�� �(�431"O�|�g	ޯG<%����.����"O�[�.WT.%��/\�@����"O,�(f�F&�RK�/�$����1"O�<�B�#
���*!]�oG��Y�"OB��DO!$_���F�i/J���"O� ��"��x���;}{6�1"OPM*��e�ĭ�r�^�}���c"O�,q�EK�0��疓W�>u��"OܑqBgG�U�p9�r�#U�D�K"O�J$K��ZYLT�`c�?K��	�"O:�KPP�{��Y"�-w���8�"OYk�)A�i�
���b���P�"O���ܛ���"Q4���z�"O�M
��55�"U9�(��1x�M�"O�%�ЂP6�13��8\I&��u"O>�v��b#���b&N0ʝ�r"OJ�C�� ��U�DGI�~;��9"O&�r��	S�t�s��;ƨ��"O�����Ie̼�{e��g ��3"OP}�RP-O���''��t"Oz�����ova��E\�r<J�"Om�̆*T�f���ש+̼��"O��#�G휵��M�'����"ON��LĮh�h{A9n�����"O�M:DN.Kj�aM�f ��"OȑCEDM;��@B��u��0�"O&���D�(BI����R8iׂ�� "O�I�5�N�z�����.[��-b5"Ot-�$��,8�C��V	f��"OʔJ���o�iKs��Y���Q"O�]S�)��w}H��-f�}�@"O� IsN�er�l��Ϳ�*�K�"O@���Ǆ�5|����j�c��:�"O�x�״IZl���5(��CV"O����K�);�"�5E�tP1�"O~T�b�H�G_~�Iu�Io��jR"O^:V��z���d��</wa!t"O���E�M���5�V�Zu���"Oj����\�Rxh��*cJ��"O��0�$G7w�𠦤(�X@%"O0u!5BAf�r�d��_(,ث�"OxT�3 �dCXrCH\�0�=�"O�(���Q�~tٷ�5���"OH����,V�
�⇩��5�8y"O�� $�E8P7�Q5J�l]��l'D��;��S�6=�fcП!�D��@�%D����C#=��i�$�ν6:`�ڧB"D����+|Ƣ4�7f�Q�V,��/ D���R�b\!:ԥ��$Fd�)��1D��B�C��x��5�"�=G`P� �=D���B��.s�2X;SfI��N�q��=D�l�S��HV(02h�%-G�t`:D���@@V�;�S2�Z>D�`s58�L-k�b�Kz  �,=D����Y�[��� !e� 	�����;D�ԸdþC"�}[��!XM �B%.;D�H�!��-�r	���U�s��$��e9D��B��&6�&d�!�Q E����6D�$�*x_���@�׮h�[�!�dh���;�J8Pg������!�S<R��dŚ�.,�(��Ux�!�݁7�=�P��O��:���cU!�d9�0�r��?���XǧվY!�DXj)$0��(Y��]�ȁJ!�DK5e��t��&Μ�]S�-G�\�!�D�\�E�����D�V���G�!�!� �R=�#�2,�p,�p�ϝ=|!�['ʤ��VJ�	v}��œ�jR!�dii�j��8��B�<!�� P�[���P�>�9�)�`����"OTd3E�A3D�`1#'9����"O���b�Y��BA�ä�� �"O�y��ċ?$�&��1*Z�'����"ORQ1c˳13�xw	X6�2)�2"Oށ3�lT;���0�÷pU��v"O2<��MdxZUs%��9��q�"O֥ �!�:��r�EO�O���Jg"O`��Q�!�P)f����Mx�"O���G�<Sl2��SeY�G�80�"OT����;K	����J*��\��"O�p�R��Y <(��S�|XD�P"OnӒk�3 �|��@��79dP��"OJ!)�' x�L�O�g� �A1"OdJ4F�5e2�d`sD؜=f([�"OB�0��0Ed�م!�3l��Y"�"OM���YxpҜ�J(:I"�3�"Ot�9W`Ù'p���たX�Mw"O��R $�VG�-�f#��I6���"O�Ӓ�KeR�r��s��u��"OJi��+ŻX. �(Q�Q�C���y�"O~��KߕxDq�gF�Hmд"O�L�'CO4]�V|!�/�6]�����"O�e)���n�ܽpn����ò"O�,��b�8T�,Kǆ",oL���"OP:��@//������%��}��']��4�
�[�Hٺ��L��ez�'�(�E+Q?azʰ96��+	� ��'��ۡ�՛ImNP�mڦ���'�jP��cT�gY�\���۩	�ҝ	�'��U(5�� Q�R�)��,[��x�'���+�B+n6b�ZF���2�T��'��=S�&�� �*����V"Ĭ���'�A0s-�3rǠ�
D��2ּ�B�'?�ABR(��a;�m*Ãͩ*V����'"l͢b��c@\��⍛/_L��'�@I�cOߕ;��Ջ�G�'&T�S
�'�x�x3�?.B`��$�q�}{�'w��\G4p�J�CEf`�DB�'���Q,E+�=�QDT��Z�'���94,ƕC�b�d�3�<e;�'�J�K���%M�r\�G%8���'9�����\;x�Qq��.{R���'mL��h��S��]J (ߘ{�iK�'������#.`x0y&d�q2���'�$٢��S�v5a쐌j����
�'��(���P�3�T�pGP\�)
�'?��HE�*?�E��������'�Xm���@��L�1���"	�'����m��j�X]f�͆ IH-��'��a��̈ ����5�C���9�'��5#�J��>`��KiAȐ��']N`&k >�d�B��t(҄@�'v�I ˄��dzm�,kH��	�' v<+��a-�l�F�cWހ��'Lm SN�<r$��h�ȅ�_H4W�<Af6t�ڠ��(M,��yją`�<Q�"�!d�:����=L*Y
�FZ_�<��2�ԁA��n�~���<�����3��x�`m��RYB�k	R�<�)Ιo�R����**�a0�[h�<ǆ*<�v�
���+&�]�<��)�q<)"H8k4&M�f�_�<9@LQ��E��T�C��}�Q�N^�<� �x�����hp�t��SR� �"O �8�J�`�Б��Î]؅8�"O6\@O6hb�z1l�9V�-t"O�pq��o�L� K��n9��"O��R���M�ʔJ�
Y��"O:肐�<th]Y"�(	ࠜ� "Or���a��nȮެ�S��)D�4��#]o8p��5�̏G�tE��%D�<ken�'8Đ|���<�|�wA/D�����'i�rL� m�yB$� /.D�x8Q�����`�D
�pQ2��6D��B��ӝA���¯���(l��G3D��F��%[76yA��Z� �(4D�t)c�" �鑁�0O��!:R�2D���m�8S�
7/���=���-D�,xS�Q4$������. �h� *D���sMƙ3�|�@Y�A������<D�x�3D�16״<भ�6��ԠI9D�����zl����G�5Nq�@��f#D����n�\:��k����#����&<D��*�DY��L����ʲP�,�'E7D��C�MԺI�=�e 	�ƦP��#D�h�G� z�N@X�%�"��0[ׇ!D�$�` �d t�@�⍮#����@!D�P�!`�!�X90��=s�`th6/>D�C!g]:���uM��W�j=z :D��I§ى,�F,�u"�.&�6�R�I8D�����څM0j���E�l�2%��b5D�\QC�J�U� �ib��2\�p�2D���AfS;\\[f�O�^fb�e$1D��3D��~�©@�����	�g/D�����C��0�ĉ��<���:-D�Ty�)��>:b�˲ɔ�.�� `��*D����I�9ym����Я@-6D�`knF=X�����f�&D�� ��2D���3��?�8���$���pS//D��b�C0�.���H��'u�|�ǭ1T�@[g"¸FT��%B��;	��"OR���g4,'M��'P�!�D�"ORmɀ��CC8)��Ɲ�?$���3"O
]�%�	�D\�q���U��i"O&�h�-s���
 e�{���2"O� 2�� ��$ꃁ^2���"O,�K�n-C")h�)ρ@bVّ"OV��'�)z>d����%}jH��"O^4��hʈeHt���;s\,��"OH����R��$"�Ҿ1BJ��"O�p�a�����͋����+�"O�1�r޷A���%bf�L ��"O yI[����d&V�3�FAA��(�ybj r�@%H��[�B����rB�)�y�� *�s�%:��c"�Y�y�ǟt���p)յ$q|��g�
�y��+� j�J	'�x��A.Q�y2+�+Xy0]qsh�?���b�8�0B�� 3@6l��W��\�-�5O�jC�	%:����c�4#�la�%Asa~C�I�V+����I�G�Q�Ȟ/+�B䉋 3���c�v��M��`�G�C�	4%�	�'-��e'`e�p�"�RC�IK�`���ą}�,�qEV34�$C�c�<\p�%F W�e�GhS���C�ɏz�n]��)��,�$��G.\UظC� �����$��SM�A;�ȕ�/��C�)� ��0���5X��AƉ!�ZI�#"OZU!dc-"�r}��V�PH�=sE"O���F�d��c�ק�c`"OhݹV*R_㰠�ga�^����"O4��o(H������1n�h��"Od��a�
�
�(�9���"y�*%��"O�qb@,�:s�t��eLr��S#"O��� U1
�@rq큧q��h��"O*TR�Ƅ*BW]Ç�]�
�<��"O(e����,y4�Y6H�GqJ�"O�9�U�^>R��8U�_"	>���"O���n��C�l��� ��-p"O��@��35ﰐ#��9�R�!"O�lH�b@-I��� ]�b?�`�6"OV]�QI�)�u� ��i��9U"O����'Q���(3I�eC��ӥ"O��"r��x� N��o=x,r�"OH�x4$	�6eB��� hI�$PW"Ob ��
�r����+8;0:]Xa"Ov�!�H
}�lL�p��j��a"O�1��.�3���9nŪ"O60jW
�'@�@i��*��#"O�����[ 5p�gуL��sB"O�1���δS'���DZ2R���`�"O���A�T[@]K�D�{�ҡ�p"Op�Q�JJ�U��0P�m�y�� �"O��9���at���gÂ1�X���"O]H')��G\�%@��$b�"O��g#I?dZ���,E,9��R3"O�}���ZkB�!*3f�t,�y�7e؞� �1O��x�R��yrCI6Y?�8���Ii�ɑ����y�H�V�m�T��0F٠�H�)��y�C_�_~�zC�J�M䤩j�+��yB�_�G���,�+}����yB�Y7ڜh���y0E)FA^/�yr�S�,��Ҟܾ�xUO�y�%�Q�h�� ��	���p楟�y�d��I���ad��X���D(��y2i@;8��"��ySH�&�y�J������Uk����R`ר�yR�ڟ!N�Is�ڪxEv��ҩU��y"��:]����>r,�ͺ�*���ymZ1K��� ��)>�V�����y�M��H���jf�!!FYǥ���yba0J�u� �҉�(ǂP3�yB���T���8�ğx�Iz�	��y�( ��|��LGܢ�!�W�y�-2P��#��$>0&ʱ���yb ��H
�	���9��$ʃ&1�yR�t���#�%K4؆)�֯��y��0B_�����(T���2���yb 'op("QNRS 	#�G+�y��0�8-��K?m�5��b٫�yҬ�%@)��#lC��@\)�`	�y���;��;0���"{pM�bW#�y��.�J�`�O��LJ�a�$N��yB"�Z�
 
��֤�酇�y����z��'�A�|�T���W�yRL�_����&�s���p�P��y"��:(�ȀҶ��<�2X�'g���yRQ"_�بd�Ȭ>܄�戁�yr:c*y�G �´�O���y�!��\�~�9��Q�}��I�D��y
� �����P/�`����R�@��L��"O��B0@B�%�b��%�� �����"O�dRW�=3nH�����?y�l��"O���E-8*pIA�W2?����"O���]#4f8!��#��p�r��S"O0�b�?z�L��C�	�Ȉ���"O,u�H@�7��$b�h�=���¥"O<p��f�c2���%D�P�(w"O�QgEؿ�R���G�Y�yq"O6�;��W~0wfV�K2P[p"O������f]�m���%G�脠�"O��#�!F_���o��}w��@�"O@MZǬ��/� ���(I�UfZ��"O�8���V�@����#@y4D�"O��$���Wu����,W�eG t
7"O�q��6|��4:TL±M=��a"OtlڃO�fȂtR�b$^1�"O��f���~�̱��GI�&ДI�"OZA��.�� хg�6i/m°"O�!L��Kc�$P��X�5�q��"O:E��9nmP�20��pڣ"O�Z���P�`'��2R�� �"O�e�B�{jp�`��1M�0�"O�t�V'L�+��0�B+kZ�у"O��W`WFnV��W˙4=�X9U"O���h�_�H���*���06"O�4G ӊLUmCM�l��"O�9�`#�y�����j
�U�P�"O�Lk�Á'����Q$�i���S"O�H3�o�1[Vd��2{��Ha�"O�;�ď�Ae�dP5NG�-���5"OF���oU3l���읗Q�T��y�e-����]�X%|e�I���yR���zx>Ř��T�@{�Ls�C �y�+�91>���B0�D�cZ<�ybOŚ:�еx�ȯ
ɸHA�3�y��	
>���+�1s�t�k��E��yb��9/@N0�� ȃn+���#�-�y2K�2(��tQ@$���� 0dL1�y��4���� }
�����yb�	�r���I�e�1�斗�yBD�R��(D���Za����o�;�y�F��� ��� Z2ze�$$\��y���!M�%y!˛U\he8$�Z��yB�O�2s0Lx���\M��z�-ˢ�yr��U��1�E�P�`d��F�y≊8�ةC�[<Q��ْ��y�@�$��wM��p{�a��y�
N~�deM�d�Ҥ�ąת�y��>&P�kG�[��%�dF�y%��L%B$�P���Y�(%�Ӣ���y�^�^�mg�"�~1����ym��)�llH��")>II2Ƀ�yB�Ez�� ޝ��E�M��yRO[��*5�`S�rqǇ��y��ٌ�$�����i�5�y��Og��A�ŊA��%�M�y��o��QV��!u�r�J�jА'�!�G�ph�U�F<o�YJriN�!�$�	�2���R������Ww!򤋸K�,�2��Y%t�<�@R�*?Y!򄒧� |�@��0*���ȇi[A !�	�\`�{Ć݉k_42��!�$#~�v=�'�{ 4�MJ��!�� �6�v�4�{�`�)U��5�D"Oܸ��MT�˸)�2�2.�n4B$"Oб�����{��ٶ��=�zZ�"OPXH�ǋl�y��놙n�h�C�"O& u�J_}��S`�
:H�����"O䁂�$�<fn��:7� �8��D"O�ēE�ȦE)D���͏:o|Hg"O�eѐ��F	A5�
� @��B"OHH*�)�\Ѣ9h$H�΅D�!���phB͚\g�Ģ�N�8�!�E�D��@D�8HvQ�E#Z��!�d��g�Ձ/�6l���HD��B�!�ą<b"����I!h�*ԩwA�!�ɚ�h��bV*�v�P��ԇ"~!򤗖���f扥FP<݈�茷c!�� �i��ŐF�A#$4��rv�զj&!���r#��(�3w�Ƞ��ǝ!��/vВ��f4$���*�f�'!�+ٌ�X��.%�\��R�E�7!�P*i�����gI(u�Q�5A�!��R�Vpe��fӾ����N�!�T&���#� Ud���8���5�!��F)j}�t	8kS:TB�ݸr�!���}���]��Y2͠%w!��{ɮtqn)M��2��<?!�$[�'St|��f_33Մ�b�N�>!�Ć�^5�m�%ET3d!�e�L�90!��'E�Uғ��,x/d�qKîa!�DǙTn
5F��O(�dx0�!�D�=<= A��rt���fE_�F!���N�>XJr��$Dh4�$&� �!��i�+Ş(n����fcN��x�ȓ:�L2Peڦp�	 �KN8�Tt��+�\Ԃ�ア��������b���1rΈ�U�� ��Wŗ�dy���]2@ c� ,hF�kVb[
L썇�#g<�B�ɣJ��qk`���FH��8ט�`�������"��j����ȓ��b����V��A�A�0�N�ȓS��T	��T��l�[gZ9
��#6�X�`�N��ǫ��N���ȓ`�N��c�?W�jH���ۮ��,�ȓ1�D$s"�)
fx!��� ˆ���Y�]��
-C��dA4Z;�Y��`mfi���*'J��䤕0�
�ȓgq�6a��X� N*8s�U�ȓ*��m0�%V f�:�J���)�Tx��~*t�)'�S\��!�*����ȓ+z���oE'9���2U�^ @�Tm��FP��B��~�b�"`
�N�����&�)��GY�d4��C\*I����OذQ@����"��� ��`�����G"��*��0N_����W�.�-�ȓmw�HyL6F�N�cJfd�ȓd'���A��2��򪗗4o���9"���d��6�$��+ݑ)���ȓ4J��C��>j8ʸ���Ҵq�ԅȓ%�xSX#�����i�ȓ%��(�<�����WRy�ȓ>Y�Pj[�r�	�q@S�t�ȓ;�Q1,��
�
k�nزP��ȓE�E���6N��l;�Kī\�����O�h��K��Nk�!�֤��h�:<�ȓXkf��g�;iP0ؒB(A,&�t��S�? ��3��\'}zvdxE
�e���Q"O8���EE$�x̱t�k���[�"OX#�C��H�b�@-˦��]pS"O��z�K�3��XT�U����w"O:�8���
:�ܨ���Y�c��"O�i����2�*Y)ዏW�t�"O�!kBݻH���̕	O��&"OD���Ea&��8��;E�°"Oڀ�Ƣ<>��X�U�]*b�t5P"Oʹ{2���`�����������x�"O\��� M����P�Y�\�R"O�}�$!pO���%׊�"On�ǩU?�䔣`�I�L��̡�"O��8�D��c�0Y�&B��~�.��w"Of�ؓD�B?$P0@ěI�NH�5"O2X�s�Rn~��n����f"O�\a�l�6> �<y#W"O���I�?���Ak�zӞQ��"O���pk� �x!`ʒ8Z��sd"O�\��dJ�6ބd�!Î]B���"OL���×s�|���u;X|�""O(���OD-���j��!�T{�"O�1iD��>�q���x)8t�R"O��أOQ��Ȕ�GeWw~� h�"O>4�A�� �����x�3lJ��y��S�>/hҒƝ; $�%�"��"�y¢���D���&?ƍY�ŋ�yrD�.>È�B�)V�^�hQfjE�yr$Q,�ɰ2� Y�DyL��y"��U(n���\�~P������yĒ�=  �8E� �C'@x���ܿ�y�ǅ5�]����80��6E��yR�� j+(ԨV�Y,�^a�$MZ�yҥ��uܽ��؇"o2���J���y�4��pP�Óm\���y�pl��2h���������y�)¹d4Ex��Y��X� SH���y��)K#}��\I���;�N��y�)�͜tA���@	:@b�%�y��6F����FM
9-���B��y�bȣ1~N��ӹ-;�,�G��y�$�"XJ�!sq�,�� ��E��yB��1�����*��"���H�#�y�.�y�������&��b�9�yb�Қ?;* ���`�\󂈛�yR������aD	u��d�R���y�EHT�����6@#��ٻ�y�◞[��S�K4hx"x"mS9�y���*	�1{Ga�f�������y�!L3?���Do@'X�ȌC�"�yb�}`"i��*U�P�<�����y%�ؼ�g�H	S�&u����?�y�ϭ(��h3���D?¸���y��Y�%\̓�g�5Q(ujSo��y���#l�BS!n2w��q�EC��y�fӻWC� ��3h9�(c�W��yB��r���ǆ�f�x�@%I9�y�g�#X܄`Q� ��haHM����y��8�D�pЃ��`5�B�B��y���<���2P0��`AmA#�y��2s|ec�<@��@���yJ��_K���E�.������>�y���^ P����3�"�p-��y2&KafZ��J�23�����֑�y
� 6X�H<8.ZQA����T���4"O��EN�M҈��v�֛R!�!H�"O,u���0HQ�q���;5B�#�"O����I��!JrN��@(�U��"Oqh!�$eB-�vL��h	�Ĭ[�<a3Y2-�o#c��xw���ybfG�����I0M��vm\��y2�֪!xJ��8{��� �@���y��A%Q����t��vE�qD J��yL��T�� �q	�4�S�K$�y��R� 9�4K�%d}��HBm7�y�℩R�	a#���H�V��a͉%�y�聧>Kԓ"���-��� !��y��"^�P u�ڂpj�Ѳ-��y�`��"���'�hSx䱒I���y�l�@|LP�U��3d�Zb`��yR�F�GU���V숇ae�,�����y�i?0B%2q�^��D$�ꁹ�y�`��,q���S��:�� ����y"�r-��(�BE��}�$��y�'N�P=^9Y"���V?L=�3�W6�y¡��U�h(�o^ Ѥ�a�O �y"[/72�9�b�	�:L�^*�y��4=����#�Z VҬ�'O��y��%
�����g Os�,֭��yL�"�|����_@s2豆œ�ybÓ�M�^���gɺc��9W 
�y�@
4G��3ХȵF~Y��͉�y��S �N�sӂE/y�䕢a�_"�yB�&
]r��U�ٗj�ܱ�NT:�y��5�2��ŏܓ_�"�$D�y���cՎ�I�/"�H!�bI�.�y��6�$	� 7��Q��ه�yB�1p����E֊dێ�s$���y�(�3'jK7��%�r}��e��y!T�h1@��#U�i������Ȇ�y'��0���P�O�x���!��yR�O�p�9�>q�����P��y�'�1="|bDG7lI&YC`�^��y�V������� /��ěG���yb�Zz�!P�l��ok�M)�$���y�A�0k��#D%��h��
�蜻�y��_Tp-����>c](1s�R�yBd�_���lU`!L�	�
��yɄLҘ �R��/)��a$��y"&L�E�v�IC�� Mi��a�AE�y�.^�v� C��t��*�K��yb�L�N�J�����e�2�&ϝ�y�^��� 6�c����S)�y��`h
b��]���o٣�y�%O<Jp�M�r�4kQ̏�y�&8�6d�#s�����К�yBn�3T%cO�e�*���C��y�g��V���%�*����H��y���,"�rDHD����)� ��y�O]VpI���2���g���yr G*B�~t
�KP��$��Z(�yΌ+�]�S�$6�r%��y�E�>.x���Ĝ�H�p!�Q���yR+Q�'�1���[3NRj=��J>�yRGնL����qKX�vK�����yhrQZ��I]�d���3F���y�ˤM{Q��RE5���5�˿�y��Z�}���j@��Ak�	π�y
� Tm�6$!ȱ�E���E�B�ڠ"O�u�tb�e��H�O�z��"OL�(@����yzvdG�
�Fm:�"O5R�UG�8�b�ɬ�Z�K�"OP�x���Q3���.4�E��"OZ%����Sd���]P��9�"O�a�0S�&$
�3Qw�u"O���`䊩����-	�@�w"O$���!���PeV�Q�JE"O�4d��M�@�Ɓ�=b��%��"OB��v��P��T*�6Y�be�w"OP��w.x���t�V @f�A�"O`�#3�P� CNL���U��16"O�h�ǌ�K}Z��2�;؁&"OV��"��hc�@��-��@f�y�"Ol㣔6m��p���Μ-%,���"O��!S�F��T��Ŏ�[�>M��"Or=��M�${��|��k;fm�"O,xHGGK�J]Ǡb9d�!"O@��"�r�dc� BC�E�"Ov)�c�C���D����-�4��"O�4�Ј\[�všf���N8�"O
ͣ�-K�
@���
#`�d�[t"O6���Cмc��Q��;	��pз"O$�C6�ʪ`B��e�,/ߠ��"O60{am9���S��n����"O�T#��A� xx0V��KA�X�"OTy[�I��O�йQ����y�"O�i�@�(�L#Yayc _��yR$͑gRExV,O�\ &��O���y�"�cԬ� ��2Q*=��e��y��D;V���	JO "`�Q��y2�R2RHh[-��W�(��	�y�Ǔ�V�>�!����JDm+g��)�y�hyaa�ΚU�}R1c�
3",H�
�'bA��
>(͒㠉�.�t��'M�	7��~|�bXw���'c��2mҧ���qk���y�A×�b�#A-�(�V(�pL��y"$�'k.�o@3VDA)��B/�y�ǂ�vMԵ�V�S+IR�u{"%ڳ�y�G�T�ęb��70�x����۲�y�,��w�8��g�֥&N�53�ӏ�y�e�/[���F���r7�@	����y"BE>L&��4�?���E��:�yb ���b��2͓E	���ꝡ�y2☂ÀIؖJO�6�,Y"����y�j�� �S5j��}&rr���y��%(��жB�q?B�+֠�5�y�O������=mA��2u�Z�yRI9G
1r����b�Z8����y��R(�kD�߰F��q�ra��y҅!"J���S�O8����ҏ�y��w�B�8�Ұz@�L����yr�І&>�݉�CT�y�n�U(�6�y�� 5Yu��k[?A` �^0�ybdY�W�j���<9{�h��m ��y�Qmbj���ɨ_4`�"���yE��	m� �h�QC�L��� �yRM��K*[�ҸI(x��B��y�	�C��T���a0�8�k���y��8P��h�bJ�|<�h���yr�Q���D�M$oyn	P᥅�yR�\�0\���� A�H`@����y
� @P�+��6�<���/ɥL��ͳ$"OU�2��2�,9F���T�Tp"O��jd�B�f~V��m�+_튕��"O^��bA�!o�����lN�?��t� "Oڬ�E�݃q�PIڌn���Z "O��95h����щM8x���X1"OL8�1Βm����qJ� z.X��"O�M�G�^�;Q�M붨M�^	�""O�H�d O=����4�	9X�^�B"O��`E�(�8�x1�?I>�P�"O ��鞀-�NY�c��� �6�ȵ"O�[�#�A�f�BV��#>{,ɢ�"O2���F؞
ܢ���B��gd]��"OB�ࢯ^��P���!��$U��$"Oy����
�J�M�y���yrm�R�h����A��P;բ��y��@
�(B�a�1�L�yBk>"� �P%Ըm�2ab��y���X�PfŜ[T��e�:�y��W�H��]�"%ԗ8��������yB*F8f���
D�2��! ME��y"$�.zK~|���K�(ܐ���ޔ�y�猗<:���h�,N�.Y��&��y��ɱ6y ]���F(D�N���W��yr�]�t�����,>�` �/K&�y�����"�gũ5l��D$Y��y��72� '��4 K��$�y��P�tmRM�-Z���˷i��y2%5UL�-���EZ��b����yA�?M�6|��dIu���Չ���yr,KY9�i+@ꚚoA� ��`�#�y��A�1<f�ǎ��b#�i�  ��y�+ν(�,�2���F}j�sP�'�y"��T�3�!?�L''J�y�F�,¼<Ғ"O�7<hTR3��4�y�+Ǔ"�R���)��Ed�s�"S��y� HZjV�*�G�9�Hg�T��y������%:�����,Mmad���';6	��(� FvX}�b�Qj�I	�'K�����݈[��ʤ�J1l��' �ܰ���V*�=��HX2Keta�'>8���!�N��,R;0e8���'�$e�E }�V�ɵ�20��d:�'���� �q�¼�H��+MXh�'�ʄ�X�cZ<I
�������J�'�͐���8"�h��9c�'����h٫ �h�b� |9�@
�'��(P�MX����E�5n�T��	�'�� ��,�v���m[_u�1��'�F�c5cK�=�LD��U����'Dt��ܔD8�qde��O�Q��')��f������:�P98�0�'�J��6$�-N�.=���԰,�P���'���Ȑ!�)p��"G\"��'�*1
�
ө2/�4゠�i�� �'�+�:L
h����� ?�2Ȃ�2D�1��M?X!a�ܝu�q*")$D�D��D$Dl���E�?�Mץ D��ǡ�&�:��D#��\�(�C>D�ty ��[f�(J#�~R���
0D�$��Mi���x����q,�A�E)D�����ߡ�bt���I+N)qL&D����a*{Z)�cE;|��l�D�0D�C�#X�]R����x3�0D�� ��BP��8-3hA#�a���p"O��9�#ħ^��$h�OI^Bʔ"OZ���
=�$�� �"L(��S�*O�,�E��@��K�b������'��%���J�&u���6�»��	�'��uC☰lyά����w��2	�'?D�[a���*!#$�]�pz4Y+�'!z�x�b� o��K�]�N<��'�Z�I���B5Y�[5HKlH��'��(��,GG�����l�����'o0�2�U�<���x�iǘsy�(��'�>�2�*J6yOH�@5%U�6b�q�'� �P�B��X�����&�T���'��jR�ߏ���3�]9U:5@�'��PA��S�MP��h&���"�3�'���0����8���&$8H��'��Xa������V��6]��'\vM�zN�Ivi�+�@��'��U c��uTCuF�A�\��'�H���̋�@�`�Kn5H�池�'P��� �I}lyঊ��Oè�z	�'�Z�ǁ�-�X�&�ϼDr��	�'� �R׮H��
��� >^%�	�'�����ge��"�I50���!�'7�Ջ��B�Gj��SoUm����'��u0d ��r!�ip���H�����'y<zR͑��f���?���B�'�,��gG�}��ѐn�D��	"�')�lK!��������KA4v>D*�'�<eI�������I!MԀͣ�'|���L
v�6E�f�D�m7� ��'y`�ǣ�AG������X�h�X�'}Fm	��FJ�{���<�H�3�'�ȕ⍗;��H�DHQ�<��U	�'|*3"Ã�!��h�d.D�<��	�'i�Pr"�]$����1�r
�'�Z,�qE��f� ���!�|$b�'�l���U4����e�I�n��'��8� �.Da�uLeM��'��b%�B�v�:�)tA�n��'�"-�`�KtT�qXC�T7W��8�'��iߚ�ނ=�"O�\< �'֜)knb�=�d�t��'V�]�I�lX�貅��`ɦ���'�䉴�T�e�)"�F!`l�	
�'��q���S�"����]c���	�'	�}H%k���'
�a�����'v!�Pe��"K7��S:�Ւ�'N��CV�P�b��)�f�E� �ȓ96PxA�^f���H�;����O�T1���#Sn��5B׶L�\Ѕ�#
<�16N�?⤈:4#��)�n܄ȓ%�5{�B�4pd���Bjϸ!���ȓy�hZ�mɬU~8#A�ʲ?����9�ԑRG�=H�* �3[�M�ȓc��������NspP�D�d?�x�ȓ]i, ��WŸ1̇�Z)�Յȓ�"�z������࣒G��V�ԅ�1� ��#׷~�`�EOp�u��'A�#S��@GR�;��V�/����<�>ᐦ؛7�ԣ���(ɒ��ȓ.���)�kH�_�`�k�+�"D}VU��C�ހ���R"�����Z�H�x�ȓĀ��I�?~T�"��c�a��S�? �U��A`����
ã@���"O�1�ܢe���� ۆ"�!j"O�a�׏S�T��L�ƮU-L��!"O�@1Rn6p�"yS�]��2�+"OB !�E�o@npbTc�,�� Ò"O���&46���#֡�8y���
�"O�БU���|�L5o�*	�:��+:D�`:b`�xf29�s�Z�bw��	e$.D�4x�+W��, �K��P�U�!D��"�"
L�ڀA��*�P�I5D���R*�����d��Z
��a�3D���f�0�l6��6�UZ��c�<rjQ;+��mrQ��+#��y�e�h�<�f*u�>	j4-*_T�l��
Dh�<AR@ޝS+Z��Щs�Zm�MLe�<���Z<N����&�`%�-y�<���3�����]��ȰtQ�<9jK�{�\2�$p�8A(�M}�<q7o�
]�pӐ�W�B�����Od�<�!�__|��K��w�㱀[�<��k�~�jP)��(��'�JV�<i�/�/)M:�X���$AfA��U�<��`w��iG�\�E)�C h�O�<�BJB#7�A�Ďم�L��R.UO�<I�A�$��qGA� 6ԋ���_�<	�+˿<����_�26D@MH_�<�U�H#"�6����eBz��7��O�<�S�B^�M�p�Җ9�ly�i�J�<��M�z�0��M�a�`Be��k�<餆X�T'�8;Pa�#T�����	h�<!�$��,�v!"Cm\�9d��ص�l�<)����b(e�ǘa�ڥ v��<17IX4U��x�M��{�hS�x�<Sm��UY܅���?(�,��E~�<iA�ڧ W2��1���4�0Y���O�<I�	�/���!�"-2aYR��O�<f+��c԰ ����	Z��a�L�<)j�V��M�C 	Pl�q��K�<�&3q���R��\� �O�q�<AҌ	#kb��!
�O[`%��cFm�< ��szz� RK��(��u��c�g�<1t��l�\0w��".p�{4�`�<)pE��f�(sH�1Ld����TZ�<�hK>xu�t����]m��r�_K�<х��j.��h�ɕI$��&˕F�<�*�*�TYD�ãK�L��,D�@�F,ϴ<��� �����&D�K�ޅ����cD�6�� �Q+!�Od��M�EϬj�^��L}�h����E�<)�яB'E�U��*+
M1`�3D�t�R�� i��%�d��	n1D��i�AQ�&%"D	�����׀-D�Hɑ(�Vۼ�h��ȭ'���#�i)D�t;��Y2;���6���$D�Ԩs,�\W�(qq��gM�]p�E"D�H�ѭ��x��)��Z�Y��#5D��##d�"$�Q�O�^	؈؁4D�@H%dȣpLt��ƈ#���7D�Y��J,V&~�I�I�V��B�`5D�\�@� �E�b�W��x� ��*6D��� �G�,P�F�̨(��]���4D��zR��y��i����y�y��4D��Q�6X���y�EL9 A�ux�j4D��R+�0&��·l)(� ���=D�� ��q7"R&_|����@�\�b"OŹ��K5�E��E�m�.��u�iJ�'A�)��|¤:Eg��ˢ!����B�����O�㞼�O\j�(D�|�@�� ��7���'Xr�!r%B=��5����+�NX�	�'����̔J>�b�����j���'�~����C� �h�!2��x�0�_|�<iǋ4%��������ޘ�6�T�<I@Ǌ6||Ը9�N3	��K�x�<��o�� �ӄs�:MI�C�[�<A�+ŵ^	 -�V��'}Ԉ���L��p=Q O�+�+'қ��Tj��EE�<A��[�5� �!gh�0:(�iF�<iѩ�2w�ȼҶ�+I�X�Q &IE���0=������U��Kǁf~�X�#cA�<��d�#.�iz� �s���r��V}��)�'��e�ЃL�mL�A��f"�ȓ%���r�];��E	ɳ(ϰC剰��WFM�������'xBB�;��1�'^$:��h`��$6�B�I!���BG�'$��1�&lSA$�y��I�7����UE)E��-��H#��C�	'��󔅒�+��z���r
B�	Yc����

\�q,�%W�C�	-F�`A�G�0g�b�	�@!n�B��n���%��Q�*
6�Z�p��B�	�B��%E�`� �?�R%��&/D�8��X� ����u�A-F]�])�e������'�����9"�H�c`L#�=
�#D� k%`M�'=Ba�ࠍ�Dx�cc�}��O��S�3�M�}�A,IrȀk���9;�!�䏏5�d�v�ȓl��R��X�!�`�<���aW	3k��A5�Y��!�ϳ	J|e��(AexD�X)q�!���7ѤmRě "N"Y9����C�ɈC58F�!4(����<^C�	fT�Hd/E=�D�@�I�+�dC�	�U�P!�A�n�p�������B�	�#�*��2HPVp(��?��B�ɴ0g����ˍ~�dl�BU�w$�B��<$Δmu�YI:,�%S�I�vB�IUe��(@��lS\<s@H\�z@&B��t
0K��\*�
���ٸC��B�	/1�bp�ҁ�����n�`��B�	�uI�q(�#��,��šَ/�NB� ,Z<r3*J�A����#��?�JB�I�eR��{a?~E��@=(�B�I�U��Pڤō D�`�g-y�B�I�j�|��7�O���Ц�\�DB�	��d�ڒh� ��Q��I�
B�<�>=����{L A�%@(w��B�	�� ��C�X ��P�����^C�	�:��A�8$���!gݢ`�2C�I�P&�p���@C�T3�<`�B�	�dXpm:�E�7/�r����	YtC�I�oZU�,O��T[�c�&5"�B䉦/����̟85��s7׺x	C�ɶl֦��7DS5� �U�E�C�jՈ��b�Z�^�K��Q$6�B�ɺ?�\�3��] '$Pm��J��jB䉸�my �V�h�0�{���ev�C�	u�FA�E̳o��Ъg�6S�<C�I$����:�v�St(��[� C��CS���N�;+��4�"�'�%"O� ^��vȘ�^�,QVcӟj)��Q"O�͂4���wX���hZ�Z�,y�"O��{VkھMB���D�u:����"O=!Q�gg�$�禀2I:�8�f"OL�3c��P�F
DTu��"Oz�P�H��I(�,C�IQ e\�Ы�"OL17�9p6p��Nu9D��"O"p�"�ӺT�]�lA�-`(�"O�!����c��A�Q�X7AH,D"O8��cnGR�V�h��=5��X�u"O���fԯ:��|��!�
 0P"O�h����<�8��M<AO���s"O�Dҁ��`�t� 4'�:�b݀a"O<!Ai�;	��A�s�h�W"O"L��@��D��
7���� ۣ"Of�%f ��r�k'A�8_4zp�b"O���hӍ�.%��P+H�t6"O�l@T�W�h3HU�&���9(��""O�����г>,�<`#%. D`�"O<�jTb�a`���C��H�j"O>�z��'|�Θ�`MH�]��@c"O� ��&/c-�y
s�8ax8h��"O9��i�EXcBn��H8B	�'�~�Q5e=�� ҧ�K�g�
�'�-���^�t�ʱ�扥,�Z@
�'��#�I��V�6��I�;k�ec	�'�6i8�W�h5Fd�iz�	�'�`��I>_=��` Z�u}b�@�'��DkR��"�� �V��>U@y�'�@q[ ����8��Ht�h�'��y�O^Y�y)�k �I��ȸ�'S��"S���h��СZ�6)�42�'��M�dL�5�H��D�G�x.t��'�0��\�3�$8�	��q�Z!��'��I�o�=B\��k�c�Ԁ��'Bl$4 �2 ��1�v�B.Y��I�'[�\9��r����L؀q�,QҎ8D�D��jT'I�Ĭ�GלA�<u!��6D�d���,!��-��U�&�� 0D�t�@	��
�A�U�(9!��/D��R���I6`�iь�~��7h3D� k�,�6/��IX$݇p2
��#B3D��*u�OR
lh6N� ��1D�p ��P:;��!dM֊ud,x�B4D��{Q�I51�z�3v�Sg<�q���%D��IF�M�)�h<�􍆗P�A�$.D������P��'�#g��H# D��q.�%|2�T��lĂm��eІ->D�䱲
D�z�,qqGFC��y7�7D�L��FP8e��T1fX5����(D��;��.y2�Q�ܣm��362D������4%SriM'%�(��f�5D�ȑ@���)�}!�dM�W�<�I1�3D�8�2-����pS�	L�OhdJ�j3D��qW�;k=��!!m	��4@���1D�`�sU++���"Ǧe���r"�-D��&��}3 Ʌ�m�Ʃ��&D��c-$9\�p�u�Ȭ~&�d�C�$D����ƒ5ɜ��:2�H:�EC�9!�$�y������f,xUAe%�!�S�S�����*v�h9;�c�v$!��R)c�������aM ��$�
l!�
�I��1��rE��{��h!�DK�hY�$Z�'���P\+�]�x�!�� ���U䐳a� �[��$r9l���"O,��N��N���J*/���"O�J��?���
W?~��l*7"O|�T�ʓj(X2�
�����"O4|� $O`f|P�/
��^�Y&"OFH�㊔G�q�����H:P��"O��	A�Id�R\ 2yc�"O"L��͚wj`@�����n.:��"O�a��IwX��p�(<2&���"OX������	g�$8�Q��"O�a ."Z�u� �6�9
$"O���&_�f��}D���a�
TS�"OHJ�� m����-�&f2fj'"OL�� SRîH6��5v�Q $"O"�Z�.7�N�pƪ[�l� �"O�l�r�R�;OҌ����7�ҕP�"Op<�F��%.$uhQ!ڐ��oKb#�'�
,����<7��̱�(��c�L��	�'I��OKCȊ����V�e�(,	�'3R���	��r�ܯT�<1)	�'��+��ݛ%�����2IHz���'
��(^�xƂ�c��VN��P�'�`Dڤ���_T�P	���K�bdp�'��D�u��2/��+/ĭ9�(�B�'�P4�%�Hf�R�H��ݾ6C,5i�'�KB9w0)@�5ϒ|!&�Y�<A�ʂ�UFB�ȠFF� >���,^]�<�0�C�{P�J&��2X���KG�<�0���}���WkH�~�k���|�<��mj�9e��;�as�*D��`�a����0��2�����+D����e[�&�nYSp�$]V�@t&D�L10�V(�ts�ͥvP4��s�)D����a6j(6�ѵ,�1n��0G�3D�� ��n���6'�	q��d�Q�0D� �n֛�La`Uf&�ظs��.D���C�}|N�rЉ�d��B��,D�\0�M��:s�ʉ'��;!�-D�%kU.~?�h!��˲�8kS�+D��;gB"a�
툷���,D�lIb℔sv��D�ĉk�l���-D�\��"sIke�ǆ)X��5�I=�!��Dj0���=~�E���)z!�ޔ7��J�EW8"�"�w��~!�$_-1��Q�%��h{���ie!�P�`�dY���^|b� �p�׽Y!�C7X�L�abH�.hX�!�D�Z!��u:Izbɉ�:Xf�AF���!�ܣ.����sDһrB�$�#Ǆ�!�D�$Z2�9b��:DnpB�C�!�D"�|�3�R�'F�@�a!��.�di���Ar/����L�J�!�L�g����i����4)�"��3�!���� �7LE�Z�$|�f�zE��dI���! $-T8P����ò�y��!F B#�88	Bt���yR�V�f;�8�M��i��@�H���=�$-���-P�� ��EL"?L��R��#�.�"�"Oܨ�G�ii�0�ό �-b��ď��!z��M*~'Zy ��1�!6�aS�f�ujt}�UJ��Tu��D�15�
�E�9
��[ҭK<9r2A8���r]"��j@x?���"��/����;�b�2R�q�Mj����2��م�	D��`��V��)����WlZ���T�\�|�W �"��Y�����djˮvR��@̑��(O��;�n����X���*���ӗ�	�g���3m#h?^6�ŕNP��k�l~�� �%����K�8\ʵ��Js
�����>U$u�DJ��]za|@M+}$ zvʐ��h䓂��Mc� �C�@����O�i�7�@U
�@\w��$p�cx^�]λ3O�T�1i >8���[�A^3d0�ȓP�0)� ڐ�KѠۏ3���A�]�b�b���xc�P�W���8�Hڴ�v��s�Q*��P�W���y��QM+�O 8A��Lo�4�r+Tdl�HR�J�7.dQ:��_�*�\� �Ə&��Y[�v���S��O����d�7j)VOA{�Lɿ�2�!�� /\����$���+f��F�bl���t���Z;e�|�#aj�i�:1��N'r�{p�׿����&CS����0bW}~�m��#���%�$����R��}QT�@%�4N|�>L��*T�)�d��u�ȡ+F+��^��X:9@ ��s�����t?b��s)��e��p	��yG�Q��O�$#�0I�$�3
ÓO�����fW�%H��!T!?S������bf�ʑ�?:J�CŚ�L���ش_7V��G©@}�HK��_�p�@����G�FQ}8��C�	�lP�4�To(�z+5�,���Dt�a#P�ͷ7��(�&Hg�>b^����F&��b�Al�3N����-�%7���ӌ��?9�T�w�6Q�ʝ
)b�8K�(Ե�8]0���\�O�
�Z�b�����A^&	��i�;.�xX�rj[� �
X�`M�2�pa�I%)��qX2A�K�t`����\�R*ۆ!� D�ĀL�7��I��|�{�G_T��8hE�E9#Q��ɿ&y��i�Y�@-:	*����D�J�E6�R��9FhP� I4a�.��6�1rԀ�lZk*u��PԶ@
�Zp�'�D)����k����GL��|��M<	 �ϙ���'���
Y�Mӣ �s���20��n���n�����H�^Ԫ�KM���=��k�i���("'T�/�����Tں�9��O�tY�E�n!��޴r��h�G)��<��M���ӖSEfEjpF�1V+����X�_�#?9���(��i�(\�����@�~$��i@0�ؑA��hx1�f��O5N�bPbѳ���	�g+ P�g��X�zm*o+/t�I|T�UZ�����Y
	U1�$��%g�	�1ٓD
�m��k]�YtH�c�ݒ�M`��%	h����+rK�K��$܀^�^����R$��A�Ǵ [�	��K�;-�,Q�Q���4zD�e\ \�J��̓$盆Æ�j	��C�
^BU�f�@��z4�t�D��f8�`��k��yb���h$�0��4|j���?�Q� G�j%�d`�V٦e�S'�"%/��'{z�YR�R�8��'X:�N�|��|���K�0cd�JU�؇6�����⌼Yu.�B��'�t�j���,���.E>**�Z�+�+.�f����-�P����R�������>X�����,$�b���*-�r��%(�>��L�>�y	��ˉ8*N)�hCǦ�+��1)-�i1�'�q�Pi�9uz(�;mYB��
�*F0|B���&�\�d��Fg2�#-�!$}� a�On�q4��8��z�!R���O��8e�-�� �O�R��Q��HH
P�R<�b*%�Ll15��M���E-D�.��-Hڴ,�h9�@�Q���=�2Lج�t2B^������*��Ɇ�!f0du
e�˱b����т�E�0kD�z�a�*ۮ%���@w�N,o��fJQ�Ճ� 5�6��-���wh ��M &z$�If$F�o������7e�� �<�0B�A�2�^@q#@ѤRv�����"< �����)e�ǟh�j�ガ�qO��Q6��Y�bT��RzQ��*ʹ7��, ���1J�/KaĨ��s�6�p��(�&��fnS�a�;$V	*V"\�<2�S�,Kf\�ȓ2@hJ��r֮�5�`@2P�a��'&$&�I4(�nYx�X~���O6�I��օ6K�	�p1��"5���l��K��<$��c�'D�!V�A�n��]>��^�&�8}'hFB7���!_8�=cZ0y g��@3��GyReD�F���G��IUvAۤgH�ް=3�J.i������x��ٹ�M�T�>0�ȗ	'�VA���'���PůCCX��`b+�&��(1�N�>n�@%(-D�p� �X�,�a�폍XM� ��g(D��%�V>��#-�5.x0�p!�)D�@(r�/I����jj�<]r �&D��1���0w~���DGA;GbF@Q��3D����b��. �<����
�d�,D�ܸ�(�� ��g�9
R2�S�*D���c,�%ؾy�$d˨Grz���=D���"e;��O�vH (a�=D�t�؈�ny�V��Q
�p�#�x�<���G1R�܌�w�C��.�I6��Q�<9� V�����A�V�a�I�E�<iCԀzB�LZ�.�6K�ޜ	��B�<Ap�Q.)��4.�K~x��/[~�<1�� ��t��Vg�R�� �f�`�<��L�a�e�`e��1�'��;���n��	Q�@Q�$����':L�sC�1DU����'���'(��`@3wD�S�T�� ���'�4�d��L�l}�"E*vN���'o��&OJv�Z���鍹�:`���� �!#�*�g�j\�M�G����"O�]��$���>�ӆ��}p��"O�`���K��W�C/B<��ّ"O�xʓ&�0>$D%�� Z (^���d"O��§X	c�d�!��:V��@"O�27��J��B6  �M�:E"O�����E�L�PBa#q8�ڶ"OxL����E�t�zT��J:��j3"O����+��eA�BT�ZD"O�!9�HyTN㴀O�wm[e"O� R���_�a�O��<�J�"OT�J��M�X��`�FU?74&���"O��Д0[��t�7��� �(D���#��=+ɞ����P���$D�Tkq�S�v(��,C��4kǅ>D���r`�;���E��+Ai�XP�':D��`��8���ܣZ �wJ:D��I�}��]@2��+�$�[։8D��x�iZ�੩2�VH�pp��G9D� SS$�::
��1X�9`Pa�	Z�!�$��^p]AQCD
k��tǟ?:!��3M�p"����AQ e����6>l!���R�+�<��� ,޹�^�*�''���&4J/&�s��J�p��}:�'>:��4X-���F/]$>�����'`�%�c@ջF|�5mO>.`�1��'\���7����-�Ua��$�T���'��CEUP0՛ahU� ���)	�'�r���\85�Z��Ļ 
*�S	�'���D�ʮw�:X��؈�ruP	�'�`�r6͜U��hqw���'��	Ŭ/?������L�X��'�q�sI�-������y��9��'L���FM�0K$������rI�e�'� �c��%lMH:�.}ঐ��'j�[Q�Q�Tj:I�G�Z5]M��:�'�@-a'@�q>���&D�KO�!s�'ZMx!���VI�dǫ��Ap��[�'�  B�P�Xب�Ȍ�(s��
�'�Й�lҬ;[ ��3N٭ŖD�	�'�&��n��]hD�m�]^�	�'�|�ݜ<��q�BF'IԆ�S	�'���&̒fB~e��*�D��`��'�)�DZ�*m�����ĉT�2�A�'�T��@@�k��K�h����'�.���,϶e�A��H�
�Z՚�'��h��ը4���� ���PZ�Y�'�bE�S!X�qqM2pb�yഄr�'� ��AjہkRE�wcF1hIL�
�'u`��Gfv�����(e�~�r�'�2�򕩂�l���p +V^$�@
�'��@��ݜ6R�����bز���'zHTʖ��*G�9��(��_qnm��'d*i����4n�h��łɝU&X`*�'p�� ��Ǽ �Y��!Y�֌�
�')��3�o�e���TI�	�m��'|b����R�m�ȠcU�ɶ����'�^�t�e>p��q�C3�<x�'�pEr���rs.y���R�blY�'�h�`$����*!������'Ů��t%P�l��M�У�?����'��@�e���(y`(�5
���j�'�(��6k��QѪ��T�T(��'��	P��4N\0{��K�xy��
��� b��d�N9P� ���͒�B���u"O
M��k\�K���(���=H�
�x�"O�Ÿu�ͰVvpYƭ�Q�z(h�"O,��s��5M�@eɳk��N��X"O#O[�-���J�*'o�4��"O&�r e��M�*��V�3`~��Ia"O��	U�ӑE�P� 0ǔ�����"Of��#�%p������\��.�"O串U��y�$�s��>F�D�Q�"O��ɷk�`�0P��� Hհi��"O�X�-ǃI ����h� �v� "O4i	$L��RD�s���sIf@��"O�Ð��L�"e�a2l�"OD�i��>-�R�)�]=A����"O(���m��8"sJNP�(	��"O�؉�%�澑)��͢0ʪE`�"O��{��G�d�ݪe��pT��@�"Of<�rF�zW
�w��4C
,�"OhMr(�99Pqk�Ό
]J��Sf"O��P��]�f�N�:P&�X1��c�"O�,qR�L�4�������9��R�'44�j⊇�]�aS�h��%�dp��'������Y��e��:'@ [�'^ę�7���d[�$]�l��Z�'��0z�b̚r��܃1�O��p�k�'	���3)F��:���MZ�swX���'��-�EA4"��b�&�{1H|��'������� T�BRf�ά!?\�Q�'ֲ<�0MFf~8�`��!1���
�'PP����%�^R��
8L��q�'���b�&�*�-W)7��ݩ�'��eY�#�������x���H
�'J��v@�0p��|��8	�'#�x���.<}5�<i� ��'7&����5_y����o��H��'�nU�T��/�ɓB/82A�e��'h52ՠ�^���y2m�9 6&��'�`��ba_���x�R�+����'�\ݚ��ȗ(�m���8��!��'w�]�s�H�e2�T�$#����'�)q��E�T�K��ޣ����'��@	X�Q��d
���'�X"@��+ar�0p�z.�QI	�'�T�E��s(��ep�ɋ�'xx˖�ς%�:-PW�� �����'z|�윻6��H��6!����'���M�h�j�K%�ټ�Hs�'!���	�|�Ԅ�$��+�$u:
�'�a�&G|��-�4D5/����'t0�CT��$3�94��+6_�-��'��E(�K�pSnu�C�ݼ|!�1a�'��uh��y���s�4�&�*
�'v�0ů�(F%�eZ�c̯{L0�
�'� � ��T%c����!a��P�nX�	�'���"@�c����0�YVG*��'��{�郧D�J�^H��(�'�CgO(��s�-K/9�61��'��ڠ"C�}к���GA�=�H9��'�n��u�X+P.z8`iB�2�6Q*�'�QKk�(9�����D.���A�'�A�NI.=,�E�V@���l�
�'i ��V�L�7��-I�K�A���b�'njl
���N-Y��X8(����'@��qU�T:v���)�F����� v}����1,�%qWF�kFB������(6�����ɞ%\$��cn��wϼ)�eFZ�"a~2mI�(�"�����b��	T��Pɑ/�j�5Q@H�!wZ��P��Oju�O�Q��AEH��K+�N�M	h(�E�>ړz}X�u`R��~�i�G���듺�Hl�Ɋ�&�A0%2;�ar����ta!�B"a|BX�P�Va,�%!�˲�Mc�C�+�$���Otq�o�15=�bYwAh��'h
Y��ϻ<R��[�G8"��8X&A֐�ņ�'�}��S�v�2��eH#��Xa"@�5j�,k�)B?tT�qR��"�u�;N��i��4+E��s��aQ�1P���qW�x�r���.�Op� �f7.8Rca�:D�|��!,��q2�A1X���W=7�����x�&)���O�8���B7]XO` �&/4�Z]�JF�th,z�I;J7�I�WA[a��;1��t�7y8�h#��nȼhA��X���<R��ͷ!�ȝ�&,�E��Q��ώc8�lK��h�J��a���B$i�o����-S*5:��i��%�ݹV�P�+�.ם1p����"�*Ex��q�6}�l�)BE�cZ�
&G!@[u�WO�=9b'�;~������=[j,@�ܒ ~��#g��Ne��%�g?�)'~���#���7|���s���&��*
�L��)Ix9l�Ђ;�Op�����7�a0��!�JM+�iٍAr�=��)ξ�2��4iH,���N��M����6�UM�&f1�A����fڲP��RG�Ǉ%�j�t�:�k ����ԅ�~�dT,��M0��DI��K�;5l��!ƪ'N��@�'�p�C�Α~v�"�Ͼ�ax/�z�1T��7��-�ƭ��yBhLBwN|�'2�9�c>]�1@_7>��(����N�<�{7�Ԍ#�q��F��!�$���+a��E횵°RdmQ�(���߸�^�z��i����8�K�=ܒ�H�K�5!�d�1㬘2��3��bh݂L����v�愑�H���)�'Nq"H�ᢏ��%	 
�`�fc3D�{FE;z�}20��C��r��2}B�P&:;�|���Se�,�'ݩ-.H|��댞v�~0��o�����D�
���3?Ʉ�Yg���=���)L��}�^��,��/� �Kp!߿5��,��'�0�0��C�r���B�nC\U-S�� ��	I-,U��ՠP�4�0�)�2E�t���������������8]�G�. ̠���]E�]�@��Z��l%z���-��@E����(4����S��13�i�n8��S)��еj��9c�<��Ó�M�}�N) ьR�fDz���D��ɉ��P���H&�+b��)4h�=|�*TR��@30y����^�b�*��'¤F�,+��C���"O"}�$늕�2T�୛H��]��i�nA��W�o�}��>I�4u��	�)'���l�`h/��J��U�UK�^�L,� �,bC>A4g��U�^	��'ì��b�߄ 9
X���1C��q�lʈ,��up�C�_4\#d�4Zɢ��"K� :ll�a�8�9�m`���-_r���t
�r�J�1��'���(�������O`��[Հ�Y=u���عh?���!E�J 5��Ϧ�� �����ݩ �b�&�P������p��aյi��`��7�|�$�Rb���Ep<���5Ez��gK�-!<T1���ӋC%�Qh��ȞKRʱ�#K�3
�.�X���a|�iՒP�)����7K�L��uO���MS2�ڣ&W�l�F��O�{s�+&��-ZZw_�A��J���܌λo{���J�V��p��M�1*��ȓ{J���բ_5qUD\@�G��ɹ��_*\(�A億VԐAD�]�xO���5pQRM�P�]�
N�D�rl°�t;��Ŵ�6��D�Yf\x"� ��c�/Q�\�����K���!`�0���%���Z�<'M�3���ұ-ȺN8��Z��Lr�<�c۽�txr'i0Q��  6
Zǟ��!'v�a} Ƭ{��L�e��\��C�H��y�΀�|j´`�fs֜�૆;�y"㍌I� �#�#R�Pȇ	�>�y2B� G�N�W�1IH������yп|�(Y5fG�E�8����'�y�*:xb����8SvE����y��ݽ�uԌ�6������y���idD]�"�M�/�^��b�:�y��m�.�Z��R�/���	䄎��y�Ɖ�>r��WK��1Mp��v��,�yb*�?w�zU���N#�d�`Q�ʸ�y�1nnP�ɲ'?"� ���y����D9e-�r	^@`�*��y���(5e��/�C4�y��B��y�O������L���p���yBk��D�X�3��5N��%�w�Q�yr�3X��h��N�VTӴ���y
� �,��jT 8�N�ir��b@M��"O^ �p*W�9�4)^6x ���"O�q�㊟4(��z���-��|�"O�`��o�N��-��fG�w�8<��"OxB�Ա�а�Ę�3"P��T"O� P#��+7����)E�Af̹""O�ț�D�#(d�5HM%�y�e"O���jA�~���ilv�9�"O�8�T�]�sY�!`��L��e�"On�7h[�_=b�Q��
�P{Z�Z�"O����S�LB(�ҊE�*i^\{�"O�@a'��J�΅��*/w7��)`"O�)� k_�J���sh�i%�Y�T"O�L°�� s$ܔ��J�n��Re"O�鱠�Ð �0�#肤[J�
r"O����L��n�	��Y[���r"O�l��瞒l��H$+��-�2��!"OLZ�(���ZH�7��@ ��1"O���V���"1�0�T�5�aX�"O����hZ.\�8+���I,T��"O��{#�/�]Z�d���$���"O�fg7d��ջ��>[��)a"OV�Gjs��BT�޶8h��"O�q��HK90�B���`؃y�>�x"O�9�v#��"tD۫ �2e �"O��Jܺf��ش�@�}��9�"O��y�Ie�D8�F�J|�0p"OfqsD�����`���:W"O�˥&�3[�LQ�R$C��P["O���%錞l!@5[��>x�@�a"O���V��F��Q%�J���"O�JU痊l65`A�zZlI�"O�I{3*L9p���I3�"��-��"O�a
qI�x
�Y��AY@�Z��"O��z椛>��%yi��M�*�B"O̊SHE==kW�Z�w�0��$"O��Ӏ'w�tuXu���]r��"OH�9�酕#Mj���X�`�1"OtT��غ!Lp<��
M����"ONT�3'�L{���C[�5(�3"O>��"��
�\��r�Ʈd(&��F"Oȡ@��կs��+v)زN���zP"O������s�F�`���P��<�'"O�K��ΝL�p�R�OE����C"O��!L��9xh�'�)�-��"O���iF�7?���Tf�$G�p��"Or�*�]�0�b �����Nd"Oxhˆ儜j˞���ANtx�
a"O0dx�d
�x̊��T t|xdY�"O~����ɽ�(�K�\O̥��"O�젧��#0wLs1�I&�u��"O.�V!�1{�b+	
l�0H�"O\,HԦ>> u�*�, �|��"O~�cDQR�b���Ȕ�5�"웠"O��4���ȉBF7q�*Q�"O,�`���}���e��^ĺM٠"O���a�W���RV�M5?\n��"O�!�R	�W��ҕb�:@;��ya"O��"��T���Z� R���"Oj���E/d����L��P�"O��j!�Z�{5�� �����N�"O��BI۶FBL��2��#S����"Ob�@�l����:V�Ҽ7��Y2�"O�����@f�HxfQ�B��5�a"O� N��*�-bX���%t�¼a�"OL�b].6I��!������"O��9��V�`!�b`�މ�1D�d��́�$��� �إ6!��C�.D��U`����� �.�}SA(&D����OH
��ě�ɕ�~d�TB�$D���>��(���4´�Q� &D�<d�כm0@�3da�����#D����
ɵ�x���@ξ2��E�S�=D���SK/Ob�pd�C*EѪ�VK?D���Qʓ=}��8�Ƅ�rE�Qɖ�;D��!���\�0أ2����< �;D�L����~� ի,�![��ڒ#8D�h�f`՞W8�ܨ�MN0,~д�P�%D�l��f�&/�������9&����"D�d�I�) .!à�+lh;��2D��J���j~^U!���A�|�C�1D�Ps� <,@�f+O�!�<�Z�a*D�Y�D�-z��S���W�{�F)D�4���5@HU9�(�:Dh#�(D�|k�L�;�j]�Dh�:dʴ`�`'D�T[ãI�.��R�P:A��,a"&(D��w#O�9^�`�ÚP���7a#D�$������2��O�1̂)��/D�����g�|9�Q��x'��dG�iü� �֣��t҄}�lQl�O�09���V^��2C-ɻ`�J�1*ӓyOlO� ��O�*�Qā�t��ݹReݩn~ȍ:!�"�:S���e�?1�g�*�SB�N�3
�Mn�P�q!G�{#f�.1B����fH%p���O1��&B�B�L�aQ#NsyL�rVf�\�&���u�@9�甫gdtb�"~��Ǎ�At4'�@�8+�E�T�.}ޜ�dC�S>�	����)�C�� �#�C�q�b��+�c0�>Yi#�C���R��.pmHe@C�ĉ�plJaHS�OL��"��D�H�\T�"AD�7��A`�O����e�n1O>9�E�J�X�%C�5¼�fL~��q�D� EY0b�"~�!��#����'��ŭ�J��� 坑�����O6T��O����X��З��!lDA�V-������0�"� ���bS�ԻGh!�DZ�_�͓�%ԑMv*B,S�L]!��~a%��!Eb0!ߥi�Pza"O��S�$��n��W�ȦK�s7"O��� �9dp������-m&��u�'�qO�t�����Q�iT_�I��"O��W�ɹ�Б�%�D�	�ʭʤ"O�=����N�0��%��0ED�"A*O��2��JC�.�SFi�h� �'�z�A"Į: �˖���6�QB�'�6<9�oӓ%�$P�ՠɊ.ԼA�'u��X��V�S�F̸6'�-)�Z�j�'��Ɇ�3`*Aqfꂇ��$h�'A� ���US�XI�b��]����'��̛�剌c�`����Q<QF9p�'j�u걉@�W	��A��,Vhf�{�'ذ��/�zt��� ��zZ�r�'PD���L9,��R�a,���'U�Qr2N�/c�"y������8��'�f}�w�	>q�M���M-�r�y�'0>�j�H/i������)~&���'�8�PHB��r���LS]��'��`�Β�T�ҽ���Q!(���'�)��5���4.D2M�vk
�'�nybt�ԃ^���e��Uoʝ��'"� x�� &Y��|��V-LU%��'z��PE��XSP�z�=k�l��'���^���-�	A�s������ � 3�i�'����F�v=$�U"O>H���̤%�e��A�*@�BP"O��R"��=&@�j�F�N$�X2�"O�tqt-L�)5,Y��J*�]�e"O�dB�޹��}!�E�:m4���"Oj��g!�%^��tyTD�O;�t��"O��ŀ�96�� �H\	,.qa�"Oܴ �&��+�H�q�HYw&t	�"O�:�m�W�T��&ѹX̘�"O��K5䌙*��z����)F!�d��,�$p���$�M�����&�!�č�[�H�q&�����/j�!�$�8 �Z&�K+&ьQ��!Ԭa�!���d[�,E��`P�n����պ�'E��a[�[;H�u���x�
�'@i[�#_2o=��9���u�L%�
�'-��K���!_���D��`�>��'��L0�`ƵbP������^e6��'I<�I�&�2��ǅQ�n&1�
�'�,�JUF�+a���iS�y�(1��'��h�.n�$XvDW�c��X�
�'�*ك��@:VJN ڹ\����'�tX��?-�dq%��("�h
�'*���4�N�enZ%6Ȉ�z�X��'2������ƢF ���yk�'Ơ	�S�ܩK��-W����s�'��D�Q�Z�Dj��F*oԘ��'G����H�~�BT@�嘿mΌ��'�����m��|��@�ct�"�'���Q�4n�P�@E�`h��[
�'��q�AEٞE;~H �	�K�F��	�'�hի���5�6�A!�)�F��	�'Ϙ)���"YD�лā���9	�'��AȖ-��N`]��݂�tز	�'v�����"V�>��vE���2��	�'N
�S"��.p��ٶ��l�j	�'+�I�w@��r�H�ФI ����'c2@�q�ÓF�l��b��&�s�'���B;���Yw�Հx	�'�
x�&�݅REo��|an���'�
�xt ʼ	^4�:Ǥ���T���'�|�5��9N8��# ��� ��'��l��ZvrȀ�`@�.�J�'Ǯ5R��[BGVPIĊ�hz��	�'-FD���/:�6$#s*�lr���'�~59�C�%G�<���DV�j����'N�;�+ډ\��X��µbȂdz�'����@�5��43��D����'����C�P����re�I��t��'�4@����t�,���W"s��-Z�'�J�Z���aѰ��A��Z��ɰ�'��]���c���i0�6�2��'w�}�0��PT�6n�/��p�'L�	xpH�Up�9E��lg�m#�'�ft�j��I�\Y��jY�.70Hy�'$<�� X�&}���F�'.�2�I�'��d��A�,<����64�"� �'�� BʩFY*��f�}}�UZ�'u�B֥��x{@��+~)K�'u�l9�Lo�N�д�{�<���'�����D�"XpB�#��A�(�Q�'\�k��^Ȩ݁2��*I����'f��3�A��y�`�:󄊔m�r�+�'�|��4a�C}����'fJR����� ��	�b�����c�>\�PȲ"O�|��F��@���ˁ`Rr�h�"Of��^��\���[#J����"O�@�"��B,��s&�d��$"O��y2jɚH�ɡ�d�B��@yS"O>x�bI
XanzVmȖzӸ� "O��B�h^%	L��b,L��r���"O���)4�|���Y;�-�"O�ɰ�a��|p6BÀ/t�pB"O�i�G��]A�,�B��VHp�"OH\d� m,���1���
8��D"OΥ�Sɱ|��m�'.��Y;�0��"O �ag	JR�Ect��F F��c"O>i8��(?�pQ4o�(4,8�"O���55���B��%$@�T"O� ��w�|�An�Ȇ=��"O��@�k�SS�k!�Ļ#O°2r"OBݑsA�3��%��*��o*��u"Om��*ؑB`��(�d�(#@�e"OuG�Ά:�n�+A�ĺx�]�t"OX�+�IO"LZ,�b��a� 8�"O��2�Al�]��A��LJ���"O��e����E���1FP��"OQ
��ۜfy|g�0	��"O��!ס�%kK��R�M�����')�B�&ھ���ɇP&��
�'��]҅LƗWZ�����Z��@�	�'B\�`PiF=,��僙�S��es�'��{E��� q��q%m������'!Z�"�-��-q5���!�V�+�'_��1�+�=����%���#�tx�'M���2�J%n�R�+�j͊;��
�'�P��d�Z��na��V�\Cf�a	�'���2F@�'yEl��	�<8��'�tu��IH}(�8zS����rD��'z��g�ܗe�$1�2�ˊm�LD��'Z8�M�9
�]`7ወZ<��'شI#さ�)UXT�k˺{����'�LR�T�eⒸ�1oNp�&���'Wh�S�O8K�p�̘	>=$m��'���[���	#��yw�&A�I�'s��b�>&����6�!�X�	�'��u�P�f�f5b��!}��`Q�'�P�zT�9cR�H�!J;{A�@��'����+D;;� |���J9|W��'�nm���7u��E���{��Q�	�'5f,����+������q=���'I �;Ǆ�(�\ٳC�'cv`�'�<�H2@� #��`�&�6K��q�'���߰[x�y�'�Y�J�Z$�'��Ж �.�#�Ꞌ�|+	�'V�3E�R)~]�z�m:w|XPa�'�����߈���Y�.HkU^��'2�qʓ�G�! l�E֚c�����'���B B�2Gi��u�0fʈ�'�0�rv�˨9�4�C�"�Xc�'?<hBE�O�p�d��AL�"�Z
�'����M�s�p@�[q)62
�'t��	���Xh
ض��'�
 g'�8o� HB�-D�;r(��'+HEJ�B!A�,�1"�.�6��'�TA	�(��p�X���E&v`u��'��}���onRL�� �-%u�E�
�'2�p2�cÕ-�e��'sܹ1
��� �����m��*�	[۶T0�"O�q�e��JP���^�D{"OD�1gI�Y�`��O
�4��8��"Obр����-�Cɘy�5S�"O|Ly�aQ��c�G��m��uX�"O��!%��5,�K�-^Ɏ��"O�����Au��Zt�������"O������7G�|�����"OF��A'ɻ;z���ͩI�M�B"O��T�E��[��V���-he"O�)CA��n���H�G�r����"OLiQ�F�K���C�G�e�&A��"O�@��O�s(0���%>i���"O�`t�Lx�\���Q�h���PC"O� Iab@%bq��(��ɫC��}�"O±{eLG�*���Ht���� ��"Ol��!�
^��h!̈,I{��:�"O��(��Z�J��P˟:irP4�D"OАst��]z�� ��"n@D��"OLȃa�M;�քk�.�E!��"Or�j�(I-KOT��El��>25" "O�l�c&T�*DKu�0]nZ�"O���V�B6+|]
Ã
�݋�"O����E�v��Q� b w4<��"Opi��,�f�ɕ@ҧ19TI�"OHP�#"��� JC8�C�"O�l��X
,5��!o׭x!H�sw"O�d�A$�E��1.yX�+p"O�%�"��/���ny�|�G"O���$ ��a-�2 ,���"O�Iac[�8�&��E�s =��"O�����v��(�Q��+X<!�"O��qp�ҹx��@q��lS�0PS"O�y�"�}LŐ�B�=Om�f"O|!��k�������%O�l[�"O�T
f�Ϻa���xb�Z�N�i�"O���6�I*nL�Qqj���D�"O|m!��+i��	jD�����M�D"O��Rk�-%�>yˤ�L`z���!"O ����q��šHJ�ZzX,�"O��zU摋d�ZY�DQ�AoH!#"O>`��
�a.z,!�	X�V]�w"O.�����3����	�WUz �u"O`�+�O��m�H݈W�!9��"OL!r���#�.�I �J�"�:�"O�!�v�I�q�9���#W"O�a�&��>Mv9#`�.�0��U"O����C�N��0�ɐ)T�h-Y�"O�u"$�����2J&6�L"""O�)E$W�:*5@�eBlz�q5"O4���%S$�0�e�Ԓ����"O!�夌�>�x��[�����"O"4PЯ��	�|$��U J�,1��"OL(�x����i�+B�2��"OVm�	   ��   p  �  �#  /  �9  �D  �P  W\  ~d  �o  z  ��  ��  W�  ��  �  "�  j�  ��  �  Q�  ��  ��  �  Z�  ��  ��  !�  d�  ��  � + o � � 	" j( �. H5 &? �J hR �Z �f o Lv �| Ђ ��  `� u�	����Zv	B�'lj\�0�Jz+��D��g�2T0���OĴ��eի�?Y����?�`�҅w+*M[�!E��$,�Ph�J�"vE�̩���;X�FT�����e�l���6v���X5E�e�$oՄ^6�aP儍�P�Q�&�5P@M�t�ߒ@Q�t�.ӏW�� �;V�L��'�?锨��*��4��3G����&_-5��LS�	�H3$���(�� �Je6��&q���Of���O���E:�����P�jG�� s΅�Y2`��O:Un��̔'�ҋ%�r�'��mU% ��ޓɅZ9bQD��u�'b��'�R�'��'w�b[w�e9An�(T�t����M�I;�(T�U2qr�\�%ƧZ�Ia~+ǥZQ��YE��:g�P���9F�̵�`P5n�J��'���7����T3ǎ͟u�zE�0������Z��0�J
�l�re�'���'���'��'��_>=ϻ1 ����_�f����ܪis6��	:�Mk�i6�7m����I��M�PBHKě�
W�L�,�c#ޛzp�c���(5�Jր��#=q���9�؂��>����B�8r�O T,J���6=�>Y� �+%��p8�������'r@7��ߦq��ER���u�C>�P���h<Ь���F�3K���ʙ>x��
 Z����z��ߺ|z�m�g�Ȣ7��ۦ���4W�� ��f,�q;bM�/F��[ūUL��u�ԢI�wכF�rӆ�nzѣ�A �nY;�_%@�v�� �%?0D(1�م2�=
ԫ�V>Y��^�>cnQ������ٴ;����#7�*8���X�fذ������aNB�7X*�e�чE����y��H $_�r�d1bh�,U�4�cC�O0㟸�V�#n�8ŃE �&@p��&,ӟ0�?A��?��J����?�+uȞPz���Έz�:}��k�O�ʓ�?���?҂I�(���'P�|��tJ�陬@�JaH�c,LZp�ܱCTN-x�Ɖ�.��Dy�U��[A�(q8N�脀Ĭ� ���U�>V����?o>�@6��!d���GyBJ�>���ey2��?{F~��Q@�-�lE�pÎ8�?!��?�K>���?*O���ڗ$��=D�A�4��(#tߴ���D�O���D���=���Oz�9O����(B�L6kx`;�'��en����M�O��ݶ��6�iWB��j��rU➍;>��b���b9����O,�ğ���ܘ�+R�3{�hsU�ؔKebqj��9��ӥ+�ҠH��'m0p��))t�.u�'��Xs����<��A-���S��K�.��]�������:Uz8�y�?J������d���O�mZ��H� �8��JQ䀛w����H��O����O�D<�8��\��C5Br�q����]
��G{r�'(H7���M'�\3ŗ;D�```� �>3�PP���V��M���d:g���I�O�D�O�˓w�Z���'Y��
4�P��@�((��*�c1{D�%������� �����$6�$�9�8�6�m�X��*g�2��(O�SJN	��!K$&�X�2��ǿǊC�'m���ჭ2�l1�ҥ�[���"�iH��,����	�?���L���"���<
�cB-�^L��s��hO?C���ӌ��NX�����
��	��MK�iMɧ���O�剰7.q�0+={�j B�x���% ��$�O���<�/�����q��@ִu�� ���!O���.�Af$�T*�Z�����O 7���`��	�@}��R�G��Y�(@�F�����©87� yѢ�4�E1�̓���8��	�Y�,�l����	��	=�q����OF n�%�HO㟴x��A�w�V�s�`ٻO�ĩ�����������G{r�$��:��7KG/$9�b/2�'�7�ݦ%�'�©A�q���db�Z@����Ĥ���uW�Q��O���?��������h���+��M�Å\�x���vN�i�v�ht❐<�2�x�ҊY�ց���tWOtZ�p��^�'��1�v�*K�>���$�N��!3Ck��ç듡&z0���0��ӡQ�pӖ�n����" �6@�'���8��Ղ�Vy�i����:��O�q��ؓP��&%� q��h�jl[��4���O�˧}����{#�9�#�^�@�X��
��6��OĨo��Oצe��_=C���'��tq����K��pA� �)f��y��L<>���OB��a��`� h�}���HQ&	���O)��1���b�ݻ�\�bL̤����D� 6�D�a���4Yf$C��B!I�l%J3��1`E�S�a�d�:c�m�J9C4h	�
����|��I��M����d�IC Xf:�8d��~N\(�s%`j�'|R�|2�'Y_��뒅@��P���1�S�J<�����Ƛn�ߟT9�4�?	�&Ui=j�19A�!##��?dn�&�'��'�@�3%O�� ���'��'��=YX�uP�ꓪg��-��C	zhD�T�3��ӵ��/f����Q>��S�L>|H��į��!1�I*ș3�,�3{5��PjO� CB@`�تS��qR�c���TP�b�E��i�z_�$Әw(|�9��[�Y�,u�ㅟ�H�� �i�˓.����	y�����tz��������W`D�[�B�p��P���O�� 17)V8-t��s�C�yfap��?���i�B7�>�������<9�7a�t0"��
*�D��Q�I�l9r�iGR�'Y2X�(�O8��7p�d=
���PY\��F�(M���a�A��	D�IZ4��(��C�id}k��d~ut3@�?+*vlX�b�+g΍� 'Y:��c2B��\���P�>�ɠC��%M6�iJ>�s�զ3ոm3��p�D�K5�F�l�.��ɜ�M�N�'.RĘ�2���i�L������?I����<�d�8h~m9�-��}�|1#��v��d�צ��I-�M;�i�� �Z�4�?��x�H� K�;o@�j��#V�����?���ĭ�?	���?��*:I�\z��2j�X�`ϙ-�� ��[&m�6E��@4�T�x��c��#U��u��$қ5(X17��O�F5R�f��g�>ز3#�4~��@#n��h"��LN�]�2��/3r� i�B�'�| �p �~X��FD��0 �9�H>i���'�r�'�`��^�4bEL�6#��[�
,��2	~�n��ھX#:S��P��s��o��<y۴�]9��m�㟬���<��C��	��7I���b:(�PtA���s���I�� I�bt,��2�S�r�X$�0�F&���("�,5 ��B������y~�-`����I��E&`��?��{��ԬvU�����"�N("s��8H'��O���#�'�?i�ǜ5��[�c�*��)9�k_��y�_9�SFK�DQ��C�2�ҏ��K[�O�@XRdJU�8��P�ŵ���'�i�"U��������O��D�O�˓E�bP�
D�|��X��،!�p<�+R؜�Q3��5dZ�2mG���I� hՅ�.*/�kO�a�o�>�Isf��?����f�� �f|��F7r�����~��,��b���/���2gU��j� z�b�l@�+&7��Dy����?q�'���|�C�.����h'H6؛���2$B�'���������O�����	J~����<	@�x5�'z2�dӞ�o�޴���� �'W�Y* F�5#)�q֓u7��CG�T�c���'6��'��Y��>��9���3}�>ȹ�A�M0l(��������Wnͅ{5� �c
v��q�B��'�(O���'Vi�C�
(4mx�ŀ�V��I���1<V�$�'��w6ʌj��*vơ��'��|M�Y���Y�f�R��Z}���W��꟠��4Y���DxҮ�%0�zЋ�N�U���#��?yϓ��'Xu"D��j~8,[w���V���O>� �i6��<I�=NS�V�'�"ʟ*NlX"�,ϝ ``e��3���'�(���'�r?���hO$e��w(Z�3�$�
"'|Y��)7L1���I��ӴV�6�?)�!��^N����@3x�Z��ǩ�e}mp�)ֹ� ]8�c�O2����e\�	�!m�[̓�	ןt�'�2�uA&'��,p�jVw2]�J>A�R�HB�X�&��9��Q4[B0�?���4�f��	�-�|9U�����2N�T���Ģ<a��ʪgٛ��'/�\>���b�ן 6+ד*3��	"	�U�
5�A��ş��	�	���XEH�/	 �!&-W39x!)�E��|z���X�^0¦�Kn>p3�����݌�p4���
�<R�P+ޑt���P YƊH�!���:�X!��	����Ju��9�T91��O�\mڃ�H���Ӭ��t`G�V�<�Q�j�Id���+�S�OB��%ƴAd@M�HR�.�tLɁ��<q�4n����DE�Z ��J�/]y��+�ꅬe�T7M�O���O�e��֑R�"��O2�D�O 睸bA���ӄN�0� �C׀��*w ��mL��R���r4T�!��#據EU�����e�hQ���=F�s�jތ0��L��e�d�xp'й�4�xa�\"!��u	�'Րi:⌛q���'�xU�b�|b��?q���yR �0��@:u�^
A���P7�y�%ڣ_*�� M�8μmȧmU��$�}����|��TD��h�"�2w*&4�%��>�j�(u
U 9��'�b�'����'z">��p��LI�
K�h��* *�x�-;_T���B�Mp"%Cq�i�Z��D�m5Q�ԡ�ɠt(�h����IY�P8�#�6q�BgF�Bt���q甼��)v�������u�T��
�m��I��a�׆ex����8��I�' ��jt�V_H�"��׺1���+|O@b�Б��<�l���N�+z�f�"C�'��CԦ���Iy��B��'�?��Ȝy�F�xd��~X0�*L��?����|���?�O��9��-=�>�`��,Hд�Z)]B$2���;��;�ON?dv�r���z�'{$}zq*޳0�Z� ���
�E;�KCgҸC��ŘJc�%�iH�:��dp��  t>�(�G�|�� ��?����W�uG�A%ϊ%M�B� ��ʲO6�'�a|�@ �W2L0Un��>�ʴ��]���'Qў���?��ċ�3�t�ꁅ�&1b������,�'S {�bk�N���O�˧B7Lȹ�E(T\�
�.��y�L�D������?ѐʝs���9�E�F�\����9���b�D"������3EÊ4�cL�����]�X�h4� �d��5*��������˧1D
�����q���	�:J���'Е���?1��In��ѧ��=_>0�a�׍8��ly�G"D�$�$�
c��ˢ�h) ��!"���>U p�Ƴ8����ֲs��];v�Ŧ��	֟x�I�n�~|�bHCɟ��������������������MⅭ �K0��bMՑm-�!�!b�&]ٖ��|�"B��i�J�����tS �7�Ā��n�'&�a�`�/3��Lq�J	���y�敲)�x�O0$d����y���t��(�a��Ǣ��!o��?��O�I���'���I:Z�v� �@K���cB9P�~$��
�`�Qf�� ��hĆ�:�F���۟���4���<)�� $��ir1+Lo��$k�]$�&i�Rhϥ�?����?1�����O��d>U���L&K��Kk@�+�ԶS���0ũҔ��;��M$r
�m��I�i���Dyb*��� ^���^ p�5���I�έ9 J�|�&�H�'ШG�2T�DLP3ֆ����K���)�(1��K�7_�����'�r�'��O#|�#-�
Z޾h��W-��,�.�n�<q��ǭ�~�{�	����u��m�	��M�����d��Z0�O�b���fi�q�[,/�L�;�� �R�'{$ݘ��'��<���h"�_�9��<{�/��I��
�M-����6n��u���+�nIG~� :Pwj�3G����M�;"�2!I$	�7M�9�sm���	 4�>�J{���	џ��'N}����ANh�î	4f4"K>�X������2#��31�/z@������?�E'l������*�lP$�V̟�'9�Q(Qaq�v�$�O�ʧS�(���K���@��4�@��ŀ�\����?1��ٷ]Q��K���#� !����'Ԝ��A�d.L���a�Kc���`�� ��$��B���V�h�Q8s�[R��~�gۗ,J8`��*9������w~2�֗�?��|��)F_.Z�YE	��&@E-!��.}~�`DJR ߚ-)���v�џ��	HBe��֢Ԟ�:YÖ�!+-B�'r�'z�ph����Dt��'���'$�.{;2a��&�?�HYj�Ad�����;����LS>H� ��^�,q�Xq�'��EСDO�2�I¡j�1C�lQ�)^�/+,�Y��Ѿ+�HD�PDH��~��R>�#!��{J�]:r�t˕�ސ:��1��T�i�&?�f���'ўr`��"�p�T�@�N��D�'��e�<)�(��e����`�fcM�^^�	t���4�����<	7N�\]F�Ѳe�0b7�E�5��<�'"_��?���?��U\�n�O���w>��ЧجVs$�a`�>��7�)`i�Z�)}�ys�叫WϨ8:p
9�F�BH ��9\Nl�W�9K����
@9Vs�$�g�D�(�Z�cG&��OV���HQ��lYۥ�?�rQ�U'�>H�"�'��D �'6����D���.��Kč��E�ȓ1��@Z��ɂ�]�,D�pS��s��M;����T�`D�O�"e�cp؋QT)W�H�rt�ޱj�2�'��I��'b=��d*���A�1B&gӪz�܄�S��66���`@�7,Vm��È1���j���(OАA𦊡'C��n[�<|ÓA�g��$`��.�֐���ۖ$�>tx%���(O���'��6�Nwy2�S(���SAU84�&IP H��䓽0>1���^�*��EX�7����e�a������T�r����W�:�0��U�y1$��I\y"K)Y��7��O����|����?q���琰#�!��:�dB桑��?���ZZ氡���X{�'��Sr��*	?j	��)Y�0@��u����[,"A���I�#l�j��%�~U橂�qȨ��GS�?���4�e���?yܴ�?	��I�]~~�1d+��5�V�+4kNX@�'�X��E{��4�H4JCi׶K������B�џ���4z����|���tX=F�Q�g,�@��
�Mt�7��O�$�O�(@�[&7��$�O�D�O��ݡ\Q�T�D-V�u��z�k��$�����Ծ�[�FG"0���"CM1�iK90�([��O� ����`�������pA�#�+(\�-�e/��^��!�Lst1����bρ��$C3���{t
M|y$� !E��?�һi��oϤ���Y���ɀ3&��C�Z�0� �4��u�'Ia~"�T�wk6\	!=\�D�%�Q����}�8l�o�	&'���SMy��Q�h%,l��W",�:uPW�T!2f�=�4M���b�'�b�'w.�]��럜���YU�l�V��& `�kŬ�R-ЇG�;W��@{��dӦy)�)�?�.PDy�MN�L�H�!!,D�Ѓ�ą�n��ۡ��&�!�S� ~-0��i�8v��1S1O�8b�QD��H�~��XQr	פ�/d�BMm���t�'�2�'��'���u��V�Z���$d� Mxq�'O1O�Y�N�2E2ڭ���G�t¸h��|bEX�t۾6m�<��"6#��N�O����w�f@�&J��v�f%�ߢ�d�Oz�I�OB�$v>Ur������ �� ����4pP`H1�CS��pV��	@��P��	�u"<�3��BȜ�Ơ��Mc匟rҮ�q4bޅ&Դ�ã�f���v��O>ymZ���Y_�ԣ2!J�o)�l�"��t��'$a|r�
���|�fM�72mw����?Q��'�.�p�M�Pu���끔v��lq���$#i����O����|JfϞ��?�`�^&\9���J�.1��L�V�8�?���9��8[��\cj�z��R��M�R��mR1�q�?MI�
��FO$�
f��v�<�bW�$?��J�4�2�	���hV�n�2�^�K�f�5�qIB�OI��9�#�=؆<�c��D0�(�O�y��'7r���<Q�f�#�0DrtE$���G�<��+��p�����6|Ɔ��5i&��?���11Kx9S�Y�a%��z��.7? �۴�?.O���s�埄�$�O��$�<y���f-����ڻ"��Lui3_ � �d��,Dzi�	7Y���8(����9��]D�O�t�G����E�@�>x��[b-ƛHh%"S��@_n$��O>%�N̉�&�|��n�<�Z��{�? ©1B�\4Z��t�vD(fT���@|����'�FAP��jɟ�'4�ђ��j%09Я3L5���	l���(^�^ipq��+� $ي�#�O���HҦ�Bش���|��'�򤑥=2L�.�|�(�� ��O�C�������d�O��D�O L���?Y����t�:����@(
���V�J!1��E��nvJ<)a���E�x���s�8hDybl�<}
�* �"��b����A���qE�8eg�d�QE'o^L���͐m}�9Fy��#f�I��j"v%��L%pR�z��g���D,!"jh��5W���J�� �y2&
!@e��a^��ҤY�O���{���|�.�b~*�'�?�ɼƱ�`G�{�<��KL��?��Bdfa2���?Y�OAah��.D�|�p�m@�eZN|�����-��'ڕ6d�U�	l�4Pb�PY�'��E�`��zVP��	|���l��$�buQ��L2za<$�U���!��L�'ź�h��?��O���#�U=N�R��So��q������|2�'l�@�`@90jHAԅ؟J�P���3��nK$�0�O�%�
�s��M �?)(O�������I��ȟ�O���c��'�ɗ��+`��`�C̠*�T���'I�F@_Ĵ�@$E�?�-ȶ!G� *0i�d�++��-5�x8����=��֨[g��Y��{�Bɶb�B��F��=�mۀ�_=S,�O�blP��D�]��Q��FO�NXꜪ�OTݣ��'��O>��pEB�O�~-�'�+.f9B�`>D���A�}s�3��V�4�el;�y�>��G̘Rf|b��$b�{r�ަ��I�����'iL�8j��Oڟ���ӟ<��̼��_�"��| �R�4�sKӑ#<j"Q/G�q��i1��R4����|w�^�9�t��$d��iW�7zJ	�0	(��@ÂU�@�R䢗抙%.���`��	N�O \4���y�n؍x���rE�:q� ���^���'v� ����Ϙ'枅�G�9_FAQ�ղú��	�'���@dF�@9�FѩN��i���?��i>%�TA�+˲w�xY@��+x�v42�(M�! B�
���ӟp�	��$���u��'��;�&���K�]��i"�.$>��ʡ�ln���ʇ���X���&�(D~r˻c��\1��%o��A�W�<m  �Ɲ��}�S�LR Q�  -�c5R�1ↁ12��H�$)�S%�?a���hO�"<Q�bX�Q\T�3�'��s�|�c�[�<I�%�����\	���q�
U��M[���dƞU���OC�3/O>��5@�Bےq����V��'�J�B��'�b3��PPfH	1T�^�Â�7X�1�"T7���8�a�<-�1K�(�/LǞUy��œ�(O���3�_'=�ʱ�ôx�PU13N�?����+ل�Cǈ���A*����q�4�d�*�R�'N��M��A��
�/(�`u�0m�vF�Of��D�)Q"��-�j�D���"m�O��=�'I��)�����(ľ3]�bB���?))OkJ��?��?9,�| h5h�O`���(V;>���Pq�]�:�P�:a��O��$�!��`�X���i�A�">�,l!bK*�R˧h1��P(��iv���ݶx�L��OHh
�+�^ј=[�lȓ.�̥�TjB'g�� ���ͬ�ilf�L���"$ʆQ#C#M�
��IDH����ڦEa��	r>���P=_�qB�,D�@*��3 /��ʈ� � �V� ��$��B [E�Lh���ޟ�s�4&{���|�|��LE�C���؃횋 �r7m�O����OBkq�3u�$���O��$�O��]�����C�θ
��@B
�ۆ�9�m��6Z���$����Q�5�Ӟ�XQ���O Q*`E	�I�V��2G3o�L�be��&3V�����*����	*q���c���|�1J�;�eλg����B��L�֙)RiɭN�� N>iI���|�<���F,;>j$��,��=P�gJ�<��	�U�I��^.�p�%��ş��I��HO�	$��K�!u�U����8HhK�_�f�*|2�
(?�l�$�O����O�Q���?�������ŗF�X�qw��}q �E͋jb<x#��@ܑ��ߴn����招��Ey�r�t���Ǚ�	8lA�F�if�)�*G>Hl ��p�STE�Ɗ�XǬ\����1;p�'��\��~��\�p�y�P@�&X��?I��'{�A�c�;�8���.��?������'c��2�hG2+�̡��˖�3��JL>ya�if�'��MPc¨~��j9>��5&��4�6 �&��7,�h�{���?)�S��?A����4Ùv��yE����9
��1l(��˩e��)���*6�`�6�B�cGn$GyrK/Q�n����%W
ĠE�TL*l��GJ!6n���e�ݸ�v��#���ez�c�!��h!�'|�c���?9�O6(��gײoA��`��&bJ��Օ|R�'*B�H/}���e��{��i��i>ɪ�rS���͎�2�dtℬ�6Q@�I}y�IK�X�z6-�O���|���Z�<�cBllW��
�v�˅X#?�f���O^��s�ڢf8\����H�?%�7*X<���5+��S�=�y�� [�det���$W�i�*�6� X너�������к8�Br���H�D�O(L�nY�)�^�:���Q��YC�O`�"��'87]X�O�� <��䇿R�R �E�V�B�
 B�|"�'�b�'K?Q	K����=iu&ҁ
82�h�:���B�i�1�4�Ӎ��jҺ�*�X�5dV�5csӸ�D�O��� CͬT;���O����O�Dw�Y�ǈ�t*�H��*���Z�@�a4F<(4�F���4�fŷ"-zc>��K<#�"^Bp(E��d�R	iR�P?�ص��"�aTh찷��
;HI�|�T�xB��i�B���싵'P�bA�1�?�O@����'��46�h��.�8�RHI�Nv���ȓn��l���3+��h�`��1S�ԕ'1R#=�'�?�*O�����
�L���hM�\n�����(H�P|����Ov���O8���N�d�O��Ӽ�Z\j���>�^����v��A���q�tb�H�$,a'L� ��OP1�C޻2��gj�0���	����&�:��E̱_��j�/u�
�<�M�"���T%'��@'혆U6@��v&��L�	C�'������R���I�B!-u��A�-D������8T 3 �\ j�ɑ�8��V�����wyR-N�<����?���eK�+��V6}�$�ʰ�?���0̲Q����?i�O�r �=,���w�-b�2�hG�s\�hWKA<x�4���0<�d��lf�%���=3(nB�I�@1�Y!?BQ��h�B��9��E)�ў[V��O*�$<?)@�C!*�E$��*�ܸ��l�E�������I�)�2��n�)(4�L�g�c�,D{*�>��	�bx.�J�m�pw�as%͞'Ȗ�ĩ<!��0�?��N�a��]>i��H�h��ɂ,�L[2�úV���I�@��.�|Z��װxԺ���S�OZL��#�_�:z�u�uJơ0��j�OT8J��S^�T��`��J�}rNV�	m&� /�*g�&́&��B~2!^.�?	��h��I�ބx�eL3�ָq�%�7$�!�DP ̱��O>����m��=�џ�ˈ�)Χq�:�:G���Y�ĵ9��vmBA���	�	1�����?5���D�'��÷%ʸ�� �4/�-qN�(�!1X>`<�.�O�p�Y�2v1�1OҴ��S2`��	��N}#��A�h��J���OtL`B!+rW1�1OxD÷	��{2�r�-�d�VȻ#�'����q�>��O0�=�D�]
v��""ī�t81�._��yB �d��P2Q%ˋC��:sn��$�j����<��oʁx@2�+Ua�*n������W�\�.j@��A0��$J�.���9��U���@HȦ��W�ȣX���b��
.�zY��/�?����?a��?�l��R���a����黢~��|0�� @��}`�X�ah()����0�@�.0�p��*��T޽ʮ��|3S���g�؉0�S�Mg�I��	nf�������pL~��^�x��5I�lۤ��]�Q(�[y�'VH�c�dM�6:���93�L0�	�L=剀��ԛ�C�(c�U��L�&=��&V�u B�i���'�S
-����	џ���B�K��0@��/\)l	Xc�QП�0�Ś4*�E���zν����y�p�y�b�o̧R�͚��I%)�������;I,E̓1bv���|i:(�g��a�~���E��,�Zw�G���)AO�UՍ�:C�S쎝.��d��Q��'��)�I8?q��-�)B-��bj�1w�<yUe��%�������vl�j�J���?��i>'��?�`�����'D>�Ze�Fɟx��� �!�	�r�r�������	���P]w$bn��L�N�JuR���8��Rt؃7�O~�&L��s 6�aǗ?#<D�!ZC�4[����>>�i��Z�q�����=d�̒��ǇE�8A��O �cU�Y��"��Q�A/�0���0E��O:�$<��y�A��-m(����U=9N43��Q�y"�U6R�2�� �9c���z��Λ�?ق�i>Q��wy.�2S�q�h�`�'�� N6�i�K��!��'���'�ם�t�I�|B��"p)܀C#K�,:d�M@5�Z�P$�dȑn�4��X���U�gCre��D(���<P�/1��䲣���C�b�H�͋�""&� �e�:�3��w�d�(�DN�46*�<qS��ڟ$���Q"A���#�G�n�aq�՟���x���h�vEs3Ʊ&�@�!5FC4&0���f>D��h�����cde��EL]��ʾ<�3�i_�4]���_:���$x>5p�Nё~�ݢ�AS8h���bE�O\��� �O���O�u	��X�)E�feݣX�Y�����}J�ċ1�@æ�2!y�B�=#%Q��J�F�b���Ёx�&#DT,��0-��In	�m5D��:��Hp@DWE�I9;����O�b>i0���m��ag�G�d��x��<��Dpԭr@��L*؈��.
��'��D{�OG��茍�aE�N�؜yrG��[ؼ\�'�}KB�i�&��Oʧ�*|��?�/C&�(�*�b��;��4!@ϣ�?1mO0EJx��N� `,���)û1��P�1���O��3��T\89c��)(9���'��83Ì@����%Ӂ8��`�k��qF�g>�ʧؐ�'�F�P�fE�B`��r�̓{�jd��؟p����� ��{�(�:Z��:$��&X�<�Q"O���˂�(��sCX�!�~չ��$�OLDz�O����(�L)����/2H��'���'	�}�р��WYR�'I��')���'�� ��^�D22��ӀƳH�X��k@�K�&��G�:3d8��>��S2C�l	�>��͒
�H��r�kT
���Q?�,i�-�5� ��Veفg�V)�+� w%��Rv�F2�պ�eAi3P;���<5��䐟� v��O�D'��y�Ɏ?�
�d(_p<�#XD���Ɠ<"��fmŃPD̡� �II@�i��)����4�'�օ�m��2�\�*e�!d�]�Bк0�'�B�'�bFm�����P�'^V�<( E�]��i�%�xÕ�лB 醉G!�V̅�ɝ1URȲ�A4>ADЃ�!)6 1�b#P�!��C�`��AS`A؈�3��-��'����8�L`��	�+�X����3n^��p��hO�#>��/�L�j@�d#'T�8�c[A�<���< N��p�!�0���|y�M}��d�<��LҲh�������'�����>��0�'L�$�����+rt�	ן����*�@�i�%Ü�"�`4�C����O�H���̐�{��Uz�	ǌ$�a�����ID�3�i�a��e���o�􅄵iB 	�� X��Z&fM1�O�����'��6@�@���tMd�z�8�oY��*ʓ�0?)e-��%��Y�%�]�\�� -�yx�A/O�
%HG�v��t����e��	�F[����ɟ���`yB[>����<鶧K�(����e!���"x��
�s}�>O���<�eU��>}�C=<���E�\H�\,X�"��ʦ�'�#E��F��w:���Q�Z�l�� ��U��7��OF�+C�y�0˴��O���។�l���ݴ9gJ��G'	d����h�R)m��H��������!p�h��ם�m��diލ�b��a�4T	�k�9:&,�a��,���'�&��3O���͟$���?��	�<�֪֑-3ziҤG�\&Mڧ�
 �h������EQ埈͓,5|�����4a�D=T�����V�Ul������_���Dj�ş��'fz�����Od�I�OY�d�1��Ń�L�>,*����6�ğ��ɮCm������?��aYwnڋ]���k�!8,;�	�2�!!q�
�MS$�'-�=���?q��֦��d��:���O�ɑ�,�h0CN-���4��;T�$�B�v���� �O������yr#����4[*x���B9<8�ԁQ"[�'3��(�,÷]��7ONPsс`��AnZ�,��	ɺ������Eɥ$��a���fʁW��6���C <z6�_�y�S�����\���O���$/��E�0L<m~8Y�4t�������C�?Qoڤ��(O�T�\�E��`�a�;k�ް����){��C�	�q�� �S$�F�QE)B|�r7��O�ʓ�?!�[?�	ԟ�����{����k%V�ѳ�ɂ�l�I���D�<�����$�O����O ��*�`U�����W�LX:��ݾF6��O����O���O��$�|���?	KA&���"Z1[
�p��O�����'��'6�)�>QS��08|�LPV�˸$��P�'l}}2�'��@�VH�,a$ ��ѩ�ZO<��?�Ǔqi����|ҜQr@�O�t G~���(Ir�,���^fB��"�J�0vC䉳tVYV��((��D�O�&C�ɧ/�*x ��P�D��/�7��B�	C`�L�����
lz8{ƣ�$r�B䉱y�������=<�R ��.+��B�	"z��历�|_n��*܌Z��"?��?���?9��=�=r M3<LP9�*A �^�rU�i>��'!b�'�"�'\2�'32�'3�i8d�!u>4!��V`�Uz�E�>�D�O2�$�Op���O��$�O��D�O�����Ÿ�Y�֬%9¬`U�XӦ-������I۟���֟4�I���	���G��";r����4�	�p�Ć�M����?Q���?q���?9��?����?�g'��Wa��� �A%��肊�-����'3��'��'���'�B�'2+�:!��'HҀ�,�(���9�$7M�O���O>�D�O.��O����O��F)�������2I@Չ�"Ԑ�mZ��,�����ԟ`�	����֟X��~D�ZE<H��A֘0d���4�?����?1��?9���?A���?��u^yh�$�L>H"�F��I�zM�%�i���'b�'���'���'���'��4Ȓɓ�>�j�2ঋ��Z����o�$�D�O��d�OD���O
���O����OPyaNԟH"�q�ѫ�W� ��G�צ�����������	ퟤ���t�	ϟ���Ɂ�-���M�=ٚ� ����M+���?9���?i��?���?���?��e	|����J�oĄS2�C�a��������ty��u�N�H�N��Pe�4j�kW�Y�m�&�c���I򓻍M�w��挔%$&�ZB@Y�����i�7�k��'V�O~:4�!�i��D��{.��5K�4^�S �7B㒣_� Q�"#E,Uў��<����� ����kzs�%��RyB�|�t�d��e�d)� <��5�z�Ė-]X]9B��d}�pӠ�o��<�,�D�!�)$)��8z0,���@�W�HS�@��L���>?ͧ�A�^w���I�A}Fu1�M_%K�<�YV�ʓ���O�}��Z�{qB	�%��x�+�78�|���=�M��B�V~2�a���擽����2���5�R<�I��M�i���#8m�f��h�+�$����ᕨZ�~��}aJ٢�bt���Iן �'�1�6��@)%l��{󏟕5�Ȕ{T�dyڴg�2��<i����7��"=��}� �K#	6<�v ��x�j�	G�Ov���l���"�jf�vg��"zT��O�-A��N�6�0�%
>��A,OH�x�1k���D�6i+ �U5e*��F!D��cD�I�l�ak��-�� � %�
-��(��ŽbK"]��nȲ��)q2�܆|d�����-iw
�a7�� �^�qWJT�26&Bx�(���j�AɌ��6G�7]� �̀ǮH��M
`o�-s� =߸��1	�zx )жWG��+�k�,�D��AU$�.MK5$8Ϝ隱I�{|R�iѳ^W�ћ���<��3t�V�d��� �wl�B�Ʉ��}�OQ�p�f)������o�V�r���'^���#S�g��e�D�)	�D<�0c��j#T��9r����I�yY��L)0�g
H	�Bdk�`�{��M`ׅ�#N�XD0 �F�8Ρ
�`q��r§O0JId���#�m�V��Ӄ�)`�t���^T�QP/�5Hd$Q�a�)~ ��S��Mk��?!�axz��F�ܪ�����ی�?����?��a�BY�=��ʞ�
$�B�V6X�,hr��� ��؟`�'��p�'�bӌʧ�?!�w(���	T�u�,�ɕ��Cl������O����>�;(:��	�n8�n��7���	ay2�l�6M�|����"�V�H"��R�x<C�쇅y���.�O"���O���<�O=�L����l�(�0���:���$$�Oy �`�Ӧ�IٟH�I�?�`J<�'Xx �ZV��"��m�5,�,f�9��H]B(�(O����O����O�	����x�Ј�5�V�Q���Z��V��Iڟ��I�ڊqN<�'�?���u]�a�B��>�i@5oЩ���[*O��$�O���"�d�O����O�H���'R�f�*g'Si]�X��O$���*y�%�����IRyr���t\�j�ij��J�����'n�q��yR�'V��'��'K�T �*Ժ4T���0�Lbl��EUD7�O���O@���h�4_���I�/��� ��Ө����^�y�B�B B{�������b�����$��j����Z�4מ9�׋Ǯ�P�S�C�LU�����?����?I��?�/O��D�~���_ F,�e33�I��Zd��.F3Z���O���O����O��d��[��ilZ�����3Q$�i�&Ż_t������" i�0��Ɵ���̟ԕ'�"�%����'�B�Et��jwΐ�z�,������ �'�2�'Z�f�n�7��O�D�OZ��{.쥈d��5�65���L�n���O���?A��U�|����?7�L�|�g ��N��HJ��U�V�� ��?���?���Â�V�'��'��t�O�"F[�+��P���Ƴrw�9i���b��	��h���<&�����Z�#��)�2��� �꼚���?I��I�I �6�'�R�'���Or��'o�X_*|q�NN%Up�յ%���9L��O��$�OPAD�=r>$�7��/A���%���M��ş��-|����ğ��	ӟX�I�L�S���_`px��d���)J#Hz4�X�l)��ߟ��I�L�S�L:2~^,�w������y!�C؟���#E����ٴ�?���?q�<��<i��4�XIy2M�Z�e���_yʎ�y�U���	���IWyB�Y�wx����͜;��0����`l� (�>�-O��d�<���?a��v��Yi(�� �F�� '"r��녨��<!���?����?���?��p	�����i�Va��C:��#@�*�J0	��'h��'_��'�rY�x�ɷ8���'s��Y%�]�vx ��w>��IП`+"��ϟD��ڟ �IƖ�;۴�?�$#>a��M�� ��a1�[�1^����?����?�,O���G2t/�I3?Q�����l�c�˅t�<��5�ԟ,���X���4���� �M���?Q���ڷdZGl�!���7r�͛��Ļ�?y����D�O.�7�2�ĭ<�'�"����[iHE��[2J�FEB��?��Q:�c�iY��'�b�O����'����PCb@I>x��&U���	�=|����Vy��Z�����?�ʇ�_� "D=���[�⌃q�O�8�ע���Iޟ �I�?��S��<�IП;��
#�������a#�|���ɟ�hǠޟ�Iן`��x>�%?y��!W�)����>^@sR��!X�ڴ�?!��?����(�B��?���?���D=��ٷf	?
sʜ1�뇒31ꑀ��?�(O����>���O��$�O��)ye�s�f��&ና��O�DT�e�l���I���ɰ���o�|�4j��JC��if�A-h�}R�<Yg�<Q,O����O��'�?�"�Ğ3�̐T��/*����rdQ�j�&���i�"�'TB�'�<ꧮ��O6�c�*N<�����C��Y�v��wk��b���Op���O��ħ|ΓKD��Z�Op2��ť�-r̆�+U睄+�,4�(O����O��O����O������O~����"D'�m[�0o댌�Ƞ<����?�����N�T'>���UL��!�č	X��� �GBß��	]�	ß���	�4� �iG *���!�w�����O�D�O��f�}�&���'���� j8ZaD�f��U���0~Xՠ!�|��'�R�;gr�|�O�ұ([#�0����1^��!����d�E�*uma���'W��ƫ<��N�����&#�-薑١�\ߟ��I��l�,��%�t�|Z��E(rĜ��g"��.���U��� '?�M����?���"�xb�'���8�gX=(���EΛ�^^��'P�����'��'~�Z�$�0^��8��N�C��p��<A�o�̟�����pr�	���?���y2Ƈ2!��)�v-Ү`�8���Ԯ�?!J>!7�T����?���?� �6yRv��4P<4�/�?I���\jv�x��'ҝ|�B��JAz��.V�R3��.e,�I$q_��IAy��'���'��j�P��H��(�j�)�|zu�S�D���'�B�|��'��GR9R��f'Hm��#�KV�>�ܰ��'t�	�P�	ȟԕ'��1�����Z�k���mEX`qS`��N}�\��	ٟ$'��Iٟ��g��,SL�"|�>��
VS�XЇ�b�I�,�x=�����Dh�e:T/~f�j2K��|��g[#_�JQ�T� ����w�����?)���?1O>�����I�����W��"iC �$dsA�\����I�4$��I�9���p�ͨ+��@�_켍�s��-$2�Ƃ�4g�C��310 	""�J�[��5�g:Nx���ЕC���[��M,q���
�D$&980��ʟ�:>L)��&^=�q�� ,��y
�bƟd�20B� 2h��Ȕ�D�,��<jUHуP�y�x�b�]�@cr�9�*>xe8��'(¸e�u�ґE�x���ԁP�$,"D|6��ȗ/I&-L��	��=C�A�EN< ��%��H2R��1��'��j`�'�"�'0�������T�"`N0��ƕ���ڛ;l���a�0�Z-�q�� Ȉ�D�:k��E�*7����P��?`x��#%�4(&a��MR�~��,�u�B&��:��dI����s������h�Q�ۘ 
��`�ӄ'�>8��OџL��H�S�ORҔ `F�8(bș�)��M��	,�Ğ�]f�ZA�V� zE�a -z��!�'��x�f�|���O�˧BE�4���M��,E�)1��2A��(����\�X��T0%P8р��݂i���ԏ�6W
;�^�OB����صh�����L�<p�,��O �҄j��Lnd�a�.1$6�� K֯K�$̺N~:f��c@�-
 �[:$Y����EBp}"�Q �?a%�|���Qc�����˖8s�%��R�!�*^���c���@@e�>h�Q�T���3C�L����%�J��RJD���I�����#D��"o������x����Ձ	>��� o���e�e�'&��tf�x��Ξ+X�"}A��HN�S&��'bx�0s`�	�>U*�h��I�tJ #�	q�ؐ#�^/b羙x�F����'i�1O�} ���'I��0w̓=-C|�铗xn�'�?Y��'�t�Z%���,��Y5gY�	��	�'j��t�^V(�5�ϯJ��)B�'
�#=ͧ��8��{BiZ(b�ĉx��/[�&9��ʷxQ�b���?���?�R����O��S��t��נW�4�XC%hX�5��D�Q���G0��`��0b�Z�X#��+Dp|��ɤ@,daA ��C_x�I1�L	=�r�����^0pb�Ŗ�"*ѳ��+'���v�=q3��%���veh�0��u`Q�)9����A��{�ڟ�&���Iޟ �?��2e�f�c� �$���	�I�C V���#��+h� %*FN�8�)z��1k�R�'�66��O>˓V�F餱i)"�'͛fȘq��<���(�$��C�OV��D����d�O��$�Kќ�8#�[�����G�z#lh�oV[��,���� }b���i��t����F�I�U�N�SI��`�N:M�DqP����:m��[f�\�J�-!J� V[��0��d�6V��'�r�O,�Q�f$A�oլX;���/�����O>�)�	��|�	��'#�=KeK��>8���%~���{��i>��ش=�RMp�I�	9{�i �.#��)�iф��dT�p��nȟ���[��ᘬc-°i5��%I̾Hi��#�"6#���Vc�O䠒�� Tn�aRfƲT]��en¥H\Z;�)^ {߄�dcבW�n�Z���68a�I�*�P�w�Y��lE��)P�o6@���m�1}��O� %���%5�iq1߾{8l��OJ!�!�'�7���(���b�>�G��}�>�!�� ��kT"O|�1�OƠ1@���W�Z����c�	��h��勓�|3d����V� ��Cے8#��'��̗	�^I�#�'g��'�"b�ҼK�"�9c�\�Ơ�;p�Psh�DEp$
�+X�[m���@���$>	�=�'�N3:�\�qH|^��TM�8��*M�b��d�E�
�ء$>u�=����(�#GW��,��j�L�I�����l8��j�$��4����-x&�9s�I(D�ȳ���X�`�������11���8�����-*� �m��-u����:_N��A�D�<�����I��H�_w��'f�	�?���ru�%lK ��ŮO�u�.��O�pDЂ�"̀i�4��dJ���5p��qlDh��@J��r����x�j88��`h�z#	�u�@a d

S,Z�ъ�D�-d��@D	=f�耔�
�1�Ţ"�˧!���T4�H��a�j0D̒�a��q�`��M�S�? �p�gȅ\�h�f�HU��iu�>)ײi�'�b����e�4���O<6�F�^v���Ǉc�D� ��9kh���WybP��ʟ�I?,1��pe�JJ��9a�U�7�,���2�0��4fV�`�p"�	�nC��
��.��4�ĠZ�Z���.�WCV%#`�e��E1 �-ʶ�9�`�c�d�~NQ�����O�%�}2���-���/03��E�<q�W=d/��:E/X.Qxu)d��~ܓ�hO�)�d?�Ca��U�L�� �BE�CeNnk��'@�Mn� t'��gy����m�tA��K�� ���/�M[���s�vL� Ρ-��=В��*@p��P��>P�>R����Q���AD�|����A����=>L�!ز�K�Yk�цȓvH�mCt�н'�x�j�w.켆��Yc�ռhk"�yq�!GbL��&�>�[���$Zz|�`�P�&�T�ȓ-�m�F��4~L95#T�Hh�	�ȓC�Z%EfЮ<)''Y��4-�ȓx�b�d��'|�P@�CKҌ��ȓA����CR�-�:%�ǭF�<�n�ȓp[
@p@^�Joȁ1nH����ȓ1��Zwώ!2���LY"!�T-����zP��9*�ԴqG'\�,�J��+Tl�3�X�|�.Mi��J�l`�ȓk�8tsbEƪN0n�h6,Y��%h(D���G�;"yrt:� ¤*������)D�0C�.O z�ĉk��JC$#��&D����͔0J�� 1�C�)4%��'D���@.H��z��.��/�6���9D���� M�'ˌ鋠jڂ=	eᣫ9D�LK��ۗ`LB}��d��b��}jJ"D�PJ���rrqQ��Y&���6D��:��//'�)y�̂OU�AK�N D�<9r.^�"�����K�IŒ\)0D�hd�:E���#ÀsR(�r�1D�DI��f�EZ�˷�H5)�d3D��A�$nq*����g+*1�bo.D�p(��ݼ;Jɋ��>q�>�k'6D��k��I�4�� a7��7s��H��!D�:�b[3 َ�Da�2[����e*?D�LZQ����Ԑ����1I�Bd�?D�@�u%�"s�*�Pw'{6�"�=D�8*�JԿq@��b&̜Ba�bF8D��kRF�z�j���K΍|�Hhi<D��!ee��� 1ۀ*;\ѹ��)D��0�J�s�8��e��En"��W�$�DߊDl&�{������P�楋F�x�a�bC��yDј|��A.
~�@�J�L�'/C�H�����Y�N]q��'�����n��I�!�v�g ��	�'������	R��y�)ܻ�NH�e� ���5�v��}�`���P��QI�Ę��Qā
��O�[q�Ǽ'.K��Ƒ����#�����E���\�2L� {!�D�	_4�y��¤7�&��&iΟM�	����ېf��=x:$�D���N�aPr�K2*�r��#��-ce�C�ɰ<j�����Q�z)K��ه8�d)[�F�K~2�3fێY�37����!�H��[�z�
�)+C�.�a�%Ҥ@�����cW�R$�S�i�X����t�n�s��ɠD��|� �3��"P �9o�ʡ:���,��O$�Q�D�u�M#���b�S�Vh@���qY��HF	Z5OXC�I#R�H��A�	;(x%���5o.�#Mr�a�P�Q���8	ѩ����
_�|�jeM���$��9]���zӬR=R�Ā� X�y2	�xb�d2���U��0G�?j�Q�w��� S�J	t�X��v��y`�	*UI���*^���� �j���`ҫN'�6p�C�v؟�&CA� �@聵�D�^.��3.�]�PԈU��^�TpK�Œ퟈�%�Ō[�V���E�[(c�$c�cCd�p�4b֣1T�Y�1��4;V������N��Ms��ÐS�XeŦ	$��`C쐥uM��AEI�RQ^p�0��7��zRd�� c:�ڕ�i�Č�# �6��$�6ji�ES�"��3݄I�41l����6hkT�Y�fZ�!�B � �h#���77&����	Vj ��"O�9p�ǔF�&�R�	�<V���Ń�EH�m�� Q�a{�`�+@�N�7���� �}�\��kg޵#VE��v��BENIb`��e%��3f�4V�;VZ:0>��xcJ)�a�aļgM��3���5�
%�R�\�\�fD�?c�<�F��>�VH����"|���1v 8O��JƧ2��u��'M���T했�<�$�Cy�F܁���&c�x��@l �I]$��Ǭ��0=�s&ō,��i�Lzt�85gA/9fP�-��6����i){���@��4T�`�N�5Ty3 ��j�JX��$ѥs������'�RuP@^+l�B��u�Wm'���3��b��▫*_�|���̎<�v�X�-�k�D�ҍ�	Y������˔�m�Z��b���l�j��P��ʟyCX�bFV>�h�FՆx����T�ҌZzI��afJQ���O�Oa*���E׆cvb>c�D��BQ ��l�үvC�U��E>-% "�O�-&�RG$�$<vTH���i��<��D4���x��2	�	S� �M@�d(�+���5 ��'W �3��Bc�0
�m�~�Zl���?`*.�F�Ӡ3�����������b�(!bc���^`��оcJ�ę0O^�Q�A���
8�N�1�E���#D�pB����i���Œ�S3�\��I��;�� � +Y�:�>� N��?�f���)���S�Nܧ]hܝX`���&��'fEKWb$�>IaCR�d�9�B@� ��@P��]2 M��ObJH���σ�b���Zb&���PFD5+n� �aNϦY�D>q��'�긓���*\zŲaτ!g\���I�9<U�������R$
����J���~b�Br���ӑ
��z�f�C��z�MցL�:����$ljA?lO�}�*�j^�0�4��rt�,`�h�%x��}�VK JDC��Q��q���ٖnW����@5v�  U��O,��q�ή^ƚ�� !PDi1�'Ĝ��` ��[^Us�'<8��Q�FK4 �������9.GF�8�@۟cb�hKRK-����R$ԍ��16��b>�1�&��L��AX���_�h�ٕi+����� ��3��8�b�Թ��P�A��4�0�3q�D 7DPY:(3�n��B�ɺLaYD���!�a�8?����B[�Ē�i $��C�;M�O ��3�q�5�"愰7�H��*2��h�i,$��!ł�2�F�Z���9\J�,���ѻ7S,�R�-2D���$�n��;C%�)7�\#=!`�6#�x+��l������\X�<���X�:	{��<?^��v��D���/�.9a�x����!�lpq��H��}�L�'-��q��$�@$هl����]MV� ��HJޠ@�D R8 l��$�%��S�_S��w.�N 	��(�iRB�	�ZԨ�cÏ��G�\�b�o�]ܕеm˹0�Z�B
�+u����Q�<���o�pP�!ֈmңEV$󺱲��;3��H��c��yزe�3�����P�M��2�\)P ��@�-$���Ю ȣ?������*�`���M0��VEX�\ȡ��'�z�IB��.>h��CU j`KR R	R꺌�""Tj:pY�':�Y��f�2Cj)C���*~�АO<Y���Q� �ѯ��x��2m�'$4����
��K5ҐqtZ5u��ȓ'�<4c$�Պ1tz)��X�ph#�h��A�L�H�G�#�"թ�t�g�ɁF��ma1
���(qoʨ!FVB�	�h��Z��ӘGd�hX���"���3��,@&��ͅC�~���>,O�p�5
�>F�;�\�;5P+'�'�8�N;xt�`��͖J�Jݩf�A�k�x\��똌GoAaD���x�8�����Άfs�1���,�ē��i҈��^W܌Y��>j��~zr ٹ6�ҝ+��� �X�0�&�j�<A�[�]�t`X��ކ)��칆�L�r�ɡ�F C�u��
˟h/܈�~&���ǆ��ɲ�����+0�tT�;$�����
�4*�BR�M�p����4[j>��`!� %!:Y�$)��t��d^�?�>p°%��;or��4m�e_ay��˫~�И1�?Ť����,E��p�L��8xlpIP!X�v�f�B�'Ѻḳ�Υ9$<�Q��P�6��m3I<Q�,M `f���z���TG�'<ԌlJ�]���֦-6�tT��+�����X�����V�"�(a"ޏ>e������.8;jU�A@�g�I�=��}
�|��`E�A�a��C�I�htR�P�ؾLѴq��͐��8(ǅP1�ٳ�횅��q��C�#sX��O.���(l��L	bLh%�	1L�f�/?�D�'3� �dh��l���I��>Oj����+d���{� �g.��!'o�<m���b��]�<a�b�p����N~&�Da���r�;j1.ኍ��(8�$�1,���y	���:q�3K|��Z�h��5���Y�X�P�t� �}W� ��Iݒ{���լU�@a{�P�}��CR���YB�K�K0q!'ɿ!?P�	�k{��d��O-� ��DƉ9#vu��$�N�z��BL)Sh˃�÷Sv�
'��8�!�$�,^���ɞ1m�D:�A��K���҅_���5�� N�.��TI�/Y���!i_2k�`��j��	�{A,%qoە*�j�0)�0=��-��E>�H����!}G~�� p*��� d�4ع�*i.� c�"g*%f��)]�|���7�x�OV���eGyrF: �V��G�..$|�����'&t��B��+zh��k@HԪt��'P��T��B�/�1k� �<L4�� #�+c�48p!BZ0 ����C�)4���+C�'��*g��3	oFah!>dy�p)U�/t۲ �@FՇ&X7m�-��.V8hQ�e�ꂈ����&ʪ�h��BOQ�b�t�m���x����\�*����*�OH�����:L���aZ�"+���#�T�[�n��3$Q�i�-i""�*<mT��u�י;N��&�� /���Oa���S ]�n1$a#�
Mj��
�����#� :�aQcD� 'py(bFV<�GEY����S��V%kr9����~X���)��#%�ӅNE�M&.��f������q�x�r�.=Zf,�`ǚ<E�1Ob �0Z�A��`�톟"����O��9:�`��m
�A�e$P8gF`t���Z::TpDK���ZJ���/0��˓��6`�u���1�`�M�%'S+N�ȗ.��Rh��:!�Z}�i%Ď~�b�1���`�Q��GؐV TȰg�ǘTc��z���J"�D� ��� äԒz�z�����D:�)�)(|O=1�?zl$���� 7��x�E�����A.���0�rN�h���>yj4Ђ������݇8��9"��`Ѧ��?^�����G�R/ay�-��qw�a�c�]�D�j7�^%����&�2���-��v��p�PK��F��1�((o�&�HW�����擓$�<��6�Cq��D�Xc5�9Jg�G$DR�;����Q+D�#L<i7���A�N���G�@�zܐ��J���A<�2W
���4� ��A����J�i�V�k�j��v� psqA#|!�(��T<�*�x����I�<�����if|�Q�	v�щU$�͹D�.8b�� �=�H]��ܝH�>��r�G~~���4�dx#p� )M �p�з'�H�1�G��.��!lO吐�PWt��k\Q�)*@K>
~2�q�e�j��m�q� '��������iU�2R���|�,ۥqJ8����%}��1d�bX�x��݅!F�P��h� Cېy��oè^��L+�(��i�a�HC�n�(���/�7T����N�֟����é����j�
Uyr�h�2֘6�bL�CΏw� D�4c��O M�D���m�Ekr���lqF���^?I�ۓ3�x�RA�ܫ���GM��Q��5�s,��ȍ�0,�y�"�`����<�܅2�)��#<A&d#bX����D	�2�KV�y��["�P�(Jr`Z�x��U�wLO� �1��dǦ#@"���-'~��{b-�=I�>x��-&��qz"a�\����y2<�R2
:|O � ��R��z��D پt청�W�� �$M�Џ<M
��3��;y�V�8`S�
�b�˄��=r⤹�g�e>1�!�$M,�9g� �[���`'LO6@L�یex�#ɍ*���ge�s�b9�(Ƣ�ԤU�h��A�T""\�Ҩ���-OCDQ�v�Ubf��`Vz]R�jb޹T �$�h�ˢÛ�$#�]c�i"����!�tAݡ u"e O~�A��wb� @m�)���%.M*��aA� F��"��X�ܸ���ۗgn�( ��(O����EY5��P��U�]���I/_Z^�ucK~�"����c+����:��R2,��+��� �Cէ�=����1H[�*�ɂ<Wx�$���Zmi�o� Ԛ`��	��'@�=�B�~���t��1*-�����(�, b�3 X�D��MR?a�E"�"O i(V�B4Ѩ�y�fŪsI��[���fEM5)R�[�MH��0|��Dw�4Q�Sftnѕ�Rj�<YU��5"1lDp���B(��@5�h�ȓk��Q)qd@8Dyt�х�4G��k$.٩M�`��7�z�ȓ6�x�ê5H�H�q�ڥ[=���1���gɒ3�z�9����<8x�ȓTh�8 N�?��3a�6*:dt��7a��k�5
%�ɰ>�
���jn��W#��G��U��L�@)%�ȓ�¸i-��?9�����wՎ$�ȓUچq"���'���8 �[�H��4�ްCQ���<\rIе	ԩ9B9���~t�[�T��XP�@ =e a�ȓ�\ĩ3�P�B 8cʙ�N�}�ȓ3f���c�;+��{qJ�8�a��kM�$K4mY�J��v��i)�L��k���S��ɓ���t��I����L�D��僿b�])�¸��!�ȓP�S����Q��uрM�9�ꘆ��i�K��w�`!�!&��KM*Շȓx�*m��'�)Z@d��H�	=�0�ȓl �RVD��z�8�s(��0(���ȓ��0at��/O�v��QbU�<��O%.bf)��/S3�Mc#��U�<	�GL(פHq� �%M2��T�_�<�̒�Pk4����!g�X���L�c�<�0*��|���z�_�-�:�PfX[�<�vO�'c��P���f�v�qaQW�<� <�G�Ra�����<AY~��1"O�� TI�5�ЬB�"A�,.Ra�"O
�j���z(�*��-�U��"OR�*$�P6;Z)���ܑh֠I�"O0D`r$F�NI�\{E�7���b"O�}�π�R1iDe
�uzP"O�X�ɑ��š&���B�M�G"O�AX��G?�����Él�f���"O~,��M׸"�Z	��ʜ��y�"O��r��Z)�&��a��(�����"O���d'[�,���#�
���{""O���!�!Qg䊀#S�3�BCE"OꐨOF�����$X�^D�{��>��$�3e�(��Ύ�����d#�{��H������Q�kmĤ`��m��1�ȓQ%��9��؁p>�l�s�B���0�ȓ9����Fp�e�V�	Lfl��b�|�f���c��X�o `�l�ȓ%�4��Bb����$�@�_{ڬ�ȓ�jqbAH)Ӽ�w�\�Q`R��ȓ
qpt��D�b� 4��(� �z�ȓg2������X.���I��|xތ�ȓc����d��v���,�8;N���ȓ6x��ǭE����
�T� 9�ȓb¸���J�r�h4󁨌0N��ȓcbD�4�o��b��-T�����0J� ��_�"��ږ��+�x�ȓ��M��ņ�"x�@��,L	Ӫ���x:�`�Aԛ$*��yǣ�O= �ȓg�PhfG_ ����"��*�R��ȓ9�<��熝�����/I=D�*���b��\`E'!��pR�N�5�f̅�C0d���l�L��,*�MS.*��<��~g1��切8��X�eU�X#�P�ȓw��c�&�UL�=�Ĩ����/�R)W�è[���zl@�.�:���d�AT-ٛ_p���O/�,(�ȓOU�����n<(�X@dŖ{a��C
|���ՂzQ p�(ӒN�y��8������AKx<˳j��d͆ȓ��-�&�)!�����Jj@H��U6�{#o_�W۸ ��6) U��/n�;�i�% �`���L-��\��xr��ϒ�Q:�(�U�T,Y�<��-o࠻UW�;��P����Ivj��g���j��[/y9�0�קA>n�ćȓ#J��M�1 �:��ф2�^�ȓ& HI"�ک'0`�3 CŵfZ��ȓ�z	���%�2(�0��h�����BIXqEvy��PSĭ+��	6�~ᢁ	Q�yB+��x��t�C#���Aթژ'+��YAAԫ^��?��T��&w�\� �.͎F̪W(!D�0Y����Y�`[�K�z�����!�
��f�Bpo�v̶��O���	�B5���'sVyyB�C>�N��Q�/����'Ͼ��u$�F����I[+F�~ܲB�Z�O"3�D��M/#��ܳ@�rӞEl�3}|�a�҂��_7���yz �ңN�'��|� ߢ:�D���F\�][3(΀~D��� ��6	��-8B���/yJ|<��n�0p��؀�(0I.n����σY*6��OB m��M��8O�������)s�Yo����|r�2�����1m �ȈE�ٽ��$�S�4� &kI��b!˘�v�R�0EZ(2 a���Q=6�7MK�Z&�I	M ,�V������)U-W���Xa�S�U/�	c@Ő�Ur�
'�U�:d[)O�T�.\����i�_��P3�'z�� �9R��Ƌ�M��G0.Ip�1%m?j�y��I3%l��ң�*/�\A���\|��>�)yc�2^(��A���E�֢}be�=n�)q$}l�z2�V��0=��v�<T��k[��a�V����A� ��RXVpha)a���0'�`\P+ʟ=�i^ E@0��RL�ugPM�Cn�1�h���m]�*7Z슊}�ڭV;��C1�Y��U�U�O�5��6mO�Sh&�� ":d��"w>��4O�2!�z�yq%
�cfH)#r�Ýs$(f�׽Wע9b��b���|r��|F�4
�K��j(�[��Wg���c�X� >d٩���u�(y]�?1�$�y6*���2�^����ZW�DEv��!)�O�,n�Bx�q�Yp��bCc�2{t��Ē�S֐x&�˰U�@�yW�U�7,�9a�O���īr�z%��O�
�7%��j�L�����$�y�ǀ�K��P��ɼG��� ��*zL��➂x*6A��O<^T<�$���(��'H���G�K	`��O��������R@$��A�՝M�61ZRM[~РSt H�D>d�?ɒ�اl�l`���n6��C���,)��&v(�2�,TH��Tc��#a,��f�
?3��9�����o�-j|�-,Bb��0�D��"P��",�8q~�=�f��Q�$�*FE/iB����̳)6�6-�<i�_'��H"@B*wp�t��D��N�$���"�$�p/\�Y����;\O���h��gK���.ֶel���1���x����'�Fӧ�S�[D��~�� 8�`Ԛ�:�(r8�8�D`��4H���ʾ!:����}�jiqr��x�$�P�'ö@�gLm��x�S�=�tisP('v�La�t��J��+sm2ʓrW&hqT 6_L`�p��O���'
�#�'QJ�0SCꁍ��0I>QG⑭Ww�2���"�$��Sܓ�>E׎ �~���K���$^WpUz5�C0m���ۛT:��IEy�g?���N?)ۤK֔4�Ec����P�*��b��L�`EY����8U�>\O�zBC�.r�l��);v��5���I�F$��=yB�@���Xץ�$�����/Y�|��{��ΟM|���C�8 8Ų�"ً�Ą`�ҡs�$�p4O��*��AƱO
�f�1�k���11�rr
K�qV�I���
����u�'�@�����Vc��Q�`���������4�� ѡɨ$�� ��,;�OH��*�}�vա�.�!\�:5���J�M�B�9ׅѐ�B�a��݇m�aHug�1�B�{�r�S��O���!ײ�]�p�a"ǆG� T���4(f�H	rapmz`RyY�z�@��m9*`����|JD�D|�󄀃B&l���gz����@��B��?	�;U$���H�2ވ���T?󤡅��.}P͑�N�f�Z�D�Ha��U��EA�R����3�����Q�O�Z��+�	y���8ڧ.@B �1���@����ܵdJ\�Dy��Ūn�B�5�
�F.@��|z���(�(�:�#Z�_������Բ'��� ��fdwcW���X^w�D�3�	�;��Q�B�� �h���(�pA�W�?E�Ĉ���6>��T?��|���u�c�9Y�^�yE� �$�r��j�v����ջ��@d�'��qfMVo,e�B�
s��b�P�օb�>9�4d�P��O��|Z� ��KG��(�!ƺ��� ��Ur����D��*p�Z$Y��7�� cK�H���Qn
�� ��Q쟘�p�^�^e��Ӻ�M?7�Ρ* ����16X�*F�6)��mJc�Y��d�<)�i�#���Q�H,�r��ȟ�-S1N��a%��j`��q,C�~r�������O0u�P�]��y�R4����&�F�hQ��(U!§@,�B��.�l��ʬ�"}�>�O��nڰ8_<H�AoN�<A��r1+�K��͓�Xt���'�]E�*K����+V=I&�S#��E�Iu��i�(,�F����F���-e����N��{q����jo�9��JTF�7�G���$S�@�H-��_զ�j�h�ӂeH )?�3}Bb��_x��\w�z����/, ��Κ 9;>�J��d�'I����,�XA"DC�A��	�H�����B��4�d�j� I�bݸl�'J�.�6Ep�D�T����ޚA��0q�Q�/�l	�3'��"j��'3wPT����0ysҩ(��i�á�J�$�P!�l7Pv��/�1\ڪeXE�5BL������ Kvݓ�JZ������(\HY�Y	��䎬R1Okl�%Q���0�܏_+Z���)]�L�����Ո)�4�@��e��urqX�*B6�B�^���S�'}2���Ƙ'Մm��'��Z5����� YPi�9:����@�"[ۮ�#��P��}�����T�tq�����6�\�O���h��y����$�f�<$���>9S�$��c�0,	�ɘs�?��r�P�Z�DI�Ok�<"B�C��"�U�U̔�����b�:Eb՗x�>�w��e¤�5eH��7�\��hLz@aYW��8q�{�-� "�|��6�KP�"�fCX�D|B,��wY��OGLC�s�@�Xş+�h�ۃ���P�{����}���HS�3Hu�u��\������ Y8�R�p{v Ξ�ē���'�e�$H(�jP�]0$�ȸ;�f��)�X%ۀI�m��$�0����� �&�ss$�s�f��O��貂�_�l���E4%�`�#Ln?�`�]m}�b\�붊�7�(Or$$��� �UBvp�C휼"	r% �����%�vq�G匜��ԟqOmˑ.��
j$�N��*� ��і\i2 �գ���M��8��@�@<z��5J��Ct$�cy�c&����q�8�¡ܶ9*�裦K݊�Դj���I��i��E�%<Le�TfK�]z>�c�(�-9�dA� R<�D�D�K<IrC	��$�;MjD$ۡ�$v���[�+��Q�p� �'b
.l��gח��4!E��Ӻ;�̛Ky�P�W��/������#K��@�&'P}=M�;/�,䯻<(�� 6�;P�LY�����ӿ�xq�FlÛCe�Ð틝_<�)4������4lD�$П~�D�v�׎_���s�gҐ#O����Q�)~���e�p=9c��l�hr�^0k(���0�V�s�(˓;A��n�7ɧ����~� *�"�ĸh�o�=״���Ŗ1Q��{rEKk�l�$��ɓREƝKT�9�"Έ=v'xd8V΁i��'�xe:*O.P�㈚cv��Sǿ��e��J�����ϚUv Q��m=�O�����$yj�!�'+�A��W�֝[X|��jN�j&! �*)^���'�^��D�X |+�y�&�6_D0����D��;�{�Fiu��0�n]me���7g�@he��'o��VN|��s��u�e�'Z�$Ԣk"��sBZh�8ɤ���B,�"���x'�D��	4F�P���*@8/�]A���1�^Aaش��ƛ .כ���83/��u���<y�O~�S��>H�R��cd�=3@�X
�s��Yv�W5��ܠ��B$*U @�rAޗo��$ش[��$�.�m�A�	u��틡vI�^cz�uj�	��\�� 3g��QU�$ ����>)�x��%� wH�ě&jD�|�ɨ
�ՙ �C���Yq
�Z
��O��[u�6�����HN�I ��3��v#����ׄo㸰("���@2��Z|6m7V�D�
�%jl�ɤ��'qP���e��aS��0z`����M��!8Uie(� ��	�72āye�ۮ;���p(˵oj�Qy'K�������<��z� �C ��ʀme��8v�m��	M��!�R 5�~��1-�4�*ݪ���>�^�j
Ǔ4SD=�p��@�mx���_zt=x�-�U�d4���G��e�6I=ʓ)�<z�%�/d5���D�d�'�HIb��N�x���buK�/p �JK���ↈo��r�n		,T��G(�I�/�H$��U�
FP��$g��5�ƆT�|�PT��h�!A��Lp�@Kc�';��`�h�pU���e;&)���ۏq��P�RG�	o����)V3���d�/1��u�`�_d�`1�9�Of�Ѡ�U:�����j�DІyca�9�O@⅕�'�4�x��VC��@�[��0�bk����G?�O0����1�fc��69n�3 �L94B%���H�}=B���nӌ�HOf� V��/Z!��KS�Ҟ^��|y�1����0ǉm[��Y�ٝ8�0��+@O�ɽx@0��#P/K�p�ڲM�U��<)T��4��T�H8u[��O Q�cC�
��p���@�<)(���* �(	@�i���w��1q�bwǉ
� ś�H�/?�� �p=!]6�`�!e5s�Դ���R�w���	�]�6Q1�@]��M����u���O��KD�.�85���
�N9���94����tTtD84���ĥo^BdD ^�s����{J]��-t�d9Cʑp����e@(.�S�G�
0��Cйj�~��اM�=�S�A�BL��p�ʙ{j�0�Q>q��8 @ųԤ�*n5��"'�QD�J�@�A�/��qOѳ���'�$Ș�H���*�	R�'�.|s�C��)
�8���`�"}nK�X\��eʖ.&ĉe��'�.$؂��%Zߦm[�jR�v�Qz�Zn`2�M	-V�2�c§��Wi�0���]��`�'f�*Xx�n�|2��	S:UG��9"'ޓOc��Q�_1_���dW�>E|h�F�1`�]�[_��А�F87��}(�H��W��WG��	�O%H����~j�'�2UD0 �lъ�\���O�Y�'�5�Ei�0!�d��N\��-���Pa*׀s�(�q(I��,��3�.U&r:C���d6�g?)�8ܚ�ڗeM�bN�e*�k�p�I�"Ξd*�cސ��ء!�]�Y��x!DL��Qt �8��'2���'"����	(�i��yU�ARC��2��,�	+�M�|��^�@oZM�;ɆSz�BK�>/ C�I���熛+�,` �g��C��;�`aa�]�24N��!�50�*C�IbfF���
�<{�$<1D��v!�+
<:1)���c�	�c!��5Y�W��4ނCǮN�CQ!��5�Z@H 	#g��j�#Z�TM!�D_�����V�ڈA�F"�0%!�O۲�4Ĝ[���:D��#!�D��n6�bw 	a����`(U�!�Q�H�X��X�a�|�Csm��!򤑒M�E(2�U�y�hm�J�Y�!򄝻t�J��TPqB��7�#F!�d
87�l�P��G�IY2U��ޗT!�$ԑ��I"$A�!U�y�S5H[!�K'D�d�x��BOQ$] hGA�!�dE�(�r��o�c��� D-�N�!��F�	L�!� ��}�R�r�-O�u�!�$ۭ	)�@�'�P�JYX`:���,\�!�� ����a
)���E��|�D�P�"O����J�1�\a�� %��5��"O<�x��g�<��&*R�V��s"O���r���]�\���~{jtr�"O�9;�'��U+DΚ�|w�|��"O�;B"�	`媥̘&/g���V"O>]{1���6��yK���5�,y�"O�y2�g:�����ފ��Ȧ"O!1�&\[X��3�$s_�ȳa"O���`��N@�׏ߺZ��t 0"O��FY9x���`΋d�u��"O���R�R+�,��(�۲"O��+gX
1�^�@hJ��"O�`�j�:80LR���T��Y@�"O��q��-��\���Ɨ �$��U"O"<�դE�kN�A3l_0��5�d"OV�����N�.�ч�H<���x""O�ۂ���ix�
O1c����u"O��Rgm+TJ�P�_N&��W"O ͪ�m�������uL��a�"O0ěEF�����1g�@���d"O��*p�%<�.ѹ@��`!���"Oġ���L&̊��14c�xx�"Oش���cp~�����]q�ii�"O��!�t�T4�B�� =ڰI�"O��f#?�F�G*EiO�eQ�"O $��� /^0ٺ�bQ�eKHT�W"OH�xg$�1c��m��(V<485"O���a/TFxbt��>���T"O\	2`�&#�l���Q0"O���Θ�+��9Ф��J�����"O�� ��C�u1z��W0�t0b�"O:H��
��'��H8H����U"OB-�����j���pf��m*��"O\y�ԣS�$J�<C���_�j(��"O�����)
�(��9L�|5�$"O��Hf˭[|<r��|�h� P"O��A�u�T)� bI��$��"O:�PsAX$�J�;f�ܷ6��P"O
��PW]�ܒ��E,ڤ"Oz��������um;2�3"O�4 aB�0d����>�l3u"O�}J�I�+y���п � �30"O�Z�-Qj���{!�Մ@����"O�������vYa7D^�0d1�A"O,qj��Q�<p`t"��\3$��D"O���Bt:�aY�@!�Th�"Or���%"��A�o�Z��"�"O��&n_9R ՒaL	��8��G"OBp�bˊ<�Y�J��(t�%��"O���r5� �)*�zsC������ȓ1��X����ĥ��#U U�2�ȓ"0�{b@�J���K��86��M�ȓI�b]8��U�{h��ʙg��% J���63C��Bk�]����(hKͳ5�ڰ��F��ȓE͎��&��9^@~y�3��� q�1�ȓ�@�@%�G���T
��X�=�ȓ3���vI&U <I�j�?D	�����J��!JD"��U�A�m�ȓ#�虢��	̀A*��X(��ȓzm�4c��Ո�,ȩqF������h���ئ�_+p2,���3w4A�ȓ�$b�%�>����H�H=��S�? �	9������|K�ʛ	����&�S�S3^����W�L"gqP�X��^6+/&C��Ddxm�QL�.�X��'���}zC�I�Z��Q!�
�,�`R��K�K�C�\@4�d~C���1#�C�	�Z� ���ⵣw�@�>�B�IO����_/ST��f�ȔOʮB�I�A2	 I����� D�4�pB�	3!�^0�c�
G��Y�G��.%N�C䉲ZTA ��}b��#G��!�C�	7D��LH�hJ0l�t�c�'S�E�C�	
"���&�"l�X}	�#C�B�9I��;3�"�b@RAdQ8�B�I�8S&�[�L�R�NpJG� *R&C�I["P�Rl�#R�:�.ٖq�VC�hq$�Ka�@�*�ybꖦNtC䉧
]:5j���h��S2�:C�O�6�5��_���C �M�=�C䉜&i���V&�;X�x��,ˊ`�C�ɜ~u&!��Ɓ�7��T�˙1��B�I=+tma�y�I��,͊!�PB�I<Lw�����X:H^q.T�$�qM#D��!�S�Lf����E>��6D�X��Gl�ĭ�%C�1�Bİ-?D�tz�ė:J�$)
��[�~~����<D��c�agT pr���6��[g)8D��w\hK"�q�G؂�ڽ9�C4D�̡ �V��0���<���b�<D���s �,���w��zQ�$�b9D�<��_;A�:�Z���X�p|a��8D���H����)Y��,� �5D� A�g�=Z�z]x�� ��Ea�9D��p���B&|����!;�Š��,D���1`�����������J/D���% W�(2!�̖G}�i���8D���jM;w�Z$�h^ � �dN8D�L���=$�L)�G����D�)D������j^ZAE�?m��A��'D���!L�	�VlKD��q��A�^�y���8F��`;,A/1I��p6m��y��A�2pARq�O�/��D;�yB"k��1&�h%�R��y�V-MJ���ҢM�4��-R7�I��y� DH�\-G�#��r�S�y�i7�����M6�p��ӿ�ybӰvbMs��^���`V쇠�yLP�n$QBU.������ygƛh��0sAQ���j֭=�y2���C�6���3;x�e F��y�*DIs.�R�͒�  u�ߠ�y(��֐)3G\��*$[����y���{D�s�	T�����·�y��Nxl�('��2��@s�l �yfΎD��)V	P�4��
E�B��y2��w�����,f�A�/ϰ�y�X��Z]����G�̕�����y�O*i�H�!�eO�h+��y���&�y��n�lhSn�:\)0@�S"���y���U5@x�ŋ�Z7lQ���ш�y��(a��5)�!šTT��!G��y��z�(����&P$θ��(���yRDY�,Zy�P 0C!������y򀍈STꕠQ�Т>�>Ր�*U;�y�I�-G��y5ŋ95@�E���ي�y
� ��zf �UtL$ �cTJl�@�"OL��iɾetՂ�O��@�X�g"Ov���]�U��L{6��/$�]p"O��GB\s-ZMh�OF8��+�"O �>o&���#,#���"Op�/�V�@�d�0�0$�$��;�!�d�t ��p� 3\�$���oݓ�!�� �3�@Aa�]�"��X���x�!�D�>t�%���	jk|�)T鞪�!�$�� zH�Z�TgT�#(��&!�D����Ո��ޑ~�H=j�F�(!�DK�C|J�ãOA
H�<��vQa!�?"��3�>�6���#��a!�$ִaGX}[6�������f�ˤ4v!�R>}�`��wK(��I˲+D�B�!�U�rv�����j&�4``jq�!�$�,A�"ݙB�;9��I!�H�>t!�ǳ	�L}�3��o���s��O?W�!����V"b�`$� j�L���mȐ@g!�$�	}���Ȉ�R5+����!��(+��0�"�o�T �$��5]�!�D�y�|Q�D�"�\�)p�|!�B�N0���H� %�dAд
�3K!�D�8C�X��_@��]y�.V�nP!�DS,/i��R�L�8�>Pb�M��}F!�ȗU� 1��TV�pnO�!�=j�4}
�f�</��C�잌%w!�$��NTJ=S"֯_M"]IS^�m�!��wDT��7��5���(w+M(%!�JRe���,ɆVώ���ϻe�!��#w%J|�Phʘ�5��Ȉ�2!�5��<���Zd>h��
ܩ|!�5W�{S�\$<�6\@jٔMm!���O�<eC'h�$F��r��'aa!�
a�l�c㧟���E.�[s!�$ɄF�ei"I+N���3��`!���hpD%�v��9�Lx���^�sa!���z(�a*,

�:�7��-c!�$�t��Q��3@�d�#��D.fW!򤗀-�~��uE6rn��!���+9`!��2e*�+&�9Y2\uI�F��|o!򤇤n�`���Ɔ�g,*���=3k!�d�7i��@	B����cI8`!�D4��$׃_�/A.�1 �%QS!�DI6M�ֈ�V���!xHƉL�x@!�䞢u ��s�؟f��S�i=!�d?�8��T���fE 3W!�d^4'"�8"�F��NA0�Q?G(!�ā�W�܄!�'��5ӘKG�	�9!�ĆNUJ2q�k���Iל�cU"O�yX7�6!��R�N�9T�.	��"O.@��ƃ1�vԐ �̙`�$ܣ�"O|Y�	߅,#�h#m�#{���a"Ol8�����t+��Kx4�bt"O(@"tDS�Y�VQh4qE� �"O��Sp�_8�4\H�f�	5A�Q`"O��P��
�&T kBhr���J��yRN��0���	�?&1hR
�y"�U�B�ܠzs`�.�&U�AU6�yR�ڼc�]�����d�ybT����D���V��염�y�oˍZ��P���3
(�l��F�'�yb���D&T}Rp�i#A�Dr"���'^��b`flT.�ْ�٠+,PB�)� @��^ Y[<�.�_�����"O���F���qr��2¨\�"O0L1�/V~8YPː��h�"O��pvLڊKY�L2qHE.>.�I�"OvsrN�V1��M�`���t"O�)ӣO������:�:![�"Oƹv��lC@�\;�|k�"Oʘ����q��0th!�8��v"O�8���K��� h �znB���"O��"���DA nF�(�^�q�"Oبa&���>-&P��lK=q�q"O(�3� ڭr� C,�"?_&L@�"O�X0�"[�46@-!$�W_2Y�"O@ۓH�1�T�) a�._^"�w"O,�P N�U��؉$��g(��"O�����۩J�B@i����	J�"O�A��6D
f���۶q�@�j�"O��B
70Q�TH�C��k���ا"O�Q@���.r�
U(2�V.����"O.*dèY���MJe����"O�E,��y"�����i��02"O�d#f'� �(є�U8.����"O.��։�5n���mN�k�0@��"O� B�_%{�Z[�U��|�"Or[�L L��8�v�O&F:,F"O�$�
ϖ1����*ПJ`�C"OH����(�n�ɓ]�]Y�6"Ov���'�x��ɕ�$YHQ��"O��!��9�����	�OVF���'^��vK	��Ȝao�T`���'^* �����S�^��Dٺ�' ��q�*X
'ߤipu!C48TS�',����#�@�"5�d�גt�MS�'���-hdYU<��)�ִ�y"l�1X�D��EE�I���ׁ���y2`��.n ��,C�A�ۇD���yr��l>
Pa`�"൩����y©L�δ�����$S�Jʉ�y.��6�{���#W-ذ�U���yb�Ǯt}�˗	<H��C����yb�N�\u���$9.�{V&��y+�<.,��*�3VbU�B���y���O
�0{�k� &�(I��ぷ�y�'�)-��dK�+lL����y�/!t6�r!a�|���$b_��yr��Y\��A2x1��#5�
�y�̈\��ڥ܀rnx�D�R��y�c��jMf�*�ûvx���t�̺�y���T���Ė�j��X����-�y�EQ+u�`��ɝ&d�ěbLӊ�yb�R"I�
xB�Y� ۑ����y��85)J�	a꘹'�5��U��yr��:h(.	 #�ځ'��i��Ċ�y�β��9�d���p��O�y2�Y�� �b���1����
��y�bB���*��p��,I����ȓ^��E�'H��/w�d��ǍX�f��ȓ[6n9h��_�qW>d�*/؆A���͂�A�\�����)K�V��ȓ]f�bBD�5�p�p�C
�bͬх�)2<�'"=�t�b��Lb������	���3���&�?E��@�ȓ&vl�Q��E�ɜ�'��2�u�ȓ]�|�C�C�Qy��D
�|���Ib������ �SA�ޖ5��Y��Dax�i�"O��ѣ	T�$�zmi��P��"OP]I4�3�myC��9�v���'����z�ǊB[n�z�I�6gr��c>D� ��aH�z�ZU( ��7j#h�Rf�:}��)���
I�-��B�k��j��E�ܖC�I�])��:��_�4#�}�f F�"#dC�I���)���]`й��a�sQ:C�)Q�[v D�lL�(j+s�:�¦!��2�&��_e0$#�d�6	+H���"D�H��#}j�(�ƣ^ ��!-D�L�Bb
�Cl0c�C=^O�I�#�,D� k�F	)ńq�����%x�*D�̘�O��"�؅_�Y�b��r�(D�����u6�hȊ�/e�\Z#d%D���".�/,u�쫴A�z�Id#D�pa��L�Jf> ��m³M�D���.D��$z�-��FM�2͒1F+D�<�0ĕ�^����n��i I�-D��(�8P�$���K"i�ЌX��,D��;%H	�byș ��:��P�a7D��D�77Ud��EI�?ψeQ�-(D�L��ߣ�X@Еb	�X�fa�,&D����-̮B�11�d�9�T����8D�8ef�<.��4d��E&@�@`)D�D��M��Z�۷�̔T��$#=D��af���}cԭ�]�,x:cI;D�8iV�[T�����������o8D�P�%��$AXFQtU#�(4D����I%O���@�Ym�b�Ip�0D���\�z2�k�1e`�4D�tр ��LM��BV�O
��Ũ/D�T���ӧk�T���DR�N���(f�.D�؊Vh�f�ɰ3�ݘ���cl1D��!Ш܆x�0�0��48t�!{��4D���0��Ĭ	c� =^-R'n2D�Ġ����Bc@��tM*�4cԦ"D�`Qw���ev�IX0臟W]�a3	<D� C�bS= h�⊑�~�����<D�hs7�^�q���1��[5xޞ����;D��uG՞M�|a�Y5|T~5�t�$D�<�e�(F)� !X*�t=2��!D�T�0��;� =вL�8x`1y5�>D�� ���3x#e�q<�Ȧ�>D�lag�,GE���/Y�,�
�#�l*D���B㋠M*���7��;�*��-D� ۄM��D� @�e�[$o�=���5D�9h�:f�A����h3i�g(D��!T�>�=-D�]
U��`JB���6�"RKN#:2^�ѕ�]9�8B�I	Z HQ�,<3=yX�'lxC�I ���6��DZX�9�,�8&6�<�S��M�V��d/���E�@N�&A�l�g�<�So�X2�ub�F�"dv)�u�g�<1B�X}��t���+6u�ɋ� �b�<�v��u
R��bo���"jZ�<ifU�����p�ǡl��p� M�<1�OQ�{n�Ece��_[bU�TAK�<��#�9��pG���8�ʵ&�R�<a�aǶ3�j�t�T�v�x�@�Q�<ᥥ�){��Tx�I�+3��4
Em	M�<1!/�`�L9�"�$=K�P;7�WJ�<���A-*���c���kXb5���RD�<��ܺ.��QH�86X�b�H�<�  ��[�w���$�.E|��`"O�Q���D��u��I�g,v�1�"O$�zd�J�0L9#I°t��Ћ�"O�쒶F�5�`�x��at ��C"Ó34���jjPl��F
�Fur��A"O8Q��-��\ID��)
�l�a"OF����S�UN?Z�2)S���<�S����0b �YC����r��w� ��y�B�.nلYR��S/ʰ�����yr_���H��Z�R�	�a�y�
1���A!�Tݸ4���y�@xg
t��c�L��|sd�<�y���@Y��pp��Cc��k��-�y�H0H�:D�ǔ.l�"Ii󫊗�y�'߭t/rA�DKXss�e���#�y"*�����jԇ}TK�'kX��ȓdb|�p�ВP�>�� �?����&�U3�قg�j�z4� 'Mr��k�^����=��B�ןC�h��`�2e��I�<·֝H��؆�G�t �T���9��.��D����ȓ]i !�qc��:L%�5 j��)��nT�]�@%��CO8����/\w~���G��]-Y���(uD��6t��P�2D� aw&L5]�4K6�߅
ib%�T�#D��9�!/Ҕ	�n�;?�RY�b�=D�����W;�i�g�	T�1�x�<����cH(D��lI=)��fO�O��8�'���CF��������̌����'�8��g�U'#%���D۶W",<1�'��Yx4k��WFP4����z���'˦��d@8M���##@��p$��'&����4�q�r���{�Vh�'T�]�
��@u2���+�Th{B�6�S��?	 �C)�@�`O$O��9��R�<q���2	� ���*`�(�נ�M�<	uƐ;��1�)ci�pG��H�<�`Q�q�ᑵ��D�ޥ���Lz�<	w��#׸p����W;7�]�<5�m�t0P���cE)�רEU�<��)������LmCa��T�<�c��5^����a�
�
%�`hNJ�<9�ĳ?���ōN�s������E�<�� �E;�q��+i{�
��~�<�O��H�ss$�*��}�<A��'p��{��H�ڽ�էVP�<�FeV�'����p��fc�2c�K�<�� ���*w�
���еc�K�<1 �ֽ'�v5 �ի@4�ZfN�F�<��&ѷ�>�c� �6&h[�F�g�<P�&q�T����8K�H9KC�i�<)#,̃~5lq����~��a�PE�p�<9���+2�A��E_�^�H0iSG�<���cwzE"��#Jʪ�8v�D�<�G�i��)�v�L�#��ȳu�}�<�'�>���@���,���S��N�<�ïǑHLPb�E�\H� ��M�<� ��P��+B�!y?,[���^�<1�.��^���S�����2p
_U�<����ed�1�D��0'����O�<	�(�5v�l�AGԖ4�\|�,�H�<	�e��"�� �F	=qƍ!��y�<!�C'��(���.�|qWz�<�҉Z�Xze0Ʀ�^�0��}�<� nd�B��M�"Ez�H�6t��"O��2*�%!F\i��GĪ���"O$�9G qw6����ZX۞̓"O��Au�݉0:�x&�G� l�Ѥ"O���➽UX29q+Ҥ(���"OA��%�k\�PI��X� �n�KB"O��
�GN�:2�Aj�p���c"O\q��G�*x6&^�'���"O0��W��o�����؝4�11$"Oެp��Ǽ���/S�Դ�"Oܴ����op-(C��it~ո�"O��F vdp��$��76�)�"O�(�A��2{	�T[�A��:( щ�"O���F�0;�*�K��Yt-:�"OJ�� rvH��4��Z�R�"O�@��N-�^���ٗ�XU�U"O$}���Z�ML�+�JA���"O\��lY�jO\�G]m��]�E"O�4
ď֒2��$�eD�$�8�E"O�h@F�5�R�B�	�z���v"O �"�	O�{�
=9v�"�:�;�"O��`gb�@xT �"C�UZ>吆"O����E)p�sU��0A �qe"Ohh�a..&R�Gf_�B��t"OҜ�E��?~v���ٹ�0�"O\iy�	O�E�r%�eD�A]��#�"O@<R�膉d�|@�]�J>h�u"O�ٺS���S7^ "V���"OZ�B�9^�ZtH2f�G��%��"O%���+S��%Q�	?8�\Yض"O mɓ��3]ά�tM��P��t"O¤�Td�1��P�w��C<b��U*O1#�/N=7*֡�$���4��'�x��`������ɂ��x���'lx��u#]�W.9�ƒ9���'�&��I�a��b�̝�z,����'r,��eI�Gg
)w�/r&8r�'�F�r�A΄���A1.��!3���'�0�#l�`��M
`�$P�h��'4p�#��G�\�AUO���A�'�F�e�� P�X '`ED�@h{�'���G&�*4��1�64���Y�'Xx�؀�La�R�@T��(xJ���'�\S`���-��(�����J6����'��\{R��}�2�߃G��J�'��]�!�@�:q�%�1e���9A�'�P���O�T)�r���:�|1��'�Q����l��h:q�L)3� E��'�2�	֠5�����ؽy���k�'~� � �� xn�%!0+ a���'Nu�a�1���I"�ʣY�5c�'�U"OԛS���
S�V�K�6��'P�@�$,,��/ǈ@m~�	�'�6h��3�����a�g��'���3�`��]��hæ�P�Z�\*�'��FJ�)	�x�&*_�z�K
�'T�Tj�M��v��X�ńğ[�\`�	�'S�,��EҲ"(Yre�<D����'R\a���B���r��O<� �1�'ژ�1��� ;�Ti�ɋ>�e��'��4��C]��Ã��;�$�'Of0�0-7K�����3}�	�
�'�f��@��Q}�ҭ��~��!
�'Zl��W�(c�},��-s�MK�<� >Py1O�QB���nӸCP�P�"OzE��	�sN�trT�N�z�r�"O�)3���C��]1���-!���k"O\Ԓ@�ɦL;��l���#�^�y�M(Q������ȶI3�P��y2�0�>�����Ek=Pcg��yG��s�R� �Ԯ;���Bi�5�yrf�[8�w�-S�Ey"!]-�y",���.T�C$z�t9BR��y2$�-)ԄR�/n��Qz��	>�y2�@[��4�A/�$}�$�3K�$�y��ՙ���܃h��H���yRn�ִL
�"�dX�hEBO��y�JQ%(��y*ۑH2N�0H��y��ì?�F���F�9��D�"���yi	2n���sI��|�E
5���ybM\�bX,I��j��o�Q��D�,�yRL����A�3��E �&��y*V��@Iӑ1�zH�U��yb��)����5��0��YA�����yCһD�|\�rn� ����I���y�,��,N,�`/�m�՘��Ҳ�y�!����L���]���i�yRVL��� @O" ~�٠�ȣ�y���3YTz) ���+w�:����	��y��\6p��ZR��{JF	�F�Q�y�P^[8Tc���@�d����7�yr�OgB����r�0�1�m���yr �9�N�KT�+yN��IT�	�y�kA�"-��@�N��l-���P��y���\�$�(�w�2 JAX4�y���8#��x:�k�����ُ�yR�ï�D�èVP��p��*�y�&�� �����
�"���ʣ�y�	!r^��q1�W_�����y"�49c��#�b�����f���y���.j���80&��[�`!p!o^��yR Ճm���IҮ�L�aR�A �y�<h��mc�K�GN�� 3�y�Z�k�L���їA�p]�qcM�y2e�j�b���P�8���2���yb��<������hɜ�������y�M�#g� ���Mh052D�͖�y�ؔM6P���ɗ���:V�X�y�B�;�д�`́	|�R�M�y��ɖs�4�`G��6����
[6@B�	 #>-��A2j�X�����|�B��}��������4�X���J�B��<k���ǋ�a
ӢDjy�B��#�	XVG	/4�T�c��p�jB䉜Gh4)��.@di�cR03C�ɋD@J����0V	Yu��
W��B�	<u~^-�d`�C�,y���~��B�I<-�ޡC �8f�5{bɈ I�B�	�o�̕@7�X?�܁7�ЈB�IR����گW$�ܱ#暈@�B�8}F&�9�^c��Û�B�	?G40�k �@Y�Q��N�FMJB��`X|��ĠE� ���K-[;�B�I��Z!I@O����`,��B�Ii �U�"f�a0�A�B��B䉲=�V�ٶB�3J;�C�W<�B��KnY0��Xmx�9M%hZVB�	<QTPS_�H�nye�19M�B�)� �x!�,��A�-BT��"�����"O��(s���xa4#E�*����a"Ol��#CO9]�)Z���<��*�"OJ�)�\??�*�C���>���"OZq�A⒕"XVU	�1;1M�yR��=��$ȲlD�}��R�]��'�.`����x-&��Q�+
�����'S�\j�&ޗ6����O�zs|���'��5(q�L-wt�0��Ô	(�U`�'c��8���Y�f��F��("k�a�'�	��F�0tv��b��!ž�J�'�D����ޝc��P�����H��'���BA�eQ��3@ܪ�扢�'�Un�� 4�8c �;����'����`Upn��(��Yx�P�
�'������,�Ա�d��>�`z�'� U�Rn+���`rNѽ��D��'XL�4��)��Lj�*��mz` ��'@y���e\�(��A7i%�h��'%� �ŗe&Q�@�YN�s�'{��� ðPaJ���aB7S��`��'4����)���2t�e뗧PT���'����`��
W�fe�\JĐ�H
�'�����F��R49���j� L�	�'F���#G���c@M>bX���'U�y��k݃XT6�a�%ΰI�z���'�T8��!ӌm�F9���1�8�	�'�z��cٴ)�@�Bv��y:@tZ	�'Mvm�3z  x`%��r� x�'լ�;�mʑ*�ZM���f�\��
�'ܸ���.� 8����e�p� ��	�'��D���R�S�`@.a#�hJ	�'ۜ�Z����N���4��
����yR�^'M_D`�މC��5�٢�y�HM5#��� G��=�AJ5�G�yR��aNh��Q��3.���#���y�_x"�P�|���������yrJކ P�t0D���s��mz�j�2�y�� 8e�DK�%�q��@H��y�!��i8J���h�3!���y�U s Xb�׮՚MQ2�S8�yb���sy��Z$ʆ���݃�f��yrh�0X4t!Ѯ�H�s���y2�8�5RG,�wfx�`���y�ɀDN]���Ÿ�a�j	�y��¨s�$��
ν�l<�����y2ж^���i���9r�S���y�i�"umV�����+���1�I���y�O��Mk����Ol��I2� �y�C�]旔X�p+#K�0��<��'b�b��ɠ$S���3v�*i�ȓ���S���Or3"h�=)����?�rx��9I_l4��#+�*(�ȓU���0�8����,Ч(��ȓ0T�Ր�M
3h�a���E!�H��ȓhT�"u�ݵR�~$�����oF�e��B�� !��Zj�$Q$�љ3(�p��t�4�q%�(d���T����ȓsur��nEf�V��3�p0�|��K�Z�M� yߠ5�ǀ��1g|��#�� X�D�-��P�"�:\O4�ȓ6���X�b���OPp4n��ȓ>�,K7�C%g��X&	�>h	�=�ȓ�`� ���+�� ֩[��Y��S�? 8q�pO�g��D��b��U���I5"Ov����BxT=�@��&p`�B"O�U!��5F�8��FB�O
p�%"O��f"�q�Hܱ�a�&��a)"O\���K�5�P�����~y<8
5"O��s���U�1H���+�~�`f"O�9���E�p"Vp��$�+}�!&"O�ac�e@�Ԃ�T�+]&u��"O��H#c̍Tތ���w��� "O�p�JW�.f�JR��>c�6h
�"Of��	��!�l�Bc�"p���y�皩C5�qc`)��:�za�(�y�%AIV`dC�e��&���sR
��y�D��:a
P��!�*�˦��y2��&E~�41�坾�}��4�y�h��j+��h IǖG���1&[$�y�n\��4�u'�s���pG�#�y�I�
mm�L;�Βk� x�E��y���=|�B���匲9
�P�6��0�y"�Ӆ�@ţ1J�D����E��>�y��D�THZ��ݷ4�"�9�#���y�A�w����$Ƈ�(��U��K*�yҍ,���>p;K7�y���P��a�m��Rr�-���y�U=MHR�[��F�9!�m�⭀��y�⇍}�ɻf��#1��b��2�y�K٤mv��;�ƍ�r�L	���y¦�d�f|bR���i��)���4�y�MP#F�Z��H�a�F�#
�?�y�LZ8t��]X�oΉcC�ى�B��yR�۴H#켁`�^�� ͒�h��y¨�2�tIC���=��+7��yoy�J�D] 2��6�C��y�����&��֨C�ų]�TP�ȓn�\4���ڎ$�N���:�X��jqꍹ���=T��Kd�_pM���w�R�i1m�=rb�ɂ �L	j�����w	���MD=y\\�S�3Z|��UNZqz��$d8E
��^%�	��Y�䩰�L�3j iQ�
�o��,��ee�H9&�L/ISԉ']3�i�ȓS$�(Q�	��>����ԀE�>�ȓ:$Ƹ����[�z�*Ǝ�'𲀆ȓD��)iSd��+���A��]:]P̈́�d� wn��P��A@cg64�!���H�3w	��*s�8��)؛5zH��phm�$-�w���c�_>�fq��)urh��Ya)�QA����
DP���&����J�P�xk6���Jִ��J��aNF�B���s��6�
���ź�ّ�p�$��T."��ȓo� (J��8[�`��BHZ�>�HT��FV��P��A�"ur|��G��J��q����@C��*�jEK���1��%�ȓs� IR��
QJn}�CKԓ� �ȓap�e��ʙ1hR��i��V�c�^�ȓ6	�X���+G��ɥ$�M����B� ED��L�F�Y��ՙդ���4?�0�V�*Ό!2��@�5��d0�P�'C6O�$!uU�!!�ȓeZ�Y贊Ĝw�N�RG�5q�`B�^�Py�w�S1�D����>!�VB�#6�v�XԊ�$moM�Ǧ��"�C�	�	N��c�[� u��#�:��B�)� @��ebT���tjB�1S����"O�(3 �+ צ�1'J wF4��g"Oh��D��'�� ��f��n@*u��"O��j ��2 e�I %Y53���"O�Mxb��r�0���	(�b�"Oё��V��T�b�}{�a�0"OHDH�l��+|�`��7�-x�"O�P�؃pǐ4H2��>X]zŨA"O��+�	[%ְx�Q"�=vW@�1"O�Ur2���Pu2��<C�B��"O&´q� �)9"�:�hR"OΡi3҇[����ؒp�4�!�"O��q�H�&�1���9	�u�"O�p#�+H1�¡a���-�����"O��P�&[�f�8Џ�:j��aq�"O��a�'�C;~�4�2�p<�"O��/��9i�%��M��c��	�"O���O�a�|���O�l{��W"OJܢ�I� �^�@-A
Xhjq��"O.}��A�7҄@�dA�f 8��"O�u��%53<�UF	=gw>iB	�'݆�R�*��3�n􀲂�&��P2�'����j��#C�)h�o�	0]��'t8��獽*��� 6n�}.��
�'o���g_5p�� ��:@j|��	�'� ��	h0$�СM:�R�S	�'�1�&�]�a��Q57`�p�' �P��0`���1�Z�z�>�
�'��pa�Ņ,{$���ѿs3�4(	�'��I��;{y&�����	p�Z�S�'�µ0�L w��YҒR>h�F��'in=�b�c-("��M�����'!h��)�`j �E-@��@��'cT��M�	\��:@m�
I!r�S�'�2H���Y�sF�8�	�Q� ��
�'����a&��8 �B'+R,� �
�'3R){����lBgc�I��0�	�'�е
�)��MN�����;�V,J	�'hQ+��sLYzq(X&3�@��'�<��F"L�z@`�	�#ߖ%?����'��w�
 _| �U�
)��
�'Ү5��\ �>�۵��X|��'��Uⅅ��[�.a%����X�'��pK��0�h �d��v�A�'����ΣF�D���WĘ
�'q�L*�BB<q����"�ԕu��1�	�'�
���Ƽx����s�Ҹ9!f�2�'x(\ɢG%�*}���&4��
�'"�1�5�D-@m,	w�Ի.�
�'%L����Ǆ�\��ܣp�^=�	�':&���+h�xc�ŵ^�ti
�'d�u��n�9�����"�J�*�'���a�ݖ�t��/G(D	@=p�'2~M(�b�;2Jh�"e��C�vXH�'�N�¥��C�t9�5c +7UԵ�
�'����Ӂ��A��<�$�������'"=x2���5�\���,J(}pR�b	�'�
as㫅�0�t�U�9�} 	�'��ef�3TÞB#��o2�x�'4r:�Aܸ&���5'? �b��'���)�V�n���;hH�z���'�4	S
߈J��te�u�C
�'��aY��!mp�Q@��جx �	`	�'I���DωXV�HJE?iZy���� �@vĖ�;'<0�G�#\Ԓ=�"Or��G� 2Zz���<N�ȱ�s"Oʼɂ/���@�y����|H"O��J �Wqw�q�!b��;�~�x"O�9��A���C˱Tق]��"O�(�����}P��y�BUI�"Ov���D�b�l��ֆR8;��#"O�-���wF\�{b��M��f"O:,%�;W�D�!v�/o b"Op�{C�D7٪�X@�H�4���2"O�-cFΒ�t�88�i� up��1"O�4c�@�Pڮ��c�ݦ\�!K"O�I�'I��<�������N�B��"O� �*r*�q��5Z2� �T"O<�S%��t:�ȩ��%�U��"O��E�}{^`S�lU�'���"OF�Д� Ԏ�r���A� S$"O:�j�T�A^�1�I��k%4��"O(�)E�L�c���XV�ڵ94��v"Oh�"`G�-��:��V�ݐU�A"O(|��C� ;�PT��&f�j��%"O@���JS*l=�df��8!��ض"O��t'�>:���W�_;���"O�8� "WRD�BU�����c"O������ W��s�׺L-�\�"OTX��L?L@�t�b��'J?��qq"OȨ�f��v�൛M�Y=����"O���C�����05�߮[�l�h�"O�ڥm��7&X�� Ԛ)p<��"O�+V�I<T�0���@h_��"O�9�BѵE������ ?Ep��r"O8`Y���:�
�Z��ö�B���"OX*c ܝTb�$`� �A�[��y�$d�R-{��Ā9�6Pv�Α�y���}��a1uޏ"hae W�yh��%ޘ< �c��,��œ��yB�E3dV`�tj+/��#�M��y��Ο[�N�k��Ѷǌh���D�ȓ;�h�r�>>�f�gJ�>S�b���|��R��`h"d�X�	�LP�ȓ/:e�M�0�,
��Y*Z�P��KM�-P-�TG d�%ը#��ȓ;��)�b��?&��mN$_�Pl��"��� �� �I.�R����J�y�^=c�lp�������4\`�����J�g�h�Ƶ�ȓ-8��%k�?�.�ҒKJ.2B��f���&�,{�����j�o��8��#���jĹ$�>�"0�	){�t��U��mX�� U�0b2	Bi+
��ȓ+�ȱ��%�H��tD�Y���ȓ�f�$dW(�¡�dN2W�p�ȓ.4�8��H!b�NI��nUVK̝��n��,�o<"�������Q�t����Z�j'��`u�a�G���U�����s[� D��\^�5C�T[���ȓ=m­XǭI�
G>�p�	�q��ȓ ������\"���}��u��b4ء�uc]8-���)��}�΁��o#L�ƙ?(��k�J0x�8P�ȓf5Z���Kc����GϦ(��)BTL�GB�3U�nb�jΦ#0�ɇ�&$�(ZǩW�V��0[0`G��Մȓwͪ0!R��|ʘm�!K�!Z��̈́�S�? 8l����
�b!+G�)7}R�9�"O P!���\� �)t
�d��"O<m� GM r�F��i
qr�s�"O��j��S���㒏�2Mf$�kA"O&����5�n��
 ?bdi1�"O�p��0@hl]z�*Ţ7X�m	5"O4���C�6���Oח|RRt�"OF��+N�*�ȋ�-�>wBV� �"Oص�� ڰF��h�����U��`5"Or�kA�L+<JH�ʅ�Ɗg8�z"O<��ĩS�bLT�;�.�!5R^�"O$PQ"铥b�B���lɨ	 m�Q"O|Y��Ǩ�v�K .�H�"Or�f(�l������s��Aw"O�գ�f��$(:uOJ.!�PH�"O�,��k٫��i�n�+xhv"O��zs��?|�"���9r@~M۵"O�Q���ŗ\����ю3!ƼG"O��"D���r^%K�l]9��C"O�La���S���y+L�<+�<��"O��!�V�
a
�F�d+A"O�6A�2�1'���'dnDaG�*D����ܟ3!�ب��
�>�ZH"`�-D��yG쓶,�֩耇(@p�ۤH1D�����x�d���"��l V�/D���q�љViȴ���N�l%\��6	-D�,�G׭��C�$�T0�!VB>D� ��F;S�HU�bfߚa�,Pi�'D�h��/��K�� ��J&LI�`$D�L��ꙵx ��T陧#�eJ�j&D��B�]���a)���#@��h�!D��z��>I@��B��78�����=D����Q �
�
 	��7H�9��i8D��;v�s���jC�[>��['�5D���vc�
�q�CWIz0����1D��*t�T5w���ѵ��(
��z3f1D��H�iM:7H��A�Ͽb�Ie�9D�8�GN�VI	r"��I�����6D�ܸ��#0w�pq�rZi�QM5D��bp�Y(-$��Љ� c� �8D��Ȕn]\���+��t��5D� X���m}DE�/U[Y��S�1D�8pfD��T*T�S�KΚ��/D��qM��u�l3�JC4Ά�q!d-D�H9E���K��) (C�O�"Æ�*D�T+�JB�"}8cOV�~��G(D�H��E�S�j5��Ǵ����3� D�(
b�?c��Hq)D50�p�8r� D�h`\�:�㊴<��U��ի3
�C�	�b�qp�>6���z����B�I� �b%.K0�*�`I�|�B�I�*��� 3��.6��	pe��B�	�:�(�R6n�)� ��X�B�	���	�����.���.8z��C䉣k�Hɘ�BG��i�nݾ
��1��l���A�O�~��U�j
�t[����	� 90T�Ɏ9�֙�$a�8���4t��i�Ù�v� {���th��ȓG��ź���1͸D#@�
F�i�ȓ=�Pr�$ޮ;!�2�A@�C杖�ȓC�lipcS���x뇷�ل�M-z�srfN���d�s�	T� ��ȓxjhe)���0m�x�%�� dB؆ȓS��0x$ڟA�6YZ��!o���S�? >� �·�κ����ɧ��u"O,�R��ν&�V�"�A�n	Ɣ�$"O|� �T�S�"Yj��Q�	���"O�@ �l�&
�	�q��|� ��"O��Zt,˂LH	�Ú�:�T�I�"OZ���͈[N�0��(m���[�"Of)C_e}�E�S��w�09��G_N�<Y� �N���A�Ǽt��=brFo�<�g.R>w�4�
��<@X�,J��yRhJ��� M,k,�C����yb�l4H���OM9��b�@���y2cQ(*ð!�#N�x3�8��̏�y�D(Tx��u�Ye�¨P&�^��y�@S$}���`�a{�<���B��yr�	�K��AA V�R�`a��O>�y�E�`�n�j�T��e�d�3�yrώ�E�� �d�C�^RL�QE����y�ѧ@��Ѓ嘑W�^�tb݄�y2"A�KHf=1&BРN4ͳ�	��y2��Vy��
 �B���"����y�#5BT�@r˟,j��=1�韬�y��vX����ړr��H����-�y���!0°b��F�a�DUh�.-�yb��SS*�`�U�Mf>�� ͖�yE
L%��!X��z��o�yBB�8w�� 	gn���\ P΂�ybbۿP=Dh�`�ܪc�qH�-E!�yR�� ZU�({�*F��$:$����y�@\�[$��*�#8wn���R�yҌ^"N�v�Z�r����F�W �y�	=r��5�O�@�h-I��ǥ�y��_>wL�1���)���ٖJ��yB���%���I�D �����K�y2M�-&����"T��C��A7�y�Ѷ%�bz��F�Q�PLb����y��M�x9��(I�����㔟�y��	7b�8Q�E.��Hٔ$�Ņ���yB������Gː�+pNX�Eb�y�̔�#�mq���W��Di���yR�
�/f���O�0�����	�y�L؄2Y8��M�<�+ ���y�![�:r|%�`�D1B��ǧL&�yR� !f����֎Qn�$D���ó�y�˟j~3���>l�`ᲃ��y���l'��%��6-@a��yRN֞#�j}q�\�*	x��g+է�yb�La���ץbD�(� ��y2���Sڠ%��,�!�\X��y��/�貒L0���pb�f3!�䚋>�|��r�^�fEx�!#!�[�!���J�t@�J�ǚ�H�`;�!�^�Gy0h�c�Y7w[�Mآ^�!��7��P+CKǰ @�92���<4�!�d�aUND�3�
>'���ъ�q�!�dH�bu��!��Q�Y{��9x!�z��D����_ux|��F!�^5�.u�g\;��*��):$!��Ϋ4���E��tfHP(���K!�$ŋL�P�##ɖ�sEX1��_�&�!�)�$=��G�}ֶ�)���>�!�D&{������! Z�30)�0$y!��G0�����&B ZP  ��7Cr!�䍆-����	5�l�5*^!�$ /a�� �ƽ,���b�}@!�� �1zAh'7���CVl�9A "O
��7�w�����0����4"O��0��G�'�h����2L���r"O��I��ܛϮ�y�K�u�Y�&"O�CC��w������Q�`i��"O��;ׂ[ J�pH��Xڄm�"O����&6��Q�f���p�"O�r��\I�%Җ���	���"O:����S���,��S>pԜBV"O��JST�s4�"H.z��"O��9d㟿G��QW �6(0�A��"O`�a��A"���*-�6�z�"O\��5d�,K��k�}��	� "Oܰ:ń�K�,�
5`�=g�M `"O��!U-�!��	h�d�
D�.�`"O�Tҧ�P&7��u�����D�V"Oh�!J���4�/L8�ԁW"O���E��z)��b�	!@�P�"Oԉ�%�V�8e��H�ZX�d"O�����
�.
�Q�S.�$���"O����2�l �f�7	��"O�if#��}���EQ{7"O^e��K�{b�A�*��BXr��"O�9Z��Y�3��a8iA;m �u��"O�H�6�F_�%�6�F?|��"O����N7Rn$H�D�D4g�њv"O*�� � 'j�)�$�V�j]�"O�,��J�K���r�����0�"OZ|� �Ac�}�Cj�)Z���"O��v �t�8��I��"�"O�̻�lD�u	��q���k��c�"O��ˇ ��^��V'xJ�ڧ"O�a�'�#k�X�����'*e�y�!"O X��Ŏ�_����i��{@
9��"O*\SV�R�D� �(S)�P$Dm"O\����2}��h�j�>�:	h�"OL�k�� �hQ��I��E���S`"O�U�#�-)P�]��b��	yG"O�%���cb0@����?�`�k�"O�0@�7��*B�L�)�V�;�"O&�`p.K�Yx����l�����"O�)�ЉϾ(ؘ�K��@(%J���"Oй�q@��*��0���F�	c"OD(�������A�d��	�:�J�"O�5��i7@P�!
� q#T"O �"ǉG8x������޾$���"O�̓���K�p�R�G�@ì�a	�'����-�	2D%�a�/*�~T��'�D<�JճiY��d"��r�'�Й�ǡ�8O#T-��Jק���'z �T̱pʼ�E���b���'?�84/����L�=���'��	� ���vt{���6�P
�'�Ѻ%W����5��t���
�'���P N)D��[�͌ܔ��	�'��uiU�]v���@���~��Pz	�'�~��!ڦ1��dW�?z�p��	�'bH"�a>�h"�D�{a$  	�'��+�O��ʙS��Σzy����'F�[G���\7�Z�F�v�Z���'�<��C�	�R C� ݩpX|1�'�l���*2�ʽ�dIA7�X��'���i)O?�9XH[/-�΄��'��P�M�d�hX���8<������� �}*�U�w'��ڕ�F�+��5X�"O���f̾��]�4��h��)2p"O� ��Ud�%1alK%(�6IYV"O�a`�OT�.#�%�2ɛ�|v`x'"O�A��X��"�ǅ	L
�C"O�9oQ�X���`¦�'}b�\�"O��x��#rFx9%�7��c"O>M!�g_�g��D�fm��=xz(zt"O���e�ް��( pI�~�y36"O��	��_?4+��"\7I���"O�%r5/�8G����A	�KCFɚ�"O$ѩ�*�]� q�`��2Cd��"O�i�K� ��7���0;�i�"Oȕ�W�V�B3��R�L�Ln��"O������Ul(T�A��	w����e"O*��f�̄�4xQ�ؖT`�H�"O�m˄ᗡ_V"d+�4<J��"O�ڐ��*�8 s��]4^U��"O`%k�K!i�*�;�-�7F~t��"O(`��iĢ9��Q�̄�]��sd"O, C��_	^��l��(����#"O^�;T��l"�C	A�*�P�[�"O,p����1Z�r�g'�6R�X1�"O���:kY�鑦��z���"O
���ۗ�,��C�֙f��|J�"O)A�(�9u>K��x�܉p�"O�t"o�	�:"䔘w���p�"O�(��kW�71�]�G)�$ut�,�C"O|��KS�EyR��%'1kd q"O��S�%��b8���u�]'%U�]�ȓuu��$cg۞%�a�_�bM�T�ȓ[*^\r҅�>2�4�cI:aJXx�ȓ<�0�#jNK�1 �,p�1�ȓv.5���QۡΘ~�R���N=D�Ċ�jƪ $P�⍙�0I�F1D�H��ߩmF����X&Mm(�s�9D����QU5�������,z�M�19D��ࠟ�>@�AQ!V$_���!E2D� 2���9:�����G�G��q@:D��Kü�B�S�)խz=:����7D�t�� 
J����GR�V�XQ��6D����#M	4�IA!�U9!e�U�2D�p�!��RUl!KR��:uݚ��7�/D����@@��m9���g2$��.D�����.���a�D�0����֩:D���!�Eu6�zG��7�ؑf:D���e�	#���2��k����8D��#P�B)R�6�� �G�7`��K�,D�p� ��'@q�D.V���b�)D����iJ�Y��4���Rɶ���2D�11c
,Y�.uٲ�_�)���Yc�0D�0qu�����F"�Z����i,D��w��Q�r�w�E�Ĺ��,D�88�1��,�נQ�|~�t�я*D��&����l{��'Q%xL#�c5D��@�EO!l�0e��ʜZ2�*ѣ%D�4!�k�~K4=r�F�C-j@@�I1D����v�JV�%'�z���#xx!�d�dN�����Np�y
��Q�s!�Q����J#��1f ���'�][!򄔊Lu\��C��h}x��MnQ!���58>���Rm��
ti;�%�I!��IS���g��V���xF��98�!�S4P�̠fM�f������5Yf!�� ��Ia�K{�lUSĠ2,��P�"O(a����.��̣B�S�@���"O�Ip�ą]�����ˍ-�X�r�"O��R�.����<i�LA'��y�"O�QXK��I��!����4����"O�=(e#Ѣlo�5�С����<�
�'�r��A�՚6��rW#(mll2�'c��2��ɧ!r�T��꟣��U��'�Z�oU%9I�)!/H�Dd(i�'�=�ŮH���!i�a�4z�B�'�0-9"eN!JĶaʗ!�Yč�
�'���5�D�U_V�P��Q��,h�
�'���s��ւAnh��F���1
�'l�3�e���\DJv�C�qܘ�	�'u�8P� ƀ0YՂ�|�] 	�'dt�8,�~Q8�3���_P:���'����Y�.�����V ^�f}�	�'b4���=ޔ�e�يI�2���'��!i�D���ɑ�摑60­c�'}؍*5MS�`���[�+P#.���'���X���^ʖ,j#�ٍ�fh8�'��M��dYB
����xB�$z�'�`Y��愳I&��7�2Z�h���65����*\b�קc�֕��c7:r@λ%�*U`�#@Z��ȓf����W���$�a���6g*��ȓR��\���F�4�,k�JG3$k੅ȓfm4�����!��j#��0x&6��ȓd��� ��U6��5$JI`����w�R#�CL�*k.D��m�Ć�
�������V]�Ghĳm����m�{e�U	V�����F��(/Ѕ��(�>E�b�ƺ-� �Zԥ3	����ް3�i�:w~�H�5e�r�D5�ȓv��H����l`���_i���ȓ���12M�HP<I�	r0͆ȓG8]���-u$��n�1�����
i��Ǔ/�Z�0��	�^�A�ȓ^�B4yw�G ,P�p$B�4�1��q� ����)x,Byh�cS:����Q ���2@A�����5.B%��\��sRʐ;�@�\�B0���P�"��$��:���茟L�:����m5��ȓ �9�&U�6՜�SR�7�`��3&�Ac
ò�zt��נ
�D��L�JM� �؞�t0��
n4�Єȓ;�Խ1P�ϧ.�V9pj kp��ȓI2�Ct��($��[eM�&�H��ȓ_ �8���G��Hk���]�m��L�P��K�E�BAK­�mN�H�ȓo�J�&�ƾ{�XЀ�26��7;�Q0�G�e��1 4+Ӛ��ȓB��\�я�'Әd��_��I�ȓ*��4�cB�h����*ݒcs^i��#�h�Rf%b+8U��K�
t���ȓTvȝ����6����s��
J $��ȓ4l>1�ֱ���q v�A
�'�����P&.T��$M�w��S	�'����#,��z|;2���0���'n� R@��/P��N
:��'a�3���b

1{iy�}A�'+��P�J
\����I�v> ��'GH�x�l	�M$���P�V����yR �+'�dԸ"+NH^�����y
� �ܫ���Sj8�˴�^5#�<d�$"OΝR&f�t�����Gv�0)A$"Oʀ3�Ȁ�j���AK��Ҭ��"O4�QՎR'
�H cp���&�n�`"OLa`&�=S�܈�C�]��|���"Od��GBʅ �-���w�v�b"OPEpE�>N,pڴ�ԑ!�$%�E"O(t��� �c��Ǎ;T�P��"O��3�G��
A�1��t�:�Pq"O�MQ�&�_��M�Άe� y"O�X�"�C�]p�Q����v��"O����"���N�t�دC�>8e"O����߰gTU�!-�="�"O�5)�.�2�r�l_�^�T��"O0��̙+J�x�%M�.^DyR"O*|�B�(c�(�:���=�Pc"O`8�b'X!e�Dy􈜋N:���"O����J�?�f��ħ�-�j��"O��+�	ޑE��A#6�a�*�2c"Otj"	K�F�����P�B]��"O��ˇ�_f�d�Gkc��|`�"Ot9��AݰJ����	
F� ��"Ol� ǁ�!
;Ψh@���ҝ�E"O�����'��ܸ��_�z)b�"O��P�G��L�HQ�9��*2"OکhcO:$�ĘP����7�r��C"O�}���J�wY�(U�0��E��"OrQ����	�'��r��z�"O k�ŗ;^ �����|�D�""O��&���\�NF�7�ƤRq"O�=x4��%����5���;�"O��0D�_�k�ޥi��8�"O�1��ǵ�a:���)�(s"O�M`2���g-�x��+�6��${�"O h��� {�X�p%�ȴ"�� ��"O���U씷:�ڑ�'@	���D+�"Oȵr5��91��P��Hxf���"O�gjÎ[\x�kR2Jh&U��"OÉ��k�RQ��X[X0��p"O|�!$2�LxWM��3`����"O�	`E�;I���M�,baj�˅"O*�2���5e���>M �x�"O=�g�%S1ȩ8ŧAF/�y�m��~�e+�.�	%(haR���y�+�B x�"�4
8vi�!D��yb��Ը��bN�=�=�PD��yr"ֱg��l�t�21�)��Ľ�y)�l�@%��%=�I�'�L�y�eڔ$i W��8y�6ĕ�y2*�8���/�9&A� ��W%�yrBĔ)�L!r�#��p|�ȓ��I-�y��%`]nTk%� T� :NN��y��ay�|Q����RM�lc�����y�C�虓��GHIК�	�y"a��I�������DP�ͻEo���y"͒.Z��sɖ�'B>��t�!�yB+��m�Nݩ�Z�S�X(������y��TPs����`�q�� ��y2/H�j��}�G'��W�V�1(O�y��	&���` �K� N�l�r��y���Z� i�O�%0���R����y�c@m`~��f��0_����y�EX�+ޘتqAY�g�����^��yr��:��e*����.�O��y
� �$�#D9?.�}r�F��(H"OF�r5���Fjjթ�EB�$ꐜ�"OJI��͈�� 9�&�[�xGx�P"O��y��ƨ�x����	4qP"O���&m�$Y P�K:��j"OHa8c��8/���ږ{�8I�3"O���#�z��a�ߊNe�U"OU�P�>�萛0)+~���#"O���$%�2t��")Ya��aV"O=1���`����f�$�n��"O���@��������K� ��q� "O
A��fA9&���1�'i�1`1"Ov}�T��.7-�Ċ3h�>`Rb"O��B��6x��߂|����f"O�l�:-��pc��a���"Oj��@,܈`�ly�K:�¡9�"OH��'`�(L((�Ij����#t"O����	X�;正��׆;�<�#"OD]�wn�V,�q�hM�R� �ؒ"Ov�1���4Xѐ�{vH�O{j���"O�P���E�L��C�Ǔ&
�i�"O�Kb��8��iv�E�a�Z�c"O@iR�fߕ2�
= v�	�X�"O*��5�Ӿy��;���$X(J�"O���v,b�,5a��׊N�2�"O$�#Ø��)�T�GZj�ڇ"O�Z��Ӕ)T|Lä���1LP���"O�Q��=�b̀ƨL�<�D"Oh|;���xV,�0"�1��8D"O2�H��L�u���b���	�:�"OR�q$�>~1�FL�
CHe�d"O�uؤB�	* =��kGd>���t"OP]�4�c�@�c
��n����"O�(�䇤 �L�jDj��gcf=2"ObQ��S�B�B�/��U�.�	�"O�h2�%4�쫖$�7k8^�S�"Oֱ�G�=z��!�GA�?��-*"O��$N
D���ӆ_y�d�"Oy#���:I�@G�?mQ*�"O �谡V�T��CfA�;�8�y�"O�8IUe�{:ݳ�%�(A��3�"O )�Џ��I�6 9s��J�}[�"O��YW�Y�	fe���?R�ò"OvY��]�lP�xথģb�x5��"OZ\�PD�+/�+D�!#���e(�)�yBBO�Q�B*g3=|��գ���y"�I�a ��IG>8�^�%AY��yRY��9U��6;���JN�y�퉙IY����D �5��}��C��y�g�vd ��c�9'�00#��%�y�$�7=�EA�%�"��I�!k��y�l��ifȤ�FF�������yҬ�(/���C'
D�@ �E
���yR.ĥU `\��H?�>U$[�y�? ,CcL�7�h�4�yO�*Hf ��#�2O�����yb�W�@��(؜��T��/X �yrK�5�ʝ3���҅Nɛ�y��m9t՘6N��3,m8"�D��yR��1c>3�$��\z����y�,L#&�n�;'�ہ**�Ȼ�6�yb�<���$�R}�Ī���y"�Y/�d�!���DUFxk� @�y"Uc>�AC$ϑ+?~8�[��W��y
� ���͓�L=� ��׶0�M��"O6	·���
�T�ǥI9nB8Y�A"O����E r��e��ԕO-�)�"O�dI�+�3
q�#��<-�l�"O������#n�uY��U;1*ajp"O$hB�8�]� Z<!za��"O0)�a][��b��4T��iE"O:�x�Ɛ�~R�0V��?[�|1�"O*�����5n��G���8�"O8��G�n�n9C�F�r��*O�́�d��@8�EƄ�C|ܱj	�'H�r��� �K ��I��| �'�����T%ST���b��A��
�'�&��e�Qڣ��:E:,�y�'�QB���
7�� F@�/&��|K�'p���.��*h|!�j��,UF9��'a�R!�ăX@�r@o�?"����'�����&%�.���Ϗ��$��'��u��ǀ�t⚸zW��3JL�i�'4�1��U�O�p�,�=GpM��'��(F�.KպpG$��_T�X�'��Փ��O�/��b&B�
��x;�O����G�	�q{�P�R�Ĩ�r�R0�����=�'��S�O��|a���Y�y1�B�J�2�'
 �E�7b'��H���$38��1M>Y�'{2��>��E�j괍)1l�6PY��	4D���uȆ22��M��I�Y�ވI�I2�Il؞��R,���X��Q'`���K%�=D�0�!d@2E����SI� y�l�ʃG}� B�I�(���y���/K�����SxX����%*�OPy��M3=���CU�M����1|O�\���
A-�@Aŏ�b���`"ON)�&`�,����ǒ�o���w"OL����'������b�2s"O��0g@�
��@�&0H���+4��Y?	��IW�,:ҡؕ�88�jp��!�D��5Y�A�1�ܓD��$��揍y�!�d%B��Eh<8�|p@��(!�$8uڀ{�H	1e��U���~#�Ik����l�|�P�؆�H�R�  .D��AT��q{�e!eˑ�:\���6D���f)���	�v��'�]��C4D�iժ��`铷�:lL�!���0D� �vD��Sh�m���K�4�����/D�H٥@ �Y�piҰ�H��j�ʰ-1D����w�����T n1NHGM1D��X����i��MC�$��Pk&1D���A��,�
xaR�i��.D�����_ú��E9FѪ(���&D�,S���VlX�QK�lh���D�2D�x�  ��P�8�!t%AO�����.D�RV��v,Vex֣GC p��*D�`�u.ضC4�����I	��E:�)*D�\XQl�4ؤ�@u�S���RS,*D�t��G�]�y8���j"u;�+(D�La��\�@�P��͖T�lAB�%��hO��&I#,YC5섇2/��
���"O¥(��׫Z+���O����kf�'�ў"~��o��j8��yh��G�vdC�b���yb�T�6��I���
�L3jAIf�Q����2�O��%ԱSĴ�SBIϐ�� sW"O��F��1�T\3�h�/*���ˀ"O�A"�_�ZI�l��ܭl.��*��']��3��>P"jqB���?�81��)���C�)� b�n�2�"I:k��wvi �"O�1�C�ٯ70u�6�_�U}���"O�Q�T��]����K�v�B�K��O�����
6$(Q���;Ru��	b��wDa}RL6?ɂ�P�l���J3��A3��I�<i�D�;������� ��w�B�'����Mc����ɉ6�vܻ4bע c��(�m?�y�����e�sh�
����Bs �<�}�Ƶ�@�	���fB��AަM�v>�G�	g���s*�j���%��m��p=	�bƆA���@C�Z��[C�[�<Y$H$7��h� �_
C��O���hOޣ?Ѡls1�O�e�<��"�xX�$Dy"�_s�N�`�ڃJtX�Sm��yr\)#4�1����#�ԉ〈��>1N���F�Ӓ)����c�@�
�`�; �9D��S'��Cw����]&z>E2��7ғ�hO��#%�LiY�0^UZX)�JS6�,C�	�{�T��1���k�H�ZjĎe��B䉦Ј�)��S�>��%xs�L��B�	)�*Y	6 �"w@��c�K?!�܁���s�A�SՂX� h��Q��Z��)�����(�H_�;�T�h�*+�B���"O����G8yV��9�Z�T��lX�R�H���|�ɾ ZN!I7�K�CN�l����144B�	�%�0�=d[t�%�����S���Y������6sݼ����"򓥨��M�c*�6)�����S�ʛC�,D�
��D6mP� G��|�~!"�h��F{��))/,�0���o`X�b��?dT!�d��F�t�iŭ��I�2�!��G�}{�
!-�Gg��WB�fk!�L�a�X�e��i����2"�g�qOT�=%?9�D�+�~�� �P�'^@ Cc�/D��e
�>$�NЂD�L�^"\i�
-D�Tc���*qRxS��'K�`1�H5D��+7c�
��Q��"H|g�I��`8D������cF�U�!.��!�+D����hݥ��L�|T¬��(D�pB�OL��B�r�mJ�[?�,!bh"D��Ir�`E^����QJ� AwL5D�xI��c �h�e�&1�b�Rt����q�)ڧj�V� �쒓R��s�V�CR"����hO�>Ea�+V0P6�T���ߜo�T���1?���,�j�a�@�f��cCX �"Յ�	}}�� ��z�`��l�&%K����y�&V!����-D�l���ibC1�ēM�Li���0<�dLB�J��B���3/�� j�\x�$��MC�E�b5ġ�I�b��q-OX�<1�V�"�Xe:��%ȋW�~�b��hO���>A�Ā�"Rp�#����!*䝰ǄFn�<9�`�� �ґI�}А�
���g�'>���O�ޝy���?0¼�"ӕH<:H8�'7���ł>Z!�7�K�jTqp㶟ܤO��<�O�+ ���j������D~�<���QSV�XD��.\V���z}��'��X2�޾���3�O�!�����'u��x��F��q�a��A��'��	ڗ#�]w��+t`�9���H��Ms.O�a*�o��eE�S�EZ`�+"O��H���L����w_.�b��f�O�����V@���%��
'�����Ol�8�)�2��e(���v5�t�S"O�C�I�$o�����F4/��+&"O� � h'C�q��U�a ��ؤ"O͂�ُ,$I��J�7E�� V"O�uKV�9 �e	c�W[&���"O��õ/ɘ��`���h����E���)U7!�T	��]2R*��� �-O7az���	^��Q�*�hU�0��n�-�!�ě�B+�uc� ]!=`Td��6�!�X�z�鷅��"zօ����h!�ޙM����U�7QqB|��FS�=X!�X<��M�5�C&d�l[`��tH!��Ҽ��Վ��@�ڤ#Sj	�!0!�d3-�8�CB�N�:uc�
�6�!�D� JN�ůǦ
���C`'t!���}
����(mJ�� �e]!�
�^|��J#C9j!g I��!�։��ThH��D�����!��ƃ���Qr���h�y��+��!!�12���&�2���Q0��+A�!�C�K��;�皸�"���-F!��UW��s����j�P���ˎ�,�!��4v�´!T�)\����
^�Bx!�Ȕ�=�7	�7,V)fL؎e!���@z�^J�}c&��"�!򄚍|V��Xf�T}��R��c!���4n�PCp�Z8I�\�2R!��]&j��1'J���=x�U�z�!�$3#���SBɘ ;�9�K-U:!��
*6�A�B�ݞQ��	�R,BB!�K�|�o&-\�1�MB�T&!��J�"]�SL�:?�����!��Ǻ��pXa�
&kx��4j��}`!�d�@��q�Ū]�6���GX�[!�$�~|+�\�Z:P��FO�;��U��[�rk�*�|������O�%s��ȓ#aZ�6�_7�p�;�,L&L<b��ȓ�q���� >��+A������ȓ�*�veWVk��g�A�ȓ3ːX�Û�&�٣��rT���Hq R�#l��u�>����!2:eS�M&AS�J�t͆ȓi�؉a��L�d1��6oW�a�ƙ�ȓX��ؒ���D(�;�P����ȓ�r��֭��{����P�<�d��ȓN%$���%�.`��L�O���ȓ 7�%x!�N�T���P���x�~]�ȓh�| (O&�⸒�n�K�x��
��������7Í!I�z!��>������V	�A�o� m#���ȓb�ҵ9djJ"
WԱ���0"O�QA�N�-	DT��$�� A�"O`i�w!ֽE.H�ѵ�n���"O��0�Ə�s;�E&���+��B�"O�8�%ζ��9b��$X�TI��"Op���
ܪJTh��B)�#u�&9�G"OHHʳH��6�]�F-|�`C�"O�aN�K��Ȳ�B9e�t��"O���p�+LY<�����b"O�m)���]Rҝ[��:8���#�"O��u^7R�*��7��	�� �&"O�i�dɈf���i��.7o9��"O�IZ��=�eB���9_U���"O����Wp�p���@m&�qr"O��;u
��3ڐ����gt��"OX����&/D�a�n�L � "O� �A�s�L|!���-hС8G"O@�)F���d1�TA��*#�V�`�"OJ �c�җi�;�T���=�"Ov�8�mڃf��YƇ�T�0�;r"O>0��řW`H8;ӦH=v�	"O����6�j�Q�ϥ\�J-�4"OTQ8��KeLҡ2္5�����"O00%g[<�̨�qbD2��E{�"O�Тf��1�n-��Տ$u8<	`"O��FÝ�&�6y[���	sea�@"OFA%�6n~i�c`Q�Ga:Pk�"O�+d�[�Jo�0� �/	 ��6"O���-�>�.�e��~�4���"O��F�3%\l��AM^+���"On��'֊4�DTk	n5����"O�����E�?���6�ù�h1�"OV�Hd�A?'��K'ě� �t�ڗ"O�p�_�)�|�!��Q�_J<��"O
-{Qc�h68I�GC�z8h�P"O�$sC!��G��P�d���u%����"O����ߛS��<:t�z�
�"O�U3��C&9!���4s�~���"Oh��֭�*�b�Tll\At"Ob������u3�k��r�"O���)��F��MAuK�:�0�c2"OX�X�E�����
&T��q�3"O~�K��0�4�7
�&u�n�"��Ic�OV�рD�]�hB�֙CjX�9�'�*�J��ב>�l#�a�A�H`�J<��4�O����6�*:^�I��W�.h�,�7"O�4�ۃ.p���@�S�|]��"O������L�^�d�./	*F"OZ�9#�()���5��;$����"O�|�F��'|(�P τ�P�R�q�"OT���'����"Wi�@�J0"O؀�S�Hi~�TR��j���"Oj5B``��d�^��TG[�~�h"O � ��U�4ż] &�R�� �"O�`���U�+خ�3�d��h��@"O5 �"	�`N�\�#�������"O�@�G���j��٧��=���)�S�7�B�`� ���T���B�	>=~��1�)���ch�<7iB�'Qў�?w&3%�(+$m��-aK���!�DB>f���1Y��y����>_�!�D�S3�ۥ$�F�rD���^	Hў����=N�HZR���z�p�y�N�!3LC�I;=�}Q!C� h��LX,C�ɱx`�q�Q�T=`)`bd
�	�,C�	�7�pajF�'�,��� �dk�C�I�N�zH:�E�N�RŁ�ĻT�nC�7�X5�DEЇ]*���"�;7>C� '�XaP��P"u��J_�_C`C�ɞ+Y�X��'ы (
7ƌ>@�0dFxb3,O���#�JP���keG3D��"O� A�'*)<�b獜{�yaG` �PxR*؏A��й5"<YA�mH�# �y�d�?�$��g�#Vrb�HY�yB`�=�ޝ��ϸ9��H[1ϖ��y¥�.�¹3ӣ��+�؍�d�y�)��̍� f	7 MH�j�fH��y���2Ve��q$B��,0'J��yR����"�� �H�ԏ�.�y�!^�̄��UT�Q�`�ԍ��y
� ~���4�(��!��r7RA�0"OL1)`��W �tZP��(���A2"O���0hNh�X`�a(�9}��-�#"Oą�6�_�31=0�f0�6]hs�'}ў"~P�6H�Z&@ �_H�B����'�ў��xi�B��>�NY;�bD9s��Z�"O�,���	4 ���7K����T�ɥ�p<Q'��	�d��hR�tI�&]L�<a� U��X���R)zx��mV̦i���i0�"Z�=��[���L��|��yڇN��i��Pe�(�pP��'tP"�@_Fe`��pê,�d���Y(ԃ�6uqTuS6ŗ'Cn�̄ȓ%i��)u�N\Ơ5����"?9Dyr�|z���CqZ� `$NxT�L�C�<Y�.�?�"���	�P4&YJ$��B�<)S�׊l�8K���%`���'��<I@��0���*B%ٚ�d,P�(�D?���S�_�$�� @G^�����TT��B�ɨ$���3�Iv<&�¬���B�I�S<Y���v(���OL�>�B�Q��icg$��^D�s�닞|l�B�I�\)ʀ� +��!�����:6B�4��8�+ˎ���G�U5 B�ɮ��1�fb�1[����똞T��C�fD��$$�� 朔�4�U>ڊC��7[���$b �w�ĉ��
U�B�ɒ>vY���"���Z���C��B�ɷ�0�S�
f`AQ�ǚ�l��j�|k�K� `�� x�`1D�0G�َj����Ϩ_��g�0w����A\Ȩ��u��@�T쓴5&���ȓ^'���VA �i�NU�V.N6Z�Ё��)��<Ib�3�rk�ҭe���Sw�H\�<���T+G��5#P�Ţc1zT��&\X�|�OHUx%i�*5̮-ˀ�P�/�x"OD��"��ux�0j�O�0�h�"O�(�P�Z@g�|�b��V���A"O�Æj����q�#�N�\��"O.���l��[e�׶X�: "O�9H�e��bF�l��Oi�X�@�"O�����	�)�t<Bg��$����"O\�r�e Z&��cF�o�TXI�"O.@y�E�"*��\9R�;+�P���"O
�+t��?��-�vgl�b���"OV`��b�0ub�1���- �� P"O"�Aa�
v	��͗B�2�pF"O�iP�c�uF
�X���H�T���"O������;��CΛ k����"OB{�̅�w�,�IУ�GAV�ʔ"O`�RG�M�лB@K����\������=�v�X�;} @7�]�1�	;R� u�<�0&�n���I�HN;/��a�f��z�<qW*�:T��)�V�8B�P�0DN_�<I ٰ}��0�u���W����[�<yr��Ez����+T��I�kOV�ӂ+ItX�����	�d^�p�iT�l����l6�d�ٴ2�H@�	�>:@@")�Ac����B�Z����H0/ �)z�Cاs�Y��K����G+ex@��#�_�F���&�X����G+��|YB�P��Y��c�P̑rF0]]�c�`�oJ����?9٤?�p D#�#���@g��y���B�f�p _%�����E��y
� ]9�%H7@�����&W�d<����8�S�ӷJ��ȶ䃵\Q� "�,X�6C�	�Q�Da#��P�G�򀛠���+ C�"�2��L��1<$�Do�8F�FB�!x�\p$ V�v�❊�$Ԝe�TC�kb^HqfaC�&��RQ�,-��C�I,d�
'�W�<P���G?
�C�	�;�8,�5�Y�]��,�Īي��C�$G��+uD>L��T��>u�C䉜n�!�ĭP�[v�(��nԲC䉷�j��A�[;�D|�B��<lLC�Ʌ�\H9�#G�1��h��EƦ?c�C�	4 `�	�l�3]��iӫ��/��C�	<I�Ĕ�f��l8�5��Cx!�C�I:ssF�UBޭZX��c����B��H�K��"p��+�-l�C�ɶn�P�j(� �0)sV�q�C�Ix�΍#Q��~36L@��	�t��B�;f���ǯ
PEf`#2�3U��B��=p�Ԣq�Y�F�F���nG�B�(��]Q��#�Z���g]#XjB�?hy#'��i|���]�C�I tO$ �O�01�>��
�:��C�I%G"�B�U�P�2�
�cˡ )�C�m{�i��ɂT��s�	0y-��$��aΑXd#� ^�:A{ÃԳ	 !�d�mR��f>j���샬T_!�DV���|ʀ�Ɛ.��i)E&Y/
�!�DF��D��p�L3Vzp5�#%�0�!��,�`�"����F��s�[�Oa!򄑩-��*p@�<&-��3g-�!�D�:=aܩsU�]�ZPl �G��8!�D<ni�HB��e�;�'�86�!�¡$�Q����`Pj��!�$U�A!��H5`]O�,�*C�A�`~!�W�t�����#O馼��]%/{!��_�(A�]��,B�,\5�ӪBj�!���
I�ɨ@d�S���pC��$�!�d����@�V8�(c�K�r�!��ʸ:�6�S�W%|���f�U!���}S#)RL�i�k_�Wg!��I�F�0��·,$RT�&��(K!���#Sx�:�H^�3+!�
5Z.�4�C!�T_t�9�×x$!�0\8h�`��*_8���wz!�� uVH��PFօa�0,0#��*:�!�D�����Pv��fQy�R�_v!��0���ju,95��\�p�Z9l�!���NAƹ�gB����� ��ɖe~�N69���*��@X'�	�p�Rt�?Q�D#�� ��]���a��L_�<�Q�K��H����,<��l�DX�<1v.�)_(l��ȝ)\�Z,I���O�<a��g�BPp ��>��y�!#_b�<Ѷfíf�
�X���vZ`A3͓b�<��-ќy)\���
�n��(]^�<�Bi�&~[�l�������+�`�Z�<1̃8�x�D�p�3��R�<��B@}jd���������)�w�<���R�6d��+�FMXn��玓z�<���)&�0��I�p�HJ�Fz�<iF)�;p��u��{�b�aeNS�<	�+˗���Jt#�<�Vq&o�q�<��&x�y���LbR%Ph�<�R$	�n��V�R�\�,51� �o�<� �Ur�)X�@@�}"���+5�x��"O��S*�|q�
/1����"O����ꇟ��:�L=:<%��"O�Q��m�:�����k��9ȅ��"O(HxF��c� �ǉƬ:� ( "OFݨa(ڔ&�q:��ݭ;�\��"O�@+�%Ʃض�L�l��	�4"O�����G�m B��f�'��*b"O��E�$?:�<
�FD�o��E�b"Od�R��e�)KƬ��kG"Ob�`c9(�MpfM�	`���f"Ox$Zg�[6�t���
� �&��S"O�u#@�C�qg
�a�P�.'�8��"O�}��e�X�6�2�����	�"O���ShB?]���H�@�},��G"O�1 )��3�a��
5oܠVS�<!�Md��-ӓ�����i��DJ�<��O)V��\)T	�`��ԋ��F�<���T
1B�$�TCP1J���1�oVK�	�J���9�����!n�8%�G�$-j%@�a!�d\
;�Ͳ�D�7.D���R�w����>�@m�%)��>�OL�ʰ�ނ"�N1����0,X�|C�ON�����,B�4�c�K�o�.m�-��\6$�
�0T�����6F�Qa��m���k��
џT��ŨlӸ%��.E�z�������	ū�>��K�B9C䉯L���9���3�Vl��FV�Gl<˓f�Lb1��]����k3�'m:��iU���A���,�ȓe�~��1ǠJr��W��ZS>�	�r�d�~PV(镥N�3�ɴV�����-\KT`��ʋ1AV��
k����n�/��=(Bo�B���;ӈW��Ԃ_ �����ܿN��(�V%N54���S'L�5��|BԧQ�/z��Q䜸b����FC���6Z��i��gO�o��	"OH,�-V;I�5�&��(-���^��Q�M4!\U���Yu!�'l��x
.*����'&�����]8x|�타@V�P6Ʉ�s��J�#Q�r��F��Lʐ�h��� 6>��\�j�2�4,�q��Z�O��Y�֩ȤcEN��R�@��"�j�>H2�d	.+� ���܄0����	�CxRI����(~eb�XU	��I��tZt�����d�W�<0��OȦFqBQ����S�*����D�Cd��G���P1��/�4j� 
94�8n�+ L��2�\2D�Y�&�H�s��D�+t�9{ \k�8(�@�zS1�Ś ���sQ/��O�ȗ'i�C�D�,.ihbo𦭀���Ewԝ���%
C�2��G��yX�������C&C+tE�C�	�ny�P��i�=�`�H��;����֧�%�M���-@�����9��ؙ����?���[�t+�ϻ�. �$��� ���� %���(0k����Ck�pD�B�a��`�ǎ����{4&D�&L
�K��rv�|B��>Ao�x�g̓4��ē1��C���`���R�̅㉼k!
i+��W'�dM�)�@U��U4e��\4+�<	s'��9gNy+��;l��]a��'˸�x� ظ�D���[�:�8�����O~�k��U��o>) VN��"bU��϶I5�0Ӧ�MkԢ�s@A�d�N�!�)��@������jЪ]أ(�:K'Tuj��D8�Ą?����D�c��,R��E�i^^p�S�[�I Q>i��/���1���T�+��!�N0��I��ʀ�eQ)��'/9 m��$��AC�Ѻv��5�ņ�3�n��%0V�S���Ϙ'k��f^�:���OL
afP���^� n��3�	0�ʸ(f��4{h�#}J�]K�`��0d3&�P�Tgűd��t�W�	N<��@'Ls^��ɖ^��t���&36���\�\�|H��+ʆ���fA�RzP�����|��S)Jj XrgĹ�����K��P�bq+���=/�4@ٷAӌ3����|8� S��T�t]��ہS��Ż�j�80�r�s��-Ŭ1`5蝽y���;s�#?.*����U��ݓ�J+��$�H$�wa�#z�u���[�d�c� �V(�~ɀ�k��z�ܙe�m�v���#��-��m�yhx�0���Ub�3n�詹��w�b��6@1���>in<cH�m(!��\>RX�����G�#���a&�x.��K��=mjb?iaó�j0��&J�r&\�@��Z4QZ�#V�,~j�,�	7��Y3�'Y2Hq��ܬ!2%�P$G���e%gm��т!
�
u
�-�*^[4XA��...��/P�B�����'9VT�eNԣV��a��oE&vN��aϓW��y�/��sC��f���^b%CFd��W�����h��Z�������bH�A�*�|�� ���)[|#�Oq����/c�S7圧/&E�J<9��J�LL`�$�HR\ -�4���%* A�g�? .L��T"���ak����"Ox���k<l�"4�:���W�V�F���c��D����S��Ip�L~��.�|O���<��[$�67���2l;d�!�d�Mm:ur���h�Ѐ��NS�J���F��p6<��A�}$�h���Nj(Y�	:v���pdȆ�3_
0��^�8��R`�8b��[�=��AWNҵ�|�0� d�E`������ĈB?:�8(Q4�O�x��Y"{��i!�Ot!��x��ވ%���J��ڕI�����>*�xҩ/���y�����	:��Y�ʘq�<�A�|^���Ŷ=V�j�^1[6`!��-�Pt�3�E)�9�~Jj���~)
j�|E)��a����[
ِx���Z��ר��(�Z<!�b������e*��y�T����-^ihP+Z�'�N���ϥ�j9 0�.;��` ˓J%t�:����[yl)���\�|Xbz,L�m�V�"�	�c� g�!�D�%{dL��E݅z�Ȉ��Ƒ=[�'�k�\.0����PES?:(�˒�"�`22�!K�
Drm���_-tE�C�ə^9ȁ�f'K�����rc[,k����Ecݛj}�jA�	*6�ъ�.�3�Dݐ&�~� �K��ZK�}���\�R`!���F �7�֭ ��1��m@f`�	W�yp�r������F$&,Obl3R��v�(YF��f����'��qi"�Y��&���d�iA�I��J�N�؀��W�C����M����xdZ�ZJ�PvB�5D��0��A�ēj�nA)�M�!�p���F �~���E�P���Y��޵Wf�P� �ZG�<I��N99б��gQ0HX��B]2W�[`�\�vs�ą	x&�9�~&�D{ �6@�x�)�z�6����<$���7�ۍrp�(av��J���q��au��p��J�ah���L�^���  ��-Z��J�D�h�BP!Y�ay��M���@u@�1M,�Sp ݮv�8d�����M�4&^� |�z�'��X�@n�2���L�t1ȁKH<B-Y��x�{g���L��[3�~�'y������0$l���F4܁��(�B�
7+\&!�x�2�%��b��X�ҍ.w��UJ�o�(AY)��Ow�g�	�W��DS�� W^yB�B� �tC�+?.\s�&;z�W�# %TY%�7RU\U�AV�z]%:@"ŐT$x+�O���hQ+�0t�D����� t` ��2)jJ��DW14
!�p� b_°B��	y��� X�PԸ���K>^e�'/K:�Y�'{���1`U�x����!ې��F�0(h	�-�6��%&����52��jbmX�lct�����$�,ч���k��5��֬�
��#bN~��Q�fI2h��D8�`�,�=o �SSBȴT���+���Cƶ��V�Q����
���k�H�5x�N(z�F�h�|���0W"�����)N�X +C�N�B䉺6_x�I��{��$�uN?<�,�K�e�!2�,���2Z�
ě��C80Qx�1#J#|����>��I�&d�l�h1Nƽ�R.]9azc� �4u��(FҳaeR{���<�/;ۚ�*��M5��#���	�����-6��H��?�r�[Zn�#jq���䎗��>H�cX�	'&b�@�p�3*8��g��J�t	ȟJ\@4O1+j������]���KN� 5��RJ�[�4%��97f�\:2cP/-g�����9h^�qJX	dB��ʧ�R�
b ��sF����P�4P��I�;6l�	C*T�Tk���k�neH�a@�5��AbOJ2-�F���gXR��c#�޴�p?���=n��5)�M��+#0�qBˆ�`)�ģ��w���RҚ"�r�pFb
�n��=	׭*-.8�Qb[?5�w�]�)��}1�߉TU�E��&LO��*�D(.�85;���=�d�q%�90'y�@M�l��c�'ǝ`^\�[��ѕ�~aЦ萺rwh��O\4@�5� @��ѱ��UZ@T�ۃj�v��*7�h��<�]6�z�!�ET�A\�%��Y?��Í�.�L	P(��h�ڬ��T�@�\؛������vK	|�TQbkľ/��aQ��Z�HO���'.|�n{hY�I�C Ot�ܺ���2��-��a_;���'��y�x$���N���	"Lp�ȓJL�
(A�h[�0�dT�"C9��9�(@��=�
ؕC�t���ꘫkk�Iz �΋-+�ED*��?�����&������Bb��G�x��Ӫ�jj���:)���'	4�`�Aׂ1 �A��O%D1���.l`3�O=�
��G/�2�cr�#:+Zp���A��Ac!�º!���C�D:&��dI^��<�k�O)Rhٓ�O?F��}�ic�![S`̊-�Ɯ��j������.�$�h<bI{�B�bd�!�T�1P�S)���9Z�����@.t2�'S7Ll��s U�/��b4@�4s,I�4�ϒ>@��R*-�����T���۔�|�A�c�'kLp=[�F.g�>�+�Fȥ9}P\�F�ײTb�2f��=ug�`�#��:�ㄮC�`A���b�ՁHi���ER�I�$ Q��I-�a{i\�@�ɚA�4mA�)��
,:�d|1�Q/]`P�6���/��ʳ��D� ���M�"��,8�`�ӤN��tI� �x��h�	2�x��A74� *�ǐ0i���D	٘�lʐ��=$T8:�T5+��	@�n#
DB���b��4L����dΧ< X$r�#�����A��5֢S�K�E�WG	�(y�Ц����ēR��-��"�LXr�	3K��,�O� 1G�R:M��H�
Ҋpb���'�"hdR����U�:�@�A�)qL���D=�
�Ej�O� �@��úN��A��C	G�%�U�P�p�,��dAJ[:�x��#Z�h��B8K��a�C��eAP�r�5p4�	�'����b��,�S���Aހp �+I�n.�{���4Df��2���r6\0��Y;,�x\sd�V)-"
�Y��U�����n4C~���"��t.h@eh�-��)֢(lB��0"צM$`AGG۫W�az�ӧ�����-U�U�IqS�V�h�
}�f��	h�!��Ȕ?MSd���jiȸ�p���-�P��4�*�����7�Hy*�;2���lr� ��%�&�	^ܓU��D>C��-��9$?=�3�J!PJ0Bt���z�
&-�\���#E7^	�Ь�(t���Y�"�<VF$b4�@�'&8qk�ovx��!�������C��˛�<b����z�t|��9�ʅ�����B���X\�MT	,�~!���	E<�cNE48�H��©7�OХk�o;S� "�\�G�Ɲ����8HL�1����:w�ޡ5j�#fƕa/�|zM����9�.�sbI�ҋ�m�<�1�H�jE��,�6Z브z �A}�fO�a#��J�%T o
��i��N��Lc�䔻Jm��� �Ҏ<�!�Dƫ4�&�@�N�tXnd3*۽�!�$�#(�6���YSK~=IF���{!�Ę'SG�Q{��6@X)C�`�xX!�d�'�"�ҁ�ў ,�yuo�=0B!򄄄%szS�l�!��Cd��|�!�d��j�҈󶢜�=p5��5�!�D��mY`�B�X�f�0�����$b��D)��U�9�L��:�y҃�"�x��Dاz��8J�׹�yB�~DzŒ���~��5�����y2�S�]�i	b&K-~�F��*���yb�3��T�&r��l9� �y".K�|��6�o�T]:0L���y"�N�0�L�ې�ߌ++h�Jpa�=�y�NQhw�q�g�SaV��)�&�y�i �OGBcW.�"o�LBa,���y��ѯ��"��g��1�� ��yR�� ����Qg��U8�`bǆߣ�y�mV�\bQ�w.�5M�b��mF��y2I@�eWR�W]�����
��y�\eԘ���X�&�r|kV�_��yb�q�1@E��:�&�y¤��)٢�[q�6.�6�!�y��?vJm��W"0��pS�/X��y��η0��ą�%ʢT�ЎO$�y2�I%�ݣ�' �w� ) ���y@;m8x��R�l(4ŀ⅖8�yR�9uA޹*�K�Y�2�N��y2֡g38@2Å�<_ih%:��'�y�#�L�VH"#F>T� p�a��yR�
x�T�Aeo��r��y�G�?��ST K�CdzC��y")\�! �tSV��`����W?�y"����\PT��et��Ӣ����y�
ӞjSPى��\Y`�Z�y�J�k�� ��%�?����j�>�yb��'��:C��)}pla�ݼ�y�a��,&nIhJ�';�XH�f��y���p�H�s�"	@pE��:C��L��
p�"m��:4�B�I/ �'�6�"m����.�fB��"��� � O��S�-��a�fB�+B��0:�Θ�)�����K�`SVB��"J�쉃�fH������A�dT�B䉷?K��p�DR	7K���hI7ELB�I�V���nP0K���Q��E�LU4B�I[nڠ0��B�)y^�`F�9��C��Y��C�(�9gR�P�c��>.C��%J�F��C$Ht�h��"�J��B䉼d����#�6Ά���Ɓ/�B�	��p��d�I���"SL��B�)� �R�GS�M��ۄ��"Ta�-��"ON�9��P�yb"�X'+��-h[�"O���w��	I�N
��9�0�"O�1X���9���)�Wq t�"O�)Ht��� �5�NQ%[X%e"O$�C�ֽ6ߚ�0�MӔO⨊�"ODx�d���vr@��K��&(h�B�"O�!�0�@�<VD����L s6�X(6"O���NN�M�o�;�(��"O��pR��|g����,�}u"O,`�Pi֫dȦ�y2���y�v��2"Ox�K��+u�-K�b�!�>�*1"O�1�/1�ͻ�Oݤ]q�d�2�'D�;�e߷_ָ��B*�G���"D��k#�Oq~�3uL��!WZlh"m-D����D�8T h�����:�0� d&D���KM%4�8P�� [��I
5�;D�4���5�qk�*�"�.]��8T����KK4���+��߈>����V"O�9`��2�R7+J�3��:�"O�$[Ë'8�|qq�eY�e���I�"O��+֦.Ty9���6J2�y �"O���`YG�D("`�B$X�U"O���P��F|����?~J\���"O*P:�KՉ3�����l��K0"OBqy��5e����*� �d"OXA���
�pf�:�b�Q!"OѺ�&�`���q��5U(���"O�y�� 
A�PW���kp�Ӓ"O�=Á����	¡Ɣil�d�A"O� r�N�Q��P0�\�<XJ���"OzEyggz�4!I6C��t/���"O��G��?-��7�ݭH�N0�0"OViZ�����ԣ�g�h�<��2"Oh���Jƶ*�0P�vf3�椑"O��R����*���d�f�P�82"OD�w(��+�䀇��8Q����0�'Yp���!(Kan`��'�l��&�O�@%	�E�St5@�'����W�Қ@@G��r
n%�M>Qw��pf5��OK`�>%k�I@4�\�#d#��+ ���A�6D�H����K��ͪ��.ਡfC�gi4��t���y"l:b?OL8s%[�x���`�?+�x�K�
O���f�3RS���U�
y�&���hZ�Pg�$E%_�\�0��'O��@#�/^�]�"H h�N���Pb'O��v��D�P���<��oE�H7����M.�I��l0'!�D	�-��EBpe���B�Y�mI���>2 �@B�/�"�ő5J�"|r�ݭ%�Zw�R+l����F�<�ƍ�8Rb�25"�k�Μ�n����E�P%:I��-�4u�|�<��
�Fe���G�p�gn�@<�V�_God��#%�j~V�(hXr#�8D懪>]���6D��̈́�	�,i��ZjB�>� foX;a�V��>1Q�^�w�
��'XoNQ  ����9���W_��#���C�h���F��H�Dز6l�J���8!�O�L(��k$BD=��L	z-�ҔN��=��Ia��|Ŏ,�'��J�R�Ë8ʧy�F��'o�2[Ŋ�[2�ؚg ֙Fz��T�W�fĻW��a��5�Ms�ԩ�gH�)�" ���#��,L�T�	v$Z )�pA��
�<������yrˏ+�b�� MMT�B��5@��D��n $�ꤤՐ+�D#D�/ҧZz�D�dE��`��E�Rꁥk�FY�YK]��a-/�|����P��`�#¡|��
���{�����J�9.�.ި��0������|��jAΑz������7= �;���1�l�!�ʳi��F�&|O�0����8c�b�k5��V
Jux��],E�=�K;�.�2���2����d�%�����Γ�W	RAn�-Dq���Ѧ��*�������A^�DQ��P W���FV��c#KJyeR�?y������vM0�/�))ݨI0��R&Kl �ׅB���4
�D�}&�����Q�<E��8F�F>irFx@���8m�
����fYr��ևń0`>����IM�5֋�Je^�aa��Z`챪'�ΗS�*(�4&� t1�UFޫ��=� ����@����Hb$��x[0B�j�.i�X8��"K���G傣#���ږ������ ��|P&("B��OFl���	 lsBiD%tdЙ���'jC2iŧqoʥ�g�5<?���������,(fU#@�|#�]?^t��m̃c`T1��13������b>9���� r�,���JɈG�j����5�dU��l�Jsبa9�-c�]&YBAQ(��2�����8!xg���s���r�T�2��B䉲h��4�%%� ���  �S�K�ӆύ�[]��c@(�.5ô��3i��O<��nx�9��o��?���a�V���	��6$���$I��/
�r�aC�-�4�)rCFS�4U�B�`(���-'<r�qE��4z#�=��)����"]�t�X�#��7,O-��-�8����� 
,= A�"i�(z�s&W�:�Bq8�*٪/�E��"׈��>aJ�&4����2��\�I�k≲g.�A��S�P�Xŀ$f�47Ě<k�b����iW^�.00��F�q DL�-#�!�Ą�:*��і�M]�\uSӋs�V��S��h�ʈ��
ն6�"�y'�	M.	p��ɦ:�����%`}:r�A����C�I�<I�M�0(�}��Q�Gw\	��ğ��L���5<,�Z4GU�~Oџ�Z���Y��01R�
 3��!<,O��Q�Ek"�I�,:Q���FO=���[���U���Q�ǈQj�Ї�}�޸�k6*�-x&-J�>8$��C��Z�)jDRP��3�lu�v ����yQ�ДL,ֱ�f*Ȍ5��C�	�IX�6mľ�L(�5)�-e�LAd"n�PěahD�_�t�
�f+�3���[\zP�P�Z>'O.u ��G<M!�Hj�� �X92u�hh�	_>�0�*햩[���xѥ�'�0]ڰ+T-ɜH!�Ӕw�<y!˓1^�%٦�$.�fE��j\$H��;/A舼B��%�<Y��H|H<y��ɄH~HG��2p����a�I�	b�!��ʹE`�� !��c?��"U�[�
5c(��\Ȯ�sj1D���j\�XeqC��E0圃j�ع��,��36Hi� .؅`X�c?O� �v LNnhu�S(vҜ�	�O���48��t
�)��o>-��A�{V�a�/�$G����`S3Xay��_52ؐ�(����EF��а<1��#��5kM��@ؓ&��W�	�]
�駧ɠS��=5�($��[aĜ�����/Lwꑡ�@)��7\���K�M@x$�����6 ��!�D��bV�KB�����"OL	�Dт%mX@aE��>#�n5�A�(N
0�D�U���#-����x2eH�n�u��C2 pxv�����x��[�f�^�k�b������tU�t��QR���9c"X5�	J:Ob^�Q���%d�H�MQ�q�Jz���1 �j��[Zg^q1C!���<)��O6!�ܐ��f�e��F�»��X3B�Ϻ9�<�C�DT�&��aj��"��承eB@d`U�{�3��wMХ�& �v��dŘ0u��'��t;f�Y�sƤ(G�+ov�%>}[�	�6��x��� �%<�D��@H$,B�Z3�
�� xk�#��ް=��7~*�
�jΕ�9��K�D5�E�w�%��H��iU�`��'n�\T!dd(~)J"E��zh�v
>m�so	�S�����ݴ�y"���`+\4S+	�'��l�QT>}���2&�D7��XXb�M��V���,	�`$By��!��p�O�~b�M��w���jW�� �J4�"�t���&i�E(�Ii�ہh�P]�@��v��٪�NӠ~F����O��3�Z,�:	��AU���mJD��.�!}R��'~��1�6e�^XJ�MH)G�1��y��ȨD���Q/��ucV�%r6�]2�p��NV<'Ԅk�G�*�h;w��K�~���L;�~��rLV0q��DE~i�$x���@��pޞM�DG�F��� R�HO
�;��y��x����|4��d��$ֹ��C�<�2��e��V	~�AuD#5�����-��(R� GVD����pr1qW ^�xm��D �)v
)q'��s
�Ż�f��H��G�~p=aw��?{g ��PĀk�DD���QZ	8z��Ĺ, ���D;���B��{����X�*bt��g!�M0�ՁP>xg�q�Ҧ�|��Z!��P�˷&�D��D|TY@D���?��G�
K�z���R����l̓S�	�Ԥ�.{Nd � ����S�$�l�KB��7u���{�O(WX&�z��]1P�nq3�I=Q��U��/1D�!c���p�������%F�.���JO�$�pV��=�D*tOÈX���r��W`�J1铋A�D�>��5*�-"�n!y�N�9�d4�H�q�#w��o�eYrd$F��pҠgѻq�6`�ߓyv0&m����S�@�\�-:��c��Xa�ܽT	H�E�!t�`HV����C���nqrԈ\�|B��%6t�K�EG�zjd@x �aX��z�*��/���� ��Dc�}���J�PH���2��%(+^�I��rudA+Z�6�a��܂��q��N�.��4�R�1��P�˟5O��X�#��� D?xޤh�4΂��^O�Y��I]e6f����؃y��'_?��&�@@�J�*�}�ͭK��1ڷ���u�lt�B��g����$H� z� |8wꇆ-�#<�.� ��E��I�*����M���q"�	�z	�-?{ߖ��A��$��y�0��2-�������!Y�?����K�S&�9%��x�ɂ��@�z�<���	1[|��i'ݭ>0%ړc�	�
t9��Hc���ӀӢ<=����u��I&W?7푈�d)�π � ��J�Ĥ1@�ҡ� 8p�'�,�q��K&E*V5p�`Ә$Z�I���Ʃ'�\tq�'ɐ!� \y!��6<�p��m��2r�9b�'�D���f>}Q�ǉ$�`�`���5&Ŋc�bШL2�9 ֋��Q$�x��`�.~Ԉ ��A�;G��Oh���F�	e�\��CߕS�J<��ˁ�x�\$hS>h�aqE��~����,�1�DŠ�f�ONyd�6T�4a�;j��s��E^DM��Ҷ��F�?8�Lu1���Q�")X�-�9n���Ch�Gd����3�I�Pm�@=��`���*j�`�i3%��{��5wl0JG%�&������Z���`"uU�����	L��t��O2zt *���>��(�[��Ʀ9D<�bF���cqV-���� �az�!�0:��r ��z1>�1r#�Hyې�>$��=�4�T�z1��:�@T�	@�+r
Z J�V��~�@���}L\eCЉ�(���Y^�(��*ɸ	3��Q���0qO��0�KC�;8�Ң%N��;:��"�Ig�^	r�aK����_"o��a!5�L�Q��C>�9�F 	e�VFy�HLۜ�dNG
"ʌ��êؑh��a����@�v�#��� [3���Pq�t\RM�!B�s�
��(���G�O���G�<t�| �p�[X�(:�S���i3�E�&_1���'?�vLN�8��<%�A��7a\L8@�C�d�s�ʡbJ�:0��"Ȩ�y�4�����m��^�$�!�̈���F�m���z�f	xgDȄ�
�a�`gؐCԂ8��䃏F�LB�	�D�X��5�v��� ��(B�"�Py�DƇ� Ԋ�[��0-B�#rpV,Y�l�����k/ر
�'�My%kY��0s���T+d��
�'��2�0�"7�P�x<T4:�'AN-@m�>ע�yGK�N9��'��0��.y�$:V��'p ��'����^n+��:�Or>\�S�'0�&S<x�v`���Y�b��
�'۬���
��:t�C%PZ����'����͗�o5r�#��I?T��͡�'��๰kT�o7�KC)�On�(��'��i��K�u�����H�B�V)h�'��]i&B��s鞰	r*SG�a��'|D�C��X�y|&�2��?6��%��'�(���!5����(��\z�K�'��%0t��i�R�C��(R�'"Ф���K�%��
v��99:�
�'�Тr�D�����T$��;����'�ꍨ�BRcL��8���?oި�'n��AG��z�X�(�MED��@��'��qYKF� ��8$��3�T�Q�'�D���		�I�l\��gN�f@�;	�'aJm��"�m1�����Vβ���'��AzSFD4�(L�W�=I?�ف�'D��b�ŝ�1��(W��/� *�'TVȑS'~"��@�����'��XGʓ�F$����D� N��9y�'E��0��
V�"AJAe޺?�h@�'���cD☃*�ԅ�Pg�{���'S
��3�
.6}tX:�׋L]2�'���#!3���)�@�@�D��'P��V@@5C��,b�<{�69X�'Δ�Cԣ�sR�y9�k�5�tD��'wr�C�u^�M�f;s� ���'m���Ï�_�%��D�hWi;�'��Q�s��bPi� g�R�"O~�+H˨0g�Qr�-f$�i��"O��K�j��C�X��'�)fp0�C"OV����n.|4��m�:t�(3�>K�r)����)z۬�j#-DL�d��uC��=� ����A��%��I���
db^�1�� �"`܄LBDʊ�^I��A���#Z��!A�nȤD�������t��9�5([�4��.i}����ZKtp�Ddݷ�!��ĞZe��$��R��	=��b�b?��thЕ ��j�.E�/X�I��<���:ȼd	J>E���p���
��]��ٰ��+�?7
, �ڱ�<E��+D�lDf-g&��{p��D,D�@��VD����<3�3�T?=��dn��0�G_���6���@@�*$�9�MI�O�� ���5�/76dx� �Za���>���G�r��ʒE#�9O�)�?A0j�,�d�{���?T��0�wk��`�?����>{7�FL،A��?/���#wW�<aԤ����w����禽���<�;Ʀ�R�h�?�ZĢ�+ĠpL���M�7 �<)(�"�8b�����%G�"t~���R#&�m�'����C �|ʏ���Q���Rt��� %�$˺	��h�OΑ�� X�I ����֦5;��^�X���f�4~J��꬟�zw]�[͢]�K<E�D�î{�]�)[�G�Z��Z�M�C6k�:aN>�'�(��irb���Wd��	�皝��yڵJަ'�ZpM>ѥZ>��'>�'5�P��hX�MĞibCC6A��}Z�N����l�)���&�	A�EBĩ�#�����B5/��'F��+�j_8O��~����V&Z��J��#��9�X�Ԓ�G�=��H�`F��h>,��j*]�"�*�ϵ�M�����>U\�H�k7}Zw�>�h���F�����W;�Z6E�O�%�qd�i~�L�T�L<�'s� MQ$�!4?YІ!34p�����ē�hO�O��D�����Z�K-��%{���O
dy����(����`e�N�zD�b!S0����	�MS��'唹��f�fx=A�BL�U"�A	�'�:BN�T���vL��'��1���� b^���e�/eg�M	�'��$�3�Cv�D#CH��I�P��'P< �ƀ�!K�pY2R�43�,��'��ȸeÙ�r{�ݰ�����'q6����W�!FTTc�B��"��	�'B@̣э�EL!���?>LP��''�Q��Ow��b2�ԃ@��̺�'�h)1SԀr"�j�mٱ6��Y�'RjX�Rʕ&_�4؀��_�-���'Xv���׬��j׫�s�b(q�'ln��ɘIQ���%閍w�U�'��<�!��V��LB2NE�F-�c�'�Z\��3w5���T��)�%�'�XU�϶r�D1t(��;���'ivX(���F�^@�������͸
�'e�@�#I
tA��g�4{���S	�'wU���@�)' dyhut�c�'��`&)�%���X��P]_ �y�'�&Ir�����*�N����'��-��J�����BK,���+�'8���!K2|rxqq�	��Bm��'K<5a��'sUh��聡��� �',\@�"x92�9 *�Uq>��
�'i��[�� ��h��H,M�`���'Dtp�G͊ v�y��΀����A�'�\e��ӌ6� ��BA���I�'C�I
�K��8�k䕠=���'��S�Ξ&P!:MC�$W7�Z�A�'�,����^1\|*�_Y����'��)�ba� Iښ쳥�V�z�XX��'�Ĉ�Wf��l������?��'D85 '�]�+������& �����'�Z��a�E�Y��1�B�l�	a��@�E ���eD�B��k�>�A�d�)��cp��I�
C�	�	Y�7K9)��%D����B�I 	K��[C�׺1
�����}��B�?Y�X@�W��)ǒT�2�غ=#�B�ƒ���0�Ј(�cU&�B�I1rX���M��9n
���X�VB䉑6w>�;*ǚX̼�f	G�_/$B��1��C�� =jňQ��M�C�I�S��(�*T�A�4�������C�*:X�16Ί �}��#ߙN�C�	�}Nr��¨��+#�@B  �B�)� �p�s�V�
.t��Ռ�r-� �'"O�<G��t�I2���io8�"O�r�!X���CcA�V,:�"O�M�w��v!@)lV����"O4�f��}� 1g �.z�LXd"O<0���S�l�X�9&�
�Q.Ba�r"O��C҉ �TS��[?:�(�"O�U3B�wl�� �C�dh`��"OfP0g�W�Y��84�J�zU�Tӗ"OB���L�65���9�J��,�`4"O�� �K���ŀW�+)6 �w"O"���
7��I���} �j"O8(��ܪR�,���-E+O����"O��T��*� P��S
��@y�"O"]���w���S���#��d� "OQK��T�M$�HԢ�?3�؀�T"O�a��jO82�L����T4�u
�"O�����?^������J
�JR"O����Ke+X��B�2�.��&"O6x 5�
3EBb(�2,��
y.q�"O���
"欴���V��f��"O� �A���[�(x��S��>	��"O�Uh�c]��k$/Y�p1(�`"O$Q�Aa�MxV�a�mI�@����"Oy8CJ��.Vn	�V��Fg���u"OX����P"��9���=^��u�d"O(�KE��O���)G$&A�΍�"Of,q���*�^�xUL�	�у"OT��L��$x�
�`�f�8�"O��Q�7�,�����M��q"�"O��0��e:.P�Ѧ�>�(�E"O��ZCH�P�n��3�K�B�Laq�"O ѐ�	�#pH���EM��6M8�"O�d��`��GĈx�W�J��0��"O�M��c��o1�B��2J�∃"O��vH�/�2�瀘�T����u"O�$J���g9ą��[�Xv��`"O�y��I'%�:AL'wT>��#"O��  �ˬq�p�D��dq��s"O����_9����-��oR��"OVdCW(T2L&�5Ð$&B�퀡"O���;_�~�S�5%NppbD"O����Ѳ:592�+(bK��"O6��DN�.9I�Ȱ�
�pۓ"O8 �u$��eF���3�L�yk$���"OL���2�N�ye��20a�	�5"O����;[$0T�.Ӱp��U+w"OL�r'-犑j�K��&I�Q"O���L�S��kb�:D�R�%"O2�c�$��P�*��e��$�,a!"O� R�!08�i�&u�����"O����JXՐy����ey
)�""O�D+r��%��T�W����r"ON��'Սy��K�C�-| ��"OHРA�&?�N���Ϗ.GC���"OtH1��X!�nX�M�y2��i�"O"!�u�G
q�T8:!ƐG��Ƞ"O��	�a�,cPT��'M�F���"OL��$d��$�  /V�l���"O� �b�pN��R�Cէc�r<� "O��P@(B�P�")�¤�;�^MV"OȘ���O�<�x&�;h�$qj"Oʔ�Ce�5k�X)��摩Q�R�х"O���r��'`@yq��S�Ry��"O� ���k��N�"d��n��E"O�p"ѧ@�l-�I2Tb�,��a��"ON �en�(?%n`q���N恡"O �h�E�8ƒ$
G�4~�j4��"O~�iaeC�m_�d+t*�$PO�=��"O�l�1̏�����IK�z/�!�2"OR��!A�NP9�)�a>|{�"O�%c�$"p��+`i^� �u�T"OD��c*I
�b��S(� _���#*O8y+�*$�YZ��Y<h�t�	�'Ӡ�s���GTX: A�!j��Hc�'}ؤyЂ���lR��Ĥ9Ⱦ���'�F`�b��rp4�('(�) � ���'��y�Vf]7�:�vA1H�	�'(�!�)ׯJ�u�挗����
�'ݸ���9�$��6�O	����ʓZBPS�Vu� �;�(8{��C�I�`U�i���'2��7���q�B�6�$�V2d	Je��+�q��B䉟C�������S'��B�I�Zxt��R����ф�4C�@C����s ��:t�| ւ�#GC�"80�3�k��\]pd!��:`lC�ə�l�7iD�5cd�� KS���C�)i$(h���\�b��Q�FC�I�xm:aA�&p>6ȣ��Pw��B�	 κ�2�@Z�3L�
���waB�	�.켩k�i�B8��M4��C�I2DR����#�;XCX�` d'�B�	3g5J �\\�F} �E�9��B�ɽ H�p�� ; "!*7��>f�C䉇Lh*m dF&R���&
0�rC�I	"���2� \�}҆�R�''(C�=�T}�'_�K��:�%Л|>�B�I�f��g
4v�b�CI�=,"B䉢m�B��)��b�v1�s�ʫ8�
B��l`8cҽ7�T����0n�C�ɃP��xKb�ԙ &y*1�A+%�B�I_�P���I���$���0eB�I::����c��1���#��2��C�	����C�O	P��a�qDY�NC�	S�tBI$V8�YAF&
sC䉣'�BI�E,[A�Z���O��� C�IHM��	V��0lxe���_�B�	�iFJY)����bp��"W�h�C䉖_-��!C�e���7E��"O*���&Al�Z2ӦF�67�aF"O�$U�" (�5?J�+�"OV�fG�SOj5�D��q����"O|�2q'� 5��$�!Pڌ�"O����,xj������#���x�"O�<s�oצSݨ&�5�ə�"OX�
!V�@f��PA�1��5��"O�m@7�Q3h���V-�X �C�"O�A�Έ�aؔ8#��#]��! �"O| ���|B�dh&O�e1��r"O���P�?k0��e���Y�ڇ"O�<r2��"��y	э�-e��B1"OR�rnGQO�$�-�0}f9Q�"O�����[>Ç�I!&p��J�"O��.O(!d�H����g&�i3"OPU��-L~�,��I ~��"ObM��F7yE�����	6 �u��"O6|	�d�2R^X!0�J�.�Py�"O� N���yȤ�*_)	�4%B�"Ob�&"˺;D��k�IZ||�d"OH�"d��(�0vWR@+�"O>����k�L�#�� %)�|!Q"ON����в� �j�gE�b��U"O:I��%P9��E�r��:��\0a"O��06�F[Ǵ����Ƕ�$ �"O�L�l
�0���C�/�9v��0�"O4����,xveCa�M�"1��"O(	���-A�ģ� f�$�0"O|�Bl;q�j�;2�;� �PF"O�L�`��pu�4�s���Fh�"OƄKI�?3�|I��	�%��a�1"O�5�@��	,��V�Q�K����1"O���dJ'D0��(I�wҲͩQ"Oho�1ڨ����4R�D��0*O���2��G�&W�\�Z�'�𴓢l�aG8�"7)P�VAұ�'�2}��g/7�u`F� �����
�'�<\��^--$}�$�@
_�X
�'Y.c�a�.r����8#)p��	�'X���@D���I/�d���y�nӊ<xC�0�M���i�AJ2E�W�$E�,:%�4C ��?Qt��=R� X*��D&����n�qȘX"��I�?�c�@��Z��,%3b�(:��
��'�-*q�!&\��:���S ��"E�vd�@�`�ɹ�G<}؈�Gc-A�R�`!.�ɧ����]ۦ��N|©���x�cǜ[A�����P!k2܂��X�	����)�gyB�ʳ&-�r.
�<��MJAcT%�p=��iJ"7�>&Ϗ��	����3{枡p4��,	Ą5jy���d�O��4�r�c���OP�d�O�6��{Vjp�@� �����AP3�@��4#
qj֠K�-ħylލz����O9� �O��Ĭ�������H����7.ѧ��CC���'��\wȉ@�̵;�o�1��l��H�H�4���ݯ9��K0k
¼�$��:�^T��D���P�`��N���e�&	�'��t������#�B�~���hܠbЖ�BPb#���"��?��1,�B��\��iM�Hy�%�%}�'1�7-N���	��M�������M�`��7t,jӯ��?8���(I?i!K��q���'כ&-<&����� 3�r�c$��R0S�Dگ+�̘1�ϊ�=/�E� �(2ILYá�$�fik���+Ki�h�ũ6��YI����ef�y��AG'e� `��驧OT���'D4@�m�2n����
�+^ء
CD�.�\�D[ئ�9�4�?�(O��d)�DR�>!�i��+H�S�a s�BqO���4HV��`�� d^�:���}(� aܴ��[�ܴ�����1p��;�M�oF�
0��z�㞓'6 db�Ĕ�.���'-��ڇ CB�'/£ԉ���	����� ��ng�#L
|B|�!�U Fe��A�`\�;�vܰ���r2�!��c[oJX �
�.zzT�8�K�n�	�cr�ll$ᙆ~L�u	?��h�6�d֦	��	�{d�{�-�2�`Q����*_[Q���?����?��4���3��׸~��q	7
�.s���@�d�R8��+�#Y;'�h��O�iiZ�;׆;#���r�L�D�Ԧ�r&����M+���?q���U�'�F�QF�V�?������A�m,(D����?���I�D�U�N�&��9E&�8��!
L�WE���Xw��Up��mĒX@6%�u;^��}␖m����UC�nl�2���Q	^w�|�q���EeJ���Nψ�:�f�z�� �O<�U�����45 B�O�Ӷm���á\9| ��QB��m������	m$��e�u2��)����'ip�ɮ�HOz��B˦) �4���!���e��qֺe�4+Ӂ^��S��3�M����?���|j�@��?����?!�4Q����*T"��M�v O�|U�$kf�ϑ\Ϫ�3�_$Yq�`j�c�3Q�� ��Z>���nN?J(�sT(2�P@�Cn�79�t�g�Ɲ	 �M#��ȹ(���3��$s��@��s�ur ��`l�Awb�K��a�r�L��?y�id6��O�T;��Y��u�'{�,p����M�dP�)���?�.O�=%?Q��i�)0���$/�[-<�R�-�I�M�R�i��'�Z���O�֬��m[p��b@�0���0�LM���ILX�Ĩ�/   ��     �  /  �  �+  4  |?  �H  �N  6U  ~[  �a  h  En  �t  �z  	�  J�  ��  ϓ  �  V�  ��  ۬  L�  ��  �  ��  ��  ��  s�  ��  ��  �   Q �  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p G}"���P��չ���"�:i[q ��rC�I��	8���21�A�M�:ph��SHX}��'���[V(�d�@u򁤚�P�\��'��+���8?��0�d_�
���4�yң3�O��ǫW�Qp85�U�2��v�'��O��B��\�Kΰ|ð�W#7�x�"OP�
�)ǱrR%�B�$��`!�\���iO�(h��*�Ӌ��T�` ��M�!�^�BIH��ş�o�|�ZtE�I��9���|ڋ��A#UXD�`.��B�h��U�.<1!򤊎5�0��< �H�2�A�!�@7���SmC5ymF�b  �%�!��*Yr��x$�X?3<5��� e�!�S�q�2X�R��.@�AZ�	�(V�铬~��'
mƋ�(�0�A@����5�
�'�N���Ϩ-�Ё���S�<��'À�i���OwX�n��5�"���D �'o�\0��W��yh穚Zv���ȓ#�@p(T��'��]:i(���S�? ���-7�l��`�)#�*
�"OlɂӌL.589T@Q����"OH�Gk�q8� D�'�����"O8���ƙ$Y12	pr���D�5"O`�ŀ�,#����?x��E�"O��QR�J�B�p� ��iijEh!"O�a���p�����95��A��"O�<7G*o#��ZF�R�cn,�"�"O�]r�Di���
1��j��c�"O���&G�;��j> ���0"O�,Ӕ�M�M�tA�O7	�X���"Oƥ��o��^x
����ěb���W"O�p!wnQ46-�,��KYNlpG"O�E#�'�?5�B<pIּW$�!0�"OΌ�f�&.K� �CH�'숽�e"Od!�7N��Mh�!"�gK�'�<��ҙ>Q
�f�Ja�vHY0J�<As&ų^T�y��	G?I��_�c}�H��B�gSNx:��@D�<�� A�q���C��g本�d)�u�'�? v�_��֤�v�ƾ�V�+��9D�$JŢ�/��X(rş,�n��,3D��('�"(�Z3�
�.C\	XA�$D���`�(\b]"0�U"j: �0d�ϸ'����>t`%U�V��w�ݾ6��d���5T�(�j��5�����oގɢ�;D��2���7����O�,%@\��9⓽蟊��E�i�M���ɂ_0Z�ф"Onѓw�,��d3�NL�
6��On�Gz��iT|�� %�Լb��4i�s!�d�6nJ�c�/F$wz@A�H�:vr���	����'�PMS���vo$����&��P�'n���זSr�zC~Qٴ)�^b�pF{*�H1 "��T��)��
�
�ʗ�'����%�I ����T(�qD�}iv��	fB��:�]0��m�~ز0��<v���`G{����:�-U�8v����n$w_P��l7D�K��Z�p�T�A�EF�@��JQ�?ʓְ<gd�8�py+u	[��Y�HTR�<��B3Ȏ�a%F�S�Lu�!��W?a��퓱k<n��#D?�	�𧎂|i�B䉱,�B���_>{Ӫ���I·$ʺ�'�a}"Aˇ0dX��-��k��ق�@8�y�E�n�B5[�놤<���RA�,�y�moV�ygM�	:u�ipB-R'��>ic_�<iǡ%h�<U���~��L�D�0D�@����	w߮bC��E=(�:p�#��g�� T�]�~�H�)��]�H9s4�$�Ȩ�
���߭GC�قB��a�<�6�'hў"~ZB�Z�s5�0���ɪ����4����hO:��	N�,H=��-H<5.�� �l!�8<U�]3t��x�K��Y`�p*�{��'=�1y$��p�q�"I�)nD����y"f�@b���ţ:5.�r �	�y��C9!p��9ud�(+ P�p�l�yb猁F��0a�%_�ǖD�"��yR/gUS�I4|�,KP�,�ybCڋkҴѻ��*�Θ����y�'<� S�I�K���� �%Y�P  �'�D�1��Z�+��h�.@�ar����'τ,y�^S��k`�W	�J�i�'��pF� ͂���ߢ-�����'�`�g�3r0r��f쌖gƠ 	�'��0f���P��E�ٴ@y�l��'�� ����-�F��V�I	� *��� ���A/��cG�Ջ ���X�O���ꃹ^ ��'Ij�:y��%C*b!�d�O� 34L�� b5�G,�l�a��	x�O`Q
�n
�BHjl������<��'E4m;�f<^OP�+R��7)�p��Oآ=E����[SDPd�l<��q�*�p<a3GII?�L���w����d� �mC�f�b`y$n(D��q@�ʤO����E`�'}�n��Fh�>y�'�qO�>�v�H?
�T� b��-9Jh!�b&4� K�$S�7�=
%X5����#�hO?�Ʉ	��]��!�L�+��p&B�ɱ���8&�>g�P��(�lm��Mk��D>ʓ$���@wJ�50���B�N�P��	ן���s1�D'��.�V��M7o|��"Ol�8P�2z(�Kwo�^`|y���o�O�ऊH�W�и�6�J�%a��	
�';��FX5u�z���n�E�BH��'���r �L����&B�%sg4L
�' ��"���(b�@�#��T@��ؚ'˛��)�R�^��K�
� �"A�!0�R���]4�Q��9a���w,Z(`a4��>��|�$EV
/֔��H��]x*,Gz�'6^��'�ؘ)���H�̊!Y#�2�'�~0��M���j���x���'���(�b��H�~�����$uJ���'�x�+EbjtJ�`d�(�'���P���)<�}j���
UR@��'�4!��"�x��V �j��`N�x����W����m�E�:LQ�h�$tV~�=��!\F��(�$Ivġ�-�2G�ćȓW �ms,�,�LI��c	晇�2Uh0ED���p$LE2@�E�ȓ=�(DjJ��|OFte`�RO�=��\��Ȍ }n�t!B,E&N$��Ap-Z�5I��p��%S�&�ȓy��"���c8H@�a�$K�4نȓ{�8I�4HJ�b��_�|�d�ȓ\�(��B��o.8%�؝p,>��ȓg��� �cЧ/|�Y�6E�V�n���T�A@�0�(��s�PP#���`�Ld����x��� �B�N��*[ ���{l����
-�|��ȓ;����A�	�9��2���>؄�Y�$ꁣ'B l�R�� f%�ȓ;8tH���+��Y��I�	[�)��gE��L���æ��v����z�JH��G�0��S�fW�e��ȓ6�#	&M�Pళ�9ZP���$n�չ�W�#�h����ǫA��Q�ʓИ	z%�Ul02���R�'��B�	�q*�S�Ӆ5�J�{�	�Ga�B�ɡ^28rd�D#q�>,�@$�#~B�	�ogL��F��=~���� �.B�	�iIx�z#U�k�t�Z0�+}�bB�I Y��&s1�Q��ǌ�W��C�	/2b�X
�R>f�tY��
L�_h�B�	�8�2a3��Y�6�3Ĕ�H��C�I�k�3#���$�L4�P��9�\C�&I�\@����d� e�2F�JC䉊Q �+@��;<z�;���w��C�=�v{c�Ǜ�Dy96!�&�C�I�E�$�)慔�S��DQ�ڃʰC䉘99��t��F1ac�ܼ|�~C�	�po*��s�ϼl1��+��C�)� ~��jѫH�,��d�V�#�<=�u"O~@s�N/���P��"�n2�"O��b��2����D��o,2"O
�;5��9NY̬H���TQ�I��"Oް�ዎ�0� ��nߘ@b�����'�r�'���'Br�'�r�'}R�'�( :ҪF�T��)�(�<%s4Y��'�b�'���'�"�'n�'K��'ˤy��H�Gl��� kHy� �'���'���'r��'y��'8��'�����V3D�>�@�+�&k8as��'kR�'�b�'r��'�r�' R�'�0�чS�i6��	4i��m/V�a��'	��'���'pr�'q��'Y�'!��	o\y�#�~�|�{�	��?i���?���?	��?���?A��?��I�
 ��gB��]��y�Uj9�?Q���?��?����?����?���?!�� ��8�`��	[�ar�oR<�?y���?i���?���?1��?!��?	 D$ "�@����[-
�A!�'�?����?a���?��?Q���?��?�7Ϝ�A�4�9���@��e�#���?���?����?Q���?����?A���?�Tn�:��%�<!z��t.��?Q��?���?����?���?���?!�BA89$L SE'�?	����-�?i���?I��?���?���?I��?�'b�*�c��[YL%���K��?���?a��?!��?y�X�6�'�����x驆h C!N�"n�'!���?1-O1�����M�CN�x)�dcG }h��b�"���'pP6-�O��O�9O
�om4����+�%'���T+1����4�?U�5�MS�O�e�`㝑n��U"O?�(���`�,��㦛wB����m>��Ο��'��>���S�q�z�!�X�`e~��NX��M�5RN���O%7=��	� �շBӰY�K�-^1�4��+�Ц��޴�yB[�b>Q	�Oܦ)�A�&��K�'���k&R�^(�X���1�͢UgP�(��4��$˄/�� ���1Y~zyˆ�,y��<�M>�S�i���Ӌy�'! 0�e�K��6�*���h�B}�O��'��7-��uΓ��d�-��Pb�$|UP�жņx\�I3HX�욂KO6��b>�"K�ĺ{��'B�-x��0�0�AmE%�"C�Izy2������Tz��ȁ�%nU�)�b�b��צa�4)*?iѶiA�O��C��9��M`I)P�ʰ���V٦�Bڴ�?��[��M�OI)��Ųz��h�i�&<`;q��^H�ZwJǪ�H�ۃ��*+GV���晫�Lܺ�V�7\�'b���&�}�`e�	�N�������3�h0D�0&�^�4�����* ��\rO�d	��:���4w��@+�"/��D����%�Ԝ��"� ���R�H�x1�u`�	V]��T�^�%�N�h7�E��p���+{��u�og�=�Q�@=t�ٱIX�o��4{���.
YPd�'E��<�-�V��Qf��%	,'0
0��UȰ��%���M{���?���|"��Y���'[��tx�hOE�D�Q�*n��D�O)�s�i>��O��hfCjq�e��Ry,Q���i��IR'm�"���Oj����:�%��!s��B1hp����`�~��2�4��Qk(Oz�t����?c���I<��I��R�7H�G�5�2�۴�?���?��o�V���D�'�"n3.��F
�Y�Ҹ�@�N���?!� �zH�<y��?����Y�wN�+N���bN�^uƼi�N��^O�)�OR���<�wnN�we��E
m tIcA��p����'2 H�yB�',b�'-�ɴ{��A��L��Z-����Qs�������ē�?���?9.O����O�,�c�Q�E�Pl�#Bf���Tg1O^��O&�D�<�FJ·'"󩟿v8��Dd�l�x{�bO�dw�	矬�I� �'���'�
�ҩ����lA�5ɠ@;3�)�L�\�@��ן0��ޟ����~��=��4�?��˸�S%�V�Q.�!3��:7,u�S}�'�R�'�����(l>e��ݟ�h��̇Z�Б�`f��0��d�E3c$2m�����I������=�M+��?����zPk�MM�j��--c&�d��)���'����Dp�#i>��	Vy��M��K�4e~6E`Fl�=a\�2q ������柘���͠�M����?�������?)6��uY̜�Cd�!N�Zđ铠��	ݟ,����ğH�I��,��"o>M��d�s��@���7gg.�0�i�Xq�4�a�����O��V�)�O`���O�\����E�Z�r��O� 6�!�L�ݦ�#m���I��K��v>�&?��/T;X�����<�Y�6���A�ڴ�?���?�%et���4�?1���?���?���"P#S��ks�L�Ճ��DmE�I�4B�)���?A����fO�"}y&,��.�[;�,Qҳi��	/��7��O~���O���[{��O��'$�-h	h|b��9�D�2WR�����8��@��ߟ�����\���G��(�A�X(7of%�PJ6VD@ljܴ�?���?���E��jy��'x������11m��]�&�x�S�Ә'���'\�'�b�$�<7͍G��I���B�#��mƅK
y>��lZɟx���0�	��h�'������MҊ�n��oZ�:F�ȑ���$5B��?���?�)O��ʠ�UU���'�nx3��lV��C�na+ux���<mf���d�O@�g5O�����\���3G��B��҃0�d6i�~��O�$�O��Ǡ��������?5zUV4�J����3sa���>�,7��O���?�%��|����?ɔk��|n:� ���A�7$��h�[* (b1�i3��'0F�1�le���d�Oj����b�)�O���jC[6�*f���ku#�v}��'�
"��'�ɧ���~�'یGT��g��8?l��M�A�cˇ�M+��?���:�'�?A���?7�O�/0a�V'�Q���dZ;q�6Q'��'��i>A'?��	^���BȆ#N���� I79�X���4�?���?ɐ ��'[���'�R�'x���uש�RG���@Ŕ0i�`�5H_��M�*Oz�H O�#��?��Sş\�I�R���)%��{�޴0JQ	L~@;ٴ�?!�(�jśF�'&��'%R��~��'��U�i 0���E�С nF��4u�ȰK�L�<y��?a���?���?9��X&X�䊖y���/�-��v;<��6�'�2�'����~�(OD�Y�\!L�!b�C"�f��Q"Y6on�xۂ3O6�$�O��d�O��D�O`��_�8aFuoډ6$h  a��
�l�䫜�X:j��۴�?����?���?,O���͍c��i� V#�m2�A�1v�<�9���4<�'c��')��'��mv�6-�O&���&x���Zb�0c�N_'�4���~�(���O���<��`4��̧�?��'��9��m:OmDL7�ڻ(�����4�?9���7��u%>��I�?y�Z�ؐU��&�\1j�c�=U��KH<i���?��(\��?QK>�O"�Y��-�pQ�Uϋ ؐ�0ش��� Q�l�����O��i@~��߆3^�q���O�ƥ{4̝��M����?��e���O�J�q�h�Gw��Cb�>o>�xߴn�z�Ըie��'"�OkO@���4���z���*M4h<�oZ�%�F���T�)§�?��.ڜ	*L��PE�5%�� ��E%r�6�'��'h8`��<�d�O����,!vN�	XfdӓÌ%1��u��y���O֭�G:O�ϟ��ܟ��0.-)&�-��$F48�Dפ�M���c�h���xR�'��|Zc�fDk�J�~���!�^�H}�aH�O���7B�O˓�?���?9,Oʔ�TF��U3V4*�Ha(ƈ�r����x��'d��|��'erC0o�n�C��ߡw�x )�jL�{f	C��'��	��I���'�����q>���R"�] �J�<麠���>��?�O>	���?�1'R-�?a@�X��TĒP!��&��bRerm�	ş��ß��'�z��Pj8�� ��%%(|R= D�?-��Asu�h���#���O�D�fS��D8}���t<�AcT8�:��cN*�M{��?�+Odى�G��8����*���f��y���c��@!%V� :H<���?A��+�?9L>�O\t#ӫ=��	�D��@�[�>�a�D9@y$���}�m�#Fܩ��Ǻ�Б�tc��y�+t�A� ��0(�	s��rB�2� m��a��$�鳇��x5R��g)���ǔ$O0i�&"S&o��0� !X�v
d��n�"�"����3fZe
d���\�� �C�rPQ�$S�ZR40Pl�(�R Yu��)�.0 ��f�k�d�.X�q%o�rd$��l	�T����'�B�'�Deݝ�����5�6#K�j$+[�||!Ѷ�K+o���S%�,E�.1��F[���S����3���֙nΜ� ��V*F��ؑG"l��	���-T���H�)����ߟ�Ѐ��>�'���`&#K�[Ⲍ���+��:�'Z�ܪ�7��6 *�D�O��D�<Y0�V�K:���Ӫ4ش���r�<� P6UE�̀��i_�(`�턈w����H�'�>�0 bӔ�U
�v���`�&[Lɑk�O��$�O��$�	0�����O��ӷ17��p@�եAs顀�ґ���p��;d9�q�G�<������!;��:u�I0d;q���,�hҁk�8�q���\�.�2�w'�;+�"L�0�_�~&���/�:�������Si�4j�"�����
'�eh�	!D�`�gS�P�:��@�cݶMz� D��s��ҵX��ĳ3�����7'��p�4��K��;�i���'M�ӅQ,t��2G�mR4u�pl[P>.��V�۟l�Iϟ�8e߳k.�1M��X'�a�c��gP���3k�|�K�kޝP�,͸ĆZ9nQ���#`�3\��5J��Rj��u����"��[7	�Z!�b�Hh�\L�r�4�(O�YSS�'�X#}ң��dU� �Ό�F�����bR�<)�)Lq�u��Ƀ,fZ�����E��(M<�ӡH{�����(H�(����<1��T"b���'��S>��#�� ��Ɵ�"͍��Piy�#
��Tq�l���8��o�s_z���Ǝd�����9*��m�|��me���v�Y�6J�ԁB[�_-кD`�1\8#��DhLf}�ւ�mn��U�$Bl�-�W	��h���HRH�#@D,v��1�'����i7���2ԉnE���'�3�@�z����wx��
#��~��*gCZ�)4BH�Q�4�������D�R�$��_���p��ϫ	@���A��<Mj���O,�V"D�3i���Ob���O�񭻁?���:�����_��X�{!+�!͊�91Q̥� ���ۤnɯ"O�D�lJ�..��!d��{!� ��� ��B��B/ր"EG*5��HbٟL�ۢ@�uܓi��HG/
�?C|��U�L�-	���{S���i�lژ���?Y����Ğ�r��lY��O)W,�#������?���?�Ϙ'�"���1�����N���4o�6�֦='���?�'&���b��q�&~���8K�4\�^�4��O����Od�d�l��t�թy>�v��Z>�p�� ��k �����r��0?ґ �+�'?H�X��,F��y�	6#!a��/�Y�n�	]j�+E�ܺ|.���e����ѵ�ʧRE$	��I�J@��d�Ʀ9��J�O�|��B	($�6�`d,�M���G*��<��\,%|ٙad����ʑd�H�<�Ǩ�0��M3�*E�~�4�ؠ,��<�$�i2��(�'<��U����>4u<���ӄC��E��<��I���Ѻ1pr@C2�m���ȓ+�	�S 5/��a��Ӽ��m��EUN�j��НBIHuQ���$����&�6���cX��@F1^d��D�\QB�Y�o�Lx��G�H��(��W$0�ƺ"X��j'*D�,�ȓF6`����9��ݣGy~��ȓbJX��w�ڟ[$e�&Nƪ��M��`��e@  �`
�U�
[)`'p=��iϢ�2�,ه���CA�׽
�����:�8��d֯*|�A[��;"��y�ȓ>x 5�����<|xЈ�4>)(���> <%Y��D�
�μi���.�t��ȓ�
a�hW�K8�ѲՔ[��ȓFP|�0㉄����c��}f��ȓ,U��▯�Q;�Uy����9�ȓ#�0�����:[��-�����Yr���$�{3,ԺĤ�8���qgP��ȓm��ܹSJ�\���if�/s�N��\I$<qD��#|��C�iH)l7�(�ȓde�U��@T$�c����@��5��}�D��O��x���`]�ȓ?��AE���<#�M�aTb}�ȓ!�^4z���S�u��盔��݅�Ӓ���0��d27�\/!�~ �R+D�h�5�
 L���:�5
���H��(D���T�U�¼�j��ۈe��u@�(D�0 !�ng.�
S�0�~
��*D�TB�@�z��6F�v����*D�dC��&�:Tyv욃Oe~�S =D���r�eo|Cv��[S���m<D�������<'�3��`x"@g;D�x� ��@\�)�c�.Q��J�'D�X�1K�]~����#aV���n&�Ovx�K�	X�y�(ɯ1�l̉v�(z
��U- �\!�F�2��=JDc_�e:�`�:�M��9�w(���O�Fqb��;J�x��T�<���'yT��"���&^LH�'�9h-O�Y�) �wތ!��i*R7���|J ��˓m�^e���L�[Ǟy�Ccۗ&����EV(<�@�Ҙ.a���+O8/��oχMt.��.�{8�b����\�>Y�$U�y��.�(9�KW�T,n?�U2�BE3�ab�L&���vO�=��:���u� ́E�4-�'���7�M��iu 6��:5�ɒ?��ЂFf��%U�X��͗TR��	r;�-�&ς�U�"H��h6������ƩT$!�\af]W����&�	�����/JD� ���8�MS��K�)�|Qv&^������XG}훒sq�̲�,� G:���ݴ�HO"���A�gw�t3ai{i&�Z Y�<�S��)� <I7a�"�h�$�s�'��A��`��h5Ҡc�U*�e(�a�6�S%�FC�'SЭ�'�p���J
�_�b��G@�҄(��*Z.���Q"���0=ͻT}Da	3'�?R��9�@8s�H�'���3H�<ͧ�D`��IR�n<|u)]w�z�3#`�q8���lą4����ǜ�1F�i�Щɳm�F�
�Y
�0����0��=�6�dg�m�3BF�`NR���I5vf���'`�¼�F�X-(�jq�FCw4pm'��0�
��Vnh���L�PH�-@ͺ'�ppa��eL�	�@
�-^8]cf�j������Y?a�H�����+LlP��Z?#<!P�F��6�Z�n�2�ʅ�dBeh��Uc��5l�\"w�,��~
%Q�@jb�X�b6��J����\��ĦIpI�:"^h��I�&����R"I�wmLɘDĸ"o4`�?S<O"}j� ��'����n�I��y����#x���<m� �Pc��2��ϳC����#)LqFР��ME p�I��hO��JBC�Q�(�{I \������;� h��̞R|"9�F�ʁd�nA���x����CIP܀fi�X�ؑG���qO���D+-��(4��: ���{�U�h��V�1�� ��lϋo�uq��%�|H��aC�Y�p�#R8�Z���,ȱ^��Y�a���EDy"7��tP)�1�K�=C<�DEw��CE��\���$W16���5x� �+ֻ����#�hO�HX����X^1��L�N�
��5��j���Aӓ
����T������"��*��{�ܦ]����������	���Ϋ/`6����D<Fnlt���ɃƜ�{���W1��)�4�)�G:q�	��ˇΌ��y�\���'B�T"a�LJ��.ՙ����O�a�TJ�0)���f�aت ���	 w2�J#d�Z����"��p@�s/��t�V����D�>ډ'�ő�"L4eh�{uo�9y]Xܚ0"A<)��EQ�Χ5���){���DZ&����,/9�Z�|I��'�Lb���!Kv��A�O�6b�D9 ʕ�A��l���'��E;$ʅ�%�m��^<��u8��F�iF6�	:�ʐ�7�N�H贛bd{�"ON!�]w�6�	F4ʑ�3�wȸ����G�\o��(`�9`"�1�#��Q]���������}ΓY�l��4��=������m_F�m�-�M3h� !"�o˷Q�f�;���t����.j*	H Ǔ��x�0#cH�Y��l⦮��D�<�	+s���s��IU��Ș�3����{@�L�u�>����ߣ0��@3��Q�Gt��X����>�­X4@Բ\�V��N��h[�Z$i\�D@%�%.��a谁��2�d���P$`��'��iڟY��`*�.]e!���l��sraz����P�FL�L�yS���Ǩ�z�U��į@���2��F��p��G�~�H�
��i&�c����LΓ~��`6�E�e����O]/]��%���GM+oݰ���b]!&����d�oN��)U2�J�Qs+U�N�F��R�Ų-S¤"��.57Rd�2��@!�#_����Ȗ{\ ��4B��5GO�y­�!"ҧ.ШqB�3H���^?r��S%�H�H�jI��'.���!�I�^x��؛{�����t��8"��5p	����O:?�uL�Oi{q뇄6��d�)[�*�� b�Z�0W4�����
fay�
�(�i:W͓UL4e�U�D�lFp�26-@�_Y� �d*���2����OL%�SnZ6p�.��(�p��0�T�!l���b�̣?FN��0�,������r�i91���(4�]�^ұOr�k4�E�Nl�ѵ�#A��a,ǘ��c���e��x�k�	I	*:�明+r i�H��+<����R�#�躵*7��~�ʁ%�k�i�A�d������́{�����fZ1D =C
��� ��+k��ؒ��5=YB$H!��Tܓl��FHZ%@�^X%?�Y9��i&�ȟD��%��w����ɿ�$��=7����	8
碄Jpj]2��8x e�A(� �t&Z�D'�$%��OqY�葴E\��O;:��a�]2zh�����1/ 	AN>���o�C����[v�$��kܓh���T�ĺ�$�ZƏ۰&7f�l�B���%|�ivk��(.��>�&�Ȗ�<��ģƂ �^��Ɏ/��mK��8�j-
V���v�I�0㐥z�D�' ���Ha�:�V,�$)^1����d �*�ʕ����	���1�h�'A�yk��yr.�w�:��V&��iP�l ES'ް<Q�\<OS�M� ��<����\�Eڈ����T7���z2D�'��@�b��)�OLt�e���g�4�{�9OD`7E�n{4H3�cO�Rj%�a�xb�׾T%�H�˄(,aF���e�&���?Ѷ�G�.!� ��Z� 6�| ��<�Z����(PiYҫ4�J����$G�-Y�AS`�O�PZ�}�P'��ܐ�� Ev��KB���yD�7% ��G�_�tTB�H�-rW
�Ix��؜kNRexQ�ҮR�R�S�U'�<#=��a��։'�^tp�Opx�4	!Dl #��,w�r���'�B��n ���.O�H1`[,��$���W�gs�e��
p�mI�����h�', H	�O�|p_wO��V_��Y����:a�	�LR4�Uqa�+�J$h��ʀ7q�SR/�a��?7-,[�z�{b��vZ
M�r�V�[ϛfH2ό0s�FK�)�n�Hr�I>�M��d�)
F�x��ԴHR*��A؊I�V�hԨGiHL� �ү�������$�<��#�5�*i"���bI��S�b Z�4�8��E�MX`XE�ʂ����Or}Fz��T�-|N~� ��UT����;�b�j��1,O.=���C�Y�zĈ�&�Tҽ��k�/LU����P�.���J��p ���L��q��i̅ ��NU>�M+�ŧZ.F��SG �N1�a�o�h�ޜ`p��� ��P�ը;���S���۳@W�!W';j*N��_�<m�7d�`CEթa�2��$�O��Gz�`@�!Hd�j1��*u64	�@� �$����i���P�ƖFyJ?�O�DN)&����)��o��#t$ \���`��ʡ�|Zc& ���B�3he�t�g�<�Xq�'��@)���}ɧ�,O�0���$W7�lx��Zˎ����Ȑ6Ȝ�8��'K�����ذvH��ΓG���Aņ�Y!���1 (^L���>��k�<YW��-j�T���OI@���jZD?�!�$0ݐ�ݹn}��0q�	z̓.���2u�Z���-9�ܜ��|n�/� �DY�◯<���o8[�`�с%M��~���%�`yf��a�=�ң?dF�0!���!�$����q��7 ��)�O�!o���M���M�#�8�M�A4O�i�<,�](#ʊ*;�^T $��1��������Y���=�̽�-�H}t�H� ���6m���MKߴ�MK�8O�!͟�	D������kEn..��Q��V~؞������{
���SGS;;�)A��\:pt`��~¢��'NΤ�}�}>m����V�����M#�b�p��5i7��4&qq�m�����A�i���q��Y�i���3�OH�n��Q-|0��CM�, ��X��S c�\�^�re$��:g��JшV���Fz�H�E����bG�b���Q@c#4Q[�4���SD�}�h��'�#=iRcݝ�]��H@N����]�f��ܛ'���>�u�Ysښ�J�*+*�ta����D-,OX���
ׁ&�}C�<d[������Y��+G�'�������-�ܔ�A�8Z���Xs�24��X����$@��ˈ��ſR��@���6k��آ�ؾ;��d�V�`$�����Q�h���+0�1Oh���#(p��j� V�o[:�1��H�9&#ţȩ}P�U�@�^�R���	^�N쁶��'Zw��x`�Ҫ\�ў�DBZ�-��i���Cz���� ���VG�v�>��5�7LO��a��h��P�c�l8���WO�<FY�M��guX�h@�xMt��т]/ ��@��g� �Ez���/Mc�N�5��x��%�Uꍨ�!�8#��z�L�:�*h
2Ƙ
q�֭pG��]:��#A���8�:TO?�$)
�'����'J����� z��ܴN�R�挰s��R�G�4��>���W(:`�@�sB�D�|�-�䱱��%�0"�y�<p�'�`)��ِPy8�Qቓ�r�Yb��$�b e�񊂱W�l���W�xR`(�@Y/(y1�'n|$��ٟ�^�M��"��X9IW(�`:�,�foN�6<p�����4R���;�O@-�uh=Z� #,�X9sĂ�Сg!rB2�┅��<�~n��5^w���r��Xn�u�Aʀ��jm�
ۓN�H�U+E�m�8�����:�z}xf�PȕRg(��iS��oZ�OO���j�7ez��[���i���#���?A�@��"�8�8x1�}�%^Nތ���Pb����/擖8jL�[���n'���Y�x�ti����%����r��A�Ċ�E�~Fz��S=N�`Њ��Jm�L�6c�TPZ�;��T-F-�)��.ؤ(�fJ���?��##}J ���Q�����¡>�090֯ ��>�T�S�7-��P+B�i��YӶ�D
5>4y�JH5"����-�L�ק���Ē�3���C�C��|+��ۃ#N~B�z�.�*>d�7-a�kq�Ɂ1����B[��< ��E'��Ozl��� P��)�{~��4�˷={���e˃�
T��ɧ��-��O���gD�|T�|Z�ԃNf�e�rA �m�Zi�� �ڟ<�`����V]����'��z3��`,h<�.�0Un0�+O��n�04I�b�"|z����e�ꀨs$F>'`R�P����qx�8�S ��<���q�m
sx�$j� <D�x��B�4���9�)D�K9�`u�:D��p���Y���%�
R�X��6D� �3��9�*���MN�Uk~��� D���YI߸\�ņ��,�2yK�(?D��l��;=��1R�L?&M �4�8D��9��g����Ae֞
7�C�,D�0���ܡw�E�jV��|"�+D��[T��	jf�s�"s1��z��*D��@U���m����G�bQ�a�'D��h�Du� :PJ�/0)b��'D�lirF��R=���H�O�(٪��:D��b�����mC3/�8�d�℅6D�t�q�PvOX��$L�?I2Px�8D� �t�ԮP�d��b�2e�L���5D����a��Q"�������O5D�왆�F�2򋍾t�e3b�?D���⣟�y}�׭�/8��)�V&3D���Q�Ր>��D���Jg���be,D�l�q+�#[�Ձ"g�v��)R�"8D�+&�ؠk�-3����;BԵA��6D��1�v���3�ϗr����2	5D�@�eE��5�8M��'�d��t%D������I{�$�a�����=D�4�鐯S�� H�'ȥB�^�r�?D�P����Mmj����'��mb@&!D�� �xcR��,:x�����
�S�}�"Od 2�M�O�<x7.Fe�����"O��`��85Ip�D�z���"O���t�ďG��(�BD��E1�"O��+A垐"��C嚝t�*AB"O؅
g�O�Bm@���#�c�~�3"O2W�V�A�5�c�B�'$| @$"O�4A��C{ĘqEC��VP��"O��`�Ä
`��5���^���Ik@"OTx��K�h�[�aPp-����"O���t�pmPoN9k��{e"O��A�/]��ɹ��Y�03#"O
�#1��E`���ь,^�e��"OhA���R�.u�u���Ջ1�A�&"O�§NL�.h����F%�"s"O�[+Z��XS�R7"���"O�I�(ؕujT�a�J��P���"O���gF�X���b�� o��"OJq���%i �z�+D�e�M�U"O�rV֖]n�)r��örc�t�B"O��lN�d<P���(#L�B�"On@c3�[AQ����=I�@S"O�����$AH���,Ć2�3�"O"YI&H@���;@�)*IL-z�"O���e�\P��̸ +L29�m�3"O���V������'7.��bW"OV��A'w������/x��5"O0͛�*ڢ'�8���)nF��k"O�%�b$C%dR�I�_.�q�E"Oܒ�l]�ڬ��(��a��+t"O�!Q�R�.�R���>���0"O(,����v]ƍ{�ʦq��H�"O�����"�L�
c� 1�F(PP"O"Y1��E��(��gC�Q����"Oy@k��,���!���k�r`�Q"O�9b"CPvR	@�g�7Z���"Od���-p��Q�a�2�%;�"O(՚"@�+>p�<��O!m�r�ʲ"O.�$���Ol�!4�ł����"O�M����UI�Qy��Y2V�NUx�"OR+gˆ�3���c�TAE��T"O\� ,D	xR�����^0H,��"O����.�|��Q����/h�� P"O�S��Q!=���k���&7�����"O1cAE�|@Ь tC� @ߞ ҅"O�u˔��$?�}*'��7)�0��5"O��b炏��@E���U�?��%�"O$�0q��&\�i��ΕBR�%"O&�ya�+'2<���B�a��I s"Ohl[�L�*G*��MW�A%u�"O�B�DW�=�65y��F ��3"O���u.@�]{�}ӹ���0�"O�QS��B)<����U�N�T�C"O$@�r&Մo��\�QE�o����D"Od�P�J0J.�!�V=.�aS1"O�izg@U�9ʠ+�.,�(��R"O�`x��O,� ��S��=^�Ds�"OR�O̺?��Y���? ���"O
\5瑠)Vΐ�a�ةN����"OT��J� �jd�  C�Wc��r"O��Y�[$��걅�_U��å��є�p=1����)TL\�K�9{KF��"��I�<���"b7��P .Y�v�y��L�<!���C�z!����,v�}��R�<� |��#�<}���X�kB�XPx 2"O�=��E��m��b�F޺!K�"O���2�C�2��(Ia�=,6���"Of��eN�2%|�pp$S�az�� "O�A����X�:,閵i��9�"O��Z��J�N��́�j��M�Aj�"O<y�l��Uhv�P����qQ&�2&"OL��e�U-��"l�tKlT"OXI3-��C6�X���@	/��2"O��J��̎f �D�_>}����"O�9S1#��	�̑3jn|��f"O�X���0=t(Pc�jI�b_^%�"O`�;VNb����F@'WD���"O��i6��)t�̡���Ξ_5h���"OP��u聿_Zft�����{�p���"OV��g�2N��x9���zrr�k�"O:t�え�tHQ�X/\���u"Ov�XĨ�3,�ц�^�`.U{0"O��@ mA�K��%�"s�<S"O�I P� e}sFC�:r���s"Of�ہ��={��`jt#_�}ô"OV�	�H�GG��P�?h�;0"O�8�6��!3�����̓!V���&"O�1@���8z6L�r��8� "OB,�d��o@���s��0x�)��"O&H��JO����9Mzp|i�"OZ�;Uoҷ_��Cp"��JmZ%0v"O��BD��/DB �_�La�"O
	�b�T�n���2Ǔ��5��"O"��d%�#YIp���%��t�-"OLX�d����
��DV�y "Oru'd��V8bk@&Y���jG"O�L��,Ԣ&,R�q *ܗ��X�&"O}��铧�60h%BՎH�x�"OʭS$W�mlZ��B���F�H�"P"O$A��O�:i���� V�F���"O�|�%c��s`�J�� E���q�"O��S3i��])��:���#�r� "OrقE�.g8��Gƞ�����"O�0���[� �k@�Hp�Ze����%�S��<B8�(��a��}(J���Ӂ}�2B��C'Ҍ�*21�~��sKԂ&\B䉒4e��k��0��k�K��m=�C�4L���@���*�ص	ah۶[C\C�	t���KR!6YפaS�?@�C�I�v�̋s�L�\�i ��̎-ŸC�	�]R��B!��$��6�^{e�C�	�T��t"1L�-Z��l�Ǆ�*O#�C�	 a4�uC�jE�e�|8DI1\5~C䉀$l�;��ľ8'���q��F_rC�	.r{�Uh���z2H�zת^�@�8C䉶^�LT+e�S�Cz���\,e�$C�ɛ�H"��O�;��X�f�G�^U�B�IoA
�)&#w����3�Y�D��B䉿!��d[�(0y7�P�vc��6/�B�ɛs�ҭ��I"'���{CV�4��B䉖p��)�ŉ��#s~���@ b�B�I�L�rc�5H����%{�.B�	�5
�E� ��
�T�3���6CAd���5y6�*�M�{���Lkc���ȓ��1&@3x�uB��@$��m�ȓx�<��bC�� ?�ZCeܵd����"�2q�ϛ��!���3%�����6� ;�m\�,�'�S*+?h���S�? @H[��-%y>�h��-T���
F"O����:Z~8�`���==����"Ol�I�{(LB�h��O�Z�Ȣ"O��D֟U�=(���6R���P'"OqPA�M!!�b����èU��@X�"O��[�O0��ah�*��V�B�#"O��iѤ@�	�n)�U��y��"O��%dd"����l�"TVm��"O�U!��L0�*��(��2G��bR"O,i�EE�~jje�vH@�2<�xe"O�1$��	m�b�ԧ�>0Ƙs�"O������-��r~�d��]�<	r���!*������M=����ŊX�<Ag
��s��#�[=��e*%P�<A���%.�-�1��,����a�<��B���J��0d
0p�h�-Q[�<�,S!:���#��?K#|����]�<a��/���2Fe����1��)� ��ȓ:�@c�   �H��wn���44�ȓE;1@�D[4%���	3�!C ��Bgƌ�w�ѿaҪq�gϿ�Ⰴ� f�XdȚ�h\X��
�<�:�<ي��	��/�\`�qR�U���)$!�d�#0�}
�F��%bX ��nąȓz��(�
�WU�pr�@�w�<��ȓi�>� s���}�Z�H�Dѧ�Ʉȓna�3m��[پ�ӯK!Sc�!��+����&�E)h�p�ˁ�o��Q��zm=u�O%tQ��g���ڌ��~�>�QL�?rB"��g��$A�$�ȓj��hRg�P�o�Ʃ�hvV�ȓpVh�A��ќǼp�a�ؖw��ȓ]%`Yh���Bk�{g!J8!�ȓ"�Z�`E��b�^��NKOA��`(�T	ކz0D�f,E$? \����4hs	J(� !���
R�.P��-,�9����i0Hёq���ȓ>aniX�/�a�d�H*�(O�t���TE��cܴDu��� �	$؅�ȓ6��l qNơ@wQi��r�>H�ȓ`��4����2u<0�����+���~��T�*Y�D`��d�܅�F����Wb�z��cϼg�*�ȓ2���!�	�U+�Re^<�6���4H΁��`ڢ7h�9P�l:o��"OX9�u&��j��IAJ���"O�ͺ������ ��� ��C"O@��bk�.��H�5�V:v64�G"ObxBAP%
z�i�l��]���s"O~X��k��A�|��w��\	�"O�����$���$C�ZkLTӡ"OT	'�ױ���``f� hl�"OT��7jt��yX%\;`"eHR"Of�0��F�pj�чF�+�us�"Oĩ@"[�^{�eR�v�V��%"O�r�Ƈi�B�ѷ��` w"Ol�Q�B7:>�Rw��N��Q"O��A�� �l�zQ+&�D�WC��"O��$ "�ҰB�&G�N���ڴ"O�!D l�j�PV�^�=�N�!�"O��j�Q8Yb:<K'�_$hHi��*O�es�&L8]ؔ��bK6�"��'lN�D��1(C�$ Sf��,xԍs	�'H�(v`,#����*�"�}�	��� ��h��Q�>�J�1׃\�'"���"O�1�	����%1�a1	�"Oʜ�b	�9\�>��"b�3a2��U"Oh|�b(F�� �d�@9"D88��"O�;�e�	{���.Y�5��"O֭@��2!4��@�Ϳvk����"O�]h,���XRa-]w�Nš�"O��
���jH��1�N=H<$�"O�m֌\�b�<I
5E�$&Q���"O�h�t��D���b�꛻�:p f"OF8(Cd��9�
�[��?A�2�I�"O��R`�V�x�pJ��ȏd��!�D"O���T�
�	G���e צj��X3"O>Y9�@�:CΨͺ�s�r\Z�"O����EJ�:G�	a�.�"���"O�9���-m�Ȱ�w@&'��"O ��v���@E�1J6Q�)�H�'"OЅ:�^"^��i{����,	�P"O<yW�]cč�O��s���U"O8X�F*�w���˔!Q����"O�uh'̀'}W
��A N�s���F"O��[+��A�8�)��P9h�x���"O�W��8��	5S�VL�"O�Tǝ+otT%�fV�H���"OXK��C�J�&ͥQ1��Ч"O�,xD��*��Te�(@�����<��O3>��4�K�u�تQ�Sb�<�q���������M��凃c�<Q�˂0
CH!#mXZ!dGND�<Q4M
<E��{CA�y�T��R�j�<�k��j۰�Ѷ�H7-[�mX7n�<d(��-�f.gu =��O�<i��>I�H�;���������G�<�t�S��K�U�b�~5�RC�<1&�Y2/�*1��A@N���LU�<A��ңC���[r�ݩ_�R��eYN�<���9����nS�Vi�����t�<�ь �Ӥ��N�Z����v��y�<F�D�/j��G�j������@�<q7�#&p�3KK���j2��f�<���
iT���ڊ8�Z8IS�_e�<��?xݾ�"���/Z��Q�i�<�b�~q̤;rƖ�Z����g�<�1.��mF�%�7�UEv��Bb�<q���_����EFըO*��0�Fw�<�0,�6.�b�I�"��((!�D��H�<��/ш%५࣑8#��m;$Ín�<��k�5Mc�P��88�X#4d�i�<a�bħU�JQ���U> �0{QO�N�<q"�J,x�X@�Rŕ?W�N��b�KQ�<�eG�V)� ����1�];a�FM�<����8h	n�Y%���z�z%+p�<I���7�V�	�9� �bЫS�<A�վ]>ܜW�R�f���O�<��.��N^����ȟ�Y+���I�<��O2(}�Q�͌1� �C�M�<�uF��a@�@e-����Ul�P�<A�K�hl���
�k:�=�"�FM�<���HQ� r'\k�p�hQ�P�<)�'#�h��ȱ`
�L�t�L�<	-�d6d�@g�.T��lJbN�G�<�MN^��J �* �\z��E�<9���!�i{�N�d/�ĪS�G�<y�I�"�<XCGŷJN�`Xb�C�)� f�����2;11FG��8 Z�"O���eAH+d��1�悇 ���0B"OT��E��Sa��"ʀX�q5"Ol�K(���ؤK���3�����"OĽʔ�Ϡ6�2i�E۸L����"Ov�)�#U)=B��c�E�آ"O�+�� 8�L"`� 2A���"O�Q�"�+4�UZѮ͓O���7"O����`��q%8	�%+�&2�U�"O�����,"���� �=A��"Ox�dJW�	>��\ᧀ�V�!�$ P�����['�w C)�!�$�r�]��G��)'D��eΝ��!�W�IU�(�_9���	$bƴe����ȓu4��1�O����.�%V�^��vƢy#��9���
=Z
����M�8�AA��%j2�ׂ�4�ȓ:�L�ȅ��i.�	4/SWH*܇ȓf	<pp��ȑf�$���l�;;�T��	��A� ^$$p�,�A� ;E���ȓb�2ɳ7���D��b�I5�L�ȓ	�͊#[3a& Q@b!��8O
���0 ⇝�0*�D�a~����܉�C>���#'���R0�t�� ����0�ׯtjiK�` �嬭�ȓBPr ���1	�r�ڴ �<{�$��C�
�r&[�*��^<��T��ytM#���#�uS��T<3��ȓYRܬ*4%K�-���h!��0]��x���D���ϊ$`�EȀi�q����ȓ	�.Y��11�>Q(R��2�*��ȓ/�� �H�e4�1�1�A�il����9��!�`92&i��$�ȓk����Q%֐_}�]tk�$�@��ȓ T�����*h��p�E	�sb��ȓT�щ�QN�4�i�AX�ȓA�p��g�
Xl��A�F�aB�؄ȓ	F(�q,xvS�.=q�.L��:�l���J�jk)�%�Ȇ�/����0���R�*�?2��ȓ	 �h���vs�5��gɆ}�bĆ�V"n	�R-%-�h:Q�K��Y�ȓB)�$q�F�2Z��Y␀_=+���ȓ~i"8��S�� Y ��H]�ȓ�Z!��T�S (��%dD>F8����W����ÓG\�(��	;:I���X�Z`��l����T��ȓ5l`˔����F*X$j�:���x|�	�Z>��`5�S��ԇȓ?�>���
O���HWT� ��w�(�� C
. ���g�E���ȓT�I�_6?P�94�Q�I�BL�ȓ6��D�b�Ƨ}4�X����x>$��ȓ>�$� �κ�5c�d¶xzA�ȓ���+3�ոU�2pC�Y�t���ȓ{�x� D:J���qԸ8E�`�ȓX�Xu�$��	3&��쑎B���S�UZ"�� �fdo�R�ȓq�DZ�o�r�j���K3^\��H�t��&�Ÿa�Qr�0q������Ӳ$q��22(�>jV���,���g;R�<���Y�L5�ȓE}P��E�*����Ց��x��vlŃ�jE!ua�-���>� x��S�? �}8p�Ю=�!�E��?N��Չ�"Oti��"�.A�ĸvdE.v���*&"O�5*��I8r���A�
F��Q1�"O�P�ud�lx�A��94�. 	�"O����6-�uߨ�F%�q"O�� �D�L�ك�Q0A����"O��˱��.A���h ̨r�"O�@�e�51GdQ�B�^�b��ȩ�"O8)Ԉ�~�rBiG9\�.�g"O�$0�H�`#����G\�v�D��"O& !r�ga�q����s��x{�"On	0��	;�+�BߑR���1&"O�����YW�2u�fB@4)	t��"O�`��d�60�R !�f�>� �"O��)���=��ժ"EN*G�|9i�"O��!��*C�Ċ��Z�]����"OV�an �4�V���ȥ���ڶ"O����!�;5L�2��I�Ny�`RB"OJ��Q�S"�#��	}�p�C"O���-�p���7늎0e�0��"O$E��,.����4j��n"���"O��j��E9ow`�Jd��4W�C*O��:ul�hV}(�ѭ!�Z=�'�d5�r ؗ(D>��������'B4�cMY{1� ���� ��ə�'O��Y�N;`���흃(&�xH�')z��a�'x�5;�	E�t�� ��'�D�i��u�]BR-ƅaO�}0�'�Ќ��m���{!K��}P�B�+r0��VHɤ2x�E�Ҙ��B�-B�� P�G�@G,�����8M��B�	�>��SDO�$���)ef�5f]�B�r#�!a`��+�%y@g�*ZS^B�6*oJ�n2#�|��f�-C�	�L�0�Ц1CJ=y���C�I Ej�!'畇Z�"��<��C�!�f<""ʉ�B�
�jaۏ��C䉱A3�La��'|�\���[�ތC�ɐ@Yj��&�Ρ(Q2�k�Η�K�!���-jxQ�G	Hm�ұ�' 
*o�!�d@z��I2�

���}2���|�!�dPn���0� k}.L�� �5iN!�D%\�6��@J	v�u3�O�6!���7g&5��!&N�<*��E.VO!�Ҝa3�Ub�ƀdJ��y)K>=3!�J^h�! ��  TG���H�>�!�$�*up�urp-��F�yc�$�0U�!�$���,�w�D !24�x"��%�!���T�t���F��R��	�k!�$fR��0v'��8�V��B�!򄆿>r.=c�ђf>��C�_!򄒅�.ٷMAxQ��p�4=W!�d��Ěd�U�Ԍ��Ǭז;W!�dC�_|V�P��N>j˸�QˇOD!�Dߢ)�8��u�C�S�V����U1!�䄢-@�8M
z�hD��E�#V�!�$J1d]̠$+?\<:���-˵r�!�$�/c2}�b	Ūj9di�m\�!�$ǵn�Q"��M:(�=aw̄�;+!���P�����9A/�@��+4bD!���@�0��U�R!*e��ꊾr\!�C<���Ɂ�\�:F�Ht�RZ!�d\4O:�(��M֮���!�T!�$�~����a*ȨT�4��զ-�!�� r���#
�8���	>e��P@"O��`�ث�%�Wgрf�>H�"ONya���z�ui�hذdL�� "Oj�ʓ%ЉVY�DㆮJtX��ca"O��U	����H�#̊0]r)��"OX
��سt��	���15�\��`"O¥#j�
�Lu"��������"O t�wJM�A�<$�����M�"O،�E.^Z�N�v�L�!�0�v"O�LRPd�:_��9��\�0�}��"Ou36�ݲs��GMI�^�[%"O�@HT�A�_faraA^)H��Q"O��2��ʮ9��p�7��*r��"O\�$���3Hz�z�Y�&�x��"O@��s�E�0=V!`Ì�q	����"O�7�)[�2d�Ta��[ʶ��"Ot��EG� ���U_X�3�"O^0�`C�5�H�УCW�*Q���"O����-[k����bH@�ǥ�y��(���6$G�lm4$��y��E�5�b��^#
�H��a�<�yaΩm�:���-o�Y�C�a��B��9W̈�AUp=F�j���4��B�I=a4�*���?	��m����X��B�	���$"�ΕZ��)"sO�$�rC�I)T[~�C5��B�jA(�/� ��C�	�=|:�q �ғg-0Ap!�֢dR�C��1-W��H�䉤O�L��ā�-U">C�I���jfBI�X�nYJ�g�s�8C�I�~��z�ʂ�|��	b����C�ɲHd2 �V�M�9|j)�1iD�\�fB䉵r���B�:B@i��B,F��Ą�p�aC�C.vsƬ� W !�G��]Yr�79i^q;���7/�!�|nR��T��0GZ���=�!�D�����1-�;72��p�R?,�!�D� 0�ɐc�
!.K��R4HS�k!���8A-�у��;Z��
4h�!�$H�$��{�
��F�����ٍ�!�$^���#�?l�m	���Z	!�$�
-��+tf�>IZ���k�|�!�d�>Wc�0NM2�}j+0?�!�/@d�,�c-ˣp&�y�kU�|�!�ԁE�����M
&�E�ꝺ�!�$^~cd9;rJ;O�.,�*�!��.:��5��E]�
�<�f	M>(4!򤎴������
4��!*Q	�=!��F�Q�Z��kN4�&��1���!���ti�&Nk:%�CB���)k}!�D'U�A&�Ȇwsn��+�xD!�䁘lҢ��fe�O��h� �R3!�D�\�`��rlB�e\���N� &?!�S�Dl�`0�cC<KFQ�1Ά6E!�$3q�0�5E�OP��sQ�{�!�$J�o��hV��8<_�%�4oB�!�	�ٮy�7�ԑ�x�(N��6�!��A�><|4z5L�g�(90,r?!�x�y� n��	*������!�V	�R�zee��~x�a��7R�!�D ��y���ĝ�H�f�̴4.!�D`�q ��J�4l�t��I!�ޚ-]��BA�<7X޼�Cn��!�рf�y�-�2OW��˔�&�!��^�T��r�o�;`SDM�w���!�� ����iɐ2i+��n����"O"Y"ՃS�L�q�&A�&D�v��f"O������@��@��Z�v`����"O�a���Ef��St�Xx}#R"O�[�.�=:n���@���J8*�*�"Ob�0��{���X���"O��AO�8!�j��с��H���{�"O`�3R&��Y`������]��"Ozi$��)�]�� �!j \�P"ODp9���TI�e�9X�m�T"O����G�*@`�k��-d�vV"O|���Ǌ1
4��_��5#����y��<��� X0�[@*�yB�!\=�B�����1N���yB�%�`|��X�X�p᪑��y*�|�>m��B�(���)6�V��yr��7ʨ��)�FA������y�/V �00#&@
\�����-�y"�1.�4�j��+�9������ybK����6��fQ���$�_��y�D��y ɨ�ɋ�LU0�G�@�yR�D-,JA4 ^�2(�X��Q��y"�X�|കJb��I��VjJ$�y�Ϙ�$�\)��@ی}�)���?�y��р �����@Vڌ���kM��yr#�:C(��� Ñi����y,jw\,�+���r�jT����yB(�z�� �tD��$x�� aC��y2#B( �h�x�d�#1��Y�e�
�yr� Ϭ	�ؼ/t�ؒ�\�y򈌈��x��#)-Lى���;�y����.�� Y���
u�ӽ�y"m�0+W�8���#�j���NO��y�� @��+q�C	"��9�.�yB��D���'��:'�<�{V\��yK̿KX���ެ$V���b�ya�/~�6eb�<"U�-[0k���y��Z�D�J0p%�ƚC�	��aW�y�e�q^b]he�q�(1��a��y�g��)76�Su��%@ �V����y��Y%���P`���<��D�%�y�!�8ib@���K�H�����	
�y�	S�0�a�M�kǆ,�`�Y��y�+@C���3mո-,�ipN���yr�I�	/U�9"~���*�4�y"�DO�"TQ�@���`n���%��\�毕� j*L��O�SQd��ʓ(�a;%��2 �P5)��%0�B�#OӞ�
A�ԛVS,QZ �x��B�I=Ӛ�Ztc�+B�*Q�'�e�B�	�gڮ	��B��N�N�j�	�'Q��B�I�E�T�%$�'$"d��%א��C�	/NPQ3ZX0H����v��Z"=D�X�HY�B���jK~ �L�#�=D�D�aFE.)�ܑ��)T�4���g�<D�\�ţZ�cÄ���o�|�� -D���]�3���E��\؞\*��+D���U���S51Xr�ؔˌtE.*D���3&+L���Ҿ��92p 'D��c�NA(_bVq�bo)I�2!*Op�����5e�t���2�B�S�"O�@)ڂL>�]�dH
�"N�y�"O04 ��2/�0�3u�ߍ{����"Ov�p"�.Z+ �j�IVMѺՒ�"O� 4�͋�p�����j�ع�D"O6s�a[�0b��P��|��%��"Or)�F�;{���h����lD�v"O(2G���*耷ASx����"O��#!z����˂H� �Y�"O�� ����ZF¹��`���B�"OHE�d(�?36D���V�*�6�:"OL�[g#	;�D��C-*j��"Oz�"$U*y00�LO 8L�1�f"OBq�@R�����1lE=C.)%"Ot�"FK,lTl(	�=Y(ԡat"O=Q΀�5�4Yeu�#g"Of5���K���y�Ko�=�s"O�q"S	���%p3� �}����c"O�q��&�$�#3�M/�6��"O����)Y�|!.ʱ�$/��1�"O�*��k�)�6��/�	�"O��R@�O�f�)�B'��`��2"O2U���MX*�PF��h�P�9�"OD\� ���$wz��+� rԎE��"O���
%o3��)�K2� 4�S"O�9s�$�5���_2C����"O�p;@�W�'+|���-[����"O؁��sPZ�3��{I"��"O�p�'�݅#t6����
)E^�&"O*�A"�֒ L	�@&nHA�"O�u����ʴx�jY�V�x]q""Odݱ�#S[I�i�e��C�"O��xU�X���r��J���E"Or5�DC޹h�n�c�&�2lo\�IC"O�l���I)��{�F@3rV,�"O�˅�'��mz�%�<�͐@"O��h'%he�"�$X�C"Oj	7͘?�x/�n�q�G2!�
�/�@�e���0b�7t !�d=}����3���R������>a!�dؤ"�45��� �dgE�<g+!�䉺A���kc���`�z]��ċZ!��:��E�J�
��&l�,a"OX� V�23}�Q���_���x#"O$L��$¹ii>��b*=K��\��"O��wO^�,j,1au
شj�\HB7"O,��I[2W�4}3S(I$:h���w"O��C� �s���M~u�&"O@|�v@J�I�>�(�ٷ0a;2"O<T@��&��I	`$F?YV]�"O^+�A�U{���G�˄^/N�"O�c@�O��49��ČP�D"O.�x�(��l]�L�W!V;�T5Q�"O��;��֢p������
��$�"O\��1�I��h�1�M�x`� "O|��!���}*D�WrL�[6"O,���6!:���J��t�P"O�ȀE��pެb��ݤwݘ9c"Oj��Y.E^���e�G�e� ��"O(��0�P�[��1e��$S���D"O$��n��-Bp!�%�6�A��"O��PL��j�:mR�$�8���[E"O�X��%á>20�0��&@�y�"O^PK����o���g�C����%"O��#�]}�����`-�=
�"O�!���(2_:��/��&�d�"O��q�.�0h���_#oUp���"O�1��G���DC%�:)>�I"O� �ʦ�[bv��Ra��7�l�4"Of�j�E�,Z�1BF A�l �"O���lǜ�.T�RIڅ"�}�S"O$X���֮tw���I	�����"O���K�URb�Ic	�8G�&�;�"O.�:��C��P��Ș~�੺w"O
�R�&˹C(~�R�]���m�a"O4U��a%��S��_�W�l%�*O	٥�9J���� �^����	�'+�u�RD�� ��V!UG<���'���PwB2Z؊ �vǆRs�0i�'f���d	H
��1��.�$X`��1�'����� �4R�%Q�-���
�'�D�C@o��h	E�Ƽ��a�
�'�.-�� �@8����S��'bt��#�I'o�IHf%�	Kg8��'?LȂe�:~��5J��J�L3�'Y+��:��Y�B�&.�f�a�'�:[6�� 6�	a�]%�����'W��� eC��(�,<T���'��5Z\�f�d-)��4=k�\�'���K�fĐ1r�aIJ��9
�'ӨEU�G�*[�����E�,0���
�'��Zv�O=o�H1ʒ��7b�Q�'�� ���*�����X+�'�
��0B
�!�i��I�x��q�'M(�jp�Z��ʀd]� ➩Q�';0<��G��J��Db�m�O���'�h1�DhAF�s����E�&Q��'?hq����'*쐍����@�
]��'�Е�B�*p�Q� D\%b�Jt�
�'$��H���T��A^�أ	�';P����Іm���R@� ]�H���'=�L!s�
YE�Ҳ�=*�V��	�'[��&��9��J�ę�2숱�'��I��HU:K(�1�h�%�f�9�'�(�r��'��
�"P�.���'�@mS7�A/{^��#��H����'h�X�OA�\(5���&L�'y�DZL�x��ŕL䘼H
�'�� B�Z�T:�04/��Y $�B	�'j����.�;���Q��J���#	�'K�u��o�f��aA�J�.���y�'�Y�QI&8yy��+-,�i�'��Ԑ��+2��y�0	�((����'r����H),<����˹ 8���'�lăэԣ-��4�ĬO8Pyrp�'�pH���_M���:G��e2
�'�8�I�mϘ�vp��fǠ;��!�'��iz�(ˈ8X��r��0:���'NT��2�RlրĘ�Ň�Vv���'t8���e҆%�>{���M�ĕ�'��xP��C�J�����!!?�t�X�'��	2d"�QE�1���$D�ZL��'òV��g@Tha�P� '���/D���E�� ^�r,�rC��0��.D�hz�JC�0�`i��S0Gԝ+�g6D�����w�"�� O����&:D��r)�J��(H&+�mby��8D�t�W%T�("f�S#I�% f2Q��k!D����lX�lR((��0B��Ջ+D��q�d֐8����ś�v��ْV*D� ����'�q��%g{��	Xt�'D��1/hѐ��ޔ��w�*D�� ��(vd�ɒ9:2�D%qg8H�Q"Oz���c̙>.B9I��[O�`2"O.a i�R��u��PB�ы�"Ovl�F��]VQ#c`Ρ!=\�cf"O�4�����K�2e��k	�"O*!�ŊL5o�9�u/H�hM�"O���F�A�2r.<A�d���yq"OhajD�Ϸ̨"�#ܯ?�^9�"Oj�!�h��iØ)��3G���"p"O�dk!>k�b���ڋK�.[u"O8e���E)�����fH�1�ʽ
Q"O"} �BC.ˑ��-s~4*s"O��F"I�-�()���M��d`b"O���Ǣ
�T�Ѐ��Q��=*�"O����\�/�^qr��w� Y�g"O4@��a�c}��"�,L�;�8*2"OhC^-�`A ��)J�lM�R"O�d�	5¤��ꃐr�D��"O�H�& <Xd��q�ؙN>p�"O��	u'�S :��R� W�fQ"O����LO\��4��=]�ډې"O�)Sac͉*�C랒K�����"O 	k2��$j��� �;&�fh2A"O��;e�v?��1!V N�~A�S"O�p
ŋY���%9D��	,���K "O��)����1.���U��j|Q�"OL]XwJ��I�)P�-j�X���"OL��aş�{��x0�`߉e�]�P"OQ�P�1Q���Oŷ��m�"O�YZ�`8�=��ӧ�T�2�"Ohu���M�s��4!S�b����"OtȐ�卼(T&X�F�W���kR"O��fO	>Lӷ�8�Z��T"O2(AE�(7�@�� L�6	�"OM�c�_��jh��A��Ah�"O�;)��"����t% � ܑ�"O�d�#��}>B4RfǶMPHV"O@L�!Q�@JJ�:gD��i� �q"O��p �ܚpG�_�t�H0;�"O��*�L1v �ՑBN�>j�,��"O�= ��Z^!U�q��b�"OdiR�)=V�(��
�, "OԠY �S,lS�kJ1��%W"OB��uC��u%��	�ׄx�I#"OX�`�ӨJT�=�dn�#s�$�"O ��7	)L����ٌ
m�Y"O�-kP
�{��u)�A[}R�xڡ"O���([�n�t����u3�u�"Ov�C��Gr6��3hV$G,
���"O΄rjY�7��A�]n�e��"O�Bb��3��3(�_�k�"Oؕ�0�	��M�&X�f�0�"O.�Z1\�>i���E="D�H�u"O�A��_�_�l=K7�\�O��l,�y��~�Si�b�0�
�c���y���;}�`���U�T���Y���y���3��ȱ�F�i貂ڻ�yR��L�9���=�T� ���yB�/#V���I:``�C�8�y���`1Ej@�*���reJ��y2gϝ�X����8���V��&�yҁ��Gc�U�$
�$t��V�Z��y,�w���hV���7��)�6�N��y�W�:�Ty+N� �LB欟��y
� �$�4�B�BL�6�T�dR�u��"O�A���# Ry��O�+J4�
�"O�<�2%��cSI!է���"L1�"O\]�`$�6D�,	�&G�3-Ԥ"5"ON��1���d�  m�� .��"Oցr��ǖ[t�ghb�"Oh����H�����d�C��]cs"O!�G�
&T
$#Y�:�j�3�"O��{ 또}��$�����:9K�"O��qN�5p���w�ٷ �v1��"O���Eb�X��	�"C�d���@�"OV|#2.� 6H�#h�2@��qZ�"O5x��	�Y8$��s'�b���4"O�5+u�Y��yv� ,��=Sv"O��g�֥1��-"E�;��̊�"Oΰ�r��|0B�:Ճ]=g��)�T"O�P��AϺxn`Yjr�W?X����"O�A��^� ��,U�0�"OZS���:���x���"O<X��D�8A8�� G���1`"O�|��
��!���Q$ �Pm��"O��F������� 3{�!( "OR�P�P�/�z����;�B4{"Oy��BV���=�7�\ X�����"O���T�����G��%�N%�y"���wU�y;0*V?<��i�"�yr,�)T��ǜ�ܬzI�6�y"#M�r�S�-BzM�,hK���y�aV �b@�N�@����(ė�y��	�~���H�.5L%���R�y2��VG�hI���&Ɛ�*LO1�y�*e�F��h��sba�ׅ��yңߚ;+LUAgb�X7�ǀEI!򄁚�q�ҏz�� ��P�?!��3S���ٵ�Q�J}�tJZ��!��	Ҕ��4�[5��2�;|!�	'0�D oˢ_��#�	<�����g�P5y�"ζKrʑhs�C��yB"R�V�^]�@��K��I��̲�y"��4�  �@`�	p�^l�1�ٶ�y��H�ۮ��A�ǡmT��FKԄ�y *��J�n�;~��)���і�ybǈ���iK⋅�^����B��y���.%|Yc"�C�VV�]������y"+�B����F�S�6��[��y2M!+�.����P�K��tX�֑�y�N�'R�9sB�4�K�,�by���d����A-����B<<|�ȓfP��aW(5^d�Ct�$�X��HL@􆃿t�P�S3Ċ"w�±��
&`(3�*A�B�Ry[Ƭ�XB܇ȓ�ؼ�D��iFN�7Ɖ%B���	b(���.����aO'�f��ȓ'9,%Qf�[�Ps���.G�����`]0�.��*����#� d�T�ȓ���ʁ�Ǣ �!�%¦s�\��ޒX"aFL�/�n����[�KӐx��"J�؛��59J�)F��ivj�ȓQ��#_�8��p��g���?)��Cqc	�w�ܺ��L�s���ȓmn�|�*�q$t��o)�x܆��p)YS+�G~
l2s�>� ��71$�B'O �z-��KھN:I��L�$)Rqg�.��!���A8�0��S�? ����b�y�""�]?.mCQ"O}�nQsx,���
2E\ڸ��"O ���b�pT2aش.#O?�|["OHM�C��FRXL@�޵gP�P"Od��s�

g��|� *]&Zl<kt"O������֬9���
ir�KS"OFI�7�F�~����aʄbI<�k�"O=��'n�tt��� <p�0 "OHEK�� iD�셦��:�"O����I
 SMx])�j{��e"OࠩC �2nz8�*WC^4��6"OfI:����0jÌ��E3��)�"O8�	�.˰0�F�rЩ�6+��Y"O�y #iر2dI[��f"O�QЗKՌz�Ȩ�&�)6�-�"OP��W�8\L��(3��3���@w"O&��'�Ky䮄��a�D�nt��"O|5���&�8�c�.�{D|��"Oɢ��C(Az��N  � 0��"O����P�T�lc2�-6�`"O�0��O"�Ec�@Ԓ\�tu�"Oؠ q�[$|�4\0��H�rĥ�"OX�SdB1|����r �[�Ν�"O��B�	��h���	�h)(v�@8A"O6 XNʺ^z4���T�yd-A�"O�Y���N�4#e!��F�["O�%���B�t:>`[�a�<
���"O�����(P5hU�v�gH�.�ybiW�^�Ⴈ)H @������y�K��*��0�R�b^z��7�y���J~"��EI�F-�}�g���y�ŐD��(�K�<��A���ڃ�yBg@C��t�V�Q�.\��a�	��y2k /j��<��b�)"h�]:��yr��z�{��0l	�(�a���yH[��y��N<f�j� ���+�y"P�d�@:�Ƃ�_E�TK�9�y�$��Y��'I�X�����\6�yBō�-�2a��@�Q�,�Ys.T�yrIW�\�D��Gc��A+�,�2��y�	\ r��K�J�:�`H��ƴ�yb�E�V��ka���/�%�&"��y��n~<�Tf[����R��y2DC�:�a�W�
ΞyC5D���y�E�px:�!��V;�X�S�JT8�y�+X�Z�����hߑD���'�(�yr���Zݦ�I!�CC��y�WL���y©��n���dْ�����P;�y2-�8,_h�PE
X�	i�"�y�n�$$���X��M�(P83��yRaB}��>5� =��(���y��N'>6��P
�/46�
�ڪ�y2���9FY����$�Z��U8�y�hM#| ���0e�0�X�*�y"!Q���x��IC�74V	�w�Q,�y2��.Si��G�0/k�����P��y��~�0 ��ʞ"N�� ��yRjS��F}ڥE :��c��y�Ҫ1h��r�^=C����D%�y�^�%�(���h\6�V�0�¿�y��^9Oqf]j��ٜ+e摁薄�y�JNᢱ���u�<��%�@��y�EA���0�"Փ��iCE-�y��)�6�b��~U,8�5aO�y
� b�g�ݕo�5�q�����D"OV�4e��3�骕'N�H�`���"O@�U+�!F}(Й�,G���T"O�ј�*I�� |j�bR5Pb�G"O�)r`�L#s����9-�ڑ+�"ODu"&Г�X䪃^�&�;A"OX��Y�r�����$�� "O���5j�c��(цԼv���c"O ��W�AdD���-b�P��"OBY�ud��wAf-ض%�/HL\s2"ONЃ�'���9�DйIV�&"O4�2��K�lDlz�D�4:$�ɀ"OB��2+W�'1��Rsc�h&�5�3"O�$���݉<�����DQt��"O���j\�v�F��$Y ��x3"O��2�c3@|�DR6`m4�"O�)�voI�\U�	��%K6��2�"OZ}[vj*8ժ)���886$ �E"O6M��gV�N����Ӣ�$.
��8"O���6"ۢh��+��җP�d!#"O���EʧU(j �I!�p5�"O���<�l�Ɇ�_?&�4�rv"Ona3pK� j3f�������Ҷ"OL��JM2*ꪝ�Dm\�Z�-��"OZ!����8�BPA���H��Q"OR5Zt@�	b���B�M�|u�Y�$"O���@%��pdHBтK'E��1�"O������.���#���wj4)�T"O� 9�>W�t �-V�1�u"O0�x���)�Z�
!/�<�Z�"O��1 \�0�]�0ǔ�4�*�"O�<RG��6�aٔg�:|ܭ{�"O�1�R!P߆%!�芏g"�l��"O΁B�����|��Ųn�h"OtUxg�͕1pXM�� F w\�1w"O��-��w
, �`F�2x��d"OV��
E t��I�]�
$i�"O���2��3`\ж� Ff�
�"O����#2�ڀ� �Ԙl*,��"OD�3��v�r@E�K~�mA�"O\���k�PD*�k�h[�)[e"O��s�h]TT��/�/[�S`"O�\��	��a���;�[�BHTs�"Or�8���Q�r���m�0!fr���"O�����\qz�|�n�(@�EÄ"O|���L2v�)ҭ�W8� �q"O�ŉ��G
�`�E�]#r�q�"O�E�Rd� q��y"�ƌ
ڀ��"O
���%_&�B]*r�_�H�G"O�(�#ū߶Q��g�F;n�c�"O��#�wA��B�	�8�p|��"O��q�ˏnY��b�ϒ"�Ju`�"OLU�g@�.I@y@�� G��r"O<���c��p�@��F`��}�F�KE"Oj����Z�L�u��"�9i"O~@xq�G� ���3�.�{&�I�"O֠��LJ<�f�a�N��_��h�"O��֛֭}1@M����E"O�Q�4�Dc�+�xЌ���"O��S��֡G�t�T-\%e���)�"O^��G\e��\;-W��4PQ�"OU�ӫ�U|�Yвm�S�^�H@"Oj�$KYFj�jdL�h� ���"ONi�噚����
H� �|EX"O� �ٰ����u�\�qdQ-r{�2 "O��JG!IrJ�{��	�Ye���B"O��%b�a(T�q*��IO譙7"O�%�b��>sY��і�Ǒ!���"O�`����,�ޭ1V莻�A�"O��c��Z $#Ei��^D6"O�i1��N����i�*jݴ�S�"O�Y���t��q����^X��"OБ���sf�$h�
33��� "O�9�p��	��L#@L�u��"O
�Zv�!j��Q��9@���"O�D��szx�.�'P+��"O^(#�S�8��]ye��=�P�"OUhҩ�&P���أ�J%6���"O��Î:�5j�(X.�Љ��"O�h�Ň���,�)�G�k�:�PV"O������nD�	�5f�j�v� �"O�uʕ랶5��ʱZ+\�j,��"Oh�0�+�7w�P�F9�XL W"O�2���"(�%� 0� �;�"OĔ�W�΃z��AR�M۝'���B�"O0����v�<@Xƚ+��H�"Oʈ�EN�3���R���]�2(�"O��g�3B�����o��(��"O��S�G{	^=+�a�*{��l!#"Oذ#�f��k!�\�#�+��P'"O�UY}�����̒S�����"Op�{7�ڠ_̸���������"O����L�uj�%��|�f5c�"O8E�`D�l�����C8sq��"O��*�i5Dw���'bL/ m
}�g"O��C��	0֑�#�աHżM��"OR9ہ��T@X��GU-|M���"OhY�fd��UAC&��/�<�s"O�ݨT#��|T4|8@Fˁ*,�c"O��R�Ĳ"�$� C��u���"O^�e�͵w e���̢���i�"O����$�2���C�6�D���"O�u ���*Q��r`�"O��( "O���"�
�*�B��"/S	ym����"OZ���F��eٕ2T8��"O\P�R�os�сTLI:^J"O��ӣJ�i�2���%�3Dj-C"Ob-z�f��[��yR���--����"O(�j���AZMH�@�7|4\q1d"O�8@QK�; �1;����F3�s�"O�T�V'Ӂ���AΜ<dv�Q�P"OIxT(F8�
x�M�U`�ͣS"O�;�h��0����.�'qyP�� "O}��H[4&��kF��b�ذ�R"O�݉bL�Rk\TA�JC4|�f�"O4u(b��$� p;F�ܿ�T��p"O$�J'�[3Yr���HK��p"O\,�X�WA���]�*"���Q"Oh| �C�1	��a��
f���H�"O@lz���FƎ��0�K$	��"O�՘�H	hJ5��(��{kx�q"O6�BuaZ�8���i��Y5j`X��"O���dO)0Z���Mׇ`�4D�f"O��u
_��0�8��� q`�Q0"Oz1+��!�p����Lp�"On��3���c��r5ڑҢ"O�)�D�(��TX'��5|(��"O���J�^&�(fO�:H��Z�"O� ��I��m�xX��޴U*���"O����_�����A��Gp����"On��҅M6`\H��:NP���"Ov�҆��{8
Etę�52B*O:Y�UiA/l<�Kт��7��
�'����fkA�d��:QlW%|�,�x	�'�X�mG	�������u|����'?� FHZ/��b�
N�}hi��'�֙cs j^`b��	������'wP��f��#��� Ј J�؈�'�R��aoOAkT�c�ה|3nY��'4�8`/:n�D��L�o���a�'�Y�%��d%< KR�B*m[���
�'�T]9��]�9$�f��5��S�'N��b��T����*���
:�"X��'�x���� "l��lX�5�A)�'�:8Ǫ�d��WC��3,1"�'�nt�Vg״s����Um[� /��	�'�v�3dA\�Zk$��3�p���'�i2�K�"b>X#/˛_��M9�'�j��W/E1	���q�D�`Dɨ�'[~Q9R R�H�P8U�ټ,��%0�':D3��\�.�a{�FT1'���	�'�m�M�)}:�s��@,5|�	�'d}b�B��Zט
c�	�(�hl��'�t�$���mg|Xxw�;�ƭ��'c������H8��'A�'΀Q��'�H[��X8s�D� 7�\�z���'Ԋ�iN��.1wG�pZp�
�'�^=�J�u��-r�Dɯ9vx��
�'Y\5����}f�{�`����	�'��9�ʍU��;T��wu��'�:D��?BYc��yI���'�+�ՀzR9X�lBn6V���'���a<S�E"��T:j)��T�<�`B#?�pI�v>b���̇j�<ёb�S~XX
���9հ̂R��c�<��F�1a&���/ԴHPN�B�_�<a#��4�P�b�%J�d���s�<) g�_P���� oݶ=�j�k�<��J?�.��pdM%d�ɑ� h�<�S���M>DeB@�.X�0p�e�<Q'��Nw�qS��y:�J���d�<)����U���;&��ã&ӀA�C�	?�x������
��A�K���C䉀0�$ei2��	|o��H%MN+%�B�I�qB��Q�L�SV�ԑ�NU�C�	]ȥ(�J����3�ƭX�ZC�Iu���w�ޘ�!@�aGB��I��I["-y���̵h%HC��(�t�q�gK�B��R��-%fC�?L|§���mDM]:P�C䉶y!���6�D&nq��S�,�vC�Id@�b�a[,6C�m�W���0m�B�I3�Z��JMXW�Q�Tj�I-lB�ɓ���aa��'��<�A$�U��C���D�Qɝ*OΜ��f�=)�C�	��"�a�M��@���iz��C�I�	p���
�*�D Te�B�I53�HE�VʚԹc�0i�B�I?Q�(Ң�1W<�;6�T,fB�(�0��&\��D��b�P=�C�O�M���\�w�H��gkETC�I$Yl,c&/ΫT��
�C�"#�B�)� :�eJ�1�
�p0�Y�o���"O���E����icqk�&Y`��A"O��P���C>L�6*�w"�ؒS"O��'B�;Dv]��I~8�m�"O�0��Q�<�p]���1m����"O��2�	+Dz�Aa�G�o�.H0"O�tI��#ҹ�,j��"Ol �d�C�N%S�땘�d��"O.��%D��l'�AC \�8�� S"ORCD.T�F<�%!�1"<*�"O�8@
�0wv�z"`��ʴ�'.�'Blm2���#{��I(�O�����'an�����?k�(��ǳv�T���zӞ�}��ֵtvz�K�i ��h9p�KR�<��͎hi~��u��M�U�1,YK�<v���&�2�h�/'����G�<����� �H&	g:�G�YB�<e��b�f����, `�B�/@D�<QP��&+�����U�&c�DY�
@�<)4��yq��> < ���v�<�`D�Ql�Y����=pN q�F�X�<$#�+���2A���l��1�U\�<Y5��-2�n��W��@�� ��BX�<��$Z�|��URC�� !w��07�T�<�$�
8I��"�*�I��IT�'Lp���=N�a�Wi"ZҨC�'���A�L�3~�yW�ӥZ�)��D4�'|�^M�D'�ZNv�(&R��ȓV�� [0�<f��x����B7@���$��)B�_O�4�J�)@�^��ه�IY�k6�����J�Zm��Nז�`���1s��!R�,|�0G,p��B���QW�۸g���j���
7���ȓx�~D�t��a���:�J��t��ȓ�HHIт�6�n�����+K,:��ȓC�b=�$e��i+�,J�,�D�H�������&��^�� Fްņȓ��i��
�-BS�$;a�o49�'��#=E�t�J�:��&L��b{N0@� ��y"�T5|��PX�*YG����"�
��'>J���L,c�������w�J��	�:�!�$��
]�H�矢)O��j̦/�!�ۢ���+@�5K����({$!�$�v/b�r�׆{^"�[`(.�!�Ē�hQ ����Í-K���3��`�!�@}��� $v:X���fL�R�!��~���M���2��+oȁ�4"O�d�D͏RkbTr#�&n���2"O�s�؀C��4���
�Q�G"O�=A��ЇS�h�ek�����"O�-��-�#\L���*� -t^�'"O,E��U�V��`��s?��R��3�S⓾j��a�.��[,�ӧ(�e����D&�X�X�`a�Z�!�i0ħ�l"L�ȓ9�Ԕ�D�M2�F���GշP|��'�#=E��e]� ;�y�\�%�B����yRH5��@0	��ib�O����'�a{ީpi�0�ぱ���)sG��yr�0;��`�Ø2�����	+�y2	ϑ��5It��VkVȒ�"B��y�a�J�1�k�b�-�s���y�D�`.iS��Pq���6-Z��0=)��VcX񘖊J�g'"�����y�?���˝,�J:R���y
� f�J�j�^W�t1 �$�����"O����F�>0�+����B�O���	��D,Dd���8((���ҩ�$�!�d��f릤�v�SJ,��_�$�!�$�	I��1�  p���֏�!�d֨'��it�>	\ �q���R�!��߬����,!,�q�D!���l�KX$#�9�㜖;!�?6u��pɍ�~�2EIsA�2�!��_�'�Н@pe�(ܚm��	{(!�Ğ�J�r]5��5\1tH1F�JC!�dѸxਗ਼�������Q:$�!�R�<�<\����L��1R%�%�!���E�J0�*Նt����#��a*�Iy��h9FO	�9�&e�0���0<O̕�?y4ܷ&��E��(zy�$Z�<�/��g����H ,=�I���V�	�HOq�X�K%�,
��*�.��a;����"O���� f��Ty�N��_"�X'"O&��n|3|����۷�n�2-���x�bI$'[��B2H��
ɣխ&�y��֒m��Y��Y�d�Z�����y�9G(���0ME���=H��y�M�*� ݀��� ���v��yb)��%�t=�!F����I����yҍ��!�J�s�d�셲�y��
a��i�*�t�A���(�yaźR�z(�
f��}�����y�������� �P�Lκ�y��R� `eZg�@����� � �yB��C�6���Y	u�1QǏ�y�Ɂ �Z�A�懌t��p#�+�yBa�=D8��-_�n����jI��y���8}�TY��PmQ �Q����yrD�
"�4Ȥ P]5�����?y�{B�O��剞]f��!��]9���
���p�C䉢R6�pi��H.S�n,���X!Cg�B�I�G�ZE�+���d	W�7��B�I�ZԴ�@�K5X��Y3�Wi8C�I�����Q�N�,�׍[�(0��I� ��"<E�D$̙(�l]����+�P�{g耕�y�X�j�*6`0ST������d[x�8� lP�p%2Hf�R�,%��
#)D�� NI3spxY�2g� g N�s�)D�PڣF�!"]`)�D�P<= �ѣE#D�H��� DTuC`P���9�'�Iz��x���	Z�\�������M�0%D��p�e�5QN=ZQ/ǎ-��A�v*(D�0j�ǚ5C��/�8yk�G�T��D ғE^����,
<Gb$�*� _�9�}��=� �Q�Br���,$r���D�V�$(R�~�{QjA�<p��ȓ�ʈ�d�{9h��/On�5��4�2(���'	wΝb��X���ȓ?�Z�AV���m��T� "��}�������ȉc  (C���f:���ȓW�K��S�Urf��a�
4Y'\��ȓ ������F�RGnR@�:|�ȓa��L�Y�2 �T±$�U��u�ȓ;��} �ݙ
������;c���� >��ї�P;Gr���,^*��\�ȓG�t׈�k�XJ��h5X��v���x	�&��i��	Ă��JV
JҒP�}Z�څ�䑅�S�? ��2��!�jY��+�<P�:�"O��W��k߸��$��4�\���"OVQ�����^A�DH� q�br""O���K��;XJ	K�G��[�r}�"O�!�7õ*%��Atg�jݼ �4"O&TKB�[��ȱq����?�����"Ol�E���	��;GX/*�nyق"Oذ���5.���˔����-bb"O������ڠ�S7Mת8�^t0�"O 8�Ɠ�JeXp��5i�(s"O�\(0�Ӆ�f1�ԩU7D�}�"O>LQU@H;D�N�(燏kMn��""On��?L^���;/3�hڠ"O4��̆�L��1 �jяZ*��'"Otu�R�u�F�0bGJ?��� "O`-2��Ȯ����倍o�*12q"O~l�Iܷ��hA�eY��)c"OT���c�~���A% 3���;�"OE0�#wP����.]|�p��"O�DB"��-&fa��AY��j�ʷ"O*	
�T:t-���ݔ~�bIa5"Ot��A� $�����ƹj0�2�"OD<�� �P�,���'ca��I�"OԨR�<
�,8�R�[$�Zm�"O|щ���
m���G��W���x�"O�A1/�+8x�a@f�RF��E��"O^$��g
���h/ C�p�a"O�ݐ��R�}%8��v��;4���k""O����7�i@w!۠r��c3"O��K�D�1���1�9+��%�"O�Q0Pg�T���I�8Jp��v"Olt��CI=��e)�"�r1"O8��DE ����4�D�oʶ5�s�Ʉ���p��5�����5Au0��-1��`w&�4Z̵��kˑM�LB��!\$v[5,FFݪ�n\��1��|x21�E¶U�� rh��\�^�ȓ� �dD�3h^��T�ƍ9p�ȓR�R���ťh���seR����ȓ�:��F�S��	s�B�"�-��u��h�6N�3Cf�5a�YҴd�� c�R��)~�������/�:���l`���sV�!��F�M�.�ȓ@��tXQA�`�x I��x�0��@/`]�r�	3(�P��aC��F%Nu�ȓ64,�����f��8ԀJ؍�ȓVw.�6�� s&�����Z j�Շȓ0�6�RA���0A����>I��ȓnS�EyV�Z$��a�1o��?�$����
�c3�]~
�`��1Z�Z��ȓc~��HR����#�+� /<��J�d�h�.C(HzE� ��L؅�-�~����'E��x�J�����ȓ4��Kӆ�!�`�  �܃/��=��93(��OF�@ZL4{A�>t�ȓv%�!�!|�R�����%��,�ȓ�x��F�8$4�rQ�N<-�hم�ej�S���2n�*���(p0���$�x�3KA�N��L�rϑ6/��݄�R<���R}R�����!sJ���+��i�S#8���%G�^E�ȓV�Y���¬-]>(B�$�ȓ5����V�G=v�¥� מRXdY�ȓf���tÓm2<�cH�7��h�ȓkԺ\IS���'�R�Y2:����S�? � �샶 ���beDJ2rI��)�"O��a�� GM�����FN`�r�"OT�ȶi�4u�ږ҅7�݊�"Op "EgB�sFҭZ����2Z��i�"O�`$�<vU�r�W@(�Z�"Oj����E)զ ��$+Q�Pa��"O��r�
C6o|�ܓt� P6)�p"O��!W�R~j8Pr�$H�`"O�:�Ssq�toW�:I�0��"On�i�'9���3�)L&~ �"O�TfA��h�&�iE��?��c"O��Ck��n+�5�e�� '^��E"OP%Cf��(xB�HQ���m^@�"O����AI�hK��Y��� Q���s"O�9�V�HN@��@(C����f"O|��Z����3���W۸16"O��婅�V8�N�2ض����'����)5B��`34��M�2\��-���Y3�N��p?��I�2> ࠒ��^ �� ��'��ɰ���$��B8��'��c>�K�Ç$#EX���I�w�<9��L>h�:L�Ɔ��Z���ņ��H;��R45�p�r�/4W��T�Q��!D�#�%b���W�<ᡌ)6�D[Ղ��Y�1���D�z��i�\�Qǡ_�(?(�Yϟ����'��e\,�e�
*�L��"
%�ON��B��t ���
.Ơ��T?Xt0塐<zw�Ă�ڻA��|BᜩIӚ���b�4KPH�*D�R��hO\jS6#����������ҟ�qG,��I�����W{V��"OtP�E�
�%lڸ��MܝN��yw�'Ʀ�aRƌ(\���Q1��s�x@ȍ����q�pRA�L�#�$]:�%�O*C�	�Jz 8!I�V�)�SG��T_$��A���  Z�HQ�9z00�|Fy��WD2�w���>���p���<�?qUd�:q���=}��ĀIz�t{�Δ��X�BڣQe����	�7�p!�.�-
�|$5�I�	F��P�5|e��' 6@�p"�`���3�=��,���(�ePV�Z?���B(:rM�&E��[q���@R�$kדa��4���$��H8%�=+G
Q��ɇ�VU薅?(z@e#� \�t#(-{�<�#C#R�Y1r���<)DU�S�ֳf���"��~?*�r��)�	<"�R�*��8Rb!S��J|%�P%?�h% �6_��x��
wb c��ĎS	��S��J�d���P��G�pUV�``�?7\Q��(�'�Z�� �b�/Dxd`�Q�a{<Q�U!J�v#��
 DG�Dk��R��5 Ȏ����̎�n���0�Nߠ8�����V3-r���k�v����-|O��u��1o�n� ��Ł5�x�Z��ȄRP� ˶
�UrL4�hV�C�D E�ͱh�r���E�4�`�*`�SQ�N�1>,�RT
��]��5�%JA���x�+Q(G�f�3F`ת �`p;�,��.���j@���@SH٣�Ω#�V���
� ��`1DeT�Yg��l��*���J`�~*EYVf7M�-�Za�*�<尿�`��-��,6|�Q;��ɝWP��SŒ('c@�2�'ݵ��i˦=�ͰWj6(�Г7�[p:����~�BH˒j@�{����`gC�8������X���\��Ϟ<��r���:�Q�ȈZ�����GDt��_?��7��t���|����/F<Z�\	 �藰;@�t*����h�jԃ��U ��=�#��y��)h$#C�5�!A��Mw߈���� C?, �AّrV�X���)ۄ-p�cB3�)wL qӞ��b-Y��+рY���	��Ò�愚�l�'�� A
ea&!���+.�R�Ba���K�b��iH�!8u�T���m����-�\��h1 ��ON�Fj�N�l���?O2a!��'r�S�bӸt�
L�r�O�`���ܙc���e���P����1`�I<r!��'S��a��]�~.�hV+� er5�ߛpu��B���p=��½
C���m�5"DKںgR4���ݳ4Hh����E����O䎝!B���>��UM\1/���*9��ɉ�ϚB��,2"1�O��x\� �ǁV��{@F��c��Ā�&��U�` u��2m�	cF�J?d�]eǃS��)��0g��ذӦ_���T��:P-�u���	�QZ�$5ߨO$���#0[��t���ѧ0F�L�%��}�e blFp�T[��)����@�$�h�!W���@�7�$�6b>�'.���/WQ̐7��-S���'2v�����;6[p���ŏ�`cVcW�)gq���i� �v�Jucf��%M\��$*$Y�MԶd�Q*	ۓm�����M��KP5�9񰀊5NX\����mG�9��C_���ێ[�c�?"d���dv݈FaS=P~�̊׉V�D�x��I1X��	��A�`� `F)B�)�Д���H� �qv�Ôe�.�RIM���ܘ�n�f��R3�'9��s��&WΌ	��J1g�>�F}��_�)jA9�v�4Kj��*wA×7N�둥<\�|d  �(r0tq��$4�g?!&���6TN�P��f��� *\?�B�F�����柃Tz�0+�	[�π R��
�7>\s�m	�X4	+�"O���ሏ�t{�abKZ� dX��
��y���$�t��b^�g���x,�MC��hM����rdt���_:LT�ad�%���:%T;D["��ΔR_��#BJ,UyR�s�e"|O^}�P�H06��aCC�Ѡ-���I��0X�H�q>*8q�-~YZ�	K��1"�l�$v4I��5&!�[�L��'�d���91�����$_>2��[��
f:�����K$�>��+�ґ+��2Tj|�� �0D���T��H�$ �7EVE �BY�9|V��J~d[�Ĕ�#����'P��;��B�ʐ�����Z�����~]i'OYb���MG�v@i0�#�<�Xk��b@��F��D"v��6�<��$���/4�E�0�cp= lүH����`Y�"h���Y2 q�b���P�".���"O��sE�^7�&@�n{��ON励�I6�L�`H٠J��!����M�(����t���p���P�DB�ɚ-k��G["]�m(Dg�.�R���M2Cx�!Z��F~��r��-j��ۢ\�y`�W��nܻr�sDJǅm�v�QE�R��~�唲r�b�!����*��0���%�.����&��郪�p�h9b:)��8��P`P��'(�p��r�2E�!ۧn[�"�
�G~�+]���B���'-��u��E�S)��쓭9�r} ��b6��W����u�u'Я���R7�CG���DڦKn�O��8��iC��V�D,�	>$�Ljv�(]����IR ���2V��9ZQ����0Ȳ��	 ��H�ǉ2PS� ka��/<�� ��*�O�	��� 7F�I�Ȍ�;�hh`� ��2��߁!��H>8�~X G@Y!&R�C�C�p����#h�p��"
�x���."q��3έQU�r���PH7�(�d �"G�,���r�Z(�� �
L���EHq膱H��K����]����{L�)�N'�6�(�o:�-y�λF�. ��(�"��4DNH<)4�D;Ckr���*̒!�V��D�BrV�KD���z��q�O&���"��F��9x�@�v�,�9V�=6��'	�݋��Y�"�>x�@��1m
��3L�]� A� g��Id(ڙ'��y6��F���!���C���!2�@d��lS$�I�<�C�N99yT����(K�l�q�C#<{�����MU�R6�l8��t}�k<V�:�(ӮD~��g녱q���;f	Y*O�u
g8�X��I�X(���t%��L\10�I���8�B4L]\�( ���NEF6h�T%�FlI Oɢ��I�U/{��P��B8�!5OE(L9G2#@�BT�h�d��"m8�����j1"ߴC��S�bU�oLV�ȠjJ*/�ic�Ȏ�+Ni�Ą	��$Bߵ@���1hCH�OS�A�Ҩ�� a�Ǭ��F&X��'�^�t�C�b�nJ��%*֨d�O�%%�P�S�*y��%��SѠC1#� e��8�BG���@���<�5*F�H��0HA�LO�'�4`H��#b^+�)H��B�*1�	�:$(��eb��f�,$p��ӓ�<гb�]-�9X��o�Ȑ1�^3Y62D؀
�8� �Ze�HW�1��I�S��0��#v2�q`e!ߍ$�hI��(?�U gØW���Hcp���t0�i��#�dA�O=�M8��C�	�,��M��JVVʘW���D}r�B�H��P�w�ؠ1u���:@HG-cjH�"�����Q)�1�n�z���,@��ba+���8!��- edl��$�(���)�ɳ�88�L�sQ�`��2���;A+�����/P�6�*��U�\��Bf'�~��i̯a�T�r U�>c��#b��I�^t�to�h�����%)N��J��T���,Rl��G}��S5�9�J �CDt��̱A���a��<�  	4dֽL��<+�i�T:��S��GLxᣬ�����x*��W >��qk��:4���!J؞$11g���������}�i����wH��+f垽:.h"����0�W��:dY���� �X��l���De<9'n�Y'G/t����ᇈ14�� Q��tu|����(h�@�H��l���&"	�y���M�(Mk1)��&ߜEzb ޅX��@�d�Ҵ��!B�O�a���̗K�0a3�II�~��D[m�T�R뉡'��<X��ݏ�~��ʕYH-��A�ƳN!r�b����*�`�s4�EjA㗫`����Bz�̩�Ė=yGl�bF`
�4��q��LCv���$�)dQ� *T�ۺ	�Tـ�G��؆,�Rl�!Aⲵ��u��7�[�GV��BĈ�5q���q͏�x;�=9�%٭E��Usv�
?�,;��ΕH���P��ϥb�ε�#*�O*�'nE��>��q#�+|՚d��l��-�0� �?6���mɧ9�z��*�� �Ӂ�ΨyЖt��ܟ\����0Iա8�0�#��t�F���'��q�e��M���B�>��)�����K�=\� `B�ՅX�,���Q)J����EK�%bTM��[�DM����Y  �O,P��ءF|��z�%F�o���L<��hˌu��5 iGAܧn���� �D�*�����+�Bh�a#����(ɷ�B�?���R��0�P
��Γ~.�?�OC��\� ��ڢ#0��:���F�'F���k��~RdF<[c��`���\|��Y��C/n�J�s��ѶU���S��	��xRNC(`�t� /�6+<����(Ozd�r�(a�p� �^ܧ��z�-�*HT��aWO�@A�ȓJ�8�bG�c��e��KO>�%�ȓ)����0�	1?c�Բ��C�䜇ȓwu �7%S�A���*�k�y�n��S�? V�*�V*f6����(�.q�0\��"O���H�Q��a�w��/m�Ȕ �"Ohء��-f�X��@�]Q["x��"O1���D�}/����[Խx�"O��9���G�Bm�Ub^�EJ�h�"O�X����tO
dR�
�x%�A�"O��sg?�p ��#$1Y�"O�=����j��`a�:3N�S�"Oj��A�N~M8��ӈ��!�"O�| U�34�P e��`��8�g"O���#DD\�&��eL@ �Lc "O�KuK�<�� ��mI�U�P�B"O���I�#b����8Rh�$��"O�m�Q����B
I�R�9q"O
H�N�%"G�֙?l��ZD"O��d��Q����I"�ty�u"O�u 1�=�(1��YK�F,h�"O�	����8i b��S��s�"!SG"OR��W�Q�QW<�r4`��`�d�s3"O΅bL&Y�@�naȑ��"O�Ekb�� 1n��<	ef̚#"Ob AB�Ս9�q����2pk>�2�"O���舁B'Z0�C��4?H�=�"Oؕ�v��5o��ѓ�ԏxN�dJ�"O*YP*/d ��{#m0["�x�"O�푣�¿rb�$�G~��:f"O6�[s��-�*B�a�t���"O�Y �@��`W`��M
6�F��w"Ou#��P�;�,r�I���jC"O\ �6M�7t�哕�L/��b�"Ox����7$ښ1�� �w� �0"O�%PEF|T�7i^$�D��"O��a�CדM�:��r����j�T"Oz]����<8���ǁߪ`|��+�"O�$�p
�t��pB��=6e���"O��k���:��b��Vx$��aC"OD9��M�='P☢�lW,# %Z�"O�I�U��4\�D|[�l	�Hv ���"O8P���{7��HG�͇l��
t"O�-��gQ
m>RDc��ѩ�:���"O����X+g�|abd)����"O�	�t��&^NT�X#��Ϧ�)5"Oz1��FF-Zgxu���a�y�4"Oz`���D�
~�%bG��_���*v"OLD��툔9��*�n�%`�V��d"Ov�seɛ�$�x4À
��"�"O\���#تĀ����.���"Of���(!p�ڤ�Z�`z��"O�9�7G��*�<��&˭%g�d��"O2��Tn�@��%�R &���d"O4t�fE�)l>:q��QD0�|�v"O���5/'Nv=����"^�d,�&"O�[�'��.�t�i��O,"��s"Ov-y  �7?f�飍Z�
jE�0"O�y�u�5~B�2��/ ���"ONx�g��3[x@#b�%"�4 �"O�<��@�*L����1��t�tr"Otы�n�??1��9�+9x[��3�"O�a;q�A7m��-�5)�lF@�2B"OE	�FE�f��KCG��|<.�Y&"O��a*-\����G�Z� �"O~�))M��k�C�>[Z�ūw"O��#�A�5a��i�D�p5v8�b"O���BL�K֦*f!�:*�ʤ"O� 8a""ƴWn��I�/R����"O���wMͲW��4��j��ص"Of���A�4��l���V��X&"OJ|A��*;�tz�ꂎ�:d��"O`QQ���/�D[%D��b<�6"O���B�6%7���ȃ3�-�!"O�=i��˾T"�X�EO�_$�yYc"O\�F�T�B���*�Mx�M�2"O��:Ňݍby\���j��Bhd���"O�ͪb@�&s�1�kB&{p�Z3"OԵ��gN�c�����d�� �"O�ԃ��C���JQ̘�j�6 �g"OzŁ��P:��$��]r�ج�"OJ���˽2mf��EW�NQ:�X�"O��&��
"���D�M�)2�"O�Zq ܥ>�����s�,�Q""O�m�V@������XZ�#�"O�D20�� VH0�+�0y,!�!"O�)!�ϭ?������J����p"O�m�`�ʧ��@�@�Yaz�"O�M��o�>r��l0�%^%pV �i7�'��E�Տ��P�m)Aa��sH$��6��?�<��!��p?1QlL.i�8#�@�M�$�ӮTo�'atEC�DA3b|�Pd9�w�_�q�|���Z�Q	maq(P�<!�Ͻy(P$	��2),ళ�Mz?Q��	�s���x�/jԙF��Cw���q�B�Ol�l2�E�y�GD,:Sd�9���W�yj�j�=l}J܂f��uᖊ�L�^���?#<�����T�ڇ�sp��oInx�t�ԯ�/kT�$y���"������>�R��H%3xZ�b�oX�:�����M98�p؉ZX
@�e'Ua�ўh���S)J-[����z�a�`�?�{���2Y]<��R��0"��I��.D���E�W`����/��Y�#��Op	Au�K�N�6��͟�;��:��./~����])}i-ҳ�	�}\BԄ�g�H<󄩘�% ��0 �Z����2L��!yB�ʝ��ei�|���P�~P��1t��&j`��bb�teB�e�� �i��ħ �<�$�K�9��P�G�b�䡹�'Ѻ9f�	����@(t�	��'�v�qb��=L��\:!���O�� ��9Z��G7��i�ĉ�-d�˅��t���0�4���AD�h�2��(]�j��$Q)���s�W�Y`�в�ߔv4 p��ΝdN�`��޸m��Ai��6J���1D�%&D��ㆪ���h���0�J(3����
$=N-#��8扙%>F=�؎�ڜ
�A�:j��%?��GQ0v���Rg'�늭X���TpCW�.vq`t�g�	fV�g�'�d|��,�lol`;���(b<�3�F�Ġ��f�G4I�񸲀���OR�h��]j9P�!�A�6A�|����W�|��� gT�@Stl����=iQA�/|����K�w<�&	����w�ΐj���#��B�d�zh����|��(���˺v8�r�/G�
��஻S�>h[@,]_��s���"��T��1uMp�"@��Z����I�*	�T�k���`̎���\)�vx2�"�?��!�H��ĉ���G&p/D�o�H��]"vb�|�H4+�n��@����d��;F׀�K1��=M�P0Kpo�M�j�3L|�S��x�F26J��TXBb�\�5���<	@+/�)1��!��B S�(��2/�s��@��'x	(�2Q"�$���Hw��tCFQ�O~"ǪюwGBY�w�S��|�˒&��;$�}[� R.b�bh�J�.mtE���T�W�W$Q^8@S�V� |6�"Ng�`aJ5e·�~�s2��t��0Hv���TR$t;P�8&q(�B�O�DpA �g�0���hT�J��8�:�H-R=)��9uMՂ:�q(�@B-4d)k��b	Ҳ�\�N�bx�邔��1����&���Qԫ�N���Q
�Q�>��"_`0P����U����%�M�����¦Ix�$>)���O~�*�0
?
��9��/D����k��jUR1≘?W��{ [�����E'���k��[?1��OD4	˷�K���ɳA
��Sr�U��$���k�/*J�~�
%���1*訹�d��.V�" B/�4%�R[�L�.�*��_�P$L��ɰ��$�q+M�]8!j����:�T�>�׏����x�u�Q!sQ.I���1|��T�Ui��FȾ�*���w����t���\���$Z�:�� '�!+
.x�GG9�D�;�u9�!�;7,�!`G�,P��x���0��n�L�@4����h6�0�C�	�D�8���)r�m�a
�&ae�5m��Eh�JP�'��Uj�f:���{̓9}ЈA2����D#���&$\͆��U����� Z�ࢍ��w"2@��L�E��9A�Ԏ)��D1W��?̀�Pד
R� Ϛ9Ĥ��̕�`�F}�@ū�;�����Ni2��)��pIőE��B���$b����m�<�U@�?�)�g�ǜk��M#r�n?��=6�p�v�[n$`�p��G�O��y�v��+��PI&ő�sT�ɠ�'�n x" �_JZ9�.ֆo:���H"�Xڅ�U�P�pA�����3�ɡgG��q� :��m�aȞ<�����ǧh��1�oǥ(L��o�}���R�	l�h`�2�2t��	���')X�+��=%^-��b�=pvpd+���E�1�J����"(�[��Ƿ`+���Ɗ�@�6��6��r�!�y���:���;aԾ{�!���~��]�(��9��h�_�ri�&JS�h�x��#��!�U��9FZ�S�"O�u��n�;�Fe��I"%MJ%�ŉ�4�4���-�&h��
D�\��g�K�]�B(>Tdά��v�0��I��"�3��=����� C�'��5;��H1^c>��˹- �H��9|O��걯	7d�8��m��"ץa�'�r�SңL�(���;�KJ�vZ��'S@ZU��O�P��6��:K*e�ȓ/N�C��ʶ�8�� jǋgfr�VS���v�V4@[S��
!�)E���]�v�TI�EЎw5f���M��y2�����#CL/:��H���	�D9q'�>=3����.H#���0�͖}��#�9��ԧyѹ��t���Q�h4��\D���:W!�9@�F5�aΊ#�R������:Dd0;�b�K��hx�X�ۜg�f�ɖB/~�RW�OS��ep�	a@��z���Ȕ�݂8�b"?鳫̉ �R��-�$h��$��=�mö$Ҏ�p�aK�s� �M�{�261K4t����'۸�g�'��9CA�H�iӢ=* ��1((T*+O�]�����xڔ���=x�V���
�a!A��}�8s���N)����O@Ox�9#0 4t��bN�qka}��7n8""fF��TԉA��7�@A��� `d��*�2avdCC�*j�b�R�7����@N̙�҈�Ī7���؆'ʣH/��*@�SHE������HA⇗o~r B`F�(}���.�(fP��� j�lLt���9тFjrn$
��)��)�(��� �	�1E��ȇ_'n|�\���Č&G@�8�b�ޑ{���))��?��`C�E�x������S%ۭd 8|x4��'Ig�m�a)�)?X��S�Z	2]3-#��I�t�2�@��*piƝ��ߠL��I:,�΁A�晑x�(9#��ݼ�����&�IB&Ė9|��3A�M(pGI⢫��f��\��(A�iȠ:�P�-���H�,,O��b�!ĦBVA����<e�i�Ꙭ@Pp�a$u�p\���)5V�u��J:�����v�$Â�T�Z�>H�Po��G���@�3&LY``,�%�a~����x�6���N�!f�D��Q����+҈;�d!��N�b|aUːJ�0����א#x֏(��i�9��$�q�׀U�I:� �\���C��I�_\Q���� �h��W�&�J��:g0�Ф�2�>�
 ��23R ��f�
O(&a@���/mƁ�S!;c���� ����Cy���"5����UH��{!����K~	�'xp"Q��~5����� i���O�D�ˑgV�T5a#T�_<0ؼl�A:݆���^�,+��{s-
�N��� �	,+��)��B��'��0��c�u��q����f�M`�jI�96H�p7�ؗ=y^x3F,�4���#�E�r��A�cD�e� ]p�*	�9�5�%
#{����F�]x� Xp�B[�4��	� |�hE��X�cmUV@��IU��y�H@k�	�*1�Z�9��S��l�W�E���)QC��A�O�@XS!�@�2G�/�Q�*���.�Q����x�q�HӟV7��"�����.��$j��Ad�a�����G@E�~!	�!F$%�)1�Ov�)�
�Fz�	Z֜�rn�8K�B�cYB�ʕb;��f����-�.�$�Q�4B�-�O�z���$@�օY�A�@ Oҧ4�����M�(�y�@ق�:A23ψ�X ���b����O�8�������I� 򬵰��L�I
�LQaI	��$PЯ	o���� ͖����I����sӒ\����*�D�AF��\ߜPa��L|�}�
�Ӗ��0	<b�|b5�qr����iٵG��{@&V�&A@���	��i$g�<c�tr�w}����9���Kf.Av����3'�����gC���>i�a1l��+�؞>s��	$K	�?U�g��\g��sြ%����F�}=������<
�[2�h]H���_` ���A�? �����O<�i�62/(a0�^K|(@�u�O��Y�	M�H|��!����ؐ$Y?I��"�h��g�I�*��g"��R�$)AÀu�����ý~/4�Ae�ӡ9*88�_<M�8�>yC�^��5Z#��
3��(zL84S�9@1���=@!��F�D�	w��? '��SĦ�e\514��vd��B��x�"�#�_;�2T�C+	o*(�'Jn�pK��<"�q;��
���ѡ�<5�`�7��	�i���cC�%�MC ���ɇ��$$!m5��#S���0�L5C�MPMbXu:Ó;~���%*�l�d
�Z�ܸv�S>=�V���I43���:��،hP2���
�8I�@#�LN�P���U���q��ژdvd��'��\��NКVk��;�A �>f*��J�`�W  K�\H�4�%?e"��Rj�x^@��q�¢�V�3�ߕ7�nЙ�E�"8ꐩU>p��EI�H\џXA�/رx�~4��O�0�$�(ړ"W�V�c?a���$���� _1 ���+�%B0Y�<U;6��|��t"rN}<�� �5���"��&����/ I�'� ���@4���;�3� ��@�$�*.~���1/�"h��$��"Ox�æ��"j�$kЄ�?en8C�"O 9q�oM�$�8�6�[Rʐ�"O��	�kƒL���`b�GB&,�F"O�h�E�Z3`�~�� �6G�@"O�%83�2�p��mi�i�s"O���FA;5�@y� ��R\%ZR"O��0cޠs�FX��I�:���c3"O�A�	M�j�$i�U�G�v0��"O�����ɾQwKբ��	�l�5�y�A���0@��<ڦt�����yrn[�>1Z]��*�.�`rD�ŷ�yBe�V���$B&rג�Q�Z7�yb�t�)��ܑvo����y"��4����R:{�X�Ť�.�y�/�Sm��7c����怯�y"*��C��i��O�B�f��Ɠ�y��O$������8Ov�@ǡ�*�y�K�j!�傻4�v)��L��y��J�WF
�0�E�����)&�y�m�HT��tF$`�b�y��(_�p�ѕ�ܟt�օ��A;�yr��z�4aˠ�x���E���yBM͔=KzX�vu�a����6�y"�UBDjS"�c9�|QaB��yrō4����@j*��7�@�`j!��Zvň���aY�y��-2]!�D�.|�Y�h�aYDuINQC!��"]4:���<HA��!��<fK!�$'��\2��H�N;�ؗ"׸=2!򤉐2.REز�3l\�ؚѫɉM!�J��� �%G�e�j�4<!�d�)��J AU�[V c�I]5W!�Q?b��t�e��^����/�� _!��O;n�t�j���B���	4"&8!�$ �=y�aQ�B��D����tLˏ`:!��Z��v�&����e��yR��(Ba`=�@n\<N�<ҴcO��yb��1T�,�I�Չ�U%�yү��FlhՁ(�&D��n���yrֈ|�p��#�7��\ش葟��O��bb�	�d�[f��3OR҇F�$s/<<��C:<������'��P㗪о4�$P������cs%�'Bc�	�r�%J�	]ڵ��S!1ǆU��R�	�g}��i����W�4� С�ׅ2���!�L�}TE+�{*�B�?�"TD�>Z�ЪE��8��A2-G�B�BP�y�~ڊ�����b��*�	��=<��<�.Ƚa�@�Zx p�%AҧZ�<14�@��O�tprH�ē��Y�<BC�܉!���!���[ �Ya亟Q$߈	�ئO�#~j�Kٙb1 ��c�˟\�P�f@	���!#P8>w�ҧ�� � �,�(��}�I7@Y?�X	`�|"�O��i�i����5u������_y׸M�U��V���<���^I��?�u��5�����d(�c��,x[F�p�雁�M۟'aNܑO�ϛv�]gy��i��u�D��Lܚݫ�k�`��7m@fL�ԍ��j���S�n��'�Ȩ���l�\�١��#z����
�j��6-�K}
�'@j�� Eċ�x[d�I�|���*QD��(O&e��S>ӧ���,Le������L��@W1=
j�&�H��`�=Q>�O��	h��
<b��)���� q���O��[������%��O��d�)!�2��3�7}Fh n�7_�f�n�z|��V������S�O��D����D�T���-b��T�$)Ъ\B$jE`�S�3��Ou�qwN�$k\���Њ`p�U�F'^�q��L&�����S\�ԁY�ޱ	tȗ/DCƀX���e��%��	��K�
��t����?��#��Y`4=���P8?�0&�O5��Pp��~��1���pF�*��j2@J3�~�.�<L<I��d�������D�K'v,b�G20��,%��P,O��Mk��|� ��a��d2 c#D_� �	:w�|2d�0���	�+��jԯ�9Ln᳣�1e��C�I���4�$�X��ʑ�w �C��=qM�8�r�e %�5�S�	v�C�	/.�
\�7H�z7�9c �l�B�I�<��!�� �( ��4!�M�{�nC䉪(�{iާm4��[�KT��B䉿?�i6_0����$Kh(C��KDI�d�K�J!�Ez'j�C`$C�I~�ثu�F�v4l��E�'`$�C�	�u]R�a��H�"m�i@C��!qVB�	z���s��߿&"�{�g�vp
B�	#d�8�7�](���(�m�+& C�I�&[�ٷ���G(�����4A�B�I�z��hr��	�Z(Q��14�B�	-e�����8V�d�ڣ1,B�ɹ/��8���[8�'ge�C�	�;m ��T�N=k�(�UdإSZPB�	003�}r�jEP�^� AH��E�B�	eO��j���u�P�heNа �B�ɱZrM`v��<TT�R���AL�B�	xG��#��!;�ڰ�S� 54�B�I|�ʔ{�Z"0{l`G�c��C�I,���"2��%n���c�*��C䉕�l��%�ȧ?T���1lA�'��C�	;1@�,�A��o�%	r퓙f}�C�ɴ. � ��ۢyX��9�����C�� ]愭�ӀY5�r�5!�r�B�I�8���S@NM�ml0!�'4��B�	Z�tyc��ȶu.!R���"h��B�ɥV-F��db֑l����v��;��B䉢T=�鈢��$1�|���̕wfB�Ʉ�f�գ�tOzeKR���'I@B�<PQ��ǂ��T�v)�D�*�xB�I�1׆-�fa�'hR��!Z�H�DB�I�nG0�	��W.t"*53*B�*jC�I�^@�bF
?.@��	��7C�	�/�Z񋣌�P�$��î�&pNB�I!lD�����W��5���R�M�.B��g|L�biA�m���3��]�S% B��?FDRE��l�`�XEj�H���M�ȓ
�"U
�`.j���ۊ0��1����[2��	0��8�2N�+��m��\�"�i��+G�q1��κx@X�����Q�e��zڅ �.�SZ�ȓ�v�{Æ�12�)@��4j��ȓ�l�pF�>>v�Y�/��h&ʴ�ȓK2`�l���[�-֍�-��E���zUO�(V���T�Fjh0�ȓc��E�n��v�0Ҩ��~U�̄�M�n��F�m���ա���H�ȓK��I���:@�n�TH56)t݆ȓ$����Rˁn`�8u�/CZ8��u�VŠǣض/̀x�oŀ*n��ȓam`�W�ڀ3>(�	;(g�ȇȓؘ XG�I�u��s��O7'_�Ʌ�xvC�f�!l��,̴%\A�ȓJ
�	Rt�J�>���[���.#La�ȓ G���Nb��=� Lԧ)�ԅ����z�N�(���)���dH�ȓP+�\#���X��BQ��	\34�ȓZ�ޘ2C�#=l���@�^����e4�E�؋7ɤ�2����Նȓ+�p��F��}5"ybRG��f���S�? ���!X��x���<��"Oj�R��-��P��@�,�����"OZM[�M
*M��eJ oبm����'"O]�f���҉pchO��A0�"O�`���̬}b˷Fի����"O�"G	o5J鑅�4���!!"O;��4,J��� #��y�z�"O��i3�?
@�@3��.fj���"O2�8�(ܘw��X���Rr��"O� Y�)�'iʠ�
"
�,U��"Oz��d*� 6H�{�P`��"O�!ZS��#l"���HߩZ���b1"O��@��@1� �N�^@�"ONb�c�W=�� ��*���i@"Or�3��GR�疣`�l�X�"O�E�0AP[~��X�W %���YF"O��1�N� ����%аM���p�"OTm�%ɖ3r�
Y��X�e(�TB"O��&�J�bsF"4����@iV"O�Lqg��Z_NP�6��#C�v�"O����J�%�qde��0��"O�0kפ�f}\�3w��-TD��"O�P�^�H�X쩅�Z;�DA�A"O��8pG�gj(<�@Z+'Pf%H&"O��ᕩQ?W�����>,<>�s�"O���t�Ǎ\���B�B[:��b"O>�@���� ���y�T�F"O0����&��a�����C"O&��N�^�(�.)����
�y��H�y��Aa�J�5�4Y���M��y2A�	"�%� LЃ3���ŉ���y P�0�F�8łU�W���z&`E��y��Η��|3v_T�`t;&��y�^d�<�	Y�5}d�V���yB�̖[{^h��>5�u�en�3�yR'�rr��a@D�;�H�� �y�R�-e�qq���2*:��U�-�y2���M���b����:]{�b^��y�D�%I��*���D�&�y��ZW�0�'���\��$h��y�9DT��R�d��$�� ��y�&��x-�%M��"����ݰ�y�@��z%Jeٍ�. J�]��y��:R̄ja��=Ͱ�s�e_�ybd���UiJ�|Dx�R�ߨ�yҮ��DD�E�s��Nj���T��y���(f�p�❇:� a됁�yR`Tb"rĎ�|��eBЊ *�y҇�S`��2��{�f�`(��y�hZ�f�����}��&���y�@f���bU�%z�*�)��y"˘�R���S�| !O��Y{�-���Dt�w��:\0�����$I-����KV�w`|	cuȞ?��ȓT�!������jF!4�����'j� 0� 8���c�/6��<H�'�1��$P�t�#/�G����'՞M��o�&�!�dQC���'.����ada��mՏgJ��
�'��Գc�+U����) #[��(��'SF�s3(7�D�P�Y�V�����'l��RI�&j��ʷn^9w�\���'�(���R�b��l�2'XX�fِ�'^���'.J� ^pɹ�	��`��
��� ���p��h���é��\:�"O�͉��܆��Q�(�0$���3"O(�G
y �=�q�U�$���"O|��&��4����QÞ�3�<��w"O�����O�c&�ȕ�FGu�\	�"O~L1����<t��ޅfh��!"O� Å�Q��XU�	����"O��d S�{�M�㦋�����"Ox4 �.S�L��q�QF�	E��IE"O��[��B22K����$��
�� +E"O�ī�o��-�Z�i6%�Y���*�"O0��ȯ&�n!C&�6d��-�v"O:T �N�`�T	{4 ���j �C"O��[$	�u���Ѣ(Q*���S�"O����Ɯ�x�|9A��=[��8j7"O���3�*Y�e�e�Hň "OH�BPL��9�=�1�
j5���"O��J���ZP㭊�&&)�4"O��P'F~]8�z�oN=7z�b�"OE�A��-Rf�yG���T)<Ey�"O �:�O�+1��3��U�@.��r"O"01��Ƥ{� �(D\^��%("O���TKǜ;�lC���O�&�+"O��#��pިXc�T?����'"O�����*&p܌0C/ s=��À"O���5-È]�� ��m���:�#T"O�QM�Q"�dQ&��2�<|{"O��#g	p?B�g���%�>�{"O�� 5�~�2���k]��B��`"OR��'cvw��3
�_�f9��"O���5�����K	�+Q�8Q"OH��N��H[�ZB��`"OHY�P�	�TB@�C!� ry4Ȩ"O�l1��ۘ ��A�jaшU3"OV`�����-}*"���|��횲"O��2���=�0i�Uh��t� `H"O� Zd�O4^&{2��E��1@"O(� $�*P���<:���"OJ��Qg� YR����e��"O�5�WE [�du������S*O&�qM�=w��,�����N��41�'�*�m>�@0C�"BT �'=�@ѯ�'$�����]�2��+�'#������<JĀ{���'	�I8�'p4����/��(K�X�V&U�'�.�@&é�����+F����'B(�`A��S	�q0Ԋ�M����'����r�ռv�`;p.�$-t�`�'d���	��F����b���h̘��'z� ��'G,'�8�
^j���2�'����3k^5o�V��R�_;����'����J�2b`�-���؋(���s�'��u��EA!h!��+���#L��U��'���ݹ"��亗�"Crd,p�'�>�&��vZ�}Kgf1h��
�'�tK��@�N���i�[���j	�'#�T���>Ӷ���Pi���'�l���ʟ"`������4U�0y�')t��Q.V�1"��!%�,Y�T1C�'`b9�ƮS-/������P#h9+�'��"g=wy�;�g
"C��9c�'řJV/o����!/9�Ȉ9
�'�D(�Ra.~fU�4ŏ*\�&(
�'�N�p��3R�fO��I�	��� r���ڮ9�u�Ӭ�=�"e�f"O��r�[c��q�H��nU��"O!*#
��
|���A�L~���"O�X�"�&a(���j_�Qm�A�g"OJ��Հ\#o%n�� ���.��hw"Ov�K��ZK��Tp�*Cj���"O��r 
  ��     u  �  A  !+  �6  �B  �N  �Z  _e  op  �x  Q�  ��  ��  K�  ��  ١  �  `�  �  ;�  ��  ��  H�  ��  �  b�  ��  ��  ��  9�  � 	 n � � 5$ u* �1 �7 > �@  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG,�!��}�:O��J��T"�o��S.�i�c�)o;�|�ȓn���ca�Q�]�T��	�9�D�Ey��'"f��d�;ɰ��d凸U���
��'R��T���D!P�A�i���<!�A)$�`�$D��;���v��b�xJ���OB�r��h��%@���I;� xs���Jyy	#D�x9Ɔэ[�.	3$�Y|T�X��s�T�E�'�]��QTĬY"R�ʑCppa+��~�Ьm�����RI�� !a�T��y�jԬGI��jRb#@���7$� �HO�	{�O�F�
a�D+5��$��~~�uK	�'W쀚a.D�w��)˷![-�=�B�)� <L��`
&s�L���m�4!���"O^��v&"~�s�ʊD���"O������SW4D����0d�,A"OT`��<0g�<k& �-�r5�%"O�]�c�8`0j���o�%�<���	�O� 
〗�:H���vG~���'%����(@#{�� ���BhP��a�'bў�}G�� {�h�"E�ju�� #HP}�<���ğK�nx����
Ud�Z��	W�'�axB%i��a�(���Tx3���>�K���'��o�VMZ�"�vČU0��/D��Q O���mHaf�c�,{C/��ȟ��5e��R��JB�ӎ'VPA�"O�X��d̵`�0� OE�e�¬��"O2%٢�7Ңq��.)���6"OƑK�cH&,����-P�6p'"O�2ϟ2R|>`J���_����"O�� GN_�JQ$�ٳ3y�5�#"Od}b��ؗ==X�C��
k�$���'w��8�j�bD��B�/��Y�-��KD�0K�U2붉�fK{�Gy���e>i�u�P��P\��ŚfT���rj;D�8���3C2X	c�C��D���G#&D��ʥ(�C�|�i���)r�Չ��?D����!Ƅg���*W,x�4D���;�d;�OTuK�D�wg �+Q�I�W�횰"Oܐz�*�C�l���ɐ����"OHy���I�F_|]��$�p��H҆"O���i�{���`�l��N�ْ�"O�(�rA����Kuf�-Y^p�Z�"O43s�_8`>��a	!G��I�d"O���R�)}.Jd�۾{E�]�	�'Bht� ����PH[��^���'�v��0�� ��3l��#�l(�'���0�A�b���Q�C^�^�I�'(����Α�0(Ұ�C!1;��	�'
�j��D�]�x���R?��s	�'��pq���K�n	K��ЈJ���C�'�F�0t��g&�(��e�'D.�83�'/YpԀ��xF�W�ȲK��0��'�^��d� @rP"�#��E�����'���2�ƎH"0�S��7��ȑ�'��/ʴ5@�̢���=@��i�'zpR�i� {�T �Gc�7��q�'��q�5M
1"��h�L=3ʜ��')�0�H�?z�|ó���UP8�'�r@Àd?���]
K��y�':�I1HA
�Ȭ��C	?R�Ⱥ�'$4 p��A�s�^��KZ��'JL�1��>:I��Ԅ
�RX0�'B���C�җN����'Cgv�Z�'aft�Bn]��,S�E�$���`�'��U�$F!;�~��1dW&j�<!��'��(�h��9p�� ���b'nu(�'�bi��T+4�!��]8$��'G^	���v�P�ٕ�	��X0��'�\��&#N��2i*���"Q���
�'�l�91E��]y��[��Н n�H
�'�H@r`J79*.hAQ�F+��4�	�'�`�EG:,�|xZ���s7�I
	�'U<��-_ 4aZ�P p���2�'��dh�k�U�E1m�<}C
�'^��r"�ݔ.�HA��M�*e؝c�'�0 '��?(D�s�O3^���X	��� ���L�W!PY2��9�b��2"O�I�OD;m���R&�7�V-Y�"Op�+��������E֝x,���"OF���-�&%Ȭ�MWꔈ�"O言�ӀG�P���+��<n�)�"OLd�w� Y� 𠄛����)""O�zJ�(��1�C�	�H��"O�����M��vա��[�=��("O����)Ē@�@8���'��݈�"O���&�C�]�,��jE�tB� ��"O�ЛƇ=7��|��ksERb(_~�<��f��\K�.P%5�B��pOA�<�AG�)�h����p��4���AV�<	�
�9	�hd����,?�P�E��R�<�5S�D94�B��WP����QQ�<I'Y�1j�1��MI�T�0w��r�<	5ȋ/fή����)`0b��J�<����p�^���*���FPA�,�D�<B�T����th� IRv=�D��<� j��u!b8��4AY+�� �<�a��SD�\�")3\={u��v�<�&a�ltJ�30ꉇI��M�1n�t�<�%D��\&�a�1�Ax�t �'�IJ�<ɦaW��ڭ��&�S��9����D�<q��Z6:�x���50�5*�
�U�<�f�u�DyW��8	�*Ƨ	L�<I5hM 'Ė�3�l��~3�I�F�E�<��p�oC�'�R�s���6n�ȓAe��c� e��43��I
�)�ȓ>*�z��H�Sy.��e��L���&H��lõ8�e#���l~<%��m�v���'�7OP`;v#�7+�؄ȓj��@�%�){̙c�L@=<��ȓzμĒ�iN4Vc<s׭�Qd���e�R���2V�=�0"D�8$
t�ȓJ�v ��X�n��%;��\�?�䱇ȓg���S'�ދa+�]�c�>�,Ѕȓ|4�u�#��=<��a]�G��=��P�:����Y;R�p)�r�ִ9��1��e��4�?]�\(���:���ȓI�؃p��!���r֤������ȓ�����  0[ =�#J����B�
��P��t^�����6!��|�ȓ&daۗ��wDΐ�q���l�����b�N� JCРY��G�n��ȓ	?�4�"��}�ZP"r�OJW`)�ȓ!G��s�.��6���� �rI�Նȓxs�Su�ҬY��E�$���<܇�D���(ABʄJ���J�[��P��Zw$�����3p�X��
�9��(��KŤp�)�+"���zslM�`�x���W8�Pi.�F��V"�;`5х�.�,ؐ��2�L���4P�
���V�8=�ըW 'ᐄyL]�d�ͅȓJ/��
6�6cNh1�m� ���ȓwi����ĥz��S�����ȓS���TnՅS��%� [�T��&�@��Ba~$pS�$Y�w�X�ȓ]�6h%���sa��<Z��E�ȓ&��E�tiM2<�A�0��*�e��_je�׋�� {���L��e��j;*5C����z�Z�j ʜ5XS���1Ȫ�#�.
lY0ÇQt�h�ʓ9gz�I��B�W���ʷ �&ߚC�)� |�I�o�C�F��AH�>?1�쀶"OB�b�L��G�8�P�C�PL�iS�"O�9�g$H	z�}p�߄-L,
�"O��˕C�6 b1���U.�T;�"Oҝ��Mi�%;�ٷg Jј��'�"�'���'�r�'��'*�'�T1k޳��`0��Z�x��;w�'�"�'q��'���'���'"�'�[�W'�2����YSo�y�1�'���'���'���'���'e��'��X�3
S�t:I��#�ll)I��'���'&"�'���'��'�'�*d)�V�B��r��A�7kH�S��'��'���'�B�'k��'a2�'� �'�2D�~�ՅS%7%,eqQ�'e��'^�'��'�b�'/��'J����@ܫY�]ӆe�*|i�h�D�'r2�'m��'|B�')��'qR�'!�cg�3;ٴt�`�ع����'�2�'O��'I��'�"�'�B�'�$���-F�	��;#E�/�.$"��'%��'�r�'��'WB�'�2�'+�TAsD�<v�H�2/�D���`��'X��'�r�'���'`R�'�r�'V��SH��U'mJH�f�y��'�R�'���'H��'�B�'�R�'��l��GW�o;���q�|I:��F��?1��?���?a���?i���?i���?A#S#I��E�S?Y�򰀊�?i��?����?i��?Y��OX���'+�bL�g��yۥ�Ұ+��!�@�^����?.O1��I��M����}� m����y�٢�k
"K��'��6��Ob�O�9O�)m�[����l��M���}��p��4�?��`:�Mc�O ��I_�]�*P�H?�)��r�Hx��K|�bɻ�`9�	ݟ̗'��>S�@J�1�ԑ�EO�nW:y(�X9�M�1&z���O�87=�)IB�%t�\9�7�M��ܭ"��ҦY�ܴ�y2W�b>��C��˦��V7HR��J�p�S�F/!��PO �	�=����4�Z����W�~أ�]���lؠ��l��ķ<YK>ᴲi�jH�yB��6%����/O��]ô@A�Z��O�M�'�7�����ϓ��dщ�
��*X�����O����&T�	Q!ݯtFc>!X�!R���'���b����K�&̍D���{Q�0�'���9O�V
��)oP�I����ˌx8�6O�	l�6���5^�&�4�x��d�R4P�a�$�4��iv6O��lZ��M��Y�!��4����d��9�A�̪�gΠb��������n8
W�䓄�4���D�O�hӢ���Oyۃ�	N)bث����ZmsQ�<���id�q�'���'2��yB$��±`F�F�[+8��M�]���p��{�f�%�b>EA�/�-���r�XM��B�$l`� `�#[���$�l�8�JUUMH�O��!"�;�'�p�@{	�L.%r��?����?I��|r,O��nZ&��ɹgx�ܢul��4��YA򩖍Mj̙����M[���>���i��7�_�3dl�+����+8��T �ȕ1�e�J,?
��@��冝��'a�k����]�Ě-A�|��'gD���O����O4���O���9��)��$���-c�l��1���J�u�I������MSWɕ�|b�(ߛF�|"Ɯ����u&��~�A¦©Cxd�ľ>�T�i
�6���P�3Ht��	�&�Q�1��T�d��3W��<Ժ�JD'��\2�OI+9�p�$�Ա,OP���O���O�X�� �8T�цG�y	 #f��Ox�Ġ<!A�i�,(c��'��' �ӬJט���O��Hn�GÛ�d	8�P�����M��ix>��1�	�� ���q�t��%Ƿ1�I����
Z�6tb�Җ!H�ʓ�R7M��u�'�36r�	#!ʠ08���b���5e��$�O���O
��)�<��in)��>���Q�˸U7��	��V�s�B�'�6m&��8��$������@ɦo�,- B-�jM[�A�M+սi?h@x�i���OnuEm_YQ����Ȱ<�GAȇL��8��A|��qe��<�,O��O��D�O��$�OFʧ
�T�Jw�Vo2PT�Y��J��!�i���Z�$�ID��⟠c�����,W�3���Y���?fnl1G��x��v�y�b,�I[}�OA��Or6�8��i���.jD�1�)�����bθa��B'�
�c�Z.N�O��?��(�@x��J���`
�%`5���'���'DRT����4%<���?��7�!����Xw�����9yh<Yj�R!�>��ip|6��s�I/���jѪ]�[�N9¡��z���ܹEC���\�g�SIy�O��j��>���1�Hd�%쑚<�<ň�cw}��џ���˟ �	P�O\� ��w|�Ql��N�,�*4j0gBb�J����C�4���y7�	�ooJ�6_&آ��О�y��|�2�n�M;C�پ�M[�'�r��$�P��Phɦo����t&	��P���١X����$�O����O����O���Q�Zo8,��-ϰVn�p;�����d���H��??�����O�����,�i��cݻv\��c��>!��i�D7�IX�i>q�S�?�RI�-9̪���\-|��ZNǒ����+�gyRhM��&��׷�$�ȗ'4�XG�I1D�.��Ǔ�v{uض�'6��'Ob����R����4�U�=O�3B'&���c���0��;O`n�Z��k����M��i
6�!#�xT��X�g^q���]�q����c~Ӕ�	�.���K3�'U\蘄��<�ӱ4�j��=� "XۑFXju�A2$���<�́ˆ9O��D�O ���O�d�O��?m*��O0c~�J�Ե7��!k�r��	���40m~Q�'V`7�>��F?	B��$B�U��Q�Rl@ ,�NH$����4rF���O�|Hýi��d�ODpG�> b��hF� �~t��
-i��Q� ,IV�T�O�˓�?9��?��+3��S���JA���A+z�́��?I+O�uo"����۟������۝�t���c[6jƄ �(D��D�p}�m�pUn����|��'|FJm9a�N�8ϐ< t�H���3g���T��ɕl���$��$<��w�mL>1�E� *_��aYo㢕�b(��?y��?!���?�|�,O��mZ'fI̽�C�еE율��N����j�C<?¶i��ON��'}�7�6`��C��>����D[�A垤o�M�,�Mۚ'h�B׻}�H�f�'B�	$�B]�dH�T�� ��luP�IUyb�'���'��'�B[>��啯8�<,�T�BXB)`&�E�M�Ǖ�<����?	I~Γv՛�w ����y;p��g�K��bqw��l����|��'��0�#�MÙ'�����$��n��R�#�<��U؟'x���9e<n|��|�[���I柰�u��0���k�n�o��8� _� �����IUy"�`��0�t;O����O �*"b��@̝4j�T���Ҏ ��+��d񦙊�4\Ӊ'(h�fM�PT��c�?�M��'��u� E�V
xB��&����J�]$T+�!q]wLR��(Sw8	q��sѲ�� �Ʃmh��$�O^���OR�$���M��|Z��e4�P�ď�?��i�����'b$o�x���#\���5O�8x�@���>�:�ɨ�ME�i�6���R7������D�Uǖ�0VFJe�`�s��M&+�0�rvCւ-�b�)A�<��lyR�'q��'�B�'�2��r$xc㡞�<�h��FӔo��	��M�@���?9��?�H~2�D�hp*'�J:� �!%捒H��y�^���424����O�#}J�Ι7 ���"2��m�XA��� "�Ұ�f�����D�'sBj�{@ez��*J>�-O(��hL���
'π�P�C�O��D�O����O�)�<�F�i4x���'a�d���56S8�yĂ�Z�\Y9�'�,6�*�	����]ۦ���4=S�V���de�e,ҡA� �R'R.t����ҳi��ɑH�T�R ��;ZOnM&?!Zc�@Hc�DP.�̰���pcHu��'N��'���'�2�'��:=�����P���ǛB&�L[���O��d�O0m��i@������j�4��@%dݸ'�*��!�%��%��t�'��I��M[�������Ɲ��*!�N1<��X�CH�s�!���*q`а�F@�F���&�Ԕ'�b�'���'���3 
m�� ���0碈rT�'�Y��۴"�j����?Y���i�2]q�d�$`S� � �[�{��	��զ�ܴ ���¥>�p%����jz,�'�q8D\j���	G���↫<ͧ7i��[wn�O��8含���ꡫ�j��5X2b�O>���O����O1���m���SG�aqPIM�%��S惊��h�E�'�B�j�~�x�O�m2"984Z7.�+h��HQE
�G	 �شK�6��*z*PT1�OB��4�K�M��&%�<y1F��*m�e*Z�l�6L��<Q(Oj�d�Op�d�O����O�˧N��܉��%`�bˋ	FPX���i� ���'��'���y�&i���M2ҝCi�&%�Ty9�`��xamZ��MÂ�x���BA�3;���'���H�։Oz�Z�*�,���'Gj��Ao�U�8P�|b_����蟀�g*�e{�y��trDL��������?1���?A)O�o�(8���ʟ��	\��A�%#��J�9���a���\�F��I��Mcִi.�O�$��#�v���AwJ�$J����C����GS e��Y# �x�r���i�ޟr���:X�,���;4�W�ퟨ�	ޟp��ԟ�F�T�'w0�
&A�v��1�ҙZv|���'6�6�?8�	��M���w��U���J�\���H2/�dH�'*:6�NŦ�:ڴ9X�mjׯ�P~R�H���<I�L�9+��d�b�ρl�%)j�	�}��|"Z���Iß�I�t��՟<i��>6Q.�ѦN��}5BQ�SXy��~���R:O����OΒ���*BN���7mR�\C�IN	�2��'�47W䦅�I<�|��H܌4��([FfA�����u^|Ԑj����@2J���AS��)0ޔ�O��I`�ѧ��a4��@�'*�YX��?���?)��|Z(O nZ3t�$�	2Q֢��:_�̱�%�ro�ɺ�M{����>a'�i��7m[�U# �O� ��A	Q��*Y%$�0w㝺yݠ(2�<?A`�46*ht�r�<��뿋� Η0B���O90��p����<��?Q��?���?A���E�0�H���	�!T�(
3l��y"�'�	w�^M�А���۴��|��	 �ʘ$Irͪ&�X�Y7�xR�u��lz>5:ĦdY�u��<�%�?Wg6�hd�QR�� ��X�cG�Ee�'��'���'(2�'����P� �"��E%�_�Q0����'`�]�H�4g`�`�'bS>e�$�&2�U��c� 3�
ɪ�%?��^��sٴ,����,�?9Yw	,|�,���O���d0V�uQ���O�]��}����Ƈ�n/�ΛA�#�*��B٧i$F�J��K5f�� �����	��D�)�dydm�(2�ݓ,(ZM{$D�X���`�"��	��M#�r��>���iK�8���_&
[���J���p��عE�����T`Hi�V�^��WmݜI�"��*O� `��c
�"F(��˅�T0,�7O�ʓ�?)���?���?������B�T�j}�䝕_�5C���{�hToZ����	�(��G�s��q�����OL�z�@,�@�Q$`�a��
ݚ.ʛV�p� \%�b>%v$����͓|����K3eh�aPdL;O�d͓[����c�C �;H>�+O�$�O�(RNZ�����ݞ,�l��c��O���Ox�$�<��i�x!Q�'/2�'� � ��5&��L�B"O0̼Y)�d�q}�m�<�l���,�\�hD��<1T�$��M�%��M�'U���CM�.r�j�:��ĆJ;"���P֟RSI׈��i����;�t� ��柨�I������4G�d�'"J�B�nJ�Pm,Y�i�#D"�D�C�'��6���:��O��n�s�ӼS�	�����f�>i��=:t���<qB�i8`6Y��=cq$ҦA�'��}jvG�2	��h#pÜ�jKl8��F7ubL4ptl21c�'`�؟0��џ��I�����=����t��R&�њ[�-�'6�7-�2*���O��$#�9O�k�EW�$�L�@#�J=n*���{}b�`�*oZ���ŞI�M!�JT�K��	�$h��=ȴ/��P��z(O���#CD�CZN�]!����d�-���A��.xbu(�h�@���O��D�O��4���@1����y��d{B�����%��"\�y	wӆ��	�O�nZ�MK�i�����/q+V�2���[J���g�&,D�f���Y큆k<��L�l�S��Ai�6b�rI��ڇ5�\��Op�d�	�L�I��p���x��`E�.f���	3ő���p��,��<Y��?�Q�i/�]p�O)m�N�	�g�^5A�aT������戭`N<�׼ip6=�~Qk$�j�>�φH�R[]��ct�W�W�LQX��u��r��������Ot���O��䚻(�D��)�e���2s����'��R�DA۴'�Np��?1���)I8r7�4T�ܻ0�P0rdɎ->�	 ��dAߦ%8�43���)ZJR)���Ƨ�.pz �΄A6��!0��q��e���<�'J>ja�^w�,�O���g�=<&�H��P
>�J���"�O���O���O1� ˓~K�v��4��"��VHDݒ�I�+����OD�n�g��"���:�M���=�t8s��O˲d��Y8��v�g�2���oӚ� >ʁ�C�L�Td�/O{׌͡2���h�$m�1�0O���?I��?���?�����^�?�]ɀA[ڱ��ʎ ��n<+R8�����@�I}�������[7����؝K�.ݶ[��Q�CK��6�sӦ���b}�����:+��>O�`�[.���2��6R�0�(�>O���lO��$u��9�D�<i��?1T-�*kMLD����F���"d3�?����?����d[ئea�DQhyb�'@tT����T�̄��`��f|��U�D�I}�*f�^�l��?!�O�L��ě�1�t؂�FF0DHh񉐘�0��E�l�s��J�>8pPt��N~"F�+O�)���Ŵ=�`б��OM��'���'7r�ٟKrJ]-R���͒G��&AR�HB�4-�A��?�i��O��� G��F�Rl0���#��FԦ��ڴ�v ÷Z�����`G�/ ��!c��7s��I2ˤJ�\b1�LM�%�X�'F��'���'q��'�4A��F �!��	8���{�]�h�4-O�����?q����?�)v�`�Kf�N%�P-��!R��I"�M��iO>��2�'o����;i�@���P�R@�$O�^ʒ�)O�"큃�v�����򄞘C�hR��~��҆)� ҈�D�OX�D�O:�4�h���֎�k�R@M!h�|4��h��k�̸q��ʿO�d����O��lڧ�M뀶i�*���ďu���S���22��(�d�S"K��柟�ңOZ,B!�N]k��&�5�b��0�����V?��)�����y��'�2�'���'���IƄ�̱��II�X	�%+��_�O��$�O��DX������>?iE�i��'d�D� ��kj���%�.=�=Zt(�٦����|r\:��9d&<?�2$P	z�J�Xrj��Z�:�'	���`"m��&�)`I>i*OZ�d�OJ�D�O�|#ե^T����(ވ��X���OD���<Q��i����'nr�'K��2u��iS >j}�4�ww�)!?��\��ߴ���O�c? �b����'��	5X��Z���ƲX�̖���:'���y�	�Ud�-���^z4��K�T�-����@��ٟ��)��^y��p� 	3�(�'�� YvnG�$ud,����&�t���O�!n�M����	$�M����d8�p�19dD%�7nױ;���l�Z�锪sӺ�f���1C/:bh$i-O�e�Ģ4N��t,1F�څr�8ON��?���?����?�����	��Eg�P	�M�����4H� 1'��mZ�*W�������V�s�����K�ǞF��D��(:��ؑf�d��nn��$�b>�ǀȦA�R%�*�HF�#9�̈& �q0�	�)�D��w�ŤkT��K>�/O����O�}�r.ݥR�~�!7�	�OW��BU.�O����O��d�<ٷ�i��H:�'���'�T}�vaóv��u��!j>�S����a}r-e�F,oZ���n�n�SBA�*�
Ep�"ٞ:����'b�U`�.ɦF�L=�C��d�L���nO��l��䓲1��%���!�HH�G���,�	����ȟhF���'�*�ڂ�
l�X��@�1� �'�6��P��	�MS��w��t�*i��9��	':�����#1�&w��nZ�43T�m�e~�k�$S�����O��� �4e�ǴZr�R�0#o‣p�>�D�<���?���?���?QE1G�
Æ:j�|��LǺ��dTǦ�؇Ll����۟&?��*Xh�}P��jV��E
&i��1I�O<o���M[�x��ĮU�K�l���,0d����	�9�>���&W�	+ ��x��ֺC��|�Q��b #w� �`ϑ�7�^��%V柈���d����Siy�ch�<�BQ;O�U��f������ƬJ��hV:O)m�U�4S�	=�M��iN 7m^�h^���!#�.U8F�:� H%%s,��@�r�L�;��9Q2�?3~��M~���kI.���Р<Z,�g+� "�9̓�?����?Y���?�����O�H8r`�I�}�:��g[�|]8���'�R�'�7�X�����M�H>aS灞@q:IQ4�9��+%��?v�'>:7�L̦�~H�m�|~��Χ#���ê	5e��MB���b��=���̛`���R&�|�S����l��ş\Z�NR<G`-x�U������ �	Ly��}�,�d9Od��O��';��ܢ��4d��dG;HC�$�'���hv�f�qӎ�&��'7���b�N�E�PM3�U�;8�=�r��T�٣l�1��4�6����o�;L>y4�ΰA�6	Ҕl��{�$E�1R�?����?��?�|�.OZ�mZ�961*��ˢ�n��bL0l�����3?y��iC�O�E�'m�6-��X��U$��p�j�BFP�_"`l��Mc�`6�M��O�`��[f��F�<�&�74Kt�`��Q
��� /��<Q+O*���O����O��$�O6ʧ�h8��[�n<�9�rk��u��i8 �i�B���'Pb�'(��y�`t��O�<�q��@�~�6e9G��.2pIlZ��M���x����X���f2OF[�j�c3*�!V���8��݉�2OH�����I�&!0�(���<1��?���1 ��إ$�k�����W��?���?!������Zrw������4؀-	�1�Z0��*�+��9r`DA�S^�	3�McԴi'�O�R���jZ�8%�:-��h呟Xp�O����C�M�d� �կ;Ҧ�*y���@b���x��ӊQ?qSb�'h��'�2�ڟ����V�#��jgf"Q���*T����LZ�4~� <�'	�6�2�iށ� �Q���/@f����$x��:�4_&��bpӆ�Nc�(����9��Csz� z���WV@Ң��;	�L(AsɃ'������O4���O^���O��$�3;��`#�f�e��s���[��˓ J�����y��'c����'!���΋z�]���ǒRX�c�>i��i��6�J�)�=B���+��I��Cᗙ�\� Cl��A�䰖'Qn옐I��5�NNM��fy"풟d(0w$��PpЂR))��'B�'b�O�-�Ms@i��<Y�H�����5��l�x3o��<���i��O*��'Ī6���K�4U
����J�R�# ���"�\M���2�M��O���jB�)O+m���'Կ����UҎ��vb��0\��22l[�<Q���?y��?���?����ϓ6���
��0@,l�D���y��'Cr@sӨ=+C���b�4��E,�}�UF��#\� 
ũR�i]ҍ���x�{�&|lz>��_��ne~ҋ�q��,\4�11hC��	���"n���$/͝������O���O&�d�/y�%)f�W	*����m�����O�˓��� �����O"�'0�P� O^�:w�5���	\�'���i$�
}Ӧ�'��lk��3QiN
PyjI8�H&-�Ҙq�f�l��e��ǘ���4���땳��2`�|rdG �T���a��0<ړ��,ZB�'B�')��4_���ش�p]1�$^)A&��0+�3*P����T~Ou�<�\��O"xo��o�,���k�w�&����2J�����4|Л֍�7:ț���<���D�`�f����Ty��H�x����ê^�aN��SM��y�[���I����	����	ן(�On峃6".�����%!^J����t�As4O��d�OԒ��$Ϧ�]�3+
h���'$�+@�90Іd`�4m���%��i�3T΅�v5O�l���8s0�A�J�<$6�}�=Ot��� O	x��aC.�D�<����?!v.�"e��UcQ�<>���9Ө^�?���?	���^㦩�a�~����� BKK��|%��ߛk�~��C�C��-i�I�MKԶi|�O�|ң �6�^�ѣ�݄�P5��`B��^Y�I��Zy�5NC�y��ߟ �j�&a���Ć	�q Ec]�� ������I��LF���'�h|�����(	��އv8<�Hg�'��7�E�	��M��wQ��zc%�,n�d�㡮Ҕk_��'�6-�ݦ��4G�����$�^~���0u�X\�vŉ�7���*0mݫI�d���'F�v�h��B�|�W�T�I�h��ٟ ��ҟ��d�τS���c��vq���SM_yb�j��;@=O����On���D�B��#�g�c�^�aN
��'hP7m�Φ��M<�|���d)	���.by�K
���� -�����R/u)^�j��5Y^ �OZ�x�l-bD�H�!����Я�m�~y���?����?��|�,ONDo�cI��	k����X�d�ҁ�+Q��I��M�b�>�$�i��7mJ����"���H��`0-��SS ϺBۀ���=?��R�Mq(�Sb���'���GK�KI�d��X>`�r5Γ�?q���?����?Q���O9�h��͙�Y��	(b���1k���'��'�6�4L�����M#H>A�����B'�(t`���ڙ]�'��6m����ӥ`q̵�t�6?��Co�? T�(�,]�T���`���3x�puE��)i���6�9�d�<i���?)���?i���#���X ��??������?����J��5�ǟ@�IޟȕO`n��rN�B�m�nؗ^-~8��OJ��'��6�������O��iҡ�+]]��I���~�j�`b��:<U�jԥ��Y�i>�j�ޖ)|z4$�,���,_�4���bƿ.�К�ן���ܟ��	�b>��').7-R[>xx�E��zD���q�:ۂ%���O�����Y�?9�_���4.�޽c'��{�d���+��}t�����i��6�2B��Ja�� ���́wԺ���K�kyb��'*�hpҀ [;葘屨,�����O����O.�$�O���|
���O���t�ʵWn���ӱA���(�C���'r����'�n7=�V��e�U+vp���F&j�(��k]ͦ�ڴ��Y�b>�P��'BpP�ɑ*3�8�H3GQ�L�[=}� �	�[�� v#D�m,��&��'���'m�t��NF4 D#M�B�0"u��'V��'��I3�M3"���?1���?��C�>s��k�AT�C!x��D�)��'v��%��(i�:���[}�R�g�nȉE�̠6s��a� �-��D��y/��@ŀ����j4�� [� ����8����A�E��c���F���O`�$�O��d,���.�,v"�0�ꐃ̮�SSA�?٣�i6^1S��'h�%����ݸm䕃���&y4�1Մ����I)�MӦ�ivH7����i`�� !��3!���VIޠ2`ڡ"u�-h������]'��'���'��'lB�'��Q��.�K�B��̔zc��;]��k�4.aJ�ϓ�?�����<���՚������V�9�{�,6-d�ɥ�M���i|�O1��$�t�ǚ ֨���h
�x�4%�d X��<��#��<i���<o���&���䓼��4�+�@9Xcr-�N�1	P�;���?���?���|�*OX4o�2��]��
pl�q��4Z2���
J�����M���ơ>���iך6m����keD{��$�k�`PbU��B�Q��	�w)*?sϋ�
�@(R/@��s�kL�V~>���O�����թ��,"���O`���O�d�OX�d6�S�o��a�r���3$,FLG%)���\�	��M�!��C~��o�R�OfP���(����ѦkT1���e�	��MS������m6|D��OP�!�hP�0�N��[��ϟ Qn�1��Վ*��Ol��?���?!��:��-9���1�3�'�7x�������?q*O�%o��j����	ҟ ��|���M��9�V�#w�8}A���D�e}B
Ӓ�nZ��?�L|���U���S��d�x	�ͨ�~��Vɞp�bU�G���d��"���?J �Oq����L��bC�F��P���O���O����O1��ʓk�f@�`9�t́
�T4K�ѭX�$�+F�'��bf���$S�Ol m�:!�����b̟J!bAR�gXP:��شpٛ6d^;r����O�e���#�,1J7��<��7y ���#�%z@]�^�t�����O����Oz���Ol���|��(ܥi����TY#���&-�*������y�'����'4�7=��9p��ȄA$MX�!R6`������Φ:ٴ@���O�,:E���yb�S�iC�e p�I4\��|x���
�yBG]���� ��G��'��	��	�k�LG�Z	i� �!Uc�W& �	ԟ���ϟ�'r�7���xx���O��,82h����8�ҝ��&���X��O�-mZ�M�W�'��I<&�����)H��=:g2C���H��mz��.~���#M~�V(0}����&1�X����6r:�%��'IF����?���?	��h�����8x�૑�7���Rd@�H�D������F�ԟ ���r�	%�i޽��è�������"��y��aڴ8��b�Ա��$��O�P�5Ym�R���!
�k>4���c�4~�����1P�
�O���?I���?���?��(�3�#�j<���̛3^z�B(O  o�"n,֐��ß����?�O�J&y�����*�����MN��e����vӶ��	v���?���:����"�*C�ܹG�_>Aޞ4Bc�l���'��j��F��h��|�W���A�"��a;�����ܟ���ܟ��	�zyrAk���`9O���e�� M���	�Sij�=);Ol��E��O��'_�6m�æ���4|��ɓA
�	E��S.�7�P����!�@H�'Y���%)4DM1�����w��9x1�C�ˬ�xf�V�����'"�'(��'���'�񟺜��!�I�`�D�����P��d�Oz��MϦёu�0?�Z �+K>�D��'W�U��?i��0�sD�!FG�'�7mWݦ��}��4	D=?AE�̝9��#��83����r��d�VDA�b�q���O>Q.O��D�O0���O�����$)YÖ'��dj����a�O2�$�<�f�i�Z�'���'���UH}A0�V�m��K�aɪx:F�5,��:�M�p�iLO�S�S�@��@�E�&�@����x8e��\�&��� oy�O�,Y�q���%�'!�=��υ/6�ً�!���8�K��'}��'`r���OV�� �M���m�x���؄+ւ9�Ѣ��g�\<�'��7-'�����Q��I;���F�P�B��!j�D�P兙��M�i>@c� ����#>g�ܑ�*��y�\˓pӔ�ؔ��j`E�ٍӄ�Γ���O����O��d�O����|���ę^�^R��H�P���[ ��J��(Z�����Oz�?�������aҏr�xpRUK!m�l��.�[\�VBr�r�&�b>5c�/ܑw�^�)� |��� B�^�feB�M��=B�?ON$k�	�-�����#�D�<���?Y!.I�Tc��0�����q�Bf�7�?����?)���d�ӦmC� c�@��؟�#�N�3n!�A˖-*�p$:�f}�7��I6�MC"�i��O���d��6��q���ɯ*��:���$��0&�	3E�Xp�Ӽ'p�u�֟({����V�<xvC�5�
]1C�U�\�	П4�	Ɵ<F���'�T���=ra�pYEM�<0�%�'�6-���	��Mc��w������k��1
�AϞ@0�J�'>�6��=�۴�q� e�[~�#�:�l�K�
"=���+��$hB���*j���C�|�Z�<��ޟP�I��D��ן��㔈 z�������Paau��~yb�vӄ��:O����O\����ǥkp!"�C��!���A4Wq�9�'jl6��u�N<�|%[�V����#uۨi��%��G�u�ˋ���ݗ`l]�	?)W(���/S�R��`u�� `U��s�$��a�T=��K[UsV��SE�J�y���V������>3A�`�C&��M�fMVa�]R�B	3$XԐeM*U�K��ܐH���Qg�O��bc�%/S��Y&"κ&�6A���(\$�,�$I1劈�A��S���`^�S���ӑ,��0 ���ɟ�8uZ��B''�Z(��gdDL8�Q�o��*G�yP��A8_�P�â�	.b>U:P��*K*"�Ո�9&D��q��:�x�%!l��h�Q�ʃ��7��;��3,O�P�8��W�TAoAy��'��I����	ҟ���/v�R���l��\P�ј� �,�4�Mk��?A���?)��?g��E2�&�'-�i~�N�A"D'jw�*$̛`���'[�	��	�@�%<�'J��)�K��iP�A�(�:��4�?���?���D�@�[�i���'��OF��R:��=�#!U�ݎ �v�nӨ�d�<���FEv%�*O&��|n����i 0��('U>1�+
*-�6M�O��:3��Hm�ʟ���֟0���?��	�w�m���?b�x��m�4p(Ƚ��O���Ä89���O4��|�N?!��c^����u��`a��(g�j��������I�?!������	� ��õ
:�|�E�=4Ѕ����M�&��?YI>�'�䧮?�WAW9|��ݠCӷn� D��۠V���'�R�'.�bT�cӼ�D�O����O�����ܐц@=� H�C��Vf�� �i:�	�M��5��fw��'�z���?���i�����"	��2&n�8<�nZ��d��@��M���?a��?��Z?]��(nh�aլ�Lb)�1Io�8�nڲCSdxj1hb���I�4���X��L����P#����o�*,�*!��'j�8�s�mm�����OV���O���O#�����1%��Q�.;�m�>A<$�!�H�Ee���H�	̟x��z��'=��H�q>�@��U*1ZVk�M�$w,V�R6��<�����O��$�O^�4O��"4h�t�4����+GQ��I}2�'�b�'�剋b�ʙa��R�D0}���N�\�rŀ�&ߚm�Z�lZ�d�'���'����y��>�����>��HP-ÑF��	���I˦E�Iʟ`�'B�p*�(�~����?��':R�\�gW�_�:1m��M��� �W������h�ɮ!}v�g~2؟�$H�N@,MU��Ƭ��R�`ݒq�i���'�v]J��p�8��O&��*���O���t�ݦcv9Z�܃]�M�V�T}��'�=(��'��^��r�)� �fL�2��,1����M�� �v�R.��6m�O0�$�O��i쟤���O��D��<F��BG�3x���P>g@P�lZ�v�"�	��$���D���'rl�.� 6�)�(;�ޅ��vӠ���O��D�EF�nZ�� �I�����̟�k�ر��cK��jI��ƥ)pt7m�Oz�$��_��Y� 4O���?	��Пlb'�(�:PQ ٺEw�p%/M��M�� �����i]2�'�'�'�~�"�OL<!8է��;L�8��آ�MfV1��͓�������D�O|�D�O���@�7I��5�K�sv���_	4uo�������t�����i�<���9������}�
����R��{3`�<�/O>���O.���OF�$Y�lZ�`�t=��߱:��<�
^)O����4�?i��?����?)(O^�Ę:g��0$����2�_.��q{�G	+l�R��'9čZ�'�R�Ш������	�O��p�?'�Qȵ�T�i�q���¦��	sy��'�R�'G��{���4dP}���78�1k3GJ#|k.�l����I|y�	
�5@���?�����-8F?^L�4�
 _~�	d�P�$�I��	��|3��w�D�'R챧ԟ.���G�p���J@Oŏa�6A��i�	�A@`�ݴ�?����?�����iݱ	���F=zaD׃tǮ ��#lӒ���OT��G9Ox���yR�	 (	�h�!��C3c���.����9��7-�Ot���O��	~}"S�����H�+40uF���i����M[�'��<�����D"�(ر�8?�<�a�ˮV�	�'�M���?���!!�x��'�"�O,���J�0%���h%�x��;"��ȫ#�1O�$�O��ă*�f<{.S��x��&GR>`m�͟���]&���?������sV�")ܞ	�@Dh�.�&@R}�JY2��'��'4bQ���ƆA�,���yR,�}!W�M�!��J<����?IJ>�*O�u�l�tzZ��&J�s~��hR��1O��$�O:���<e�ơ=:�I���,̂Џ'|�a���4c��Iş��	{�	Ey��ި��dͦ����N� � ��
��Z��I�����ٟЖ'�6x��l �E�10��W���*�� (��O,u�&n柔&�H�'�u��}2��c�����/�9y� �$"��M����?9/O<���q�������� �Y�/�����1v.�$qj���&�xr\��S6+.�S��� ��h��C)U^^�;�@��M,O���J�U���f�$����'ϔT�$�K�D}ڭHu�H�b0����4���Rm�b?�
��(u��`��K6¹;TixӺ�CV�Mצe��͟@�I�?��J<����4t��n(1�|��� ;X,<�X�i<�������tB ��N@9����$��x2hݗ�M{���?��dґ�$�x2�'Hr�O�b�kF��HÂƿ:�K��� �1O���O�����&y
w�:*�0�&��$���mßL��C��'�|Zc���c��H>-�`����V��!�O�M����Oz���O�ʓH٤C�.B�3HLk��V Y�*��2P�'�R�'��'��I,M����D̆dќ�R�(�w/b-Iq'#������h�'�t�5Je>��o
O���k`ܛ-'S�c�>����?9H>�/O|M{%^���iϷy�x���*ݝ1�yw�>����?I���Scr��'>I��I��h�R%�U��^�:��ȓ�M�������ā'��O&	�4�E�5j�h���P2d�b����i���'��W��J|R���5$ղL &���CA؈�o�-U��'1���#<�O���k���6���4-W�4
�4��$]qRdmڲ��	�O�)�V~)�|��1c�+-v�(n���M�(O����)����X:$�
�R�4�r �;4�7MW~�dUm�����	̟x���ē�?�ő�]��Y��*��CR�����J⛶���O>��	�]Ӱ�P!�U�	���r�3w/P0i۴�?!��?A���	Bn�'xZ�M#�'�
�wl�׶�Ȃ��!V\tK�} ����'&�'����N�� �I��.MN�*T�%�h7��O��&�I��?)M>�1V�9j�+۳+:NA8��&8����'9H]ًy�'n�'��I6U8�� � ��+�<�{�bʮBo|{&E_���'Dҝ|�[�L�֦��T6�:qAčM4��SL	Z'�b����ٟ��ny��ʻ7�n�S-�lX��B�g����GQzIBO"�+��<�ǂc}�C ?Ȱ�Z#l8�k@�����O����O�ʓ
&vd+����X{��V6�}��6i�b7m�O`�O������>��H8&΍��$�j���]�I��'}�ɚ��"���O��	L���H��M�*t�P�1�Fj'���'�Ǹ��T?����I>Qr��$�ِF���TOx�X�t�R�2�i���'�?���J���	|AB����W�_ZvQLגp�&7�<і������L<��b��UQ x����0M��hA���e��K��M����?����*�x��'�<�fH�EoH�(Wf�1k�r�95+o�P�[A�-�i>c���	7#�]����f��D�G��]��4�?���?��"S��'B�'?��D�dڕ g�Ì?�$3�!�#��O�(/�1O���O���]�=�So�

	����� Z�o����q�� $���?9����{k��S*��9e��.K�Iڦiw}�hޔ�'B�'��X�|��F��C'���x ���QZK��zL<Q���?�L>Y*Op�b�GP9�������V��d�ƤЧ1O��D�O<�$�<��֐6����<mt�P��c�*�H�;5*�!��IğP��a�	Dy�����S1l���"F���J�h×-���p��ȟ��'�,�B�5�i��e>�)��O�]�Ub��G9n��lџ`%���>D���q��^?�A��^�<v�7��O�ħ<RV܉O�b�Od�9��ރ:q��9 g�G}n��J7�$.�O�8�F���GZ������F����i��I:<�v���4^�����S;���:kxZ|s�F�K�����*�/wO�v
O��k�[�'�`�ǎ�=����ӱiy�ɒĎo�<�D�O�����H�%���I�u��!�U��c��������u��b�����)�'�?1K�^�,P�A�9t2�p�9Uh���'8�'c��Z'f-�����J�>� ��oB����<����>7a��?���?� � n���r�lS�A,rM+�A>�@P��h��В��'���|Zc�S[1?DYk�+���e2c̴>��Oj̓�?���?�,O8T�E 3F���k�`���ۑ��<h�=�>������D׵:���������aZ�C7�����$�O|�$�O������$?�t)��`˴��@��.��R�$ՓƞxB�'��'��'���Uɬ��M�`�2u��
��vw*�'I��'\BQ�p���[�ħ+;hY1!%؈Q���wJ��G9
��a�i�2�|�S��y��&�I�	j<xbHE�+(�+���E&f7��O��D�<���{6�OzB�O>jH��ЀA��������P��Z��6��<����U����V$k��Z��
�&�E!�!��v]���@ɋ,�M��Y?��I�?�y�O|��ġ#�,ia�}�B��!"���Y�|˓,+�S�>E��:r�əNv��؃��:U�finڤM-��"�4�?����?9�'=g�'�r�4� �uӢ�RW�6�ske�2�ZԷi��\����S�<�`"ͪArL=9Ӎ@#}�Z��o��M���?y��$12�x��'�b�O���W�y.%X�N�?���@��
�1OP���O���^	H s0E�s0�XK%K�|m���8!�臯�ē�?q�������� 11� X`��+�9���Z}��C���'>R�'x�\����'_#J�@2D�MSZ���N!&��L<���?)K>.O�ub�mV{M�8ӎ�E���)ڋh�1O��d�O��d�<9�Kݤ,�)I=MT28��!bv��T'X�@������l�tyR�C���P���R�ƉC�<p�%�L�I�l��؟d�'^����?�)�kW����]�+-�`K�Ԋ]v*�oZܟ8'�P�'�`i*�}2��1s����pD�)j��ȡ N��M{���?9-O<K��Ey�˟���9s<�ycG�� bkl�`�Zn �O<�.O��1#�~j�9ƾ��d�zZ���FĦ��'<fx��eӊ@�O���O�V�%�F�w#ӍU{0q[r�<�l��`��zhn1�?��g�I,w�����(�8��e,�ZO6mX�m�|l���Iҟ��S%���?���V3����R+
�K�ń�i͛�^8
��O
���O"���N0k@Ε&T�1�do\mh���'��'f�!�#b-������I?
s���c̏7>
f��0n�[xR���}��[��'c��':�ˏ"�0R�Ą�j�L�0Ӄ��6��6-�Oz5��LI�	Ɵp��ݟ𔧿�B��b�|����C>E��ݹ*�>Y��c��?9���?�-Op���C�B�$�SgAR,�bǉ54��>�������dN�����'ꏕȪ�+d-޵Y��(���O��O�ʓv�X	�3�8aF�6�X!��ǫɞ���R���I韀$���	��Z%�b�#a�D9��� ��b�(���-������O���O��~ƶ=qf��D�xu8�֪���fE�&6m�O�O&�D�O�|r��O��'=�Md�N&TD�� t��-��@�4�?9����ć;*��&>����?���r���rL?���pH����?���Q�� ����䓉���R?3�Дqq3?�lyBڨ�M�/Oʀ�BF릩�����$㟤��'�YI���]B�`�!I�Nx�%�ܴ�?I��-���̓�䓌�Oq\(�I-L�`98��C	2�Y��4)2ٰ�i!B�'���O�0O���I5L����1$Ԕ����I� �*En�~�0�	ryr�'��ry2�'P�Y���}�����M�7����$b�`���O��$E�"lI$�x�	ҟ��+AP���κg��F�d��mnk�I�Q���)J��?y��T� Y�կ�x�3�F��� ��i��Nt��b�h��s�i�yc�'�& "���&�� ` 
��.�>�D�?�?9)O����OT�Ĥ<��`��H�~�� +�����q�
��HS���O�OF���O�`[��	>�0���9G�D��!�b�d�ġ<!��?QM~r�oͅ��޷_؀[�/�>.�dS3���?9����?1��.�|��'#�.�DvH�`b�>�>���O����OB�ħ<�4�}�O��mqF	]�h_%R����=���}���ĩ<���?��d,hd�*������鲩����@�B� ��*YoZ͟���]y�%��`����D���itV�_˦!`��?F�9���s�I۟ �	cN���u�	m�'�
 M�����;]}�a �U���'0L���h���Ox�O���� ���AQD ���c@�L]oZğ,��
[d��c�I]ܧl\~�G��%e\T1D� y� o=X�V�۴�?����?��'"t�'n�㈳=��z����E��ā>7��6V���4�9��Ɵ��G@�l����#Eu8kR֪�M����?y�1�8��b�x��'2�O��p*��:z\1�WH��t�-9�i�'M6!雧�Ӿ�l��q ��t���5�ė%azND�)Ҋ,�!�d t�l��H����0�(I���z�D$v1F1rR�*4�=(5'>��<;!nL%RzDE�sg��D�B�ɼ֮��d�Q�/c�h�-*���{�kG3~"�%X�a��po8�AcQ+8d�� ��
@��AՁ
 ~e"���o�}�%J�B	 x`0T!,L�=�#.R�jRV��קN#d��CWǜ��(�9���M@,_��?���e.�]I��?ٝO��d՝3��m���j���E�,8���%$��$dU��p<�@f^|uԸ�S!�	eA�ћ�4�4�D ӏy�֙)����t����ɀM?������]�T2ю��#����,��i$Ցp*/�I\��8A�HZ�t��<*�-�cGL�':�ĺشIЬ	�&G�I'2�)!���>aϓ��$�:#2 �'*"\>�(������a�
�}KJ����F,���������ɽ�p��-��{�=�r�J�G2�.��ʧl�] r��:ef���/\�{?N��Ojp�"#ң|�� ��ͥ)&�D��%ܺ��H�N����%C@���gb��Oڢ}���ok��Q���)Yf�}���)h!��ȓ;�P�B(7t�ФA&lU���݇�	��HOD%Rv��#du�4ƔiU��Aw�UB}"�'�j�j���a�'�b�'���� �ea�%Z�Cv¥x�׮#k)�v`�2g�ӟ�C�\�f��c>�O؂�C�`Ġ��!o��u���4hv������P�ծ��9�q��'�Z0bI�)9J��V��:l�@�Z4�'��i-`#��|���dTA���uFKR�h����0Y!򤈐fĥRP
���xe��@�'V�ɏ�HO�Gy�#)	�) �%h�qj�	��j��b!R��'���'���П����|*3(D(�YI��^" �A���x$ ["gZ�g~Z
�#�Y��l�p�H>��X⨍,\�勔G_� XXl&%k�1���Bj��D���_���J&H�O��W'����D�O�=����� ,Ό�# 8z��M@��3�y���C�
�@bi��B���u5��y"%�>�*O�:q�Kp}��']��JF��7���O�%�u9��'T�8���'��ݗ�����-[���p0Ɩ*]*��0�3� �8 %V4C��i��ҁ9��I��$�>��9��Z<g�>�RPA� �00�,�k����iK0(rh�x���,�p� ���	 K��'@�8X*���G��<�\{�/¹Oec�P��If�5�o/1���
�#t:�"<Q��4���l��q8EF�#U��ȡI�i�,�	Ay�LU#k�7�O�D�|�r���?��!ˮk��PPWAl�d������?��}F�h�� �lY"���'�o���T���&\��-��X��"�xd��L%h��5yc�>Q�7y�.Uj#�F����L�P9���2"�ي �Xl��G2#^`[T��Y��[�dG2�yӊ���O�����P��9x& WB�T%��0=���Oz�d�O ���B���0�8`�T�1+)P%ax��7�!rj𫄢��G�x��c�L)e6�hz��i���'l���.u�><���'"�'�bem�}8cbFM�m���ʹWR��sAE�R���D\DDj4�޸#T4x�|Bף�%;��I�(氼���S��p�	�J�B �����"9$aЩ	+~�R�>���[�BG�$���:8�(kb^�*2!Y k*ȕ'��
2��Oq��'ϔ�"�HN1��9�gQgh���':��p�R(?G8؋%뎔8)��H�'��k<��|�M>y�P�g9�$J���<U�lh��G�<�`��1��p[ӌ4Ze<�qBEB�<AF�f
@4�!��~+�1@���|�<���&}�A	�셆r��Nv�<1@��� �Jٴ	�rPdY�y�"�N�H(6�.X�蓨��y2ǜ�6]���F��{���ѣ�Е�y ���ᎈ*nи���/�y����x�����k�=�����
�	�yb�8GvR�
2�:BD��G̒�yrA�;V���A$��$:�
�j��k?D�LA1/�X�9a� ;I�^��':D��(3$� �1�� vL
�7M#D��e*�b�B!��J��S�<D� ����qo�q�e�J�6��u8�F6D�̐ge �|�n4��%����1�B"D��� K�+�p	x�C�L�z	!��-D��B*�29cb}��,C5 o
���j'D��{�#9!x���ԙF��q�`$&D�����,d��=p�G 5o�U�$�"D�$Hժ@�7��a�A�C�$��E�K D�܊�"�O��	cŋ׼H6tE���<D��R@*�f���!��^2pѳ%J<D�� ��f�Q�g��aoRe���,D����!�K�l���RY&�� 0D�pȔ�R�]�� �*C8B���P�C/D����CG����_>��< @�7D�����$a�20�w!^�B��Y�6D�\*�X�`�ƜѦ�^�#l��O5D�dzB*�y2���L\�'@F؋v6D�ܹ�́0��1B�AJ\�*�2D� �� d�:��`��R:$�h��%|O�]#�KR�f�Z��u �5QC�?JXuz�":�FB䉜I\�X�R��5e��I����%~ixc��zr�O:�&p;g![�>V���&NH��X��M�L��%�A"OP�ʠ�.(n�}�CBR	I�DAt�L����Ϸ�$�� C�#}p3O� �1�@���X�V������15��)�"O��q�B;k��` H L����៴��!FT����!(8���hO���D	�$���hR��?3��:��'�
��c�������C�x������u�8j�ɐ�R9�x�sH+ZQ.]��I�Q;�"��]<`\��!!$7�c�hJG �-!}F�ZT��?6q@�s���O�<Bp�T ��ҥ\N:(S@I�6HC�I1O��H�`�7Rh����HM��Љ�� ��}!�.�.;.����S�O~��*&bTR��3j��s��ɠe�B䉾O�V���*`ز�9T�
m�����'���@%��ժ�R$mݍY�g �]	�G+Ԕ9�spL��$�����7��P�F�x: D��l�g��bRl �W�:�a�e�Ц~�F�*
�}R �����I�� AGeC_t�I�>�T�=5��hC�F��&0&(�u?���OK���'���l�y��99d�b
�'�p	�eofLJ Ӆ��+-\ �e�~Vq"¬H���ʵ������hg�A��O��j�82���N-��� ;D�L�AE�0����A��856�˓%����DZ�jm��/[�*W�8����>�#�FT�	*��S=��ѐ$��~؞t���FZ����!V
��B��-E�<��E�����d@�i�H��V��q\���	-W��3���%&VAW(С�0c�p`�4\�	rĀ&�Z%,}l	4?"j�kSʎ&����M�;�!��L�^.$q�S텥M��ɢ��P`��%��J�zU^Yؠa�J���O�O@$�?t�:�ځ�� .l)���,$�B�	l�T��-XE�6���f�s��!�J�l:'/�cfjT�;��}�$����'�TA�q��Wf�a�S��=v4�#	�,��4��Ȟ9�Ԩ��\?�|��J�VC>=�&�˞����'!�c1��3�p=�RGјw��QpR�g�4q7mR�p��L���[=����C�Y) �0�u7�;4h�P��
<�rYВ�H��y�N-F8�X�f��`��d�
@&n��`�+��+6��
�T�a �Sܧ��S:r� 0aA$\��t(��&Z�!��.g���#R50��򤓮Ya��q��Jb�0�S��a�:����	f��p@ˇ��d`tѣ�(��z𢬇�:tRN�5a�:r���4��©t�I��e�'k瘨HU��J���p�E0s�R�)5�ۉs3v�x�:�ɬ�^y��*�%WA̠H����Ņ�f�x г"d%�T�Z�w�R�r"O���6���TA�tZ�ˮ!���X ��/*IJ�]��:�Dƾ%�>-��~��X�ρVm��&��J�l���w�⸳t���dB6U�E!�Wx�p&��(�H"lC��}rc��?�>�4�[�{��If�Ñ=cԤ*�u؞|:�o��%�ᣢa���z(k�L��02��2E�~�`3���v�(P��	*:��e�׷{�:1&�ʓ+��\{v���t}i�7ta0@<�dN�.f�c�6i�,���y⁜�}ג��6��6����Qj��Ȉ�s%�.s�1k'A��|e6��O����NF��-�cj>O �s"E��!�=4e�%+	Y�i@a�E�'0��@U�H�2��Y�'� <��𙟌"��ǸK���jW���؄�"a'4��$��.3*%���6:]@XSUF4 ����4�J�H��h����ay)դ["�[rŘ��8�R#ˤ�<Y��!�<s��V�	A"��pC��@��y�!%T�AP*��5F9dDY�ēj��U�']6t8:�LJ K��'�t:3��`V�3Q��
�ɂ7��J|�`{E:5����<<CvC䉽FH�@��X'Ny�A�Q�����h2��94��t���	�]%H����0�3�dȅ_�Y:'�)�|I�k��
!��O5������([V4[g��6��S凕i騉A�mU�5f8:d�'7be6��<����߅����˓9Ѐ�'�K�K�Zx{3�V�,$�7�ܢi,�D����d��u"O�q�C&�1j1TIң�k;��C�|��,+�"�A�z�B���	pɂ�N_��ܸ3b�η� X��'��U��I���l�
"z�ܴ ��b6����S��M3s*��J
�y��GP�w�(���	Md�<�Ei[$e�鰑�C)q�1�q*�vy��VN%HŇ�!9��{�*�)�2�Pa�,��C�I�1�\�o�'fX"x*+��R�dC�	4e�:�e�f 6q��'�FC�I-�<)���D1��*��{pBC�)� T�X��-���j�p4�,�E"ON����o��� $Č���q�"O��hB'��E&���(��dZ�"O\�����7��#q(F�(��	y�"O%��)�Qܔ| �� ����h�"O�ES*+U�5�-�J��p�"O(���gHr��@���چ2*�Q"O`��iOUH�����綼I�"O���	az��
�J���=��"O�	"��5�lQ�D�׬\��V"O��(��h�h���+�,zQ"O��2&]�`��V�(ۈl�D"O�4�!.69�2|�0��2F��M v"OV`*GG�rD��c����J��u"O �2�f�+�
q�f�ݱ=�vd�"Onт�	y�,x��^_؈x�"O��s�N�}�>���I�����"O�q�.��{�4� T���y#���"O֕�FC�*CܔR"�)C<m"O����xt��
��l���T"O�h��Q�A(R���#�.���#"O4�战el4���&_��,ig"O�Y�V�]r�Xz���4n��tt"O|�� YS���u�2$�&�3�"O�e�ĩ݂��`3�*W�^a��"O�P�l� ee��
��� К4"Oz9hR���xwdXx!/S�2�z��"O`�ʹ-Fn���ݖJ��z�"O�R�J�6��Mc&�I�@�T�E"O����#j�m�b�Z/�r���"O�9��L�lmµ�T�(G�z�"O� KǠG�2��3��*4�H�Z@"O�лe%��J��xP���
!�(+�"O�q��I;6l(��?F�a��'#RS�KR�F��Coȯu�=�'W�B�X6J*(����%l���	�'� ��ѣA�����F�>c��Q+	�'	��z�-�~��ېǈ�i0�H�'
�*���Z���Ʌ&yߠ���'Ղ`�MY'"d�HpL�]Kȕ��'f*��GE�&(���F�"�X�'s&���d�j�<�G���DC�a
�'�.�J��B/ub Eඨ�ID�p��'�Թ��mϑ(L��ACC�A-!�'N��b$�K�o~����x 
�'�2D
�F(��4(!"Ⱥ�ؤ�	�'����m�8��J �Ѵ�@�)
�'r�9� �M3p��K�h�	�'x�(��i͢h�bE�W5v0�	�'2�ᡱ�_�G��ɨ�'^Rs����'�%;�N�*j"�����K�j�
�'�$��"�'��Yp��yl8�nT?H�f�S
�p��a�/O�) vj�<`��A:�N�4<xp9(r"Op墲L�iDق���v9���#�L�F����"P{��x�R�w��
���y��]4����/�p�>�r�<��e���s�d!���
"�PD� �
=͎T0��.D�4�qBҔO�p #�`C��*��ɖK�P��ɥr�X�-R*l"��з�Ʃn]�B�	l�H�(UFҸ'�v��&+C�pB䉤V�ڈ�@̜)��m��$@1K<B�ɷz�Z�XVfPB~eaTe^��C�Ɏ{�t�J3��y�cH�&��C�I.QҬH�g��h9P��p�A"w~C�)� n�(�.��Nw�́�IG.����0"O�rl��}렀�P(נ%��	�P"O�sO�$�*��UM]�&�4X�"O̼ztg�[
 �s̝ U� �"O�-��4_Cy��A�x�$<�"OnU2���X�`%�U�Cr�eb�"O�}(ᬍ�mR`�2�X�XT^�a�"Ob��r�A �-�@n_�QbŚr"Oʕ��C8Y��JӦ� WlѨ�"O�M�U��E�T�Ƥ<�Xmb�"O@e����}��l��Ňrߞ��"O
A���X�P�D��2&��h۴"O�	��g@M��ѻ5�R�ۅ"O��Ap��#$��鈖�S?V�~��Q"O��á�E�w�@��e/ �n3�Y��"O��j��/��zs�R�{!:\�"O:h3C(��#D2�9��X<x(��"O��A"_�Q�Z��5
��i�"O��*��FWr�\ZR�9n�0w"OZ�3g#��:��a	��M�0��"Ol(��a\�X��!�n�*m�Fu�t"O� �AX�imt��W�T9�С2"O�lQ0�(�K�Z
]7H��"O� ��]�H`-roͺR Iٔ"O��)��>���σe� @��"O��@T��i90�Y�U�7�(e{T"O��+�eM�@�h��P�W�Z��js"O$]�3�ބ/ �����,��<˱"O�0谆��8��1�	A�[��ٛ"O����&�k3�Bq!����0"O��1���2ET %&��^	�`"O���U⚽ �Bt)p%
-ָ$�"O��B2��*�H����ini��"O����蚀��YÃ�Qhj\5"Oz�9�l�)-������)BB�	�g"OV(�`M�es�I+ԩǢB
�pq�"O��s�X�@&��J?\aG"O.СF�_�ISh�5yM��+"O�E��HOZE�5�0c@hA5"O@��ԩW8���1�5v50��A"Ox�Pe.�~���⋤v�X��2"O����N_�R���@M�_p����"O�< F��%K~4��B�(�FP�"O���êP�Ml)arJO"c����"On���_�y�hL�u��7�n��Q"O �G�Rg��c�W-c�h�b"O��@J#������%`���a�"O ���C<h2B�����"O��S�e�(��đ/�dd�ya"O,��Q�Y$:1j��؀c�"O�8{dG f��P���	��Q@s"O��`���y,= *	����"Oب*t�E�(���V)����*�"O0��.�~d��H�Y�ֽp�"O�p�jT�"�Tj��ۗ=�lY� "O�����=KPL�P�'L �<q�w"O�a��*�e��8��ʱ?Yl�5"O�=ä��.n���Ī��)�q�e"O:��%$u�Hz��Y�!�Rqb7"O��{�d����H�I��p5�7"O╂�b��"��a���K�w/d�QA"OE
�̈́�oU��%nD7)��"O:5�
ˣ-�%��� �:~�s"O$���Mo��RS,ſ~��&"O� �H�#�<�B�t͎!x�<�"O��8�݃S��J�P�xp��Z�"O�P�L���1ɛ�0WҘx"OD��͙)}3���q3V0��"O$�3 �ؿv�^h(���La�Q"Oک(TG�V�Z(�M�!�)`"O"�C�.�'B�&��fA�m�H܊e"O�ɱ�mWp���UF�.��A�B"OD�s ��)c��u� ?����"OL�d��(L���֋�yjPhz1"OL�R ��;tRL+�ʘ�{^�1:g"OzA����:�\�Z�J�/@�\�"O��3�$��*����îO���a�"O�I�,��ejД����_�^�*�"OĽ�R'�|}�(��B���"O|� ��� �R��g��Ef24�%"Oԁ D�_{�C%�K�dN¸��"Oę@�萡M�ڝ`CN$T2:qkP"O,�YP�#L���ȋBA�09w"O"��LQ�W}t�;�FG�rP��"O�50WdU�x�ZX�`h�&m�(\S�"O^yy a��l�xd����s�����IAX�
��ۅ-��pc��T@���3�'D�`�C �!N�	#VI��{6I�'�8D��@���GmV��)܆S�]�4D��:Q�c���cR+ų�XZQ�>D�`Za��7	]V�8�����u��8D��� V0S���#�(ջ=w�]��2D��Y�'٩RGĀ����s^��'/D��q�ܢ#d��pA'�,
B`Z�,D�lb�P�n(�jfC� H�
<Y�5D�b i��cM8�Bc�ɤ""�p�m/D�(���P�^}	ԉF��ޤ��A:D���æX)�1�ↆ�t��a+D�,����~킭�6�(qW@�jb*D�Pq"�X/@:DO�� cDEK�&D��Z�dñX������R���k(D�p�DL�f����ڸ{�@���*!D�0��͎aN�|qt �D� Ƀ��;D�d#�Θ-� `�}0�[�	=D�\"t킍[Z©��W5`�(s���>	��Z3P@�m��Ι��@\����B~���+�ZZ��	�D?Dʢ���y�.
�|���S��;:�҄��Ý(�y"ʖ�2�
�� >�(����y�"2:D ���&=�l��aW�y�Zh6uҕ��"����U%��y�e���A#K�hv�xO	�y��Z�G�D)�LT���WhW�yB��FTLP�ee��* if�7�y���\�ʨ��)0g@�Rn��yrG��nK�MŌ)R��m��'���yB鐌(�,p�ЁY�B���8�J�y2-0�
��`%9a�H�%���y��'d�@�k]vX�Q�a�&��j
�'g��p�E��(��9�Qh��[�=B
�'CT���KɟD7����B���HI�	�'B�(#���!���
S��6b��	�'��I �q�Up�@>"ܜ\��'��q �(��Й4�1-F�i�'�ԅ[�d�'g2����3q��r
�'*��z0�ӳ�\*��<]��X
�'�0��7dՒ/��ݚs!ďJ1(y	�'�����	��L�Q#R�Z4���"O� ,�d,�	b��Q�3=���  "Oݘ�
��T��=�� ���%"O��@�'Hf�8 �@�����"O�ؑ�˙"?�����T�9�D�Xb"O���OR�����C�A q��D��"O�4��Cر-��};U��<~��<C5"O)�B�X�l��ZЂ����tq�"O�X�5m�TG���Ā�"O�1YT�ٞ��!�Y�T�C�A��yB��eL>�bTc@<`���-��y�*ğ?��, bHY�.��0m���y� )�Z����ff��r���y��F�.�@a��[	�0Wo��y�A	4K�����gL�[5��y�)V&M�B�d $ub��y�	X�A꜈�MR�OB:e��dL/�y�$[4.���j�<H��șB)���yBB[Up�ex�"��C.�PI�'���y�W�v��} J�6���i'�Z��y}�
lZ�˙%F��D�k��y��^�zU� ����?}n*���2�y���+p���Q��H0/9�a@�y��P�$� ��5/�5*4�ϙ�y"Ʉ�xR�R냩zq2��N���y���H����+u�mS&�yb�Α)!�V䖓\dx����y"�/e�ީ(��'U��(����yRm�"�Y�	X�D��-��'�*�yRA��*�X����K���ȃ��y2e�%�j�����*3�H�>ѴB��b�f�Ckύ-��sf�.�B�:V���u-ӟe��H�DB%
'�B��SmB�;2aT�hz\#DյepB��,}����C��}r4�"-ӆ*�:B䉄,J|�2��4E0d�h�;0B�I%R�	s��.3\�х��C䉏^VJ����%lRL+�V5%֦C�	�N�B�M=oTM�S�H��C�I�K��E����O@�� �.8C�IB��]{��{
x��B�ąS�^B�	8�.�K�'g�"}�"U�3bC�I�I"Ȥ���K�}3�Dd��#G�TC��,Bw�%d ,~�����ѕ`OBC�	�3|䝲Qc[�C����O�1�NC��0B@("3�
���P�¶q�PC�	8=��p�@��i��)�e@�K
���ȓ=�؍����:��,�wI��7K �'ў�|�K�9�v���$J�@��Ѐ L�v�<	Q��gFh�P�ɔ~@L�'ap�<ӆ6:R`
BBS:W�Nm�ȋR�<��� K@��r60OD�!f��%��x��C�!N.����<^��ӭ���y *�`�gI�U�ܹcÅ�y��G�KW`)�&��"�Ha�i���yB��aJx�������� �,�yb�8\~�H8�&\����B��S5�y�F"ʤ����Ƞ�-9�y��6{5��A��U�~��(C nR�y����30`v)�K^���J��y�M�w��Mxg�9Ԩ�S��]&�y2B8t��ك�\>���	�Y��yo�&D>��l
1<zRQȖ�C��y��8}�Ne��N̚<��lbƂ���yÄ�L՞��2&�-��Yɥ�:�y
� �t��M����Pf}��EAc"OqWf8/��Y����5\��H�v"O�x�tB������:��v"ON9+# ��'v��j H��H�zA�&"O����&>'�m
G'�
��8�"Oܬ���\<<�	�/O%�����"O�� �P�8�����oȺs���y�"O� `�0S��@�哺i���K"Oň�Ί�"¸$����t+��8C"O��Ś�W2H�;`�Q�m8X�"Ovȸ�aB�-��]	���?gt�q!"OVMc4O	2D"i����u]X�g"Oj� ���>�����cx���"O�sjٷ	^�;gŊ&E��3f"OqXv��K��i�a+^�&UεA�"O<�!@�\��L�p8�|�"O,{�M3d��{�
1Z���"OB� *J�1/�Q�T*�Bk�2V"OdJ�+��A
��y�Ɂ4\T���"O��'ID&Se����!R*�+�"O�Myg�Rq���s�P�]H�"OdD��Цl����gV>K���)"OhXcε�esv�ŏ � y�"O*�`�JM�!��&�t�2p"O�i{a�
,���A�$�I��JQ"O4��!�:�v$KE�:��I�"O
 	v��%W�4�ؠD�-�� A7"O,��W�ؠbi�����?�0@�"O������5��8uG�m��z@"O�Xc��T:_Ä�Q�L;8`�U:�"O8%�1h���tX�^<Vs��"O�<��c;�,u�r�@	jPR"O�d �	%�z���˟GS"�8�"O��@5dS5&˶! �B-wA�H�"O�����q}��	��$*R��D"O &�Y�k�4A�S.�N��p1"O���8��u�/
�H�"O"1�Rϑ�N�l80���/�i��"O�l�D��ZX�mN�Z ��@�"O��Bf�Խ���X���^ )�"O��(�*ԅ ��,U-���Y�"O����6p�Yː!exw"O����A��OA�gdF�����"O ��֠�#HZ�p@�7��Ũ"OA�Ä�-����H��z�Ȁ�1"OjH���'t�8����*6Lyq"O����[��	A�A��0��"O��TmV#�D9���]�<�z6"O�q����r��07�y�^ P"O��؂n�)��q#�U'"OT�����VE�!�'��fA�pj�"O��x�T)�T�,�4{0�@r�"O�i�#��6�n}`#D�--(�@"Ov���$o��z�#��(�Б+�"OJe��aB��݃�A
�����w"O�$Y���/��%��w%:@�w"ODؙ$	�*�tX��v��� "O��Y�a_��2)�٧+����"O��ɷ���Q��l�}�℈�"O�lBs��$y!�ԓ��7u"��u"OL|QE�"�E���� j��U"O�� е31�9�ԅ��k_��z"Op��Ck�:��D�#�R6(EH{�"O�a�Ǆ4��,S��>`2(�zr"O� ��#g"ڵ^�\��C4\�ő�"O<)�Q��'�v���AC ���Kw"O�4b��W$1'�0����*-��dC�"OP����|^����垽<4�P@�"O����ћ���T���}'����"O�)#�aJ�6T�(h�A�;)DH�b"O��Wf�K�d
t�ׇ>%.]��"O���ei�b�"ԓ�()
2| E"O�m�4ĈF	����(�9�굡�"O�����
Z�$`s�aZ�B���P�"O|t�DG	JmX�3� F�t��4�"O�$S �̻N�x��c.C�y��9�"OB�16��GB���K'^b�9�"O�����3eE�ha��Hd"O*%8��̂4(p�w�E�bU��"O��9�e����HJA�ߖj�8��"O��x�	stn���!�.��k"O�eC���F^�� ��U x��["O0y[��E6-2X�U��]�|	�"O�q(��F��a�Ä"IZ^���"Ot :b��U�
�?V�}��#Qo�<yc㔼t�$���;Z!��E�n�<���/Cg\��5�H4 �8�)1l[c�<	'�ˋ��`��3E?|��g��[�<���=<�r]�&f��c�B��ʈM�<	��@��Qh�DP�@|�)��NA�<#N��Zwi٩`����OU�<Q��߫
5v݈0��)gX{�-�P�<��
S���j�LG�
i��Bc��M�<�e�ԣ�`@��\�-�hl��/N~�<�r�J�!�z��2�M�kҖ|�R�Q�<����J�P�o٠>�P��M�<Y5m���׃��(p���m�<QS���(a�afԱse^�ۇ��S�<I��@V���甯oq��۷
�E�<i�ʜ?xX����� �i��@x�<���Z�m����揟1gn�q�2�p�<�1����}�Lͪ_]|�ygD�B�<IPL�;O�p2��.�|q�"X�<�$ �к��2��/�
ݚ-�|�<�V�J*;N�xT�[/`,Z)�eoS�<��*�
}��x�D� Ψ0R�)�F�<Y��
|B���"�t~�Y��LX�<��h�'h@!@��d&.l���KQ�<���K�fĎ��$d��F �K�`I�<��d��@Iژp���;sz"q��k�<�Ā� `���PRn�4` �m�0�L@�<!��*F��X�@��P��3��y�<��˛�j�6�����h����x�<�Ո;}�����R�q
^<z�ʕx�<��M�(���h�/X�I>�����v�<a�&��d�r��t%��8��*���u�<1� ��3WԲ�n����亰@�p�<�#!J�b�!�+�b�B�j�<��oķUi� r�'�>��QP�A�<� �ýL��� 2��S4��YӥT}�<a �53�zx�`�P�?ݢ��ƞ}�<i&�ǰCX�����l����Fe�<qc���Sm�K"*�� �.!�V��w�<�c&°q�*��N�!���i��t�<���";�>)5fG��	@��U�<�Dk���L�����euF���g�<���X�#�m`�*Փ	�t���z�<��ǆ<5�-���>p6�*#LSq�<� ��Pa�'�~����B�u��ٺt"O��0��Ԧ;��+Ae�-D>Rbq"OL§`S/uRX�eP�2����"O ���<u�*�c��_n�2��"O@qb�K�M�I��M�~q,��T"O���oҞr)�dx��).��Ra"OnM�b�7�T5Q�n+�vyx"O����,���	���yT"O����OUT�YL� E{�yXb"OXX!G)T�����+_h�Cp"OP �@��'�#W Y6A��"O����"�pғ̖6~�]�$"O�0�L��F*F�q�+�K�*�{"O��"���*��W�7��Tyg"O$}22f3k\�Q6LC�X���$"O쉐�i���2c�[�lP�"O�����F%v��#%.8�1X""O�̊�@�!sSl\�G*�/���s"O|�B�5l���q���{�i�"O�x3`�])N`�5���[;,�SC"O�X�l	8M��Ĩl�	8���YP"Of `D�>	
 !��Y>��4�"O�9���]24]�-����,��"O�� 
�!cXb��|���R"O6�G��7�L|��O �J0FѺ�"O��Q�H2�̝B��O�TN	ї"O��(���9XF�P�Ϳ[ۖ"O�I�X�s*����O�X�z1��"O:娚�;� ��D_��z3"O�}��F��&�A�dEܶzD=
"ODu� DB�C�	z"yԲ��"O\3w��*:k~4�4JS~ŀ�s'"O2�"�gK��&��2IH5x7"OfݪU�ѵy���h0�F�z�"OڍS���e�  ��A�z4�I�"O,�0��X2��P>��B"Ođ�Q6]�,��V�Ƙ
	^��"On@�"�4�,=is%��6�@`"O��îL�q���`t�6S�ā��"O:�!��+[6~�qR+8� �1"O�5�b�#u
1Q�Ȏ�o����"OhQj�/ڂaި��R���"O
l9PcS�S ��X�FB�wwP��T"O$x0�e��D:x��̏,s�$R�"O�x&�U��lX�Cʹ�P�:�"O�m��#�'p-�U�ĉ�7�8$��"Od�sBB ~Ѣ���P2�~9`F"O������0:jz$JD(��w�"O�ҨD�FHD�M.�9h�"ON�*�/��Svq�K�:W!�!r#"O~�h�gO�WBl���锉j���S"O���L��Q�ʡF>[㚸�6"O�E�@Y8������X$tј�"O| �0(�(#�м�� D�&�r I$"O-�C�/	ߜm�ŀ[>f��5�"O��01�7p�JT�_���0�"O>��k��'E�A!g.	�'�$ h�"O����nؙb� ���m[�% ���""O��!�c�#8�@IZ��M�g�]I�"O�}ZW���ֱE��
X=�q"O|������� )�e�#�
P�"O�x�ajJ.HI{d��D�"O���Ѥ��3HP�9��5��"Oʴ ��B�LDJq@V'�/cs��"O�  ic&��L���1��;(m���"O���$@�´�w䟨r�4��"O�a���tP:&-۽*R 	)�"O�A1�N�Jl��`QK
��(�"O���6KE��ۅ�Թ8�
�h�"Oh)��W�$�P;�N T����"O�Y���.\��kA���T��"O���E ɘ ���W��a�-j�'�1On�����C�PI��g|\+�Z���	_�Ț ��{�y�B���'Ѵ�:` (D��	��2D瘼!��5?��b��'�D'�Sܧx.X���%^�\�Z����8.�tńȓB�-s�F=#�zZLC��m�<�s��AvHI�)^�T�� ��N�c�<����K�DA�q��E�$�RR�cx��GxR�͋
 �`/��&�z����/��:�S�DmGTOt��Ӂ2(,܉��P^�<!E�Sj�\�{VDX�MO(�"��~�	��x��c����dĻ:�L�G�]�`�#��$c!��I��)��o�16� �ㅲP�!򄗸�Y#�%2"v�=�v�A�T�!�A+U�p+�&VV����L
3{!�	Q�l�zA�wPrC�둞m�Oj˓����pDB^�v�$����d��"O�˥��=g�����ս*$��'�Iş��?�}�r�^�1"*��a�dj�2DJ�L�<w���l���.،(����i�L�<a#`�/k�6�aE@Q�rJ��²��a�<���?f�̱V�Y&-@����`�<Q�n�GAvh��!� %o���t��R�'Ma�d(M�.��52��CP"5���ɭ�yB�:�d�zD�N�;�rqi�� �y�T�3���*v��,���ᦋ �y�
�r�ZQ��T*Ċ)�5H��yR�_()��IK�a˗�W��y�	ν}� Q�2	�	�t9��]	�yBʤ@'���a"
��@�Q�֗�y��W5���uR� uA����5�O���*�!``�D���#���"Oz��Ud�4��lA5�O�6�v���"O�M"��τC�R���N!"֚���"O<��'��;Bjt�q�C�nV� ��"O|�p��ӧl���ؗ͏3����"O�E�ޝL7���̔�4�~���"OtHQR�+?e|E����w��}I��':��p��B���+P���PG�ֲl���0'>D�ܚƭ_#^��p��dV]��T���:D�LH�NVp*bIG	g���0�`<D�Hx�[O�TrV�ĘM�2�%B9D�������u�@s�'�Ep�J
6D��{'@X$ 3������{���d�!4�0c�k�['�Y�GLםq�,D�"�Y�	Y����D%F�j<�e�߻ .�<IQ�)D���A��k��Y�G�]lN���(D�t���)k��� ހ�xD	%D��1��ҷ^�̅Q��ܲ
r����!D� *w��#l����!Ł1㬵S�.=D����J#S>�xA(��=w����9�O����n�ܹa��
<V:�P'i
=j$�d�<����	�S-�Ec�aB?P��e"��6-!�dѻb�jE�rDO�U�`�2a�H!��L�P� L�z�س��֒!���5\�R�ɐ�ɾc��蝷!��>Nh��rW�"J�Z���.9V!�� .�pbNp-f�����D���'���4��Ȅ.@�@��GBd*y���OTB�ɔ-[N]x�㛌q~P���ywB�	�u|��"���O�6P�鍄z|�C�9G�`L�b�2�ݪSC%x��C䉫m�h:�^�ĕ��∍d�B��*M���@�A�|߶�*T`��?o�B�5,���Q�
��=�'�E�B��B�I�-sHٲ��*��P��eW*\�C�I�y�6�;��5`״�s5�U�<C�I�A�\��a'\M�2��,mbB䉃"�J�A�Shl��>��B��\��#�D�@�H�*Z�s �C䉏L��x��JP	�@���X���C�I�|X��"ֶ�Zp��W�]`�B�9}	��Y���'�|-����fkC�I3!}����Q�pI��H�-�B�ɣA5��QAkЖD:���ŋO�B��;�y��C�|� �8��D���B�	6����X���id�U
[�B�	���� B��$�6�"+��C�	�^e��兊+�`�ĀԸ�"B�	�X�x�s�4W���bo�,��O��=�}�7d@�K�cѿ��]2P��X�<��^"L�|���aC�B�=rwG^S�<��/7���+�M��-��@��l�P�<�u-Ės	�(��2��d��J�H�<��-Q�MR¡2�,�*\=Z�7#DE�<1Ɓۂ?�I����5��)��@�<�E��Yt�8C܂0}�,��$��~�<Y��E��� pt*�s����|�<�2gQ�x��%�,ѥp<Ƥ#m�z�<!�
C>J����b��[b�<�b�3#��M����*�����T�<�#�@� ��Y?<�CRj�S�<A�mήD}�� ��m�\<����x�<!��>v��RET� �ԙ:{���]��k5GV�&�����g�R ���ȓ���xs��*{�t���9 ���l�]!&���a�α���J�[��X�ȓd�mׯ��[@�`y��5=*�������(��6S�T���+w���ȓH� �)l��H	���\ܾ����Je��`�4M�$��S�[�5	R��ȓ ʹ�h�މ	D��#aђU�	���l���a�X��ć�3z����ȓ;Z�I�$&Ȓ����_,&s:-�ȓOz�q��߾	(�	1��	�����m1���!�48���BR+
�1��C�ɲ-�85I�m�1�Z�+��74[rC�	�
H#�*�k�6��#GD-`S��$�2:�ȱ�#��>�U3Q@s�!��57�|�B�U�ڨQ����f�!�ǺC$�!��w�|�%c��W�!򄄊Mz.��u�9$R^�I�� �!����l<cQēG�r��b�J�!�ƖRis!� �M�"�[Ak�&j7!��ЁX��U'Gb�Z� W,��5!�d �N��^%j�T���3*�O~��d�'E�0�D�˔%�~�Z��ޤD�!�dR�%�ѳ���!y���c�_�!�d�F΅���.q������.�!��\p�8��9od���`���s�!�,#zthF�K������q�<� ��!/4��!�cP�R��:0"O�@�V�������>�p��|��)�Ӌw����]3'�9���A!6C�IXhը'#�.�p��g���}v�C�I/4����@	�c6�P�Ԉ2�C�	 U����"�:,$E0�i�3b�LC�	�!=t�� ȕ�\!�rsO�:snC�:C�yc��YE��y�hKD:�C䉿7���q��庐뉙a�����ɃZ(�;�\7H����+G(l�B�I"�m���7�y��GD�J��C�I<���"���B�u�Ъ��v�B�	�d)��*Z�r&���3)��C䉃K�"�1ц��m��	L'&�C�	=��s��6`���!�֕g�dC��6u�fxҎ$��(ҫ]��p�D(���ON�?�'^����6O��H��U�C@&$��'��8���JR�U�e螨,���P	�'�D��K�"�v����#J�	�	�'�>����@-!��A4@۹c��ȇ�3�ʥ�KJ�v�=��"X*Q�����?/��1�.8:��B����=��S`����O$�D����ޗ�$�|��I�b�@Y�G�� h8\@s��ׄ?>�C䉃'���Q1�H�3�٣0�U (C�9 ��i�5IX�U��R���)5C�B�(�.���T�r_���v�S�JS�B�f��vm��/�NeK�,�?_�B�ɜs�8%s1c�V}�R���VB�	�x�T8�7�G8&��)DX-H�C�I�	�B�����@�m���CL�C�I�X� pYъ�fȼ��!J�B�I� �z�b��C�m���i0�ވvB�B�00�T���&��Un��넭�8�^B�ɇ4��X0���"_B<�B��=�0B䉠|�pQ�5~��8*��\B�ɫ_'J�DK{b0q�0� i�B�	$l���L�}l���L^��C�	�&��2��ٍ$p@�\�,B�	�-n�i����~����([(&jB��?�و�H�)��Pɣ�Ʀ5�0C� ���Z�iA��T���I�C�)D�LP���G(e��jާ(��C�ɱ_!te� �L�I3��� [���B䉱t8Z��D�Nlqփ�80��B�	9����Ɨ�}�����;G�HC� �<Bg)��[�� �+�� w:C�	��%q1��7R9�TB��U=*�C�w�d<�EƝr	°SSbRP����-�p�D!��( U v�@͌�N���ȓ;zV�3����DɞI0�CFj�^�ȓ>��v ��UNi��0j�4Єȓd�$;rL�a���G��	���ȓ�d�[:[XYj�!�'3�d���		DL�2md���`��{;b|�ȓ:s�-��`�z���1��|�
��?I���� a�V�ZQ��KB���E�n|ў��ᓊa����&��\���5`C�\l
B�Ɇ	�*�B��$��|ң����C�/[x̠W���pG����KG"a��C䉭;^��'���r�IH��-|K�B�/V��u@S��PU��#F"M �B䉒O�4�Y��S�1x��J���O<�=�����U'��e)��	�p����K�,Y�!�� D��s-K���X7��%F��u�"O�(�h�(����e���Y�,"Oҽ1ϝ%v d9���/v��tR5"O�hq$$��* W�?�PYu"Oh	�e\�|��A@M^	
�� ��"O6-*c�A]L�yC�+O<R�(#'"Ox�@�M�.Մ��sQ���"O~�S7/\��@�$�AE����"O XӍ�5��y2���sD��D"O�,�'�\%Ӗ����X�,���"OޠiBo�:M��R푩)�R�"O:{��Q
�;�,�6uFLj"Od!R�K�_��l�q��6�PyR"O�Q�p��\�(E����4/�d�"O<Yɶ#�2~ �Q���'"O�p���i_ڑ�8u�R���"O����O"u�`	4̊&.��"O|�C�j�����+�R��2"O����UcWR�!�n�QȎ�1O�b�#�y�Bp�+�;bu�Mc��O~C�	�{iR�h�ꏫ�����g� >kFB�I��rTs�� c�*DxBc�C�	r��H�1*L9�oĆA�B�	/l����c�@��IY�I��f\XC�g���$��
I��[@@O�*C�I�(��cQ]K�Iv�ߚ(�B�		}��ɪ�D�P�J�y%�[=q."q��*!`�8S�Ã9�����'��/q@���=���像;y܌����}��Ѕ�I�&��d��:YR8�����
4�H��=���s�x�"��0���䥆�?hLtQ���64B�:�LY�p�t��ȓ�䨊�AG3>��E��W	�A�Ɠ@(���H3'b};��ڧ0
���xҋE�e��v�Ɨcr�	Q j��y�G5W:��!O^$G��9�GP��y��K����sH<�� �ڃ�yR��>=� ����44:$��C]��y�$W��|pǤ�>Czf�L4�y,ǉ%2(��-]g����Eć�y��߲>qR��iX)r��� �E� �y��I#Eu��{�Γ�hz��T���y���j��Gr������yjD�gO��q���cϨ=ʷ�O��y�DN�����nBJ�f��UDS�y2oW��z�����y��h���y��9I!J]Y%��p�X��V��ybC �|�Zdr�iP7g�n}�a���y�'��r$H�M@�W�}x� �y���i�1Z�-_�}θ`����y�NE�xԜ��7��^�V�<m4C�Ie��a���.d�q��Y*C䉏8F�%b����NuQ񅗹zy0C�����2	I$����2d7R���3?�s�^.(�R��w��V��mra
^M�<9`*�0HiBåT�E� ��O�]�<)mM�'2�iA�H�eD,�Q��]�<A�b��@������>OJ��t��T�<��Ùjd 
�d��B�(Ԙ珝T�<$��G&pA2���LH��`уE�<1�@���}�Q7|�)�F�	vx�̔'a½X����&U��(�-�1[v|
�"OKٲB&��тh�lV�$k�C�	�'[p���o��m�ve�΂Y�B�)� �� ��>Sx��e�N_x�("O$\�w \$2x\ջ��_��ʄ"O���#�&��\�v̜�U�>�җ"OT��EX�-��ۅ韤���PT�'�1O��s�NH�v�^Q���
B��:�"O
Dj�@�\�:6d��dO(��"O�YW�,���4��064�C"OF���.'m����CV�G��!@B"O��P j�1�.L �6���2�"O�)�$�&��]�f�e����"O�e`Z�k�~�`�n8l�P"O�Q��UCf���e��ai(`�"O �E��]���&db�5��"O0�Y5�ې|h:��!�9N�0XQ"O$Ę@����Qb�R�F����"O��j\�t�ʨ����0є��"O؁�D��+^S�@�v+�&�L�7"OP��.��Rk7�x�"OL��0D�rr�$Cp+\�h�"Ohؓ�
�Z�R�"װQ#l![$"Ox�P�%��%愡@�D>>t2q�v"O��`�b(y�� BVm���"Oj����!:��P��˴L�^�S"Ot-����2�����f/L����"Oh�[$�	m�%�)Zx$"W"O�2��	:6q04q��"Yӎ	+�"O$'#�­�$�=8�V�h�"O���P�	�[��l��^:�P�3�"O��dE
^�L"%D�G�<��"O"L�4-�j�*Y�$�a9�c"O&�2�ŵYfPpp%�D&K&Ӆ"O:L#"����*���S�!�6�	�"OZ�r�kZh�H�"���"On��(BP���*Q��Q@"ON�BebU�@�1qfƑ5��H�"O�I�d��Y�TI�%G�V*���"O��c���s����f�z��"OD�!#.Ж#�H�O^�ks��)�"O�}�E��=�(U���O:ٰ�"O��:w��(�z��V���
�
V�'R!�Ĝ-r��� w	��VD=!�M %!�
�k���ڷ	�0m�ΐqbmR!򄋽�V5J� u�ab�a
�
"!�$T�K���ұ+�+X�(�����!�DOk'��DK�7�$�б��Py"�Ĳ� �kVϔ0\����fӈ��x2@ۻ���W�= 
�'D�cJ��'qa~�_F��Q0�S�h2�QVDO=�y2��a�*��땨YɆ�U�	�y�������F2e��P�wb^�y�K�33��ir"]5j�@x	c���y2NӀ�r���I@
-D��Iu�%�y2'�"��`�,�)n�8�I��5�y��4)*�Y!M��<�����S;���"�O�趭�A7�Y��E�3���*U"O\��$��_!��vdݲ�(�ؒ"O����e�b�ˣ��2h}�q��"O��zF⟡3l� \�lq��kܡ�y"J�;ϰ}��V�HBa�F�T��yB�йQ��p�"�ogBI���8�y��Ll�`	�c#8� �^2�y"��E���
'��%`�"�yrIד+��i���i�^\�ĉ�"�y�nD�TΞ8+�M�26D�8t���y
� ��
�/�?O  #��NPJ�Y�"O��Y�)�����#�
��kg�T��O�Y����F�ʜ,h�p��o>��8�O�B���b ���aP�_� �u"Ob �a��ы6"��+���!d"O�;g�
	VI�#[�7��M�"O�a(wN�ep��'ㆋA�@�"O@�ZUG�OK�AA����af"Oʐ؂a+ Z4{0�(�h�c��Io�'��`�$���K�k�!i庵IY��!�$ؗ8`64�GdW�kT0�V�\j!�D�6zP�G"�rh�YȰ �i_����%,��9�׃�.SI�`�N>V���$�O����@�x�hyc��	,����&�!�Dك�� ��C�I�B�Y�ڱf�!�䚚(�\ZBY�����b횶K��O��=	��y���'�rp{��5t� �G���y��\*p��yv�ƍmKfɹ,��yҪ�2a�� ���Q��"դE-�y�a
�w��=���Jmp��q�� �?��',��*c�D�h6��Sa� -�Q�	�'E�\���<�4I��.�`�	�'��{RZ�[$⠪BZ�dg���'vɫG���,qcn�k�q�'��˲GD�k���%`C1�="�'�r���R�_;��6��'Xz��
�'خ���*��(=��mI�3^̜z	�'˼X�!k�AG<e(�0_��8K�'Æ� E��F�Rp�e��T�~���'S8�cC�1Tֈ��iİ��!�'�`�۶F^�3O�]�%I�&8������`T����j^Vs �3�y2�\D��BfEU���2L��y��	fs�8  � �^��� �'I�y�F9����1��k-$�p5����y"&	I���m#l}KV.��y�����t��D��%�R�#��x��zz$�����'~$	c���,Z�!�d�oJ�B"�΍Iؑ1�-|!�^r@�
^:F���r �X�e!�DO5'$Գ1��70����*Y�!�䊎y�@��Uk�3I�ŋ`�O* �!��
l�� ���0�,e "#N'I�!�D��M���`�i�;�H�Ѣ���!��=&
�0`�L8;ɤ�K��%�!�dj��e�D���ލ05o�/�!��)nj����K8p�l؁`N��G�!�dG�"�~|Z1.��c�VM	(F;�!���{ ����iVC�p% ևYR�!���7�D��lɸ51���F�g�!��^�@�Q-�)%��6Fy��O����F�#��9a4!�3p���R���%v!�\�N��l����6�@)r�BW)t_!�d^�$��7�c�.��p!�4v^!�D�C�L�jkB�{��|kEg�DP!�Q�/����劑9��H�o�%0�!�\�l%gfPA��-Ӣ� ��!�D�+�챣Vh�%��D��k�N�B�'��O?�g�{h"ar&�y���J��l�<)V�T; ڼ�w�_9X����hGk�<�ac2Nٮ0��#�2J�|!��,^�<YE��G/Ε��k�|���2��[�<	p�������6B���1c�l�<9q���_��a�E�1'�0P�bM�j�<� �%��S'>� (��ʂr�6h��_��G{��3Y��e�� 3|�1xq��6M!���ub�Ai�NN�Os��ФbO�P�!�dE�>�PU1��-B�Ƞ#'Ď�z��w��10�CP3 ����Fn�Y��4�h7m��yy~BG�8$���w���8F��5]φ�iV�Ƕk����D��YE�ģ?����PI�6Jm��E{�'��Ŗi�Bl�-��K��Ua�.�!�$ͅȓ��M�p�ӌ,
`9�R��x��=>���,E�=B��A�8�����23��&h#�Xۆ(�L_���m���׋�A�i���t�XЅ�=}�9�qFS���`�
�-�}��j��T�Hב�����f�%3��E��I^yr���q�0oGZ
�;e���7".D���R�ԣ�.=�7N	*���(-D��3��V-I�u�eS��4�W�7ړ�0<	�nK"^�ܨ��e�W�Ɣ���CN�<Ŋ�����Q ��-��q{@�K�<Y�O�8$��!&�3���R�_H�<�fG:e޵�ׂ_�^�>�:�˓^����}~2ŋ�fҠ���V�ƞ���☋�y�֙i���2�D�-_:�<YW�9�y��8|���(X'\~�\#2��y�������h���3��m�4�դ�yB�Ď��] 1�
J�m�ED��yBjH�\�4hX2J�Y4���cZ�yb
�@��M���>fX
c�#�6�yBL��(,����F��e�1����yr瞙Q��1���/�~��G"�y�B��k� �9�*U0~o��hR��y�'�]������ph�bG���y�ဟ"h����޲gf����3�y2ʃ�c�ވ��*��oKx\؆M��y��4l+�I�Y�n�з�Ƿ�yb���*�j+@��;X���@��y�(Y�gw�����*�p��@��y�����V�A1c?���I��y�߽�� g�^�Z�I��	��yrK\�YJ�!#b���SBL��i�+�yo�[�pP�ѽH����@��yR�L�jo&�A�1e��ۥ#C��ybX��N���յ+0JT��G���y�J��E �X$�#�f�z�@X��y�I2blP֮�&���	-�y�H��Q�a�c�P	�ԌQ]��y�E�::�T�W�SX��)ݜ�yb��8'� H�mT�I'�Q2Ŵ�yb؇m����b�'`�); ���y��!j�b�9�	գ�tșA���yr�_����Y��A z0��zf�]*�y�C��;L�����)q|� ���?�������8p �i� ��I�7��w�89�ȓp'�5`���J�b�a�jر ~��l����Ãʸ���w䛰$�D���Ib1�G�K�a��.y``�ȓ'�n ɓ��0�b��N�m�̇�fL���� 
	���q��#C�x�ȓbZAk�l��aMd�� hơ
F:�ȓ:s���V^��I���N�X�f���kx�dZ��֣R� h���jEZ���6�ԥ9E!$q' �2 �G8��@�$�#�,�h����a>RDU��S�? �(	d�^�"ʺE��m�&�hu"O�9vD5Y ��)�Q��	X�"O*}�D�.r��u��(S�NAI&"O����"�9.����*�&��!�%"O~!)���3�¹���۩v��b�"O�Y"�
[����%��(y����"O����)�C��i��GԪ:[�%�"OT�i&�ûm~YwG�n���H4"O�����м'�T�r��7i3HhH�"O -�h
�[,�����!�"O�2��J =�P��>8֡��2O>�A5gٓ�`�br(BLeB(��M< b��>8�~e�5a
33f�ȓ {aѱ@�v!����A�> ȮU�ȓ<?�����	o�搸�fӺ6{lY�ȓ����g�i��X�W�	�!��U��g�2�bB�5�F�8'\�7��`�ȓ�t1XQ#]��%!NX17����X���H�F�d#��1����r�ȓF�*9��m!!�ɜ+�Ɛ��`�P�)�2��1�cN�Q�\���\~�
-`�&�Ȃ�H�j�p��\
�y��M>	|�8%�ɑW�D-8����yҪ��z���SĂ�$���Ph���y�Ø�6㴥�$�A�"�T��'��y�ǂ%\^Z\�E��-Lu����-ӝ�y���Tڨ,�@���Zc�� �c4�y��?`a(E�7e�&C�rPQ�
����>I��?1�Eͫ3p�d�l�B�i���y2�-/��5�L6b�T�ER�yB҅I#lh!���?V��]�MP&�y�Q=vW��`�LЂM�>p҂��y"�GN���q���J�.IZ5`ږ�y����8�z��E;��hs���y�!�NK^��%iݐ2=0d�������>��O\���"^��a�jN�h��0�"O&l�Š�Q�D=hK��m)����"OD��feK�O��T#Ǫ�*?��2�"O� �����r��ܱ]��5"O��C�+��+_X�A�ŋ�@`���C"O�T��EC �T�򆥛AV�)��"O�uXciL�|�EZ�JS9�Y$"ON��ת�e�x���W;!��%"O
){�@�)(�n�ʔဣr���s"O����ʼ"!tx`�`�!^&���"Oh�J����"�x�cDoK>7%���"O� �6
ېY��!x%��#$ր�"Ory`�8x`d!�P/1�1�"Op�Sj]�zJtK �C3? ܀��"O����@�";��{ G�
�~�b�"Op�`��U'I�ń	%@fx��"O�����K]3:P�2�X�UU؍��"O�UҀ$��|T a1`"��Z*8�s"Of���L��O���qaCR��ؐq�"OH}(U�3{`P*V~\T��"O���c֗�h������K"O�TR���}�E#�oХ;�)�"O�-�b�вl�<����5֨��"O�	+���g��p�Ba�3"OP*�!�?<�f�1"h�(�h�H`"O,�"����e��,��8�(2�"OX;vcУv�JU�ˀt�>�i�"OT���ҩ[����w��'a����"OM�JVdx*��&��� ��\Ё"O� ��� �
\����(q]��"O\\�G$$r�9��ee~! 6"O�X�0JO�v�*�x �ǆ_W�f"OLl�C�<n�����Β#���b�"O��� �`���(���=�6}�"O�t��	��6-�"�!q�PMJ"O�83�#	�
�I��`:v( ��3"ObM3����mؖ��%���v+��!"O,��f��UY��Xt�P�Vn�0I�"O�S�-���|4hŮ=GC°�T"O6��Si�X�6M
��ȋN4�5�v"O�m12d���}�R'�Nd�g"O����n[7-�:,�,(M8�+P"OXTɐ�Xf�ib&`ͣ1�>�[�"O��R��J�@8��U�t��"OF�ɀbԐ �	�:.��A"O��Bȓ0�pT�&@�T�z�"O���	To,���n��`�y��"O4�(fhݕ_W�T�`�"6�pQ"O��t�q�T0�Ʀ��[R"O⌢��҅
��D��*���f��"O�D:��L	#L�!#�L׿r�}��"O���S��#'+��AdN�'�R�"O\� &k츀'N�M���Ȇ"O��3vAA �����n
4���"Ol5Y� �#z�����΄g��"O"���+�
d�L]�4IY�o�@ð"OȘP�
Ȣj�vd��H�/��0�"O��C"��5B� �n�p�"O$�����7C�mxC�"Om)c@�YT�b� 0>��3"O`l��B!$w���"ʑ��"O@�+�o�$%@<��R�4�u�"Od\�t	�b@td�B#Q�M���"OD��D��IN��hV�M�u�g�<�0������g�U"E���v.�F�<��fD3 B�Jr��#�N���W�<�����ja9���P1�`��T�<Y�#�Pf���G�o��1T@T�<Y�!Hj�D��,�
�V����Cz�<�s�D.%nMx�%Mwnܑ���n�<����(���.´0����`�j�<!E/U���9���4X�����!�h�<ٓ�")����gN/j�P�R|�<����:�0C�)/�J04Ex�<�ʾA�@J�喴9@��(�w�<Q��	H��U	c�X4�:0(�ew�<i�E�aD�=灏�p�&p��.�q�<y��<n���w##���@ �R�<�W�&�=2e�	��@�4�b�<y�e�)o�tX���!�P�|>B%�ȓ1���'Ȭ�R�����a�BɅȓ+^l���X�~ςp`��¤x�hp�ȓA�e�W��JrN}	�B� `c$m��U��0r����nD�ֆ�4O_ZX�ȓ�$�Qf �.BVDa�J�3qX}��Y2��j�;?B~Ey��I
�����鳴&͍D��T�Շ{Ip�� �Q@6�(&q�%:zu�ȓw6�<��J�f9vX��̒�&mDu�ȓrø�5,׆p�l�KǬH��a��$"�A�.�	��t��� _-�t��O����dS�3ߺ�ZV�:h\V��ȓ!��t`q]�"�*I�%�"t�n���S�? HHp-]#H�qqEO�k& qG"Odi��#�G`D�)IX�V�0��"Ob�G��	��	*�ϑ'El��&"Oʜsv,�p
-�4J�q7T}�$"O0�ن��\F�	�h˘d��a*Ox�VE�7���Z���E;�'.��PT(�9L�C�VG0% �'�" aӍ��"0��񂔭K�(���'�����R��0= `.F4��	�'������'�(�{�閸-yz�a�'S�(��	�Z��(��S$-$$��'��A��lG�S�T�eM� 1p���'Њ4�"�ΔP.z�A�#�R���'p���B���JW�s�-)�'���G��R��q�&m^Kmd�i�'�flZ�cΧ�*Q�e���@$b$��'�L��3�̻	zX��$Ӗ
���'����Қ\喕�X�q���	�'z�p�0�R�u�\�3��=���	�'H�l�c��(���7B6=x,8	�'��� bM5]�KN_�0o8�[�'���C�5!��v54� ���'&aL�6'�J��r�]44_H���'@�Ļ`�U"%��i��-+����'ZzlqJ_�8#	yan�<!|2���'�����j�~#8豢Z-�ІȓmFF!ё�(n�qh&C�
Yi��B�q	�ܩld�t��� !�Ԇ���5F�|�[�^������w̹���W�<$$+��1M�P5�ȓ0:����[�I��:��z$����c�`��Q}��aJ�Lڋ{o:���(d���b��|��U�s��"U����ȓk�\m;F'�D�L�
�&~��ȓH��	!K��9�W�F����ȓ��}H��׭A�fՉ�։F����
� p��̘'�ك$�����E�lCqfӲ�T��T��j��ȓ,#�y�@�N�%|�P�}|�t��xH�Xs�L�6�0��'
�H \H�ȓ-���x��ءq��h�(Y>V@���t���A��]�x��e\C|��ȓ�Ȱ�Ꝓ!�2��ˌ�z5����V���Y�"�3�IO3h�H��ȓ*���@��2�D�	#��'����ȓ'Adx�b���u����f���Ɩ��ȓg'��[%��j��D;�G%=�Ji��a� A�&]%� �2a'�!h�%��2<��A��Lx&lꧠS�v�ȓ-ϐ��#d�9:�)J����,8�ȓOv��s� <)��Cg�΂IB���U�\qeK~pn4�UhG�[|̹�ȓ%�*�3��"���J�Xe��ȓ!��4���%>�B�js��F� X�ȓ+<��8P�2TŚe��&M���ȓ0�;c��e�>��4 �!4	L|�ȓw��zs˓G��hB#�f�����6�P0dλ|�:�G�Jq:��/��ۆ��b]����I�LM朄ȓ@����!`�TPʸH��V������$P��A�#�"܄��+֍neҵ��Y���¦�T[�h�ҋԐ)�؇ȓG?�sH����ጐg�*��ȓ8U�TSm��0���Se瞋|@��S�? ���F�/Pޒ��D�Fe�ȑ�v"O���#��(_��y@P���T�!�"O�`���P�
T�:�HК|5��"OΰY��S#J������"�hم"O�aq�D��$�:��3f�~�]��"O�(����u[å[ lJ09v"Of�������d0Ս[�l��xC�"O*�i�iS�1�9�n�\!���"OLQ1�ӄv���0�@�J����u"O"ث6������b�'�ҍ��"O�s� �U���K�)<=����"O�lʔG@�CQ��҉�M'y�"O�8H��"�Q(	�ฒ�"Ol41Rj̱�̴k�[�!��s3"O
�{v��x���,�)�QE"O�����4X��<���Q8O��h[u"O��Z�� �Ca���T�=IH "O��9$lV�!�z%EӬL8��[7"O~�J�35(�&�Q2?#@m��"O��J��X�Dg��"��ܳ)L��F�'M��N�(Ͳ�!@p��w�O� 
C�I�-��X"��X�}�r����˖{�C�	0�̘���I1+���{�	��T\�C䉵T#̀�2���b�8��&����#=9��T?���W5s\�D��B9���ċ:D��b'�Y,1���DE+|�
g	:D��P(v�X�A4+�E��*�m6D�������B7�H�q/�	5�q�	�>�*Ov��I��'���'4�豯��5�rD��<W|VC�I(�L��D������
C*ZB�I�ٚ7a 21 ��3%ܶW�4�DG{J?-���U,
M*`�T	C�zм��e�-�:�OH�y�D�l:ر�Ag�F��\�w"O�i�A	�+v*1���
�3P� �U�'�1O��A�I�<.���%��J�%�"O���I����⁩(3:D��"O~����:tY����144�!"O��0gܛE~�Q��Q�w��h	��|�)�>#0�;V�3#�yFBC�a5 B�	8v��YP-�d��{����}���IW���	SŐ31����oQ!�<�#�/D�H�B�HP�½�'oEXf��ĉ.D��Z�T��x�+1��xX���c8D��I�"��
���aǢ�i�� 3�H���D{��IՈ];�x�,��!�"�*�!򄑦`/�����$I1�ՍN��OZ����#b�A�J�5s��[���/I�H�O,�S��y򫚀ڀR��/0��)��<�y"b_�.<���/}1@��Q-���'|ў�%��%�ŻlZ��XRMJ ��}�
&D�t�U�6Ԓ���ʆ�^1��+>D���h�5�Z�2c'E�~�F�ye
"�d&�S�'X ���̂S�p�P�(����R�M��A�A@ يd���d�Gyb�'�,q�ÎR�,���A���
0f[x�<�D �y�L�ā_�0�
��H���	\~�BV�<Z�L����(+0��C,���p=��]�|��'^\D�3%�4Tv�т����T`Pz�'�X�SE��8DtTK�$3n��{��)�i�$6D��OBc �Tb�"\����>�N��!���6�R�rA#�f�<i�#�c��	��A�)	�i���K<��XP8�G�;}"�!s�-7��uD~�7O#|�`�����Yd_�O�nU��E�<� �=�J�T�vL͛�+��`"O�ET���#���l�Z�,Ux""O����!ϒh���������C"O��!��i=Hd�q	��cbE�"O47ȓ6��HU�D2�nͳF(D���N60f�H���U�<hne�q�)D�|����TEh�0�/?���#LOޑ�>�CG�PU��h��N�hQYA���1�'�O?7��+^��Pa�d�1�#�	s�1O��Dz���P���bt"ôG���b���yb-�	}:B�S���)�mq�mA��(O����:ev����:t\�`��b�!�D�7,�ա"�Ü&Ju��K|����O@b� E{ ?$�ؑ���ϑ0v�x�#[�K$!�$)g���b:l��ہ$?Y!!�$J�zE�rl� `e����\�wi!��Z���W�� �A�ppՅ�˸H"2�ƓTX1�O-E����lU�A�Uđ��,Ń-I%8{X`��26,*�N�W����� )�~x��k%��0+�H#Dq�_{[Z1��4���g��$�¬Η'M��l�4�hR�J
IfN�"A�w&D�E|���\�PqCnD�ɦ�⊠�zB�	�M��QH�˵3 �	�lH�=)���d+�u������"9{��"u�!�ȓL���R'�3D�*	�w�_'�l��G���'��c1�ӵ]�H���K�:@��7*�00d��vE��R�E����u�P%�`ġ7]�Y��ϟS��B�I9H&A�
�5DP(����3Y�FB��10$AJ�$]5��Eq��N0-1�C�IxҊIs����n���˓�˱s|�B�I<jO������&�j9���.8�ڢ<1��T>��e��</�d��%&�P��D�*�O���F�����-�"��K��z݈6�6�4k?2_@�0��Z&2W���7*(D��l���@�(�b$��)#�%D��Rw풓T��eO�q�$"D�� D)��-��ax�H�>|����>����61��l�GQ"B����K[��C�Ɇ#����-N�n��}��	F�C�ɞ&�8tSĊ����I�@�H�<��C�IP����CbEe�f�
Vj�C�	=����C�Ͻ{0������
%�h�'�a}�dE�!�V��t� "��rm�<�x��'Ij���8?Ê���		؀`ߓ��'p�H�;39�t�g���=��'�"Ի��Ǿuؖ9���+�%��c�'ў�'l�@��CS��4��d#�*�'�ў"|���Zq�<�bRdʘj���e�AH�<��
#,�aZØ�>f��`��H�<�a�I� �8�k�*x�VX��FQB��0�OZl2��Ž:�h���O߯|����'��I����w�L��iRA��6_X�1�c7LO�7m~���'\X�i�J[ ��p��_оxx�'Ehp�3.D
ysl:�T>l��c�'V����a?'��Q�'$� �+K��E{����
1K�\�h�.d�@Mq�
�y"�H�U�~����"`��0I\��yR/G��]�E��X���"\��~2�'���Q R#M� z�kA}#ZhJ<9�yb�ĥ?1���Y2kh4�"/�y��%���(�OR��I����s�(��Nu&M��A[�XB�)� *�觥GCn��1�����)��'PўP�d��l��0��^a�dae�(D�t�H[�9�Ju�6o���V��E(|OFb� #q ��Gtdy8���j��A�3D�Ԣ$G�"szh�V�c��`���o�\�=Y���]?�D�d}���b�s�_Y'�B"O0�;��Y,+F��V  �����	MX�āfP>*NHA��΃x��`0�^��hO�O5�F��� &��)w�&����L�d���w>D�1 �T)PCn�RLx�����)D� ��]!cM��	S㞱T>����,��,�O�Y�T�ɑ$���RҭA�C�F9���i�@�=E�T�ձPV�8�Hƫy#n��F$B?!��,�� �F��h����ùN��9�OL1yt��z>�9Z'-�;� u�A\��F{���\
lJ5No�px�&hK�!�Dơ������%�\�a�X��!�ֵSd��H4�X>J�z-A�\!m��{R�'��	�9�����/v �Y����k4B䉱~�)@�>͂%:�@b��C�	< ��l� h�<y܀�j`�N�B�C�	Y�T�JT���)*ɚ�iQ [8B�
�r��#��h�F@K��O~� B�IQ�`*�ǂ�6��3֌�4F��C�	�X <��)<c�l�E��s�C䉈��� e!Dn��z0��C�CۊMk��W�oIVp��-�"J~C�]��R&��*��X��DY&O�dC��#��䛰m�3\��U��'6�B䉮S�>�r�?9�X��a��
$�B�2��ac��:�u�gO>|J�B�I�B�V@���!P޼����2o��B�	�)�����)�5i���둤xT"B�1{ۖ9#�8]��b`���9��C�	� ��(2č��;�a���C�Qg&J�#Ԛ|��E�i��Y&�C�	���Q�&\�1@�AN}�tB��/3 �D� �^��Ma���1�*B䉗p� �{1���0܆)�PXc�C�I�9���r���<7��M�G�+�C�	[����	�+t]�E�=6�C�	�w��d�/����_"f�C�I V�Z呒��7H��ݢBXC�	� �>��Vq�z0��!�:(C䉜f����bhѱZw�m	`LB�	�9r��fDyWti��I;}YfC�I�D��	��+�j59��IO_VC��Y�J]I��:�HG�"qG�B䉍	�mc��ڸ<��t�
_*5�.B�	6e�B��F�1(�����-x3�B����*P��d�
���}f�C�lt�e����
,d��s�D!fx�C��7E�p��tl�8#k��+c�z3�C�	+`@|�z�m��/FؑRN�e>rC�ɿm�$��E��\������
n��$H;'��0�U�E"a>z��%��0c!���Oބj�a��4�� zj޴s!򤟰Pfd�8Q��.9~V����D�!�B�gȰ�1���?Whp�ؕ��!��A��|�s5ːE^�-2���G!�d�@���B�O�t�7��9�!���b��0e:
�xA�.�!��Үb�<��5�\]�&�!���-L��5ρ0C�L%����(~!�� F%L��8(pT�5G�+��m��"O���7��s�����M�R9�"O����[�r��4��-؊F|�Y�"O�I�C˹1�0!�,G�#�`��"OДv	M�����1O*�Y��"O�\򠭟6!�b��ք�4�%"Onl����=&m��Y�B^nʬ�a"O�%��O�o&V@Xk�D逩�#"O��k�gʩ0`��z�_�ZƜ�I�"O~��QM	.2�X�
ĝL�`h�s"Ox� �[m���W�=Q��QZ�"Oح�͒&z:�!W�J�HHX� "O�l�Ak�~�Ȉkϊ8.���y�"O�����1`02�R���o���Q"OΕ0�O
U�&�A�NT/0���"OT�)��/%�H�a�O�
�:`�!"O��ʅnU/M��sp$Yp��
�"O"E�&��f����
$<�~��R"O�A�v��v�(镢�!��$R"O�99t��,?' �����%H0v�"O:5[� D.=D0HPÐ16�� �$"OX8�S!Q�_M9�F"�D�x0�"O�Š&�^�(�^����>��`�"O���R��0�tD� چ9���*2"Op�{LR�QV8���ŉ�^v��J�"O ��F��<�uaƊ�_w��*�"Od$��`ȅ:e�]��Ծ-WL�qG"OJ!K�l��X|����Z�0�"O4�*����Hl�1�!�7��\�"O��UK�,|H��`S)[y����"O�dKu�X9�ʥ0�iɽ\m�!�u"Oؕ�BV���ə���X&h��"O���c&�H��q�B8sj�P#"OX0)P,�g�e/eUz��צ	��y�
sLz���[�g��{rl�6�y�C[$vQ��"7, `��H�Tk�&�y����I��f�	S��ݒ����yb���	���嫔�Lt*��"�y"&P� ��*[P|B٘�)ٻ�y"��-�6z�a�,ST�$a��yR��|蘴�tOK7V��`�ҬT��y���b�^I95�\ _�\�B�P�y����)(d�K5��%���y"�G�L�lUj��:��l�CV��y�/E"�`�[���5$���@uL�!�x�"�vLX�D�k`�y0Q	��V�Qr�*G�4N ��'p����ĤORD���J�CmtUъ�$�6%"q�JT�z���?uY�BӪ%��@h�ȜN����B(D����-�<�&��D*�jŦ����?�x0r��W")5�����3��°��I�0�òC�ZVZB��,@�&��o�*gl]2��X/�t�"T���r�b�%1���R�'R�ҧ��>��Q�o��1Ś��Ŝ���>�5�\�y M��; 
����L*{h��t*0�\��c �X[Ĩ���&lO��r0G��M��ȴ�I�^���:�鉡]Jf)���Z�N�Fx��ݮFYXҥDփ9q�)�7E�P#\̚�N�TA�|��'ph�#��2m�����Iz�]�G�>��p �暾B�`����kvx�ʍ��Ͽ'�P�*Kl�s6%�����RD�<�v�N�"�p{'FҕFD�����n���ROɶwe*A���X5<<��yO��3s)*�I)�pij�O�0:�)jVH˸k����dѳCY�I�6΄�|����R'�@��L��F&Gh���m�.)|0�H��O�ubhb�� <O@ؘ��� 8�ѢƆIX�5���ɸG8���Q3Ey���͌�!��S�CY	��C'AQ�	��#�h��<�%J�ph<�2���*e;�cB+
i(=A��>(q�a�O��g72�� ��A`���Bg��,m3N~�;5C�l4Cߴ��Q�7��2xs����S�? �U�U��g���!V�C$(	<���͝^�<�h6�ޝc�,l�"@B,-���Be���֊"�d!H� y���n#,8��M�.{a|B�.n�x�#�ѦW�H�x��φ-�|Ԓ��3X�@D0�)	A&�@�bȆ,Z�!�5�'��uY"̚���8�U)QV䳊�� �~ST5�2d�lx�`S����Eճ,H��
F�DH�I�aE�@�T�r�$:4�� ��)�RQ�&o��C�>9�Ӯ�T�r-T'm��Jd.� Z�$��p�!+�TY&?�]sa��	�AZ���I�!���>bpB�I#9�~%IEn�DA�VD���: ���Q�Ba�qDѶhN� nb>-QΔ7Ce'�!!$��7Z4�)�	9c~�H�D%�OL�9���;&"��HR��+7�)r�Հ\Zp������3���%�N-���
x����$��Vz��(գ�#��鐯B�u��\�N?������FKB5Jsa�$�P�S�*"'` i�	Ҫ]^0��ǉF��(�ƓT� ���̈�
=�x�%@�=R�A�l��hςd�@�
�\�考�Z�P���֬'��缓3�\�*m #�X�J.ޙ8���L�<�.љ;���k���4yX2�14� ��3_�F�vDi�k� �*0�';���C����)\H��A鎓D��ň.��o�Ȇ�	,q�zl���*�PY��E�
'�e�!�Y�&䨁��'T�����bx�u+Nx�`�D*� d���P�B�>�N���#>�|=�q���g���rB�:�@����7L��X�`��5gHP��;U��ѳU�?D���� �h�P`em��p^Ru:�FO,?��殅7RѨ51�ŕ&m��ң�i�R�>�n,7�dѧ�$�H$�G�3{!��[�(�:��KW�.�ra螭Ȳ=�r<�tQ	 LB(��ł�\?���
@�++�l�.t�J�
c���F�p��ɜ D�`��B��5�4�󊟚��\����4��i�aΒ9��9�(K%+ a{r��H�p�`��$|p|�ؗ��;��Ol�bc�l恻ԯ�.��|b��柖��x��\��,�y��6"O�i���2[~�H�,p��K��~����e�R<	p�2ե�3��"~�§K�&�q�ě�6X``RG�H�<I��[�P�(IR�I��,�H�p��F!E�����O��Rʔ�Fn&>c��ӥQ0<	�@`ᅍ�~ $.��۵N�>g4�Z�%G75(�(�7lQ
+Q��cf��_pp��I�3���C2��,f��� GO�KbC�	�b{z��'�&�� A-A6^B��-1BX�PF���\�SF��8C�"�.+C���nF4����"{��C䉗D9$]�`S�H� t��;��C�	�pU�p�o�pg~I��Y &��C�	# �ޜ���yd����X�`B�I��ܨwǏ#z���c,߉+XB�	�a���T!Q�	9�)b$��A0B�I-D�R`�S#G�Y8F�*�(
hB�I�9�<���Ci�B���5J�B�	(f�@�R��Jv����A�?��B���F!��LI4��5��3h�DB�	��ڼH�F�K�E��N�pEB�ɘHr4���`K�F��p�`��Q�C�I;e}nت��I����O�	#�C�I-��yaD�޹=m�AxG��~�VB�>C�F`GmT0�P3-T���B�	8/.�Y�i�bQ����(X#S�fB�ɹh�����\'`�� HvC�	H]$Da�.Ĉ � ��@��B�C䉷2�5�v#�	�,uK�J%%��B�	�ed �+g �A'�ђ�"O��@���Kܺ��� $����"O~����-��]����3#�N�r�"O�5����~��0��fa�25lō�y���<ԩXA��!!H�$�ԧ&�yr <(�4}q�����px�D��y�� ��0ٛ�-��&aá�<�y�`����U,�'�IhSFމ�yBa�>K
�뒣[Jx��CG���yr��Y���/B;OؒT2#D�y����3��Se��Odn�BC����y
� 2r�۬T9�t�B�,aX6)Q "O�;GbI�R&�Hǁ[�"&��1�"O2����=L���fK<c�<C�"OP�b`G!c��t�f�Ѣ4q"�Ra"Ov�ِ@Y�>��pXW�
#e�,�C"OD���B�G� q�f)�"zA����"OV��Qv��!��G�D9pT
�"O������+3�Tk@&ֈB!tM�u"O�LQ.V�.�q3��M�2��T˷"O-��^.�R`S��(~��1�"O��0)P&uה�83�F�v���"O�E�4ʏ��1jbi�=�� AD"O��B`o�
Eo���gQv����A"O���q(B����I�&��s~Kb"O�D��+�0�(��Ѯu��1�r"O�ո7!�4c˲�`c*M#A�:�k�"O�ԃP#��H�I�`W�ѐA("O8Q%+�7����B�F�A�:�"�"OV��мc䢨S�m��+,�E�"O�@�B�(*&��s�-S�xixDJ�"O�7*�r���#nR0WE"!Y�"O��җ�������L�c��%"On�HuY�_�0��t�؍D����0"O��cp����i��5z.��"OF%�s/��y��Y�@e�8Yv"O���2�c!��!�0m�`��^�!�]-LA�C��5a�AJ�D��&5!���l~}ʶ�zW�쑡��>!��pJ`pFKȩ?5�xJ�(S�D!�N�%)V�uc�w70E�5�^3:!��L7`� ��e�8G9���g�3@!���'�FժULL�L CsƊ6b�!�12q��y͇�o>DZA�ǧOs!��(%#�mc�l�����Py!����~�T�"�oQ�{24Hd(	�I�!�7����lQp�����g7Q�!��"d�4��q� 麗&Ŋ:�!��"$�~y�/�1s��iA�Y#u�!�� \Q.dAS�2	��z5�*vp!�D��e!��A� �0U�(�2�l��n�!�DݔKJ��I�DF
&�ꜚ�kK/u�!�$1��e!����_Fl��� L�u�!�ߜQ����oLX&���M݀�!����;x8r&�_ ��%�@�+�!��ܖb�~���_
-{,�i��A)W�!�6j�~�[�
��Vi�i��0R�!��D�phJ�!��iQ��i���!���4��$4����u[�hS8b�!��]l��$	�C���Fq!LU�0�!�צ��U�[@�l�yԅU\ɊB�:mO%u#-$H���j�C�I�w��tf�W�.I���iXxC�I�(3��K ��v��ca�=�B�#���G	�!aH��(ʡGt*B�I�a
��J�ː>Q�R��֊��f��C�%K��}j#,b
�J�L^X�C�I-f�쁡mչ���;5L�#S�C�%:n���`��q�P���.�2�C��?wD0U1$�$=�t�I�Ǉ���C�ɒ`�N��G.K�Dd��X?AĺC��'z�<�(p�ɭc|3#
Y+Nl�C��.�	3&O[�~��%�iUx�
B�I�5�Й�3AK�r�J���4w�<C�	��:�:2(�a��(��.y-C�)� p�*��F%!�A���۱[���:"Oڠ�UG:`J=)�A^m/�02�"O*
E� ?����6yr�xb "O,Q��#�(�t��|fFq�"O��:�O9g�܀���Kw  ""O̤:�H��)��ݒ��@1 ���"Or5P'�+2H��â��I��
2"O�	���R`r�f ��Hy�
�"O�4!���_���*sN��ZW&��"Ox=Y�h
3{d����T]���"O�u����lG���R��m�@\�"O���իH�V)T�@��8>f�@�"O*a�#X�4�ʐ�	��|@��"O^���#�5�x��R�'��*�"O0�Z�X�64D;�ǖ�<��$
S"O�ē��9�H�����\����"O�Ջ�Ƣ�`���͂M�\�u"O�@�Eb�,�@�`vk�(L�Z%j "O�LbR�:Ո|C�)��v�a"O�����3��9�2�S(~.���"O�,��!H�I��13��Lr�!�"O�Q3�҄`W����K53h�)�"O�][�CL�����ܼ1���""O�����bgN�K!��4�d��"Od�K���:f�bYxC垚<��P�"O��`��A<>�j����ǩM��%J""O(���B�keʱ��1E�x:`"O*�����Z}t�'��6�$	T"O0q���^����G�5&W����"O�a0��Cu0.U���	�L_���"O`�8T Ԣ`��Ƅ����'"O��X�	�;���[4W��:�"O�����E�w;�쁢��F���"O���ڒ; �$�ތ.��l�"O�Y����:eXb�κN���q"O��Y*�8�ly:FF�)ݜ !�"O|�F-��J92Pez��N���y�Y<VV�@�&��A����y"==���ˣe�'ڦ�H�F�7�y��94G��K�QD�5BG���y�� ��g!�6G�>�����yBG��$�u���O��F�
5�y��#��h���G���t@
$�y�-�&nl܈`ȃ>F���To���yBg+p��e�R$^'���:2����'.�@����N��U�U3}l(P�'�T���ǁ1N*�����pU>��
�'��K�역%2զ�~N>��	�'�,L��J�R�),.q<���'�P!VH�!\��$O�\�*9�'-�*�ȃ*�I�%D����'����Y耊'�X)aX�Y��h�y"�[5Bt��IS�1^��x�@�yB��C��PvI�I4��Q����y�Z�'�-�B��^���3����y2�"S: � R<IzP(:�y2�Y�O�VHP�F��I��`:�AB�y�ʈ�+p����E�2�`]��yB��t7��q�N��b�.H��o¥�y�*�?\���� �J�VY�COC��y"�����A;���K�$#�ޅ�y��ѺC_�Y�P�_�1P��gD;�y�-�&-�R�k�kɌ��x��P$�y2c� L�3e'}8�@ voE�y
� �q��!4""e�%M�4�.��"OM9V�֥T���S
��p)P"O���)�1�*�8�B�s�"O$+�;�,�5�B9^m
���"O�;V��#$z��GZq^��"O��U�Ӏs	H�2E��L��h"O�<� ��)Al�P$ؼ6���1"OBMz�,�A.X�3'���h*�U"Oy�0�J�I�]�w�"��ͳT"OX*�O�1s|�a�1���RӚy�d"OP`�pE��L�08���T�R�uI""O�$�i���3�LD�qr�"O��S��I7'PP��=�l�Sw"OJ�B��~O
)��b�=����e"OZPهF%L���f�]&��@@�"OD`��+ѢS{ �X�σWA�\�"O���v*�]��g�*,T"O�x�.72 ��/U�ʌab"O���'�7�4E��S;P$YJ�"O� Z��9�8P�����$W���"O*x���w�Y��N��	��H'"O
����_��ٻ�O_�q��Q�"O��BTCS7O!c �?n�z���"O�H;�K��`�b��$�^�w��T�"O���W�^$I���	�S�j�1q"O"u@�ݥ+vҬ�R��S��Q
�"O4ݢ�`�����E��2  d"O����)A�r��ę�ۣ"�^��"O���XU��L"�,���6�Qt�<1�J��>U��3��_��B��i�<1��A
�������5�Gbd�<1Q�M�I��1�g\z�
'LXb�<�[$,[�y�Ƒq��Y�ve5T�8�P&B`L�sV�Ӗx��+e:D��a5-uN�2��_�;���1,&D�l��M,(1Sd����Y��$D�d��I�*����l�"Ppp �b,.D��RcUCa� ��mZ"}�HH��G*D����B�8�`�r���e�L*F�*D�4[��A�)�mP�tV<�K`
&D����(=�� �p��'K���	��'D���&֨KB.�#�	ͣ*�r����>D�̰��M�ESn�U�M�X�6�s`�(D�4+���]+�]�I�',�8#�%D���7�ދ��ɰR��B]��� D�dPA�R$�������	2���n5D��aKϞ9i	 7���"��P9��3D���->t���P�fľA
h\�RL,D����,,��٪�̼Sc���e-(D��+%D�9�����`�8`�� D&D��h!��D���sSbKN�ڑ �$D�\i�`��Y}"��c�6ܹ*%�%D�d
�i�3ei�	BB�h���0Gg<D��s��0oy���(]%s1��Y�&:D�DP��_J��Yxs
M'C�D�f@6D�L�sn�NS�a�Mޞ8,2D���.�=S�^� ���\���g*O �/K��H���-��RQ"O�Hj��N�{�"-b�\#nfq��"O�� ��Y>y"�@�`\�U"O�My���m:��#,Oz���"OJ�R&�;'�����*�xAB�"OVh
a-� � �;�C�P��l0�"Oi"�,Э>ߺT��X8|NH�A"O� vd�D"S�U��K��-�d�D"O`x��oּ]1 �ꄏ2�0@�b"O~ŉ��T3�J����ٜM��R�"Oh" ��:kB�	{�H��|{NH*�"O�D� E��j�r��qR���"O�,�1,�|6TYl\�f���p��&D��y��Y�VaXt,��9.��"&D�d8�O�MJH ���*��U`Dg&D�,;�i��hLT�1t	T$e��K6D�,��/�zð�j�$0��rb D�4��b�(;.���䏵,���o>D�����8&�����M4
0rgK<D��Rf꜖��bW
(���o�7�!�Cqu�͓�ԊC�.�iǅ��a!�d��!�&����!��U<!��>P��"�'�c�,I`�A��M<!�dh�d�PkU$�q�,��{׺�R	�'�2�8q�/;��#Q�ʳG�4�k
�'�Z�ɱ�G4L~.q(A�DE\��'&QA�;1$ļ����;5�tQ�'cҥC�	�CƁs�,̟)_��	�'���@����4Y��k��32.�A	�';^�[�a.(�D�á	
�{<� z	�'\��BC�B�7tJ�3$���b�$��'���G�9j0r$�@ƞ�XA@��'�(,ȧ"��@����?X���	�'~\0'��Hn���,N8H\��'k\Ő�*P6J��E��:���'zN(�5�=LX|j���*݈�'I�h�ҏC=D>�S� �_z�,	�'FI�k��<��L�W�T��M��'3�|�1m�9(�Jl[�e�N3DU��' r���G�)p��#�R:˴+�'̴I�S��9
 �|9B��G~���'�	���7	���A�I*:��Yi�' ���q�����[2�\�!�'��\H���&R��qx��S Q���
�'j2Ef6e��1w��J�Ě	�'��D��-͈�:tiF
Z=�REa
�'O�t� ꏲLd��̝7g�!Y	�'��e:��Fy���R����_*�I#�'�������
J�Z���㚌SM<�;�'����#uq�W��S���'����V�>|Ґ5I�d�[�$�K�'�����j�\$�=)F�^T�I��'�6`�S�y����W>��X�'�f��F¬tW���/N�X�11�'Z���
�QZR�a�N�5H�pc
�'�8 e��;H(���DL�?��DH�'6<9k ����l�F7���'�<�"Bc��?;нqDC�6j�)i�'��12�$�� �ެ8aE�f���	�'7�1�6��.&�o�6�@�x"OH�����vG2mQ�.�2N����"O�e��e�>�E��|���&"Oz؁��p4�1��y���3"Of�PP�P;,���ڀn� .tr�a"O0���g�k(��!���q� ��"O�`2�ဓ~�$��D�EMz9��"O8�S3���4� �7&["84"O�<���A4�\��K�#%�y4"OD 	�dI�zuH���Jۈ	�@esP"O��!���mYPGɕ�"��"O���A�p������ v���"O� ��R��zyLm2��E�*�ũO�)�I���?��tl3��M��p��Ǘ�@�)6���6���T�[�gy~x�'���*çc�rl���x����O��@��|3�����G�) ���O,���Ӧ��[<F������DX֢l?�!�Ϙv��tH��r>U��,A+	$\A���Jy�@:eix����`��T(���GO$S����IÝ��b�\1G7\A��%�2$�6��A`I!-g�{d�U�\^��O��e�&W�`���#��M�]�"��AoocrV��?q	_O>��Q�֊*_z�2K؈gD�p�(EDh�Ί�)J>mX�NH -PTMඊ��lvJP�AƘU��DB7Ula�C���2��s�q�������I�V��Pk"D�5a;񄖦F� %J�6���5��o��`���ɩ4~���_� ä�M�@IL��S�>E�$�ИB��ɡ��1-R%��G�;�?q1����J>E���K��(Y9�X<�!��$C�r� �p?�s'�:u���
�̔�����W��Q�<Aâ�>PNN�2�I�o{���EJ�<ɢ�U�f�(�S�K
W����c�k�<y`��'O|��d�
^�l����f�<����|�ehP��`[ڝz�cm�<	7@.�6%�6�|�&�XR�N�<����%e�pP��5Y�yX�F�< ����E�1/-M���B�<-]��e(�C�1f�!�&��q��C�"pԛ ߠ6_~��uႠd��_ �.�	ң��Kp���J�!�	7|=\��E�FF�m�� !�$F!|����&fP��쐬<,!��ùS��Z$d�[T|���s!��9�Ll)RjJ"ibF,� K�7XG!�� F����_�A^��q��8=!�ą"����R�{E��e��G~!��W
(�P|�+1D�dj�M�|{!�dNEZ���<:>M�kP�!�0g�*�;�GV�5�HI%Eի\!��\F�6l;�n��^�����b�?w�!�$1�R�5I2Mx/ۣ(�!�C�<X����AW:�9�k�!���@�T<�3,\����D
^,!� ,/H�b����eQ�!'[$!�Č�n� �����J8��:�!�_�8�N=`&��j��٠��JA!�D4L�� �ʪ9��D0T���!9!�d�74Բ���͕�E�.A�rL�'{"!�dH6� ���]�m�$��Ë�#-!�D�/����ʓ*����i�}C!�d����VCI���	G��2/V!���L�bA*�*Q,_��mC@'�{K!�$>s����T��E�$-E!�S�6��T�GGK�|���U
Q$a�!�D�}ylA �k��^_Ĝ#�HG�]�!�$�
���@�{]R@��(C��!��˾�@E��ՙe: �r�$I=|�!�$5�9�F+��C;��`CQ/io!�$��4�b��E�d�YV��-�!�d�y��B&�Bn��N.b�!�D_p)�xeP�u��eR5���q!�d��Ag�����;A��!���й0Z!��0*-���vŜ�J�D��ԣQ $!!�$;'�n�"4��r��R Õ.!�dğk4���G�W����ܔ�!�dQ�d�,���=g#<MX�%"X�!��KU��E F�	4�J���i�!��e�8��� �P�	c#S�!�D
�iphɗ�)�������!��%������#s�	3� ��a�!�� ��je&��(�,9�ƅ�e��<"OD}��f�ML>#�&��P"OX *e�Y3:�m:�N��g��9C"O �0�\�,�h��">�D�@""O�l�FÇ
����-�C��]��"O<�S�!��m��B�E�����"O2u+�J�9$�h�R"I	z��!js"O8�C0���/�}�(P�d����"O�I&�W	l�q`��I)a�8��2"O�E� Y4	>]�DD�1wAB�"O��ӓ-Ҩ`φ���E�t��hR"O|ф��7�l���L�-�6�e"O�q`��Y/��@Gl��ưHp"O�3��hE5K/�0g�p�V�\l�<Q�ؖ>z��xC�-l=(�2��C�<���p�D�1c�L�Wy�{a�@�<�1.�2��$X�%	�uv.���Q�<��=bq8C��(��ppL�<I�,��7If�
b��%w��$D�]�<ّ�m����Ƨ;"X�!���^�<�T,	�?�H͊E�[/�����X�<��-_�7�
$���6	BpA0a#�|�<a@C�v?vժ���VT��b�M{�<	"J�"9:���,U��A�w�<Y�a�33
��j��h0��oq�<! M8�:�*��
�Zh�Ah�<9�@��@Ҧ.��a�&�+�� d�<�� �S��ML=>��`�C�y�<є!J-2�4D3��=F����@c�x�<���I^rp�sH�q嬩�-Aw�<I�H�u��k��k���	Bmx�<!6��3T�eKeƏ<�5
���X�<Q#�7m������Z��l�$��S�<�lW�{N�8��ݫQ*q�@�U�<�U'ʭV�$Y!FU Q�n��3œO�<!R$0A�$��ת;sj ��XO�<AGC�yLp9��B�t��)�#&Eb�<)�hTz�Zm��.�& 	t� U�<�+fH�R�"Z!�%Ґ|��hO�O��c��#W���#A��l�q�'����ƈ����$���вs�\)�'L(2,��e ����Sp�"� �'�NE�bײ\�J�JL�/NP��`���pW�:��hjE��6sC�}���d�ԟy����숩hu��S�
:@F!�d	�#�QvhۯcϜ�fL�<#!�d�)z� �a��S��p�$+U�0!�)��pB�Ґ��`WIÄ*7!�D�9"��̪'G$s�����w!�^�Y�~D�Gk��YH,:��\��!�����j�N��q�GL!�Y7?��;�!ߴT 䍰�I�3h,!��̑1F�%{p�?G.!]�8l�'���@� ɍeLDU)���0�
���'�$d+2ř18�`A�qlű07�4q
�'��@`	A�c69���!�n���'���K �jh:q� �,	��(��'h��mV�drp�CE�0|HR�`�'!2L���_�Rh��0#,ш%�B�#	�'A��	��=1P�QrD�"��}c�'��9�� F�B��H1�� ��P
�'<�h�aڪ���ԅ�3H"��
�'�������lІh�-7�(�+
�'Z�4���̬o�8d+��Ț8pаS	��� �����5ل�Ӳ�ɮ�0t"O�p�
a�D�Pu��*adbD��"Ov=��*��{�
5���vTj\�R"O	���A���R��ipA"O�}�n�*S���
4���"O>!�ad6�4*2� ��� "Ox�.e�fz�C�:#�b�c2��
�yB���n(��2A��%��U��+���yrE�+V�n���φ�\љ�/��yRꜹG��i�r._�5�X�k'�=�yb-��`6�lX�R.��y26�!�ybb�1"�|�#6&A�^���%I	��y���:U�(���c��J��Lu�0�y� ��#1E�0,�j���k�0�y2EJbZ�m�P���"� �dJ�y�gH��l�r��nm��k�8�y2N�C}0��q�Lk'j)��ڻ�y���R� �d�:�� I�M��yBi�b�
�(�hX=(�4���ĝ��y���6^2��S�*,40p,��y��D�j(��X�阣� ��PC]��y"gw��(�E��tT0�����yiûU *��G䁝4��I�&��y*L&b�h���S3(�:��J�yR`�H\�ՉI	8���Pb��,�y�-ȕ=��m+�"?ю`��ݹ�y��P�<���@v�A�/�=av"�,�y�'_���9z���*1�� U�\��yR S.R�dLӴ�U�ҥ�ϐ��y����j��[�6N��	ch^��y� S|,]z��:(�Xm�⁎��y�,�L���1�8���%���yR!ӥOe��iE��S B!`�>�y�\�E�*�@7���_Z��i��yr�Q�iGb�ct�E�RQT�����y�Í7eȅ����7`����W;�y���q���Q�$j�y��Ƭ�y�р2�^q1&i��#�"9���yr�V�i�(A �h@��"�9$�֘�y�|�܈����y_N��db�2�y"��6V�j��k��!SQ#��y-�%+ڔ�BoH,14�ub'Ȗ�y�E4)��Zg���?BcS����yd�*�P�lήm���9�ѓ�yRG s���3�N8���r#h�(�y�e��x�p�M�5�-P�ŧ�y��� �*�B�(^&�@Ȫ��^��y"�A2@�  �P�>� ���/�y�m�%�Jxⷮ� �b�RF@��yb�ް_X���̶�I�&�&�y�J
6-���x'�¢'�����V��y��ݫg���)�
�J/I&#���y¯R*���cW��H�j���*�yR�S��<M���O�uv��C ʉ��y"��5Bި�J끂h�`�j�� �y"�ĞC�,�C�	%Y�x4�t��y�e�68��QJ��b�v��#�߅�y2M�;��j�E��T4T��j�4�y2OX�C_mb�H S�^�+�U�y������8R���D���rs��yB%�+�A`�O5��9�g��yR��H+F��0oM�:ά0#��yR<����b�?fg�	F-��y2#J�7,���`0�`����y
� `D��L�%;l�2�K#<R���"O�,K�̶	��Ca�i����"O9�� Pv7=�2� �C�Υ��"O��B���J� � 1�%җ"O���W0c�8)�N�;pyT�"O�"G�?NqB!��;zv`д"O���������rl�yS"OT�I��<4��R,�W�a�6"O*eSQ��=a�$�A�O�wLFyZ�"O�pRʃaخɐ��1٫A"O�=Yf�̏/� �S&�Ԝ/D0y�t"O^��U�ȣP���E�>�@
�"O�a�#��l)Uɐ��!"OftY�∈\4�D`�[;\��X�"O����)�\�T��7�S��� 6"OD�
׿qS4XťJ�=��)0"OV,ȖJ&��\�V���:.a95"OxI��H�~�zu��A>*QB�"OfD��(�%90u���A+�b���"O��A7�\w��s�͆Km~`��"O�L���ܜ�����6SJ�˒"O|�۷�ƭ6�p �C��G�z@A2"OT���`�)EԂ�p�Yr�($sC"O����r��v�͐=�V�C"Od4[�*�52 P�ₗ�0FH "OH1s �Չ4'N�Т��L��)2"ON�uJC�+�|�Y�ؖ�(`�"O�p����"	���d ���&�E"O�!���U�*R&,���
�@w"O�qS   ��   O  	  �  �   �+  l6  oA  J  uU  h_  �e   l  Xr  �x  �~  !�  c�  ��  �  '�  j�  ��  �  0�  r�  ��  q�  :�  ��  ��  ��  ��  ��  �  )�  � �  �  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p G}")7�7�``5�:Q,L��R�H�2��#.O ������܅kW�� ���bk[�%��Q8�(O?����4�|�z�+*�Zɨ��;���d8�SbSf��boۀ��%��R�%��<A	˓ �R��V��2)��KE�`�@�Fx2����}ʙ'�i�|r��2E�0:��L0eO|��A�cR��IV�$<t����+���<�Om���!#j�$�N�A��;M����!�ybF�:l�����F1,*�:�+<����D<�~B��$Y?}�3	��7'�<HB�K�K�v� &	.lOL�x�b�\�C�P� ��f"�!�V�7�y>Y�O4����-F�@���� 	���nW/Ĳ��i� �>a����IƄ���C��r!v�����J��p��I�u���c������Q�^�I�[�xR�|��tp��U��d@h"��?Q�'x�ə� �(C؁���lᓏy���wܓ��'K�qF��F�n��0��	��l���k��F��/��!Bz���V;7v�D�w��y�aפDB�PJ�D��`چg�1�y
� ٱ�d��X'��P�^�@��R�5O�b�`@��<qs��Se�|	��|�2¦��P}�)�'6&)�Յ�7`���貂��DoD(<I�K!	}��*� �m�㪑F��L�>Igc�{9�KnM�9~P�kP�@�'��?��ӡ��J�"�>V4��ˑ�?ғ�hO�Ӭ_����UJ�Hi�)e�;]��	u��h����dg�'�r����fG��"g"O��2oR�T���F�:R�� ��C�d�cbR�M	�����"f�A"�>�Odӧ� �n
���c�jRP�'"O2��
�H���0P'�m���IA�Oy:i��*]���xp&<Df�Ui�'=����&�(-�&�ڧAg�}�'�@�z3Ɏ�`�����B�3~4��
�'7�l�w�_l�lȒ�ͬ&��y�'�ў"~$�P>/�̉�� P������O�<A��mO o12�*���L�lt��D��,D{�'kDL�&��J���4��Mh�U���gyB�˙q&P�h���*�|�� ʛJ�"<iϓ+�~�*�ȕi�x �� ]5ڰDy�X>�pѦ2+ˤ�!#JJ�Y��]�#;D�4����>弈�,
�=� `Q�&}"�|������|b���@�$`�!�A�$R�)B)�yR���v��呠O�l�J�iFdM*���0>�`aɰ2Z�
C�^#Z SQ��I�<a�h�x�6��#��T���CD�C�<i�� ]PΡ��F�*p��P��c�<��撚�ܽ�aA�U>\ ���X�<Y�1&U���F׿HZ�|���HY�<QE�	o)5{w.�&b�qQ��V�<�v�F]|I4�ˉ%#rM*6S�<1e`��~�H�8�F�O�&�ВΆg�<y��F%����b(:18v�n�<�����8 d�Уk?&�Q�	c�<�B�Pm[��a�bל�.��.^a�<Q'���2HY �YϾ��BfE�Iy���O�q��EZ�w��M�{�\h��'Ј� �Ċ�g��Sa� �y��љ�{r�'��x��d�@�P��2o�DЁ��~��:N�LL���ˌ\l0ECfJ�!nB�I"�i�0���P���Y�j�*MW�C�	O`"�І!�?N���b�Q�u�C�I���S���r�\$�1Fx� �OZ�=�}:��#t�MKC�	
���@`��a�<�f�M�Y����G)l��U�Z�$����I�m��a�g����0�#F�MۂB�	=J�x��� �]h� �&+%'�(C�	|��������(�p�	}�6C�ɥZ	ta���.9�N� @��fB�C�	0O�,��#�47?j\4A,{�C�	�a�213����=J�o�o�C�	�q��ۦ@�Kh"a{# �C�	>5������5\�0�"��Z>XB�	!��-��'�([��ɸA!G�*B�	�w��\iS��c'(A������C䉨���Cr���%��(�&syHC�	$�Z�A`Ua��`�'��S�Lb�@�����9ҡ�?^�����Cq��	�'D�X�3jT�~,
��G�t�<<q�d� ��5�I00��EO��!PF�߳-�B�ɀb<�Y�/D�'�-Z%��6>B(C�:�ܣ�&I�2UaWE_|\��	u����(����C伉 * I�\�u�|Ƨ� �D[3ߺ
���1��%f��<`4�$;LO����P�$M�B�	A��Y�S�'��ɠ:���9E�I#!+�Qj��w]NC�I�6S$�z���0:wB�遂��k#�<�?���$A�Dj\�z�n�Z���c�T�yR���� �*OO���t�ߠ��'uў�Ohdİ�,�+d�d�;$㍘D�����)��<1�G�T�x ��DПGx�a¤��]�'{�y�Z4:]�·PiB�uxdi�'��HP#I	�^L��1��?rnQѲ젟x�P��wX���/EJJ�B�K"V����$lO�j6b���*�Yg�oy %�aC�!�hO?�Ү"^x�V�2@��l��g�[#铕y���	Ɖnm|��QHF/'�5�F�#��Y��4�u�0M/�0�G����c<D�x�ӉV��q�掇 �>���&D�4��%����55mF;�8Y�*�>)�;��철-D�{����:f(8��4&)be'lF�9"sʃ�rhh��ȓ-��]��
 &�,�aK
Q�M�'�ў"|ڶ%ɭn��I(ā<<������t�<	�ʒ �.	(ơb0��KTg�n�e8�ZT+0)NP�h���r
����6�O��I�1�bU����洛�jl0ȆȓI\Ҵ!Be����d͙�'���G}��ӭu�R0p�"Sߘ�ؗ�Q���C�I�)��a��[;�8$y'O8*��'�ў�?j��	)�
����E��� �6D��As���$D	�R�2�Z�F3D�	�����ӱj�+�!��/D��qG� �쁈C�N	���AU�/D� 2��GD�>h�&��y0�lKQ-D�([�j�W醼�`Å�C
���)D���G��lߎ�35b3cǶ�5)D��I���q��ҴkS>�P��%&D��
�h�h�H��
ѹU�0e:�!D���M�{%�@*5�MF�n03�E*D��!���~�n�ps�M?DM6,Y�(D� �I��O���F��\
J �uF&D�h�,
8DA�*�8X�s�#D�l	Cے��)��0�dp6D��#�P�Y#jUkf�J�걒��3D�x��T�
| �8��ݷK`z1b��/D����爛,�Ri���3Tb͓��.D�<��"��[~N	˰��!2�%8s�&D�h�Q��|ƚ��Ei�Ј	�@2D��(g@{HEd�\<&;|7/�Y�<A���.W[�=j�H\�e�||z���W�<Q���j��\@AE��{�EZ2RW�<ٱ&چ*���r�ͼ2���Q@c^G�<Q�l�X��S�COq�	)�Əz�<�B
�b�Vl
�G��i�PH���w�<�.%nTƥ�E�F�z��pQ��^�<��*}���v�V�=�`P@k�Y�<9�7EJͩ��M>]VA����T�<1���%L��hБ�9+��y�E_h�<W��"!������Z��`ܫ�Nc�<1�]	pThA�#Άz��\&�]�<�vᐷ\bx�����z�l����P�<�i=O�m�E!	?b����P�<ɀ�) �0[�
J�s�� !�M�<�TCQ�F1�R���(%���C��E�<��ȏ����*�N"7���+�M@�<Q�Nܧs��Q�q�ϙd�H��0Tz�<� E��GuҶ%zDG��s;��c�"O��T��gU���oZ%i�Z�I�"O�Qq c�9\Ђ)h�eD�1�^|ڤ"OJ�r� .Zzb Cʄ�SszՑ`"O>A�W�3 .@�#���H7� �s�'b�'�B�'dR�'r�'2�'d��,�Xޤ���H#lo�����'���'���'��'o��'g�w�.e)ԉ�>'���0�B��l ���'��'��'�'r�'�R�'�>�A9���aąS6r��-���'iR�'7"�'�r�'�b�'�b�'P��:�(�9
R40�m�;ٺ)1��'���'�2�'���'Z��'���'�� ��Ωho�͙`N��@�^����'��'���'��' ��'�b�'�+E� E{��]������I����I؟`�����ޟ��I�\"�JY_ Kb��r��0�����I�����ʟ���ǟL��ɟ��I�T���e��=�1�L���$mɟ��ܟ4�	쟌�	���	����˟<�S��3�̺r�� ]�*Kf�Aߟ ���d�����Iӟ��	ş ��ݟ�u��
V������XO>5k4����T��ß��	�@�	ğ��Ο�I��l��G�Q<��o4+d���'����I��,��ܟ���ϟH��������8��<Z>�cD3{����Q�0�����Iޟh�I�@�ɜ�M���?qb�A�=�8��G�%3
���}���ƟȔ����T֦͒䌃�e���2t
���d� I�0�`�v�'�ɧ��'C&7X�DYJ�92M�,s$�t  ��H� `m����Φ��'����A;.k6T���1���b~ �C��ֺ%��xV���O�ʓ�h�f��e���=p#���	�:�X������S�&'�l��>F��w#��c���!]��L`�N�0�Z1�{Ӱ�l��<��O1��d��$k�z��Ȱ�	?�~E�@�"	��手�0�C��5�L$F{�Ok�GA�u���6`�	�JE�e%�y�_��&��zش#hX�<q��\�`/���bC�&w�T9bw����'�8� .�v�f���g}2˄%V��)g��0E�*�	Am����%1�^H�d@Q�a1��`��q݅��g�����!�r`ұ�P�/�p�y.O���?E��'��q�ѹ>��t2% ^�nѼ�؝'�7mm��I��M���O<B�a��	�U!,U�7�d����v�h�4~F���'����V�i����7Rzi�sƙ��j(���7[��}˴h��_ߴ�!��G�G��"v��{�>�X�̙,$D���� t�p&mU�K��ya�B�[�5���)Zi&O��h�V�O,2hL�'K�P���:�KG�v��R 82A�x4Kz�H<9�̊Z��iS��i0���W��X�U�,G�ԑ�"�i�U-��J9D�]�$qԈ��ٰ����>��)EG�m�>]p ��r�D(	@O��j ���Um� �(��ȇ�
�\I��B�A��0�f����L�!Zi�^HК�G�<�R�c��ˤ`h�H�O27�1��n�����I��h���?M��ޟf�p�dz"�=a��vD� ���O,��Q��O
�ĭ<ͧ�?���6᪴
����ɗ(�~�@̪�i6�5{C�rӾ���O��D�����O���Ov�����h�.����R�g��R����-�������O���|�H~���p �7o�;��D颌�+�j�` �i���'U�k���6��O���O����O뮔�zJPD��
y$D����H��	`y�a���4���d�On�D��S���P��J�Co����*o�mZޟ蚦,�M#���?����?eZ?9��q�T��_�I<䨪�A�i��'���0�'�"�';��'WBY>9��˯L���0a|Y�<�s���/����4�?q��?���+��STyb�'�����lڛ�L$Y
��?iXAr�ɡ�yY�@������I䟄�I90;��pڴf���b�̺<� �;F�`�5�iz�'q��'�RX���	J�S�(^����M2:�Y#ɗ�ndM�O+���O�D�O��DW+T�(�m��h�	�9�Vh��눈�����y���Iߴ�?����?�/O��$�r\�I�O�����M�R�qRB i�0�ࢇ�9ff�#��O��$�O��^�%��m�ޟD�I�d�S1�X0����e:��S!��q:^e*ݴ�?�,O���bP�I�O���|n�/^k���%��t��R����Y�7M�<A�FX1F֛v�'b2�'��D��>���8lS���^���+�X�\N�mZǟ���\��h�qܧb��,�2nV�.h�:plz��m��r1�Up޴�?��?��v���Zy2dQ�z��R$�T?~Li��OޤAĂ6�T i��d#��1�S���Z�aAh�fa���[�H��i8���M���?��{��EC4U�`�'���O�;F�L�w�H�t�	g,b%⡱i��'�.H*�����O��d�?�s6mֆ-�̵AA9��}���cӶ�" 'xm�埰����D�	���i����A+Q�NАh��
}m��ۆA�>���M�<I��?i��?���?�����I�jR�+C~8k� Y0��(&�x��f�';��'��~".OJ�d̼',`��ݽeǂLH��/4´MR!1O���O��d�ON�D�|��@3��v˺$��|�a��*�T�x��
�1��6M�O���OV�$�O�˓�?�a/��|�1Nn��1�C����0O�!Is�	ܦ��I6i������4�����z6�L㦡�Iџ�an�fa��v�Or��Y�R%�)�Mk��?������O���E6��˓i2R�H�e���j�r[���eX@ʊ��?9��?��_�vd�i6��'"�O��Ļ�Ϝ�5�݊r`�`~�{r�r����<��W�~<�'���|n:� ����l�!j�$)�B�;�L�`�i?R�'}��|�`���O�������)�O�1����'�Μ��憈�.��DS~}b�'D��e�'��I& &�e�I�5F�Y� �k��7ʘ+t��7��'iR<lZ�<�	㟨�S�?a�IΟ�ɂ�P|�A�.j�l�8� ̂f�ikݴk�����?Q(O�i7�i�O��xB>dp�S�g�&�n@������	ן���6__���ܴ�?Q��?���?�;f����݊T �Q��5C \l�Ny�P%` �u꘧�)����Od����,6�D�7*&8�@�3����=�ɢ�XE�ܴ�?���?Q�� ��K?-_�&xq%��mfL���U4}��6�J�Γ�?i��?	���?�,���a�ʙ,wR*�J��T/�� 3I��l�n�@��џ�������<A��?�NY	Q��'7&��	"
�`�����<i��?��?��������=ΧF�[R�_���\*T�Ձ?i�'���'��'��	Y�P�J�����|����G[�D]�'_b�'2Z��PI��ħ<b^��IU�S)���V)]0����ir�|2V���m$��2~�����'֓o�����h۟[}�6m�O����<97�Լ&�O���O��H��B+��=#�"�;ƨ�+�3�D�<���_���	�8T�&��$B���u���Z�Ls``��M�Y?���?	K�O�̃�)�+�l��"���2Z@�շi��	 L�@"<�~���#6	��LT4'(�!�2�	٦M���E��M���?I����'�x��'��<����(�( ��X�p��[��w���q�)§�?��B�j5��Da�y�-��ҦP��6�'��'��壔�4�D�ON�$���	�.ۼsg����f� 4
V �5�-���YMc�,�Iɟ��ɺl ~��t��xPċ����Y۴�?��R�O��$#��Ƣ@���.Wn(59E$� nRn��EP�c�,��ڟ����t�'����C��R�P��)j�4��*�9<�O���O8�O�ʓm��i�#�24B�:�'�??Zt�+CB̓�?���?I+O��"I��|rAcݦ)S.8q@�
����Zd}B�'�r�|RQ�T:Bn�>!��J�L�+&��7u�,� �/_}"�'���'��i�C�� w�Ӆ1�Y�5��5�`�7&�� �:�4�?�I>q-O�����ǡW���V@�p��B�=y?���'eX���Q1��'�?���W���E��(!׃�u!��p�xR^�|2�"�S�ĭ��!�@���Æ����kʻ�M[+O�h�Ǧ]+��F�����q�'�~�PҎ+-��T�׉	���ݴ��+{4�b?Aڣ�/(
�&1t��	rBu�ै������Iݟ��	�?�(H<1�&e<�H�'_�98��x7��-a�T-iD�i3������� �cgϞ:��P!�J�UV�ء�͸�M����?��w��Y��x�'���O 8�)���T��i	9T| bt�D>�1Ot�$�O���æZ�\,�'�4X�nHs��3k���n˟����ݿ�ē�?������3�b�PQ�0�����M�f}R����'���'2�T�\X�Ϝ
3����J��XKĠ�G�҉+K<����?N>�.O��r�ٜRb
y���G_g�\Q&lC1O��d�O*���<Y��
L��	_�):�ԲP"���`�ܙ<`��ğ0��H��Dy�.��DW�'�\U��fܘ`��\ sI� #^��� ��͟�'��8b��5���(#-�Y)���^�ԅ��l�A���n�ҟ�&�ؗ'Fn��}�&�{}v������.U��M����?	+O��` }���@��{`&M'nօqD�S6I��^T�L<�/O�P��~bt��=I@D�a�G�O�x@Pբ妽�'OL�{wib�P�O!2�O_ ��vu�+ݗ
PB�� �܃U��Po�ny�G	�O��d�h�Y��jD1d�7��� `�i���R�kӆ���O
�����>�����@��A�N><�aa̷x�����O>�����e�٢\�>Y���3<1����U���8��<-+��#�}"�'���Y��X��� �1n�8JA숒��O�����O��d�O����?>�h%yt�_7���ڤ���	�	)�0��I<9��?�����P�ũ�>;��LA�/[�����X���,�IꟌ��˟x�'����Y�^�K2����8Q"�¶s�O��D�O��$�<A.O�� RlW*r�6�ʅ�О8�3��ކ�1O���O��D�<��oI%�J�9.�B%#�M̢�z��~����l��[��jy�����$B6fZ�۳��4TYm��'0t��	ٟ���矤�' ��D+��Yz�(�S�@�H*������DE��mZ���$�З'fh�9�}�L��&��i3W�ѯ��WC̖�M#��?�-OP 1�ŐS�����&�P�;��Pz� ���8z�6��L<	*O��j��~zt  �jp��BF�c�00�!ۦ��'A<�Z0�a�ڰ�O6��O{�H㮐Jq��9@3�,q�N�91��l�UyR���O��bЂ��v?`�P͌�
�@��A�ic�`�@�g�@���Ob���8�$���Ƀ?>.=*�hZ&O�J@�e۷F������?)U� ��(��D xjN}�g��ElhhA6�i��'�r�N�* �OF���O@�I�n�$���5�y�#���h����OD���O�����D	�, 5t>-r2����M��^:@9ఒxr�'=|ZcZ��c�u��Q-�u� �����O����O�ʓ@7
��A� jyS"�.l�T���/j�'�r�'��'�剂w34<p��%��E*���8}|�y�(�����˟�'�@���m>�ڒ$�?}#�E�3��{"V@�FC/�d�O�OD�J���'�u��n�3o<��A��\��X�O����O����<�.ʓA�O�"0��eX�G�D���Ο�tP�Q��sӺ�1�$�<!��C^�m��i��F;7݊틶��7�ZPn��\�	qyd�1������	��޻<�LE��;(<@�Bd�]yё�O�ӫ6x&����d�p<���ķiy�ɥ"�d!�4X|�˟l�S�����x>��r�U5\pI3�U�6	�_�(c�.�S�{�.����O�@Fds�&_#_Y�l�#����4�?���?��'4ٱOlġE/��g=�A�H�''؉U�JҦ�9��.�S�Ov͟?*�yI�C�8�Mۢ%�U�7�O�D�O,y�B��r�I��X��y?��i�P�,�R�':�� ao�8W}�<����?��5P�C��/X��r�ʝhd��3d�iv"�	Z�hO��D�Op�Ok̜s7�Qd�/?�A����:�ɵ,�c��I����dy�
��.�eg�
~��B�G�f-�lA�2�D�OZ��"�d�<yN{��ecPb����Qb���yj�Y�<A��?�����@ (�6��'H�䠖�Q.nJ�Y�E�cm�M�'���'
�'��I�8������A"��i몉x���`Wܼ�':r�'�V�T)�\���'G��@bao�s��bp�0g:A��i�r�|�Q� ��>��7�^M@�n�}F�P�U	'.��6��O���<A�dG;��O�B�O�^yf�Z�Zמٓ�	4o�����n*��<)�%Og����ܕQ��yTN�0I8�@�N�1�&Z��{�·�M�QQ?1�I�?�Z�O��k��.�>X�Ģ�
�4R��i���#y�#<�~��&��oQ�HI��x�����¦9k#�ˮ�M#��?����#�x��'���	$��"��$�!/��cO:�� (c�8�
��)§�?QGM���"��ꞁ#�D%�F�'���'��(�b�$��O�ļ��s#.1[9�
�#U��)�w�'�	�4�c����֟`���<���b�'�l� ����
�/=T�ܴ�?!��'>�'�R�'�P��؝�ٳr
�<a�2jI�
�d�8����<����?����$��pCn��f��O�Z��@�֍s�0�{��{�	��������'���'�Z0���ƉF_���t��7D�J�X��Й��'���'��U� 9�T<��� � T=�yb�fԞA�"�J�������?1�����O6�DK�tC���j#�)��᜘+)��y�,`t���?����?�+O�c�%�[��
cҀX�FD�1q�@{�M��k�<ѫݴ�?i�����O��d\=J��>��\ �(�ٔ@�.��P�p�⦭��ԟ�'`ny�d���'$�t/�X�< �@ ͆���a�K8uD�O�˓^~=z���x{2���*��D�����eK��W�iN�;a�A�4mU��ԟ��S�����P�"���M:E���H�#�h���'B�V�yr�|��t"[�E��`8P!�bDT�b��D��MccCTi���'�b�'x��� ��O2,���N�|�%�����1������-��+����&�"|�����0W���
�e(���i���'W�R Z�ZO����O��	 �����7w�;RHއ%[�6�0���7U^��%>��	˟L�� *�ٹ��ڴN��)5� _�R۴�?9�IDL��'wb�'�ɧ5��3|�PŊ	C��*��_��$�"qV�<A���?Y���W��H���0�Z���K�0�)#@�I�������Z������y����R�ľG�})�
Z";�f��¥k���'��'��_�<"�1���	a>��ʳ���v}
D�����O���1���O����~�0:s���@đz���꒠�L���'$��'��_�����"�ħy��)1�G�L(�s����愂ոi'��|�'&b��"e,"�>��dՅg�x��`�2J��2�����IӟH�'�L22�"���O��i�4��9�e�B4i�TpQ��%��'���I��4�e����X$��'ST�9p�h΍'mpUQfE�� v�moZ|y�됩,I"7��v��'��K2?I�`�Xh��K�������	��D1�>�S�'Lozd��.�;��1����%X�r�o�e��1��4�?y���?��'z�'8�'C&6�H�"�Ιe����O*rj7�#�֓O��F�T�'�HH�a�J:)G �'_�\�Εc��uӒ���O����DCd�&��������1�Zti��C=�B�����>?�p�nZJ�	�y���(M|2��?��]��g�0�]�����v�DIG�i�BB8,�O����On�Ok�����8e�X�DRV�#g'�f��I�D��(�	xy��'�R�'��I��� 6p� (�f|!
��"���`��$v��'CB�'��'BR�' �	K���)0�w
[�k�.a0����2o�W�����8��^y"�DC��ӧ*&�����8�������G�r꓆?������?���*�Γ�N@�E�ho6��4F"+}�Y�UR��.��R�υ�_��)�')�����C2�����L����(8R�+��Q5H�5�fjF�q��t��J��M�oQ4W:����d���Y�_�)hw��._�q�cF�D͙d$W	o�R v��,th��יCRZ%�U��[#&=�FN�lO�-X�#XS���Z���66u��7�܏o
�Ѡ��0x�%sQ��t���$"0
r�RA��/w&T�BǊ�sX�q�@�˫7���1�O�D�O�����:<{��1Ц_�Sp� �fƊ�%V�|���: $MoZ�6�&�p�Ak��w�L	*AE� 25�����A�\�����=&8l�P��6��#J�cG�
6
q��m��/0�:�NÈ'�X!�G�~�� ���'#r���	%��,����!#^M�&"˜Wv"��ik�D�ISx�t"W ��@SN�[�j��c��l�R�*�	П�K��4�8��_3
��$������v	2�'�>jK��O��@�_?zX��O"�D�OD�;�?)��1pP^
�n|�Ч؍P���+¦W1�&�ؓh˟=��6�u2���DbPb��2Z�Y�VÓ�k�v�����d����g�x���ݟ�"=�7JI�Ov`t��L�&k8����Wq?�3��ݟ���4��F�$Db����Us�Sg<[ϒ�ɞ��y��G9dNP h�De�����"6�#=�O�剰<��4E��1��śZ^
 ��N~,�����?����?�5!��?y���$J5h|>1(7�[w ���:l����V M-��y���FL�yR��yB:t��A�y�P8��SB(fȑ�.Bd�x���Dm�y�NB��?��`��1�� �Bq���<X����d>��m�� �G��4���e$ʐ�
D�ȓ-�.)C�t����(وa�$ΓN�	cy�n͇���?/����޺89H���wtZY�-��B�����O����$h��m���Q�(o�]E.Ń�M�O�䅈 �/n�$	wA١C��{��d� S�6M����'E�̐h�Ǘ��O�X�@��'֩)Ĕ�Aǁ�Q��k�O�lzI�~Jt�� Ma��٠��*l����1J��<��u[L���@�DF�`���Q�]fR|��	��ēaJ�D��K�h�r�	5%��̓O�Y��^����d�d�ĮB��'�RD�>�v)��g�,on #���
U�Q�S��L�I�� ޫ53CP�5Ȥ�����w���ѕ��-` ��Վ#7���N�g�&�����{5�]q�%��B��x�թҾ��Ͽ�B̟bq��*.Y��0�J�8P(�����?q�O�O_�'�M�g6_�ܭ��Dl�'P�=�+ǆ �*�Q�Ń!8m��y��'��"=ͧ�?ɂ�����T��k�`���*U��?Y�6�҈�ʊ	�?a��?���g��N�O��$�}�8	0�DD�	a��A=&�R���	_NI�}9o�� 
�Pb�ݟ��C��*Ϙ'R��"5E�m�fy�fJ=F`�p�c�0d7r%��W4o���j7'Z�����Įb�|��<	�T�t��ы�mFL	a�OJ��?)�k��?�i���'�B�'Y���yW,�pD�qC
T`�����y2e�9Y��) `��I@���y�h"=9"�irY�T A#��Ms �7ĥ�#�RX%ag�S��?����?��4���x��?əO��p��6�貁�ڜ(|��!ꍀ
 dJ�I�)n}H
�.�
��.�� br�3a�H�a�%��\ �@�D9v ���	�L.>��Ț�+��աUz���Z)���@��,�M[��J#��<9�m� ^���Ǡ]��a|�<AC��\-N��wZ�d�� 0�!�<1"^��'"���e�>�����I��6m,0y�^;B�x	l�l`Y�F�O��D�O>E�e+�3I�x��Ңp����|�F �rNd�u`�	QX
����x�'oH�����E($�y�	f7�O�yZ�+l DU��Mǖ{+�ɏ򄏑|B�'D��R�� ڠ�p)��x�T谠=O��$/�OLঀI^� !5�H=঵�g�'�<O�@����>y�S/IŊx�T<On�)`�����ϟ��Ok�u���'��'��q�i�����@��X�Z��A��)P�-�f]��W�uh��D���v�P�m��NKB��6�NS:=Q�t��^����w�_
#�4�B�\��p�	V�F�%qk�!'N�����w��M���C"��"�kXzX��	Z�ai��`�"d��*���'<�dB5�Ґ/!qb��ãm�B���'["�$)ړT����ߝv~�(qf��k�l��<����*s�6�O�	��DXX�.�8�<5��YlT�S��O�đA�h����O(�$z>�$�S���'��MJGkˈg��A
�3L�C�'�����i�z��c��\AR���'jDt�CnE�H�4���3R��PG�KOazR���S%�Y���,Y1��Ӣ�<G�b�%n��zӆ�n�?��?�/O��"���|<����ˀl�*m8r"O� �����?X%(�y�j�T� �&�g�'f�S[y��R�R�6��'u�Ȍ����-W��U����rf��D�O��D�Ob�$��O��dc>M�ĦK�Q2f���蕊�2 ��"/p�N���ϙ���|��&Q�N��d��A��S$���8��t:hBq�.)��ɠQ
���զ����71mr��G��sx>�0nŒ���?q������iI�'k��3�A*y�Ĝ�'��x!�d�X�42xT
�K�z�7OHa�'�'�"}�CoO�>�Ωx��+bIt�`n�[�<c-˴��ŧto>��Co�~�<agE�%eo�daQ�H+/�B���.�}�<	�@CJR5IBC��%�(Q��C}�<���3}'UY#?{t��~�<YG(T�VP�Q��E�B��e��}�<��cR�?�ܸIb�>A^�3��s�<	���m<(���ᅴm#jyXa��v�<B�'x��qy��U0ܰ�����u�<�֠7�V5ѵF˩�H��KPq�<�&J��D���e�K��,��K�i�<9bhL�'�10�f�!?���"�]z�<�� '#�
�t#N�ty mc�u�<y��P�.k`�����k(�;��V�<��c_gF�1�ɕ�qw�9K�q=�'@��0+�3`�$��@� %+����'�`�䎰f���G	]�ۮ���'��jS-̀@�B 9�i��R���'�Qb�_�i<����(Z&
���	�'���I��f���5� Ќ��'#Z()�q�>h�5��a���'S<�k��(B���D �G���'|�,@ee
"#n�[�Y6�K	�'R�6��=,�Y8�<�c	�'�T���@�?]z�S��\*Iу�'�9�V���lo�Y�L��Q5�	�'0�Ujfc(2� X�$�"P{\(!�'Vm�]�<{�8�.ҍ(�@��,$�C���	"-ΐg����!~�CQnQ�#�A��H�T	N��� ���ɓ�N/kbfy������ȓ: �Bh#\)&� �$��I��Ԗ'p����� �&��W�O�ر"L-V�*p␌�/r9Z��]���`�NIh��,O?�8/öqtAB'O�e�d-��AU�#p2m�'�*,� cA'N*���OL�z��ؼ]���3�5TږřuŤ��H�h��/��в$ތk�Q���ų�v c�a �Fx���DK�%d2��a&��h��ٽ4�\@J>��e�:��1��!�=[b���� �h-�Uo�(�b�<���b����<@h,�Q7�h��WG�	�b%`񥏈�<����&}��[?Q�x���-6y�Ƀ0	H��?%?�a��Q?u���˳"K�r��8�>q/L�U٪����X��1C�Z�'����Q��&����5H�%�K��$��D���U��OP���1@�et剬;�x�4�r�H�w�f%AC'�^�̣,�O��ؓj�;1f�M���9;�X���})6�g.�4 ��GiN�e`��<�s��Ra�K�Q;��@�C�F�[�%F��0��a��K���Z:�`��F�?` a�ٜ�(O���	�X�*�b��V��!�;b0�-��ۃn��"��ȵ���bW*F��4Lѩ4ɇ��1�C��Q:�:�P��Z��	=F刭�u`�	E&�U��K��j�l�n~r�"g��� ��$Gv2�إ��5�(O�\�v�'M�����2�ڡP�$���B�	<��ĭ'\�4�w�FZX*�˔�C:�~�оo>ax��αB6���AD�8����(����)`럨
�D劗Aʭ �iz���k���#6�9a���2JLb1�3kOzP�x�?��⥡��T�����-�zi�&���JFy��z����%mvzh�"�`����f۬\� ��_XS��2�I�o,���?��o
�Q��}��m�5Lɶ3`������Ɍ!ʶ��cԝE�0���	Ҟt6��i�5nbT�c ,(��8k'�ap]�?�$~�q��#�`@sQ�I�x��	R3���#�zK�PmR l�!���"1kϙxr�V5�)�'���',�'��r!뉎D����� �=B�y��	W2��J���(O���A��!��I�,38ѩ�P���O
q�Wi/�)�3� f\���'�4�r�-2/�Yci֕ �<��F��5��,�^7@�ż2�� ]�	��6�j����D�05]z��Ot&��X�>X&ܢ�I�R�1��;P���*(��1�ɬp�؀ &J?l�nP�?��ob��׈W���HTa����"d��C՟<�A: V�Z @�!���iL',k�O��eܾLa�0~�E�u���dP�@�m�x.DRD�
�\��J�	�-_&��*Q����aA���]�2��GFݾq���#R����=cX��C�,��<�'/UB���J�
WP��p�
7.����V-��(O��B�*����t�n���:6����.�)vŒ੒M�K��c��ON�)�O�|�\�s-(�	_u��ݑ|�`�����P�	e ٶwqV�'�X�:�*\CH����*H�E�0�h�5�ԟ֥eJK֬9��m��1���[�bM
&�˓��gj��ʊG��pyi���
�sWG�/�L�X`�ϰH*D��7����N>�O�ݔ�yg� /p�4��H�*<E1`�t���o_q��E�f�C4C �Hc���ˋ�,��1A���wf2����,���*^h�1�Ix���I6=b�.��q�O�"Y���Ѓa	̩�q��/:Δ �%j;����GC�QQ�N�}�t�+!�w��`j�Z�o�F!�ҊU�āg�ªZ��Ńc�&��T��f2@� ���t#�K'8U�����@�3�6ys$Y������N������	⺐�ŭ|����'7V��i�rJ_�w^y1D�Ӌ�p��z�]��z^E��D�Ot剞y�z�j��֫9�Ar�^A���S�ǈ69h��'i�;dw�(O�I�~P�nލ� X�I��hqC�Z�M,p����(,��d����6w���I���/��">ͻǺ�iU��X����	Q���O.�a%$�)�ӛ#*�m��"J��p�����#M}��;��'4�;��3��`��J�Y
葪2	�k�(�!�{�E�?��cC����PD�D����O��+ #�����w@�$�dYP�	,'d
�
��T� �\� �������Ñ�L�{x�!�d۪P~xq���O�e���	"�����)�����	�z�p��	��MFfeX'LXK6�"n6�Ҵ�،Lk�id�P#u�'�K��1	�OW����o��2��ճ�A
�x$�s	�Z�r�zFÛ�u:�s@�V�8h���Q%��'��d/�S�������뎦C ����o�Y�j��S^X�����|Qt��0��P/BD�� �2E����,����'X����BE��(�+���$��9C�K�'n�*-ѫO8i;Q��"\+�HOZ0ѡ��5���/��](ly�O��r0�A"�Y��F��]	���!�����ҝtZ�HD,/	�f8�wE3ړn���Y�,�'P�"m�'G+Qg$�nڛz��D� �I�mzd�j!✄]��g�'��=�ǤZ��̙��DB�TQ�|P%��38̪h��'I���$���P>2��a��d����_�����	>a�Q��2���;F�~�����]��M�ЧB�J���ēo>��eaƥs�d�h�%}��'�i�@��4��;2j�b �|b��	ƾM˶�&(j�J��<ɲ�?�)h �Z"vB-� U��)�ԭA�@��9@���M�"�E�4*�Ѱv�az BsPr���%y��k
�HO�a ����~bA��<c�ŖO��iR)P�/m�m37L�~p�M��'-�4$�3e�r@Ȗ�34�&�ri���R9Q2�O���'t^&諞w����3,��O�µP����u�^Q�'{���ɏ�Yʩ�-Z�\�kVi2ғ
�y��O�Ce����)�$��U��M f�^-D_b1��ω�:�ў��%k�0����S���(�q&��O�N_�]	�h�bIQ�#���E
�!1��d��n�8F�^?ڤK_���dv�Zk��}���`�r���D`�.]	eE��O�b��DO.Q�	�2�O�#<1���� d�6�,�H%9�B�C��|"�P6��>Q��=��](�Ǎ�.4H9����8u�:�a�O�=�Ok8��;
D�X`��8R��Q��Q%+P�}��	�
֠=�&K��]�jYk�٩=:z�P��P�	�)��'��������ا��0K� S��	)��S92}��e9HG~���N�>�HO���Eȕ�\��ö��c?\�x#�OL�"u�8?qLh����z�<| rF����gJÞP�������s"\�8P,ړ\�x�R)[���t�ԭɛb:$%l�c�*d�IǵN�4{WD��D9p�I~�'����%�Լ}X@.�1/��\���-J̙��'�7cV8�c��lt��h��1�f4��>x�Q��'I:M�;]�n<���ķA�H��g
�=t���ɢ^:L�q�ɦ��d�/l�� ��ָFt㞐PBcL:�!J2��3�yc�N�?a�?�^1!M�,A���
ܱ>�xa�'3P;��[0G�����ߟW�LI�}�'`�����6���8�%E��B�D��8`�1�~�j���c���'^<	��P�v�"I���X3Fz��S�@��jc#��8�(Q�1k�<�|�i�uceh�Ւ�X�8ɣ���0!R��0��֯*�v.[�P��C�0i]Q���wp��%�lB$�рZ�x~����]M?1*ɯFTb����ǟ�ӄV��y�F!_>��F�ل@��םL\`������N�7BY�A��ǽ���	� 4�A�a҇h��L���1k��ja�
+<�heA?$�&|��c�j���4 �+�*\t`�0��Ԁn�ԸZ���!4&u��֝��܋�fκ�O�S/!��IhS$ÿ$���A�Ƒg�&b�d�d�)��	��v�2�I��[=�u']����J�I�>�(��$;ZkӣS�\��u���C��2I>�OqO��˚:���F� q���xf��`a����K[
+ĀӆM�'v��<���p��&cz�XkP����#_��pd�Q-l�8��'���%d'�y�X
�uxEm��{������SAQ��ɛ�^�tzAe��;*����S��$�aO�u�*0�d "`^Ь�K<aB� @��[��D��|2 -,aSح`�H��<e�A�ç�Q����'�|�+�=~�����o��ilV�Cش���|r�MԡЬ�#�5��ܪPM�wYD�O�7����:�j�5�d9�N͚���9��JDB(~�R�b�O���:�5N��$�����Ƀ5fؘ��SL�R��}p�G��^<Xa��I�zEy#Q#�'G�dI�Q�3��?�n�� �M�%������L�s�\(����)*Mہ�Qp8y󥦕K	�AÔ��*Lم�A-^�8x񡮅!�yg�y$)� �/F��=��aF���'@�a�4�ԟZ-2�띜:����M��j�ʁ�/@�a���'�T�QĦ8�����]=�����'������:w�:Y�f�v$ �sD����u�$�DָQ��k ���'Z�ݺ��	L����P��zM���ύ+�ؐ�b?�)ڧ66��J�i�	3�2�X��G��B jcK��D�27"ӨUl��%��(O���m�g�#�"��9X�(�ODT9�)��؟L�Eۣ���Z���/[�Q^~,
lL�]:��Ey��G2Z���'K��~-d\��M�Ԥ�<:} ��5 KR����"�m�#�jyP���d��̆�!�H784k#'Ϣb̾�[�$�t����a�::(��gY�I����N���C�oA&_�"=Qc�D˚�
�����A�'�<I��A�@jhi�D�:ȂB�5<@,iV#�*z�Z=���<��̏�ez�H�8����1*K�IY��A�$ha}�͙�up8b�#�/[�={E( |����T��2��ClÃ7D�Aá�	�y'��/T(�s�nE�o+�U��^���>	��V�GBZ�C�ᆃD�Ӱ�/cB�q�:l��9KB剓dD�Ѵ�
"o�B�u�,]�6D'a~)Ae�XI������9&@��0  ������Ш��H��X��3`��9�/��� Y1Հ�/6����w�*��Ě�F|~����U�#�T����ߣ ���XL��<�oZ�r h��f� ����7$Qrm"BoU -T���8l��x �)�F4��,Oʕ2D�L�h`�2-�p,i:W�L	�̵l�FX�8�󏔩GBN ���@(�Rǘ~H�x ��<0h�B2m�O�8FyR�p�ѠRhU�N���K�j#S/h��s!)���#?yC��+	�ph6N��jꌈF���rQ��
�����6ʓJQj��B���2�P��*AA��mZ2FF䙧��Z��j���A$D%�OV���PȉI���X;DXCSg����'�)2��&����-�y�h�'Ծ1�0�O.9p̙#H�.Fj��t�O�����.Ț�pIg�X�$���@%[-���B���H𭑿��O�>�4q�VC���h!�C�	ք,@�� ��~BQ�]BN9�"l1��$�+TB�M��(X��`����	��xY�D!�0O��ۓ�ɾd.P����VD�s�Ȁ%2t�9j�@���|1jqHTZx�8h�L��ok|0�%TI@�Ik4N@gt(��Ri,��D���`���
���-
�l��'Y�IZ@]�ȓ�5�ӇW�qC������r�ąȓ!���@i͸w�0��5!�*�vȄȓ1���9%NW� (��� M#5�R܅ȓ9=�����*6�����f,N�ȓ"�,����+T��&�<`��Q�ȓ3>�A2���LU@�!R�L"��ȓN�y�D�91<�ɡ�R��v��u
�I)�@\��I�lo&ՄȓNș��ͻ%=`jp$V�{���ȓ\�ֽ���.����%�DH��M�8��d��.y�Z �����v�T��pl��)Jd(��%�a��H�ȓ2^���<V^���+_�����ȓW���b_Qz����:,�`��ȓ3v�AŮ��`p�0���X ^�N��ȓK��Q��7O:�2@E��}���ȓ5��9!�Y��-#�v�n@s	�'��`��RQ��{���b��	�'�v��@͍i �����>"V���')��Y&�ۧ�xp��.I�qZ�(S�'� �� � ��<�� ǡZ��� ��� �p�/ŚA����Ī�`���"O���FS V-�\�v��'�� J"O�Tf�' �Y��h��r��[!"O�8p���j���h���{��	�r"O���H�=$�P4�î(�����"O��
7HX�[V����kF��*��
�'��6b�?��5Y
M*g����'��yۀ�Ln��DK�,K��5 �'�U�4	���8�%(>6|2�'m	Q���hmQ��]?&���	�'ܚX��DJ��%�4@�)&��9�'�d�S����iVı��G���h�'��y�� ьz ����
��I�'���@E��0�~��h���
�'�V���#�PJ�آѥ0(؈B
�'c��c� �Q��̚��/����	�'mz�K�/��w_���qNV�
����'�
鲆�>c6�A�W�nn�3�'��P��M�q�iS1��1;����'��d@����|I.�J��/�L���'�B�X���4qԽ+ǀٻ+y�u��'�P;�D$Dv���>&T^q@�'�^a�v�J��مk�8!|��R�'�	���nۨ8r�C�vHa	�'��p tO
�H�|a�a�j|��i�'g�8��ј�T��*�d��Q�'���5=Tq�wHd��8H�'
�d��f֛6M ���	?�:���'d|�	����Jyfآ�[;V)c�'�,��%�Tі���|��z�'U4�Âh ���W�y`���'^䌢4��/+�=�@�q�
-p�'���* N@x�Gd�zЬȲ�'�)2�W~WL��w�G z��(�'�Vh�҃��<��8"�s.(�x�'j
M��ڏy��@7L��_����'�>��cϒ�w7���7��9(6����'�Ȥ�U��x
"qG��i1tȲ�'�Ȱ����x��HVDa�@�j�'��Š�GM�E&XR�ԄZ�'j��AB#�)�@h1EjW�Oe,�K�'���ц
@���-X��B��a��'\4-�Q��R�s��?x`���'Ol$8h��	����͎'9o��j�'?tm�e(]6eǴ4�"I�(1�pa��'�2Bdl�_Jl�A���$�8B�'%N�x���y�f�q�^����'Q���,��~�&�2D%_4�%3�'�2��n�16%�hT��a�^[�'� x��e�/v���4��k�dq��'#l�赇џ4�F�z���-9XC	�'���pEZ`1D�G �.��'Ȯ�h lҬ6���0K�v4�	�'6�b̖�&`x��N�w��
�'+�0��$��\���@�I�-��'~��W)������$��'�� `��Q"9�ı�2޾w�>�z�'zqj�o�/3!��##Y t����	�'��<�K>d�:a�E��6똝�	�'���9T)\�#��`*�#X�i�'=����O}T8ऌ�"�Bp��'hT!��Y9�C�lV66���'� sъ�?�|����8t��}J�'
JMZ!�>9��s�i��sDNia	��� <QB�-�z�����U�9��<:A"O�%����
a�dH.O8����"Oh̸@����؋W�6F���"O���R�P�L�DІ� 7� $ґ"O�,��*S��={�)Ֆ��\��"O��׉��z���i.�i�	^�����)M�5�b�A��[�B�#O�!�d]�u����&Z��H� �'�!�d"l����cN�\��}�o��Q]!�D�<h* Y(%�ǥ8��!w	GF�!��>y�DHlC�9 [�+�!�$ y�0��ê��)� �X�wZ!�$��{-^��7HY�n& �E(�xR!��2<��g �a�8D�V�_7!��`�l�x���=ʾ��S��)s3!�"t|$"V�ҩ/��}�U12�!��Tx��-E�F���i7Cşao!���X��ݥ5�r 8�BT�!��]�C����p0�/\={�ay"�#k�� �J�z^Q��	��p4C�<2^��Ac �f,XyAwg��O��=�}�Wmύ6��f"S%@{J<9�%�`�<a!g5"WH�ڤ�^"<,"Iɠ��f�<��̓KjJ�1�K��nlsM�z�<a�I�<q�r�a�H�J	K!��P�<I�e�C�.���.�^<��7c�M�<�+��e����*�H!B����<�¡K�8͖	� ��i!z��Cs�<��؁O���� q���	pi�Z�<Il�-LAq@�P>S���W�<� �"�ȓ�@հhܱ��i�V�<Q���Od�p�B��L9l��ue�z�<aƤ*x��� ��1��!�r�<���L&R�8�AV��X7�I��m�<')��*���M�0p��]�<I����ٳ��67~a���\�<�un�'rE��c�N
;b� 	[�<�CbKoJ��cC!�o��:���[�<qVØuB|��V. �0s"�*`�r�<��ʗ�,�c�䐟bԼ�0Ŋz�<���۷S�D��i%�0q��t�<����&I@�@yר{9t��n�<����eę���<0S�$`�<���M(E��k�E
9P  ��[�<�#��+<��դ�Q��D��{�<�RfX���2VL�g��]ʢϑ}�<)���f$�^�J��|�<���#6��D��Q������Zd�<A�j���;#��t��J%Ȉ]�<�t&F4=@��B���-�H\����U�<9�@p�DI�B\9�6��I\�<�5��L��=��I��g��%$%�_�<�E#��?!XH"qGB42l�@��� C�<���"�,�aOI�ZP}	$�N�<��gտ~��=@� r�i�ɆP�<�ΐ�ggvIY��
t�b��
�@���͓�TY�G�d�J���l�K����ȓ�����]d\@�JF��Lun�G{��Oo"a2�k�4�,Ɉ���$m�M�'���G�+x��Xd��{.��k�'�b���M�,88�K�F�&^S�!I�'d:�OL�p�ɲs�

K���'�2|A��Y3&pq�jH0u�N��
�'w���r�	8ޒx�F�V9aƾ4�
��� P��vC��zt����
;�ڄ3e"O��	�W>>|F�p�X%8�)A"O��2b��
N���叿X@���"O�6���P&�ȡ�Y�\c�"OZ�� N�/�lx��"Z���Ѱ%"O�8K!�۫�s��6v� ��a"O�MYWEˉ�h�H#�.�d �"O�U��t���s @�Cu$,�"O�9��#�@���aR�tbj-`�"ORHlI����f��s�e��"O��@��u��j�(R�Ba��"O��P�`�B���+��_�Rn�[��)�S⓶O�@lB��Úx�݈�cƎFی��hOQ>�1��Wo<|�����tXRh�$�7?��ᓿ)�h@cC,Y� �bj�:I`C�I4����R�D��I�Y.G�B�ɉ{ڜ��	@�%��%*u�֓HPC�Ɏ3�=BkM�O��E`�e�t	B��+(d�����h��9FaR4�C�I�\j���҅ɄDg^`��Q;<�C�ɝS�F��\<`A%�v�
Q��B�4z6�1�N�(&�sD���UiB�	/	�M�o,a)��a%F�$V��C�	3]o51@LՇV�v���1�=�ç,��B�J���xS��*��}��|�����876���늷9R���'��\9a@jl�lz��	�"�Z�'�f�I�k�`��3�h��'�( �����=%��
�%I�~*���j,�S��?�6���u撈�3G�q��T��ʏX�<���?pq��$O�h?�ؙ0�U�<�&ݻ<�r�!3�/ny������G�<��-���𥠢H�=[f�\k�-D��h�c֌x�\Z��TOv��jPD0D�|"WJ6N��Vu�����*0D��#��Pz�
���j��n-Jk��0D��j�D�)��ƓpS9Z0� D�4�� a�yƆؼG8��sp�Ƕ�y�G��VҀy���R\ Eq�-X�y�̓
E��l��hG)P��1�E�yre�(\{h�Ο*Z�� ��&�yrH��&E]cR'I���\B�)ҝ�y¢��n�^l�u�|����	���3CI<4���spR
�M��y��ͥ^-6L�d�Y*f;����J�y�-A#�l��5bn�l�rfg���ybŅ,Nέh�ei.���
�y��~����ƙ7\������y��͹r=��RB
]��q���yr`.v�虗��l���#�"�yB�^IF���"h���ʢL��yb��2j���b%��[&f��a���y�∅I� ���1S��PсE��y2��f}��^��8�=�y�mD�~w5Y4��c����sL"�y"'_�H7�����	��`cG��y�����;���-v�)�SJ��yB��>4��$���V ���&����y���%ع�M��N�l=*���1�y��/��B%��Dܠ0gÔ��y"���m����E�ΠM�\�ZfB��y�)�!g�ȨZ4���v-��3)�.�y2����qE���" ��GZ��y��V>ϐ]��ŀ�x�"��Q�+�y
� "U(�
���hL���1�򰛖"O�!	�@,O�R)"�	�JT�Ё�"OP�[7N�6ς�x�%T�-�A"OBU����,����#�кd,t9[�"O&�p@���/�L�c�����"O�T�m�Z����xv��`Q"O���v���A�0�N�ygV��q"O��PC�9{��	�m�&k\����"ON��n$$��(C���0F��"O�\���ׯs�2����)_�Bd[�"O�0C�Z:R��sIG�y�敩w"O�}0t��43ѤHQ���?���9P"O�M9�M�<9
#)ߤOK��%"O�x�����5^����'!�6��g"O�Й5�_1GL�0�jؿn ,d"OV-���h>�]�*�@U� �"O&�zc˞CIQ $���ZC,���"Of`#b��u��R"�	p�8�K"O,����3�De��#�P�"O�Uc&��'�ēÀ޺X~X("OH� `ł0�x%�q͓k=�	�"Or9ҁL�F+��hl�[!��x�"O�!�ucө5��X��j�>m��ٶ"O^dQ�b[#f����"�.n�@��!"O*q��.܉e4b��&���'��q�"O6��(Ψ zZ�� �9����a"Oz*EFM�:��i��������CW"O��ГaD� ����L���3d"O
u����2`TJ3��'|<�"O\����XpĲ�Wc� y�\�u"OUb��īz&���$&CZ�m�"OҠk�@���e� C��
�"O�Y���#�%�V�=�.�!t�S8�y��.�����\�*�ܩ�skU�y�&�<aE�T�c�;��b3D��y� ��H�N䂀 ���0�CԾ�yR�1�~i�D�1��]��,�ybO�>z`,z�OZkp�5i�cQ/�y�GW�Db<q�7���j�aS����yr��86P�j��C�[L���B$�yK��;���b�@��(q��S�eE�y�	D:x���s�N׫l�=�`��y��O?%�e
�M�8w�=���y��Cc|@x.4�AS�H�gf]�'�D����8��M�M�Y�r���' R�J�i�	\0$�p)�>�
�'����#O�?s�E��_�ԍ;�' d�$I�)_<��C�V�X��� �'|�IB+�+H�t$J3�Ɂ"²���'�@�1�2H��؀񥖇8t�
�'Ty�L��*B��7v�̱��'Nv)ȓ�G�|l��q�)(�'V IG��9zy��HP�X����'B�(C�-P�j�aˊ!L��8��'g�}��E��'HL�"QGDHQ2�C�'8�@����r�V�� ,U:P!ze�
�'qd-�MV�&����͛H���	�'$(,Y�nU�4?����qRV�	�'�н3�����MR� ;�ѣ�'�:��Ũ�V9hTk�̄w�����'��`V�ۃu������P�k𪥳�'�D�G��A��`E�_��	�'ߴ��P/P�ؤ�����c&y�'9ީ[&f��3���(2���T������� �({ ���'M&i�TcO�K�b��V"O0m�R�t(D���n��$"O `��,�	 ��h���>����A"O(���<6�֌�pF|.(��"O��c��ɓlL��a�D4T�D�r"O�}��N�*��L��W�h��p�"O����� t`0J�`��!"Oz%��m8jŻ��)�q1p"Onٓ��Ǆ6J`-��m��Z�lMXD"O\�)NO
Ѐ�+棃�=6���"OΠ�f.�F^I��a-?/lE[d"O$<c�c�!e�p@Q�elİq"O%@Ҡ"�"��c��7�,�g"O��b�jT�b`��=�xtð"O���F��2W�D��A��9����"O<���Dܽp���� �T�u#�"Of@)׋��f�>m[W/�$U��m�S"OD��D���bLpT%�B�6�x�"O���
�W�
{0�	(P��mX�"O~�
��Y1@��Bː=���!�"O:���Q�p�������!	���"O��ˤͅ�5^tc��^�j\��u"OP�ȅG��[N��q��D�z�#�"OuZ�Ϟw#B�+ЪS�Q��� �"O&�a���]{�k
d�n�b"OyEb�0CJ��RW:��lh�"O4E�� & ����7?8�E�g"O�a�1�X E��|У-W>|2��#"O��ek�\�"<i��&u��R"Oԋ"��/`�^Q�)C}24Z�"O�brS+�I�e��7���U1D��BD]�Zd�9�T%R��`�C0D��;4�p��!׬L�ML��)$D�T��#K'oVa!����lx�&0D��Ⓞ	�W��D�6�B'G���!�@2D��N)8����K��5=�X�6�+D����Ɉ+V�@Dj���::�)��I(D���ʃ��8��,�+�����3D���E�C
[O<�	�/�77�Α
�3D�P3̏7Q��P4�J�U�5;m1D��I$�Ԍ0޲�idCӴj(�q�aj1D��JP��1AAz�H&�9C�Xa��&%D� A�)o�X�!3-��=�@ZǪ=D��1��A�w�������`�&��$:D���EB�(*v�P�]�6���8D����l�+�D<���(�o�$B�	�+��� Dàc�� [��B(8?�C�I�2̮��(�2�z����$b~B�:lm4�j2��%���cl�9^��B��5~�0)���c�+�#��X)�N:D���aLڳ2Ln����]����I9D���bi�$5FQҶL��s��AG`8D�ܠ��c�\Zvd�@��+�/6D�T� C9Q/�WOYi^�@���/D��S�@�A��t�P� ��!��B�	�F�8�6�Y%�&�Qg�͘a%�B�	+]��3�̀�HKYH%�J#�LB䉲�8ˤH�+���p�� Q�B�	�)B$�A'�w��+�j_{�JB��,B�t�A�K��움#ܠ��C�I�=g�������I�>�bB�I9���0pg�>rP��'܃�$B�ɹ�z%ە�����b�>��C�I! �݃�l�k�5r�dY+ ��C�)� ����k՘�p��"�ry8d"O�A�G �+�:أW�x�M �"O@Q!�I��i����-("O�K�f#�:���AN�:>��A"O���A�6�h�`@C*����"O��)#g�0u?-J�=?-���"O�xE ��c*U���'<�BU�r"O|�T!�������9u��e��"O�=R�lJ�Q6]��P�`�R��"O4|�qи3L�X3�.ǒ�$�1"O��� T<OX�4��Y+#�2�"O�i�d�-N��+t��$��"O��)��KX�y��.��\��"Oz� �k 3y��
H����q3�"O�p��.^<���G?!MJEJp"O���P�\=3L��rT0�pW"O�(�6n�#���FT#5�j�1""O��J���&���A���j�iE"O��R�
@�h)�dG��,<�5{�"O޹��GƳ!^*$@�C�H2��"O��p��X9g<q��z!� #�"O̥�f$�L�4p���.���#"Oʄ*��+=�]�$�.4ppj�"O�`I��ȚI82X����34"O�d���5��9�֬@!,���f"Ol�0�U�S�z� �
�j�h�"Op(�a�2}I��` ��uy"O0�q1�׃9Hlv,��`(9��"O�50�)Ъ;`ye��.jLy�"ON�0D��de��WX��� ��y�i�$nh �[��:$�@I&�y�'�;O4V �S��6�T������y2���*��H���@�2d�/F��y�d�)*��
��눩����y��wq�XK�	}�����HD��y2Ϗ�u�^���Ǟ�����#0�y���t���mیl@� �S�I��y2@�_f\���O�j�-Q��\��yң �-��IP������ O
�yR�_�n(
��󌜞5\��ܸ�y"���Z:��jtjH�c(��.�ybDR	[i �PA����"����y�A�WF����$۫S�Ƥb0͞�y��Z���9s�ޥF'�!�Ȑ�y�@#Z�,Q�W��Xb���y�\�(ĳ&M�$$*�2 �y�c$=T�����=|�D��pfC��y��B/	x��g��oP��P1@Q��yRm�}�R�Zq��bfRd��B���yB�
�l��U��.ڦS.�d�4�y�LV a��c��e����W��yoR"����S"��Y���ֺ�yb�6#����)�!k���e��yrM�?o�y tI\1I�U��֍�y�c�,b��#Q�3�B�ρ�y�aG�	+��;樝���%�C�ِ�ye87��,S3H@�׼�a"����y��3A��RqEK'kv����H4�y�c��i����-�#�����ؽ�y$R;)�&���,�
!�,�! ͖�y�WgK�Pr�j��F9�t+т�y��J�n�\ �����h㐍�y"I��_D��W���:�e�!�yr��3p�2	B���QV�Kef�&�y
� dSc�D�>��u��40�Z���"O�h5��x�8]�$�-0t�\Iu"O�-��	�욥dQ�3�|U:r"O���J�;�mR�Z�L:P�"O,щ���7<�`H��6qiE�w"O���֦��9�ТCD�*
Z؝�@"OP����Q;�X
�3AL�a"O�)÷��~��U�qA7"6���t"O:��îR#`Gp ��Ư&)���W"OX��-Ip���c��G�5	���"O���ϜV�^�Ȱ.M�O����"OrI��_z�P����g��X�!���=�.u�G�L
�!��L,i|!�D�=�H4+�B��R���H"��R�!��IK�j�c���ZG��8AF^�;�!�$�"V�=3f�I#
nP���4U�!��
Y��ytɇ�9�8)b�dm!�d�q��˶�5Sn��ڐ�x4j�'����!�e�И�lτtT�ػ�'7�(BQ㓫.�qh��\��`�
�'�`+PGʭ���m�V�Y�'��mҐ$ԋK�|A6��[ұ�
�'�}�F.3���E�IY��J
�'�(����;��B�ۙQ3h���'E�[k�4�DA�VM�NBn��'��l�Q��h7�ʐ�I"R
Y��'5�(��;9��i��E0}oHLh�'�Hd+�L2Ʉx0�Ǆ!;�Eh�'��Ա��\�̍Х�ї����	�'��Peۓd��!A���~��'�8q`�.J����jzkA��'|t��׉ȍ#�]J���3�԰�'O4��ǐ�^0��FL�b�̤Z�'���j��U#``�	p��X�\�j�'�veȒ/ĩhĐ"�Q�>�f�
�'u�U���%'�bi%��=.���'��0�g��h p�!-�0h#�'!�P[���_#�8�v�P!+���K�'�d���ݑ�I�����%F%��'ؾ3�K �2HB-^W��9�'��E;P�7/�`I@-ЃN����
�'^RIzBO�8EY����`����
�'d�y#�'�cG���/7��x�� [��cf^�m�t��Q^�+�"}��&Ŝ5�6��3�\,���ʋ@�F���e ���됮\�Q�%�, X��>��h�qc
;��di��P !�2$�ȓ3��I��[w�y�*ޖӜ��/�`dh�|���pc�_J�:d��7�����O�����v���B�����e	9,A䱈2����u��[�.!B�kP��:ă���,�^ͅ�c��[� X�J"�l˄bέ�T�ȓB����o�g�2Y�Ceϥ$���ȓ7q&�A]L���Y-2&b@�r1D��Cp��Z��Z��ØV�2xRp�;D����ҍR�MsCL*Hk�+<D�|
2.�)[ܒ8
�a��Dm����M/D��W�K��+�cJI�$S�2D���@CD� 1�"hF�SwV�� �&D��`W�Z�X�R�#CAZ敩J$D�|���S ������M�Ԉ)�զ&D� A��1�,�K�(M'=Ѥ��b(D��QR�84�P�'Xnל��U�%D�� \	1�h�� �zU�c��2����p*O��!shߟB^�iC �7�l��'��R��[��1��mݵC��5	�'�0� W�I<r�R�z'�1>މ9�'�pq��I�!P�=���  �`��'�>M�&a�ZO�	�&�
�'Q��#�܄=���ha�h&�#
�'�Th�ү��<܈�ph#�7"O�	���ޫ	�&,�G��"^�+4"O��kF*��X�))Ď ���F"O���A�'9R�cB�F�1����"O�HQ��?>�����J�Y:�"O��R�ɳf=����BI-Ѱ"O
	�E	A��>|��+̦X,,
�"O9g��G���"*�.=��	�6"O*R�*�.!U9��&��<|�X*%"O�R�����j�N�"Co��v"O��"���J�r�P��%q:�h�"O�<QWõ[��P�D�'i9М"�"O\��� <%>�a�ǁC�$��w"O�,BE�GVp�K�G�r�pZ'"Oj KDD�=��u��C�G�~5�v"O:�)`͹S� ��Rh�"��U"O@eh��R�N\��Ӗ�v��5A�"O���b��w
13C��1���ȇ"Ox}0� ���c�գY�\|��"Oĺ��Q�J'Z<9�l� }2�s�"OHh0�E�P[T��@�t���"OæNX*�^@Q�-is:	�u"O�`�p���M�v��k�(Hg���
�'�8�����$40�=+���&3L ��'\���)U���y�\l�'L����F�8�k��D%��
�'o���Ĩ� R"�x��
C��@�	�'h�#d�3(�ʹ4�Xc�X�'�*(:7IE�Cb���6K]�U�p�C�'��p,	!!��e$­Tܭ��'zx��+`R�ӳ��1!�)��'��]a @�N&�X��=p��l��'�LĚWe	�5��c��ʞiJp$�
�'D��)�o��$D�,Fe�i��()	�'4�e�t�k�Ћ�K^Y 98�'����fɯ`�6(��R1]_�|h�'a�� �˲&���0�/C-Z ���'�~����R,҈��D�R�  �
�'7:�j�Ι-�tY�F�z�uh
�'�^��t܂9<�H��@�
�V�
�'�)R��6JZiz�U�U�"�0	�'\��Y��8�V���.��c�����'��Xq���	pG�#X;g�07"O���$Q�p7�=�E�����"O�	�&������V�\���"Oإ*���0�U��!� %"O>$�F�ޘ|C�9�J��1`�"O�l &�+z\��7*�0<���!E"OvQ	qZ �!�ɘ7�`�@"O�P�`�+i½[p&�b��Qp"O���0��do��0�
XJ�Ce"OV��97��ӄ/L��$�[@"O>t�6�T;$0qkG�f�#d�Jx�<���y��-P�a�?�9tN�g�< C�O<�r�B��*�ʤ�FVc�<�g�͞#!t�"V��\�P�X�\a�<�RX�I!�ä*�r�3P�s�<� ��r�a��0lL`�m�O�T��"O�Y��w�z|��+�:�Ł�"O�	���<�h���j�$6��ݒ�"OfH�,܋oo��yW��5&& hh"O�����$B��J��Όl
��A"OT�B�i�G�-�����L����"OJ`�CƣM��� �x��A	"OT��튣@^����J;	 *�1"O0�X��5$�������mNA�'"O�E��f��{�lp����=(5"O6�B�#'�Y����4{�\���"O�I�p�Z�D��]�%.Ef���KB"Oh�$dڅJaE���r(K�"O���CM<�AS�����i3�"OU
�D��~v�r䮙"d���!�"O�t����B�d\ C���lx�"O�5�e$.�eh�ϟ�x|�	�"OɃ������A��	��"O�T�s�Z8="8�Jc�їX�V$�q"O����\2��Ɂ��+Q���p��-D�xᵮS�!���T���Ń D��҇�X�ʉ�GG=�\��B?D��@�\�?����f�'�x4!�<D���w!��J��fL���3=�C�	]i�-[��K+C(�is*�q|B�I��h2f��9h�J)Zq���k�$C�	 3�ˡŋ�}�j%�U��"O������&/�d��_�4�N��!"O���E�+��ĲT�+��*�"O��A���1j^Zma���4����"O��k�ED0V����Пf�HEx�"O�pv遤B,��~�F��"O����F�D)I��A�+�DL{�"O
;"# D`ҵ�Fd�ŹE"O��#��ʺ>�|�{�b@B�nqx�"O0y�`f��V�,�9B�] u����"O,d�"倂6�>��/G�M�Y�"O�I��S }�����PO�ذ8�"Oސ*��>|m�}�f�Q�4��Q��"O椢�^J@�i�

]�zU��"Oj	3@Q�*]�i
�	�H�|��"O&�8F��l"��C�)?m��0 "O��B56�e�Ite�ܒT"O��9w��W�L��N`�`C�"O8�$��R�
Pm�:B"O��Pm�b�"�����nƄ��"O2��D�*`N�I�����"O6}�EF�	@�W�P���!�"O�åŖ�1��]2$��N'V��T"O ��~���f��b5��"O�Թd	�	����tKњI*���"Oj��q΁%��2 �vF���"O�e�%�Ů�����L��u<��z6"O8�b��H�\Ũ�lS3(M�"O�����>ֽQ��V4[$�8h5"O♪c���B�dh��;Jq[�"O$̘�� #2��x�K������"O81�b		� ��1ZFI9%�643�"Oբ����~m�$o�)����"O�fHͤ-�ФR� !!{: /�!�$�itH��,G�B�k"���k�!��ϤS�+	Ad�J {��8~�B��ȓv����X���!,EV�܄�2�,�p%k�2
�n`j2KJ�x�Ą�S�? �x��j�;A��+Ũ�LK40�7"O`���-�o�v��h@�~B��@3"Oȫ5�ܘjy�@c�՗?=L�"Oh���M� �L�9r)��	+:"O�s��:m�� 	�8�E)�"O*yp0��;�<-ɃBD 6��@�"O>��D�ڻS�^�QcC�qfb�J�"O���̧6F�X� �.�E3�"O�|�Do�7D7���e�[��c4"O�O�%^�%�� ��0%"O�XT�U�,�����-�m�V(ڲ"O>��$�&g`}�E�P�6�ڽ�'"OFE
!@TV��0�M'P�����"O�9t�"r�U���+|��hZ2"Or(�Q��".'�������3"O��S.CWX�ѱ,طD��)Qp"O��0�/�7k�	 �lN������"O�XJQ��%7����H�V~5��"O @�g���F�&�*Y:89 �� "Od袷�L}�(��(��;���"O��J�|��:�B���rv"O����ו@�*��ɋ	�6���"O�8apĞ ���Ke�ƅit�Z "O��a�h�`��ꍨKt�۰"O>|�����n��̋ �|��"O�ݨ��B�9�s*S +Pݲ�"O` ��`��q~5q���!t�l�U"O�EPj��0"�@�ZM��"O0�4E����r�\;aF b"O��%TsE����D�OG���"O.!H���;=A}ذ�� v0�l��"OV��
T'���(�_�:)|��"O���Ē#6\��P!M�)�'"OH�{�/(YL����@�
O��"O&�X4��P�<tiS��A
���4"O��I'��.�4�v�U�p�"O ���`�lk���1��v�[�"O�,����`G�<SuG�> �j�"O2�cv&$-��I�T�tLY"OJ�@Jf�h��r)QZ��,�"O�h�ꖂFtS&�޸�z���"OP���І`���c܆j (��"O�u���n�b��g���B�"O�e�B�մf@(��7����F"O
q�A6�������^RvE��"Or�"tE�6	�+K�:|̺�"O��+a�	d��rC��+%��[�"O9����/��g�Q:IĒ��"OX�`�4Jn���!2�d�Bc"O���0B4i��Y�/�X�b,G"O���ο/���HZ�l��"OnM�B�K#�.ac!G�$Q?^��"OB��$D�@T�W��7��q�"OvYY
=�� 'LܠwB�"V"O2�Jdɕ(����bh��P_r���"O>�1wiڿ#�)���!bLƠ�w"O�As��ë/�}�񨖚%5���"O�Чa/uZ,$��̛{�Fu�"O�E ���9c2�k@"iE�0i�"O2E��H�薕�!hLe����P"O���EL��S�$��C�Ux��x0"O��đ7����5ʒrt"}�"O�����f�vL{�$�=;^��@D"O&|��MY)�(�zQcF�Pt��"O� ��y׎$ �X����1���6"OB��檃6s��� U!N+.;"O��b��� �;�&�-)����"O�]���J�M,���;7�����"O��!�L�m��HVi^�K����"O���e@�c���sH��z��h"O�8�藮l�`�qwf7��Y"O����F�	�b��:pxI�"O� j��"\V�`-Đ*�`%"O,�<,��m��O��*�F��0KH\�<�D��l{6�떒o�NłAN�Y�<�$�S�y�
�8�ń<GB�KvdX�<��$֤C uai�D�YbA��R�<a䣓�W/ڴГh^�xPZ���M�<Q��9,�1L�Q��:�Ur�<��*`.���0�DB,����XH�<����=%�8C�A.y��QA�C�<��jN�oK>�l®6e�� f�A�<qfG�X�T�B���0K��kF�b�<��[<{��B���u�@�4��Y�<�k�9|D�E��x򸨂Bi�^�<���	�6U �Μ�hBpN�\�<Q%H
W���SA挎>1v���B�<q����V���1���>⨨�%&�A�<a� U>X��$�g��,a�IA�<)�T8S�tę`[,�L�(m�D�<	�� �adI�d� Tx�b+@�<�b�¥5�ڌJg��?�~�����z�<�����BC�5r���'%� "��Nu�<YB���c 3�"��[L�s��o�<qկ8O�F� a�R�@��7Ȉo�<AU�H��fA�p@[ _���э�m�<Y!*�uo&a$EN���Xp�0D�#�H]�h���²�f����5�,D�ܒ֧5r��L�dA\�;��p0�C,D��#���aI2�U�!�zX�B�(D�,2��#G�,	2G&Y�R��E��i%D�4�[?�lPi`-a�l��"D������ W��y��존.D��XTƇ�}�H�H�"P$a�4��+,D��B���)�v%��Nn���+#o(D��A�.'��)�`�gK�0c�`9D���;\�~M§��\OB4"�7D�����w���'ZE��)��6D�@*(@l�6���W��%���3D�r�k�U����I��]�J1� +0D��Ki�/1��4^�[1^<"W.,D��(RC��9�*��ƩZk�x�AE<D���DJ/X��L�RpZd�u;D���K8�F�X�lU�\���;D�T#�	,N�9#SN,>,���-D��2�9H���H�� T8x=�0D�Xq^�k&0���&~�D��� D���ʫj�z����BE��?D�4�7�)�(�P�!
�'���i��"D����"����ì�0T��n"D��J�	�v�"�I���~�.��>D������%?-�������� U�`
>D��`�/\�� 9e�	�v�@�U�!D�pp�A¨*�-�J��	3�(��2D���ӡ:! ����DFX�A��2D�0��B"�5��%�g����0D�8���P�����E�\�
Ov���,D�d:���!�<���\kAJ(D�� ��j�m�r���1�"ޮ��e�"O�Y��Ѱu~L�vB�Gl���G"O哧˺nˢ�D�D¾�z�"O���îpZP n����zd"OV�+� ߡRG,pq�l��8�2r"O�h�`�-L. �V�b������v�<�rb	߼=i�f���t���ŗv�<��֣P*�혧�\!<5$ԙ�	U}�<A3�	u2z ���9ɖ�11�B�<��퓞,R��I$Ƃ�v<M9��{�<a��̞^w!�p�#���6�N�<q�L� U� �:�-����8у�J�<)�g��?m>��VC#\��lP�_k�<�hGRa�����5P�]0�h�<�`CT�	 �\��`N�c"��bBc�<I@����	�̛�`����Cg�<	ыB�Q�����@�ܝ�w�XJ�<�C�ɠ �bx�@�c�<k h`�<AgU�n� �22a�Ld �PÂ_�<9Z#�<�1�#N� ᆉZ��f�<�3N�o�2�	�ǐ'.�ȵ��_�<Y�I�?��iG�uV��aV@`�<AbJ+�dl��N�o&�`��EV�<���G	Pl� 1�R�)%p����U�<����� !FӏJ^1��/�H�<qwj ����6#ևD� ��%z�<!!�� s��J��L�R �Y��oIx�<���̮S�ƙ2��<J�t���t�<���A-lx"��θfp��9�*u�<���U"\9�dP�AF~ʀA+Qf�<T"�3n��)�F�v�&PA�N�<��hH;b� ���K�o-�1����u�<���['<�����!m=����W�<���Z�/��|��I�V�eY���x�<�QN	1.@�L0W��	\5MY�c�M�<�3���X����,ݝy��YA��_J�<��Ԓn
,ʳ�(T�0%�p�<!!L15ލ�����	fY�M_o�<�2G4C�pZ�'�$U�(�7�Lh�<Y�ܗ'�����t\y��c�<��(�4"^�s����MP2i�c�<���86ٺ�1�JY<�\U@�u�<Ap��,�L}j��Ț��$DEL�<!G�G/_���F`�LU =d��N�<�A4q�����J+V��� �]d�<iP�l2x�q�C_�$m��͌_�<!�IL�U���f�pa���[�<��P�C*$q#eo�l	4!zE�KO�<����N�Ȫ���*H86@�ǫYO�<�"��,1�a���I=h� ���C�<�#dX4J��Lр��xN��ؠ,�C�<Y$��)���`��m�rL2�iQU�<�BD�(,�X��G�K��YՠBP�<�s�%EǤ}����q=�P���a�<!ԃ�.�v@`�-���i"�\�<	�+ɢ<���Rg��	��Y�OXt�<���N��J���f�q�Ze�<��Ø�UH$��.��A
Yj�<�A���lɔl�d#��9�𘙠�[�<�S��oD��Q�>($����Q�<�t�Гs�hY@��ڔ�l�d�<���������Rh��8�q`Be�<aѭ�� �t5 1m���)uy�<9$@A�J�[lܮ.���Ώs�<�  Y �WN�3 �+H�P�"O�l��ȗ6*s�)��6)�$�"OHP4	��Bj@�]�^
�1"OF�R�Ǆ% �{OӃ:���!"ON�����Q1�`8!�x�+pI���yR��	ͬ��G�Üv���EW�y��0.U��6�	tQZ��D_��yRo�e�V����3`T<���M6�y"���rʣ��)-����e^��yҁعm�XK&)~`hم�T'�y⩎�>��	��6�:����y2i�KX����/�$	���+�b	 �y2�THEr"j��y��Q��C��y2�Կs���C��@{���O���y���	8��1��[@]��qF��yR@S�u,dx(����D�tUy4l�0�y�a�"��@�ԏ����# ��y��P�,<���vb�|�C�:�yrA7$�I�큓醬k�-�y�`�$Y��y���5`���F��y��#~�ʵ�S���!ɔ�	�/�v�<�D��K\���
xt(4��_s�<	����r``eq�"�	k:���̈S�<�2Ec��qm�2"���N>!�DR�Ֆ ��^ �\ʷ�R��!��*�40:�'ڍt���yL�W�!�P�802U���L�)�rXd�ю�!���yƦyHQkH�\�>��i�9�!�ͺ|�F��t	���@��(��C�!�d�-�]��d�'�P�btIĻG�!�D-�|(#�E?l`�b �!��7��R#��?c`�� A�?�!�h�lѻp�ژ&D|}y2OZ��!�dM�d���(�H���T�!��D ��m0Ԯ�(sj�7LI�!���vh^(�2�ɒo��*���
2�!��zk|Mz]>~iX�y�<V�!�_�V�)듪�0� �S��8Mw!��O <���0�f�0�b��=g!�$ǲ7	����Dk颩K��cb"O����HІ.��� ��n�"���"OΤ�OI�����b]�Z�j%��"O��a�I[t�� H��ʾ7�ѐ"O���#� Z��uX��E '
��y"O`��.�1k�)��Ud�$�d"O��92�O�JF�p'$��Z�Hҁ"OT�@�����Qr	I� (P"O�9q&�0*�X���"p_�4[�"O�1茻( :�dXL홢"O��Q�¨&ê塤bڠ
�)��"O�`���8]|U��(��k8�Ez�"O�i�V$��!فGү '�Ibv"O$5@�%�*K�!�'�V%#�` g"ON]�G�].X
�x�̡��c�"O��E_�mg�`A��I��lS�"O�P�"�Vf�cV�U�%��"O|��p�u%�ڐu��9���O�<�paXc�"}���0��\���s�<����2����ꊬO~�Dhx�<�`��/V�8�
�B�,����Y�<A6�͙RԚ q�K<���E�X�<9�hO$������,6��B#�Q�<��'��j�Ss�C'?�,Q�e�@K�<��-�~�2C7C��=Z��9��\�<� |L 5bE��,���EV.u�<��"O"1a�c+,�hSg%ɽ8�9
"O����g��ܡxA��PV8"O@!�P	��V��(SeE!-V@�F"O�)ru�-Q�̽[F$F:�ڑA'"O�ٔ��l��s��?��(yD"O B��s�HM+��[�=��Y1"O�U��h�ua��� +�vD� "O�D�uL�1&(� ��/sXV��6"O��
���;�z�$)�8H����"O�\��o�^�2QE�� �!�"O@�����NάT
��y}r@�s"O�Y��E�	s3T����ח)�ڕ2"Oڥ[��P�|�Uم��.��<"R"O���#c�5�J����H�1X  "Ov�����1*|(p��x��h�"O��BU.DR1���4 ��>� "O~,����5u�xH��)-�,Aj�"OZ,��� ��x�E���`�HQz�"O��S�f�n�(��!ʙ:,��aY�"Od�0g ��g�L��W]�L�C�"O����`B�h�*�����Ye�p�g"O.�i��3c�T4�#( �_K�;�"O�)��HD:~��q���"h3� �C"O4�����]S�x@$#K�n��T"O�yq�u�����4\�l""O�Bf�S8<��Ht��b��L�Q"O,<�6��'$�*�/S)����"Op��6(O)]l�c�6��;F"OX�a�CF�Q��ߊ��(�"ODa�B����T�z�.ˤ;���B"O\��b��4���`�M�^gN̋%"O��;EğR�t(#M�rE\`h�"Ovԩ,P	ciRX�T+юl�6e��"Ot�'�
>�q�E��7@��2u"O`���	Y�v	�$�ώ����"O4�[����:�*���H�#f�^X�"OؑX�#G�W�Q�D�q�z	��"OL�E��d�� Y V�Eִ$��"Otp�EA�  \u٦� %N1�,-$!�D��h��ѹ ��T�
�aϦ3!���z��X�'�Gxht�`��4�!�D�� ���8Z�u\ö�K>%p!��#�h@�D�� _���QaJ�pR!�D,x����ts��	VE�yG!��%v���Ic�%:k�DR��ݻjA!�D�|r����^0}^�(c����!�d��{)x<��
�B��ʁ�P%�!�$�W�@�JV��*˞Ȁ�ĂIf!��߿si01���: ��S2�2uf!�D!g�J�����D���0e!�N#D��u�PA	lc:��'�$(U!�$��n�Q"�&M ͩ�A�!U!��͛�mMh�m>��	S��4[!��()!BC�:t�D&E
xS!򤙥�Е����+l�Ƽ����e�!����x<P'�z�(�l��!���c���lҥf:������!��7y��:@�%  qFc�!m�!�D�f`5�� oR�@P�fo!��	�K�>YPTKJ�2$[��ߛ�!�Ěb�2a'�֛3�d8+��<7u!��u��	U#�\�b���H�;h�!��+!:��S㐚W�j��Bg�%WX!�� j�R�ǘ!�dP2f�h>�S!"O~H��Kվf?F=q�N �
zF��"O�}�Fa�����1N%vJ![�"O��Б
RAh|��,љ�� 0"O�����H����Ʈ�Y]:͂`"O���n� [���sE�ғD�$�3�"O��
�J� `Yf8�� $i�͡2"O�y���]3����&[q�@R�"OV����$?hF�3�Tu�@�w"O����O�p�%��9f�"�"O��8W�.{ʐ�xӪ_�d1d��"Op=[T��!ud0
0��/Dr%�"O�M�#g�i:��Bև��q08`v"O(}�
Q�R����`MҺ~搳�"O������20�&��P��3x���q�"O�ݻ�� 3Mɐz�v *3��!��Q$S]����Z�����4~!�ĉI�7NX=h�&ޏ�!�$�^���qB�����#�%h!򤂺d>"���D/T�rf���[�!��4gB����Xi��f��h2!��A�y��P�B��f��a�1�!�^B0��n��@�a�G�v.!��
�PS�J�W��0 �<`#!�$�Zt����� w�|c&�Y l!�DߜS�H��ܧsZ�ѳ�`A�W!�D�Ws���hʹ@�,P`�P�S�!���l,���,�XE�G�hT!�$U�bhl�E�Z?F�3��oJ!�^�<�qbe&�vtz<B��-!򄁃�H��D�b�(&l�".!�d��[_���D�ßKH�4j�K�&M !��3�4�) �ז;&X� �O
!�$ޙU��C�ل���´��r�!�ā�t��6/��r�p	�%+H�q�!�dT$����$��(q���>\!�]W�}��G�2���	�Z"q>!��C+Z�a�FZ$$��`A��7f+!��=`C� ��B�	�$�W�U�H�!�CiO�Z����-w�I���x!��O�v(X6)Ȝd`��!� |!��V��"aP@O�QJn��SJY18�!�ĝ:U�
��ck�s̼\��H��!�$�E�L�Pt^+"x��afP>i!�$C�|��%a�a7V��ѹ���V!��?�^����	ܼe��ʾU�!�Dí�IKf�Ǆ>8�<�&�8�!��يG!�ћ5E���d�a��T.x}!��O�����ͪY�D���X%?m!�E,bԹ��Bн./zܲ!k�+W?!���w�"!�P���!����K�*�!�W!)�`�1��R$�U���R�'�(���O���{��F�v�L��'�܅J��ӆ[5ґDw((��	�'��K��±kJ>x b��n��}
�'b*�@��x�,�
�틩lL�y 	�'�j[P�I9��r�ꔛ]�ԡ�'�hY���d���8@�¢6.�(	�'�p聢�� u p���V��z�s�'���	���h��@����+Y�u!�'�u�P��#c�Qrj�[��UJ�'j��y�˔�5��bO)YX�| �'���)a�է.e�鐄�w�N1�g"OF�z GŬ�.2�h'>�(i"O� @mҴf-n� E�B�ЄxA"O ��1���_w^ej5�O��u"O����A ��s���#�)1"O�Y� �K����I��D�s"O�)�A�-��P�,@a~~q�7"O64+*26����L3XY�k�"O�T�� �ƽ[�Z�Q�nP{D"O��i�!|�x�oQ�Dd��"O`����6�T����!:1NȲ�"O:�b�a\�!�����,�w����"Of�h�C�1L.��t��"O�x��f̳�8DS�m.,�t��"O�mP�O�"���5l�lr� ��"O��cr�G#Lԛ��܍bI��PP"O�0bG��5w��ĘS�U
z����"O�yt�B)8f�A���Dp��h@"O^uc6\���q��3}��<(3"O���&L��H��6��w��A"O|yQ���'X���%靅��)yC"O���)P��Dh�n��C�"O��ʔ���ur<yR倆=��x��"O��P�b�s��c�PyT� �"O����.$쎭��M��t��@g"O���N�v�Nɡ�c6��A"Oz�!T�����EL��|`p"O�-��wTf�1��S��〘�y�͕�b/�	A���@�����y"��>9���j�09��@���T��y��ĮV�� H�6ߒ�03�ǣ�y��������@�3[��S�Ǆ��y��c&�e�AE_/1ݤ`
�y�����a�c�H. �B�:�+���y� ��cބ5b�CF���yRO��`h����<���G���ybCC��%�fJ��T������y"]�t^U��җQ����yBJ�q *u�VO��F� ���yҌݸ����v�'n.Q3��ك�y���{V!Ehc�q��֞�yR�qr��SS �6f?6����/�y̀?��ѣ��^�hR&�%�y�P<L�k�߽h��!�ř�yR�Ǻ5���igN�7z��r� ��yr��6T��ը�y:�J]!�yB��\t0#��E���bQC�&�y"�6u��0�˚-n����ʸ�y"�Z��ر��X�h�d���I��y�:8�:���/PxX�=c��A �y�W8��� Ŷ����c.ח�yb��x8a���ڂ���*ȉ�y��"^�tQ� V/�dqq`��'�yr㝰&�`�G�9u�By�Fڏ�y���<N9V�r�nكhxqw�1�y(J.\��ist'݀n���J�ޯ�y�6R�dj�N��#cE��y�o��%f8x�JK�6�S���(�y`��QS�$����J IfHЋ�y�gX�kl��	�n�\c���<�y�Bҙ?p�%3 ��l~~(3���y"eגu��jW��6km�9�E��yB�>�b������t[��9�yBDݤ:楩�mA27�2�h���y�ؽ����V 4�4��)����'�ўb>1���9@M퉱�K�Tt�S��;D�� ~aHrb0^W�$�Pg�<ֶ,y`*On��'/�'vQ����W]�|���'�D�91N��4Pxd+�
Q)nl"�}�',.�)�ǋݺ��t��E��A�'5b@;��O��� �cP9�d�'�~e�5M�~�J�:j��D���1���ɪ5��Z�'��T2� ؐO΃/+�7��<�R�-|Or���� +�h�
ϭe4�Rv"Oj��qHW�Ƅ�X�Ɍ#eh���"O~ؚ&+O9����'V1)w�|��I`�O��� AD�V��x��`A�5qf��ȓ ��j�'�v�
u/2r��A�ȓV;�M�k�"�R0	�93�`��'�ў�|�ɂ
��H+���$7�T�1' f�<Q�
�0V�.]�Bw�m9r��G�<�sIY�t��<� �ZX�`5Q!gZJ�<��j�=+E�4u)��� r!Jy��'���r��wBZM㝮e�H��Ó�hO����ń7?�B�)��/W��I�"O�u+ֆ\�`�=��۪G�(	�G"O�E���9JV�ix�g��Bp<Y�"Ox�Ja��	x�&��*J�h��"O�j�iS)3�-q���+!����a�cH<��*�U��!����?g]�Y8C�EX���O��{��..7��9f	_8bk�}BO���Q{(2��W+'%��L��ޘ-��	Vx�@h�큮# n�Z���f<n����6D����^8z#(Y��@��$6B6?I��d#�I���D�$ ���cD%Z�`C�ɴ���k�\�Umd���"S�LC�I�0]�4���@�����o��km4��p?��D�5u���!@��t����w���'u�PY1�E�Vs��@�I���ȁ�'�p$���1q��0!�B��5���1��d�ƈ�����G@�qĺq[���3
y@�|2�)�'�T��ű�>d��mu_���&��$a��S=M�탄/\�Z t,��J���C䉝!Ldև��K�>��󨜸f4\�'�ў@�>�-�l��a"�� �r�n�_�<��I�;"��H�Q�&<m�`�Q�<����F�^�(���'Nr���q�'ў�' 86`a7YrGz�{ŀ���y��N�@�>�
ְ�鷣��2�,���Ζ�����ȓ>7��Q���j�����Y�L�ȓE�������MH�n[_Ά}���<,��hƒG:�p���� v�q��<ڪ�Cf���,���gF�
4ą�"j��"�ÔS�Pta��^�� ��ȓy�x�9"�1((��Ȱ�p��a��oLp(xS _(+����fb
8�u��"}b���f_�� R<"��`�5���O+�	=�0?�3�=o:	BP�5,14��I~�'&�O�X�"���~ND3m_�?~j0Y��'?��3Q$��Č�,KWn�ɢ��7B2vB�	%��HF���U�B}��`� O��p���OD�(N2E�gt����;Oz��w#�2gs��Z�c�o����"O���W.���N��㞄J��S"O����r<X�ٔ�ٵ|�|����A�O7j)#��:x��'׶o*�й�'(04
�=,�&��P�	b�tm��'���aS�k�<���	\;EQ���'.���ո����bfB;P�:���'�6�����Gu@���*��O%������ *��dfƭ'vh�#5E�.��B"O��Q` W	9���W Nʀ�X��	Hx�x��$�q43��&�X�c3e#D�,��QaJ�Te�c,�����hO?����2��i�R��
3��9XqI3va{���y���q�K���p���JN�'�|�o��18���Cže8���2��;�ybbӵ�����N'\��L��o��y���D3�0f��|&�TgH6�y����� �lD��q�J��y�ė|Gt��/�2VU�����Ƙ�yB�¡=�=�P�\+@K��`3"��ybc�R4V�A�ԏ?'v�㉁���'a{OO�My����kM1e�A×���'��	r�O��ذ��η?�JAB���H��=��'�X8r�ӢiH@�H��X�qH�'�4-Q&��)'���
�?�4��'��Ё2�S%[K@���N9���' �%�e�oJ�=�`/�z9�7�Y���)�f<j�#"�rȴ1r�%H�!�$�&��]�rJ�#X��I{���h!��Ft�`����H̽0�`> �!�U>a�Ri���}^2�SeO�s��z��d�������L# 	{���6z�!�d3\�buPԩL-����'Iy��xD{ʟ��cv`��Y|�哠�&���5��$$�S�O��<3 n[5�by��GL\(�'eVLp�a�6!�p��!�#����{��'��]���K�H�
�/(5m���'��B��0{0�`WĂ�^-�M	�y��z�`�DO�*~z
�Ĝ�p=��}�bت#>�XC����{  ����X �y�	��4�.0;a���n#���D�/�����:�)��I"�Pk�G����a�*Jx�Iæ�ϓ��S�OyRhxV��~c���Ӡ�B)��1	�'�Z��J�k	�9@�	Z4��@k�';VśǍ�.��	d'�V}��H�'a��!j0E���W7E��`�d���yB�\
K��~�;KZ��p<Q���l��KŨ�;r5��f�K^a{��Dۦ��aK�28��PFkQ�A	�O��IP��~��3l��M�ҥ�k۶8�С��'�#=���D�E?6�@Z��WZ��`"O|K��,��� ���*Bo~�*�f*�S��y�JW�8g�p�I��F���D7�yB���#� aC��R�rA�B����/�S�O,�|z焐�s�a4�Ѯ2�`l����~��4c(���O M.����2mcqO��=%>�9$�_�g]�����B�`q�:�O��v�(x��ӉK��|X�Ο9�XM���M#�� m��L��>Dp����l~��i��"|Z��H2>���P��W����ħ�i�<�U��)��A��S�>@�ኂh؞,�=��.\�'ylx�2�D�L=�uHA+�f�'�?!����H|J��(jL��"���c�<)�>L�>��DQL�@�@�J8��Fz�O[�F����Ģ'�"H��͘��y��ZC�A��� &���r&)5�M��'�:�w�ݾU�Q[�N�\S`�
�'��<�aI�f��D�s��2A���
�'F����&l�T(���ĨA���(O�$�)ʧo vm��	Vk[��S`�@�wZ2���Dx�UƄ�j�{�I��6Z�чȓЪ��τlм)�"���n)��S�? ���"y�Tiˈ*?yʙ"4"OJ�TF�m`��I�#`�|��"O<�q6��J�X�GJ `O�@0"O�����Q|is�<^���A"O��)�*s���x�ͯV^nXa�"O8�:��Z�e9a �gSޥ��"O�Ճ� /i���ܺ[s�u�v"O��+㩞,9�x���K�pI���5"O� �q��Be�+�?2$عR"Oҝ `e�'*p`H@�_�.���S"O�4��l��Ka���k�/y�N ��"O`E`'O�#L�8�P��ʷ���#"O�-ʤD����Yj���:L�<��"O쑈X�L�>��j[r�@�S"Ozx�e̛���o�-���""O�aJu�3a�nU���9~E��"O���3
��i� ����٣L(¨�d"O<e�DW�B�FEKd�7/<��E"OdQ�J�!��E2Em¸;�0}+�"O0�SfKҦFP*�Tk
���X"Oe˱B�z��aP�	��|P�"ObHQ���?,�Dq�+":Dȗ"O� �� e��;�_7O/��5"O0Ma���&�b<sw)��L(�E	"O�P���ðtEr(:���YF�̨1"O<(!Aʙ!Y@*��dx�)׌М�y"����� 1h��!-�)�y�#@%���c��>X��1(��y���`xD�!�3�[�f�
�y�L<�aX �j8�1�ٜ�y�n���|=�Kߎ[ԣ�,
��y��"J���3�\	���3��
�ybI�]*�� E�MΜ#_hM��'�x%c�)͞�% I���1娚l�<�'a�0߾���������6�H�:�X�� mf!֟24<��Q�(Y��קVh�9���V�\��ȓ��""吇iuIVF�v����'���T�Ct�����	�輆�?�j',��+��t���{?~P��Ϻ�B���u��M�6`�9c�BͅȓU:��ǝ*���b��2>� e�ȓ;҂<�t��I�7�,m�	�ȓQ;$=�t��(�>���aTF�ȓ��0%�χC\��iql$IU����q<�0`�A$��<�rC
�<��u�ȓM���(��?5����C�/V�����6�ԣz��,f��-a>4��9�z��w�C��5馎ܗMl�\�ȓN��up��	�I2&� ��ר�,��ȓ~zx�+X-{X��"�^*Sd	��,������GD ���f���V�<�T�Ņx�`�F�|L�k�B�d�<��nXDo���P��76M�H���k�<��@�0Gt�`�AG��U�u&�a�<9�2|����S@��M
�+��X�<�����;X�
��.>�l����l�<�U(X�!߼͡�IMn4�qE��k�<���Y!.�!�����9��_f�<Y�fÁ4��&��!t�zM�6� b�<�W���@�"i����6��Y���JA�<ه慶iS�0��I0��C�Jd�<y'�ƺ~BpsT(�	�� Cb�z�<)�(T>X{�L�������Gv�<�3��,�*�ۋ֠��$z�<� ��x�IƝcQ�)�.�L��`�#"O��x�#T*0K�yhB�Z(�"O�)�kW�H�,X�E��3��HE"O`h��w#�T��+�1f�Z ��"O2ػ�)("�$ajπ_�ޙ��"O�`a�����IS���t�D�0"O��صM�9/MJ z��I\��y�"O����?��m�TbI�|5��"O�(h��A?D )�a��'����"O=8�!a�]�[�@�p1��5EM!��CP�z�iҦ0{�e���ͦ$!�$J*�@k�΍ W-f�D�D!�D�2%��PA��(|����nׇ;!�$ϵ`�>\�a�%(g���U6r:!�D׊_\�·��6kAb`W�`�!��֙u	n�*�K\Mv8��v.ݨQ�!�$�;�j�+�EߏNB.%�E+Zn�!�$�iT�5�6��8�����v�!�$J����b����i� �Ub��B���<�xA��28
�q�Ua(iH`B�ɕq �Ő��B+w?���aH�;�$B��"|XHM��bX=>��5����2Z�6B�
@�< ���#	���@<B�9d���g��SL>��D+ e�C�ɩoz,d{���DLJ0��ީ4~�C�	?kDX�B�̎S�@��O��~��C�əw�Ɖ2a畜(��t�$�C�LC�	�54�TP!(�/[o��a���.v4C��'y�����&�%*VV�� fܯ
�PB�	??���F\(w $Rcڝ#��B�ɞm�"��*�If>�XR��P�B䉐my��+���H2��v��O7�C��4&Y��%*Q쑚�G�1-^dC�I�h'�� K	" !yp��vZJC�I*e��p�����w˻>TC�IZ��K4#�(7�Vub3g8c�C�ɉ0
��
@��x����J�6m�B�	���j0*Z.d2ة��E|���,ռ$�SW>�^93b�ڂC�!��X��ik��ĔB���5�!�D %6�Ҙ�r�,9�x	U�	�f�!�$BE������,q�la2�r�!���$_��嚕�K��y�W'ί!�]w�\#�E	Gh��2���F�!�Q Y��%����1��	��#@0!��L�i@2�E/Q"^���eM�5!�$ё���a����H�i� ��?y!!������'�̩R���8S�O!�W%bW��iU�F���c�"N_!���n4�)b�͖*C��H���!�DC<�$�b)	�;�b,�p/S�&�!���>r%ik���-txD{���p�<9��ڤ	���n� S��s�<�2MU9e	��;�m��.��h�<Q�"��~v��㷨��I"��2F&YB�<-�|f�W�2G՜�mG�<��Ǟ�zrɠ�A�����b`��u�<����f1����.$Y���#��n�<a�J�@	��m�.z<�����a�<)�Q�:A�	$H'$(�@iSB�t�<�ADƤi:�\�r��j�H�P'l�<��ɘ�]���� ݜ,V�� ���l�<�!F��b�}*%����@�Čk�<!���-+�cS!=� aE�b�<� H\h'�N�[܌5r���G=l]��"O��k��\(N�Рj����aI�H(g"OF����,F�0�Z�C�K����"O�})���/����E�-�&�K�"O�T{�@H)p��9�Ȏ�'����e"OV!܍��98��K�R�
Չs"O4�x�
�������fI3���1"O�pH��"~����W�J.j0�"OJ�J)�r��i�e�;�M��"OJT+�#��]	x������E6$�"O H�@аg��!��0y%���t"Or�A��V��y�VL6��;�"O�x!R�M�T�a�CP�<���	"O�k�ϑ""�1L��� ��"O�|@p��k2d�c�>t6���"O�hksD�%O���w"ѺHQ>48�"O
���G��29<�ppLV�"T2�i�"On`P��D%4%���&G�V��R!"O�@	a�I�	L�� �畷.�����"O��1��H�e�;�k̂v*H��'vr� X%Od��Z�Mʂ3�l
�'� ���!Hb��ȜNX���'Zj\hu��5�l1���G�� ��'����J,4���U`ٍ"9��a�'����߿�`��e/ԥZ�p��'Jz�k���b8�$GӦ�,h�'N�h�ǯ��5A��a���~n%p�'���r*�_�<�;��B�R �
�'z��CcJ��BA��1�>G����'z����T�kFȌb�b���L�"�'��3�A,,�����ܠuP~E�'��x:4�,hɐ��R^�c�B- �'p�b����;t��q'��U��a��'O�!�����a����A��D��'Qp9C�!J�g[�+AmB*?/	�'` -��g=#xFI�Я���`�J�'N-@uB�z�Ҍ��6M��P��'��4����&�4@�A�m��'�H��%*Z?>��-kt�ғDJ���'�1���M0�J��D1�
��'�ޱ�Ӫ%ڞ�ڷ ��.��xB�'���R��A��Q#�-��!���'��Ւ6�ۮ9{&$�f�.$����']��n��W�|13a�	�$�
|��'��A���"P�g�6c����'z���m�1s��!',��+=���
�'+�fo����V A	���N>�F@����$�U(���v�]& �
�Z�.'��~���:-7P��`�ʺ\ö0 t�O(`��1��΍4d�����Zi#���Hj-Є
6s6XG|r��+o�ZlR���D�Oذ(���T�el*R�iX8����'���� ��d��-'zwbxI��&�1�7+�a�W��"~Ұ�<3�d��N�%���Pf%���y�C�~��P��*K���piEl�!*�<���V]� �4�J)f� A��HOLt"':yy�s�?'��98
�~LnIK��K���f-W"�vP�BϬE�DH�"��l�z�(
�C��ASIJ?�f� �j��M4
HDzB  V�2����W;d�i%�~�OUt�0b�(RC�}�5�i�<ɖ�V�:�Thx�eT+#$6q�3�]�ٲG������Ťw@�K���i���"�
0&)�0B���.*��`k�'���`�LREXn���$�<"v�Pu�ȟ<I��D��K�����鉯L��P�%
�:���)Ð)�&��D�#T�e�E�����)5�TT����@�Κ��-��P�N��䐉jz]a�5�: �%�a��0#D�9��9�E��Wx��� ��B��7GNd٦#�5|v[�"OP�`��˃:l�:3��)b��̂�im�dQ @�/Sm2|y5,��X��#nZ�)4�ʗ��9k\ldZ�N�~S�C�I�q�D�$w&�8p+ĻYb�9��'� ��@�ƃ_)��"S]>�<I ,9,�x��	s�:0���kx�4��hժ����ŃD�x@�ԅ�BA�T-�
_T0X��'<��j��O���$)��4q������X���ÀQ%�֓�8�m8\d␰��\��H�$"O�YI G��JҞ�!fE���t�OF]���،0(��N��}�Ǭ�<D�m)�F��F�e��v�<ّ�5�0�[�o�=	cL	��v�	aH��'��}��F�uR|�a��&e�=��'.��3�Y�2Ӗ��J:D%T�*	�'68�k&��/�4M�!F1#�ey	�'�N��$��^0A!,1�����'f�� ����PA�*�7�@�q�'�~�qH�:����6%�v��
�'��q(�cJ)(zTP!b�opּ2	�'��h�[yH�<+�#��,
�-A�#D�T������HӈsV�� � "D�����0J�:��1O!x\T����?D�xK��4`�=svE�=>�N�R�;D�tQj�?+-2�B�H�1N�Ð/:D�����ye���I�	=�&�8D�Ȋ���-�V�� �~�!r��:D�����?�����ΛH���;`�6D��k�$S��	yq�؋K�~@c��:D���1��$B�H*@CV�b�B�d4D������?.�v"�� U�Ҝ�@0D���U%�mC(��!��]�vC��5D�P�Ҭ�6x D��8_�<=!a�3D���W`ĴZ:�8!N�7�M�.D�i���<{ΘD(0JC�"�Ɛ��M1D�$f6+ ����C�*yD��	� D���N
�z^D���(��<j��=D����ა3�$
��B�>qZ"�8D��X-E�oP-@iJ�~4Z�I;D�X�L�j�`h��gB �#�8D�L"���9�bs�\^s��A&b4D�p�(�*Dd��XGmɷY�.�[�(<D�Db�o�$^\`0y�"I���ɀ�y"g\; $���F�&k7.�W���y�HҢK4��䧇)a���2�ݵ�y���:����(�.b��3�I��y��J�ME"]�s�R�Q���WT��y�-"Y��3 É�~j�͝�yEN�vj0)Ԃ��?S��ر"��y�n-@�w�^���a� �ҷ�y�)`���I�x�X��ᅆ�y��
*��$�uH�6fZJěVi!�yBH�'gk�	r'_�޺ye��yB�Q	~����`ǳL��d���y2��$��ᓐ շ[���iTŗ�y�H����i���:X�	�k�y�nD�}?�Ђ��K��H�+���y��تp��ٱ6FJ�N4@�2�φ�y���y#q�V�Q�L	AB�6�y"�K�F?ɀ��֪e�8�s3O��yV�4<�S�ސX�A�ܤ�y"��~��!HԂl:v���E���y�ɓ�=�\X���B�X�j�����)�y"#@��D�*E�Q�BEz���g��y�+ݥieZ�cԇ��:5`�{�n���y��Q*q,��&��?b��F�σ�y
� �����F�$�r0�^Z;�p#"OFl֭(�){3(g^Y��"OPĨ�G���:fD�4	���"O�U
�7a��x���W��5("O�8���|4R����2M�0\hV"O܈{%�:*M��'J�^�Z\�1"OL9	��Ѳw�t�Iթ�5�v@`q"O�l�Dgb-Z�cC.L
T����"O4 5�X���5�̓J$aV"O��� vts#���q>��PR"O��җ'�?J��H���2���"Ov�P�L�]�X���A�M���F"O���#�t:��� MA�^�(�"Oi�� H�U$��ZV��+�:M�b"O�hs�)�;tA���5�9�N�h""O���Fl����˴�&k��Yg"Op��b��ɦ��Q
Q	I��}:�"O�)�GvɌ-c�!���11"O&i�d�;}o��k���
fs����"O�E9��GH�I��`x�K`"O���=!�p�s�E�>����A"O��[��R�U�Z�b�� "O�]+d�ݜ湸� �6[��$"O\��.�b��sl��,0�}H�"O
�d�L�o��8:fK);L�:f"O �ab�3<0���/) B���"O<�𧨒�P�4��'Ė7qL�\#"O@��cd��')B��Qa�?#����"O:y@t��4p�z%��;�S�"O�r��>AL\��&�""�Ph�3"Oʸ�%KW�r��U�r��C6"OZ��гW:
��@�,U� �"O�RDl��3�ဈ@�<�SW"O,�1�İ^�0��m�B��aB�"O\�P��_kБ�jǿ(�<1�"O�5��X��������r(�	"O
0҆�M"zJ��'M�x��"O8�ؓ�W(9Ep9)�;Q�d�0"O��,�	��L@p([�]\Jh��"O���
�8H��LE;]\��'M�E#��X�FW�,h'LR���I�'A�Lp0K�dy���i�%N�Z��' ��D Ly0u����Vg��x�'��1�͚D�2�c�A�\Z���'����.�!	��eH�CT���'N��J�]l�xp���V����'T�А(V�{LJ8�&�KC�(P�'Q��8�):&$��Q�jJ4CC����'AШ�@h]'zB~��R䄤>,���'�q!�V+!����À_�`�0u@�'Wj�aTb_*Q`�Ș��T�_A���'7��".
�} `���M$I����'��ǔ2~�`XH�O�Gp0�q�' (١�,t��e3F�RbX��'�.l���pUnЅ_$H�j���'�Șs֥ĸ���U�ݝN��%*	�'�l���'].{>	�)�6���	�'ƬT���y�I8!&��b��x	�'X�i'�\/i�>��@��t��1�'�@H���X�TmbE��k���
�'�*�R"k��*���t�ۤae��2	�'�B���)�4{�D�@j��hf��'�xQ�l�9��@�7��
�'�%��a�I�I�QW2lX	��� � �rb_��D�Y�p�E+�"O����	���
�A��ۢ"O��f�W�w�y��Z��\0�p"O6�c��
z�$-	��ϯ_���y�"O`$��$L+�0�ee�X��#w"O&Řb�åY�t1$�k#Č��"Od���$��jθ`��Ňp)��"O�P2�J��tE4H����b����"O0�SP�I�~���Q�! �)"O^] �D��{���F�#<�Tڃ"O`L1�j�6H���`. �r-�&"O�����9
$ܘ��YP "Or�NT�&��ԘiP�1�!�䐆<Z���d�)7��:�#�4j�!�ď�Z��m���0 �%�R�ۣH�!�Dޖ3L�JWMOpy[gS�7�!�Ğ�!�>Q�Ȍ6�,h�/��-�!�)pF�b-N'+�q��m 	g!��X!�H�3����g!�ė�8�:5`Ă��!xp��Zm!�^)1�m���$����vLYFX!�DL�! �Q7c1Q�B98f�wD!�DеM��ّ�̻A1��Y̘�;H!�ā*3d��ʇ�o��F]!�dA ip�f�2B<�Q$ �%�!�4��آ�CQ9$�%��E� �!�S�!|vY�0g8�����!�!�$�5@�MȔn�%�<a#��K?w�!�H�`@��E\&=�X2��5]�!�$�Gg�X#Aq$Rxڦb��i!�dF`�����Ù�e KfAL�Q!�D�����D�"<�� -P�)\!���s=I����*^a�!m��s�!��FR�!���p4yX�n�4w!�$R�A�r��`��!���6�Fi!�זD��+�jےC�f����$}r!򄄀^�b��7g]W'�2�F�i!�Đ�����S�B�*ÓC{9�|��E~�x��ɢ
t����OAWl�]�ȓ%h��W�ɠR��G�؅�M+�݉��ɮ!�<طۍ
����ȓV����hL��!�x��ȓ ��s�U�vuT�9�T�X�xنȓ~�J1A3��3\�������;m��0�ȓJ�D�&˓�i�H��s��6:~zY��'���x���F������
D�d��ȓq��U�_MnT�6Μ�_�ڽ�ȓ,���[��^:sd�{RޱF�|��ȓp�k��V�A#��k����4��c0��� �T�N�q��n[i��P�ȓz���*2�U��D��$cn�d��ȓZ�|��7��#-���� �j(��ȓ���a�4?
�X��2\@�ȓꍡA�C5����`EK�Ꙇ�q�D�cg��F��EV��0��}(�M[Ao��>@��sgW�d����O�@�M�x!<�Y����$�zɆ�f¦m9���?�P�9�����ȓ~}�Y��O>xD1�Dn)Z�цȓh����F웲Q9�e��o)D����aM�U�T\s6QT�0uӤ�+D����.�	
����Q<m��ŀ4E)D�PaĬ4Y�5�c
O	)j�x��!%D�(+�:J�.M{�d̚GK�K�""D�� ���Ԍ�P���@�X?4,�1"O0|���I�n�^��+�
^�� 2T"O|I�gA�/I󴙪�
LM���"O���Qa���|@PSIH��ڑ��"O(E9����1f��J�"O�|3&�ɳK��mJ��FQ�t"O�e��!��	��t�#�L�	�����"O���p����1ʒc�04*��hW"Oؘ�r��>G����CI4_���1P"O��n�~��!"�L�L�"O m���0SG���\I����l�!��[	J����Q�>�Q�E܄�!�dTDD� 0���s� ��ń�V�!��e�^��w� =���K��Jg�!� !t�`���ʢ\��m;u�Y]!�$� k����5'�?S��9P �@�;!�����7g��0�G5ZD!���,w�-1U�܄n`�-S��Z<%D!�d�h�@���K>\�8��` !�d�4	5\�v	[9���X�A*g&!��{/���vǆ6��L�&gc�!�DP����R�3���� ��/4v!�6o6^�[�䌨1R���D̑i�!�d� ���*M�\F��Z�a�"`!�䊥0J�@f�ܬ7kp�0�mi!�F�\�Q�EDڲAZ��j�`b!��Q�ea���Q_�+�"�9~!��1X�]�FM�Y�f��,T!�D��y�����aT5ol���	4!�d��K�8k�m����"�!�$Ҿl=���+��~L,{����R�!�B�<)�*���Y���ؕ�ݍ�!�d�#)'~�Mϝ���!i]-lO!�ĕ�}�b�����@k��3	��!��/H��5d֛KS����&^�!�DX2|����+st�񠥒'P�!�$KAF(X-/i¤KдĨ��'��p��H@&p��9"���4�5��']VD���*!����$jA��t5��'�l����	�)����`Ұ�,Hc	�'U.�Y1f]X��q �	=iq	�'�Z�"�jB�@O���$/
&S��J�'��]	5$ɸ���H�&�Ҏ����,�ޙ�@G�*;�I�[�:]�⬂)C4����I9"�8��'�y�(L�"d�ͦ5!W����M#g��ק�)#�$�E�%%Ɓ-zt�9&� �䓎hOq�N�!ҦW�8_�tk�ϑ�)!����]�xE{��	Ȕ(6���e�:$#��^V���M����DH0GD��P�Z��D~9�E��"Ota��B;ju2�t�T<n"6R7"Op�� !	-*� �%_�B@�$4ʓ��)��XX�d����H��-3�0�a���>/O��O�>��c�)d\��f#O5x����AN`��J��D:�h6&�*�)���!��4U�vCB(�剛Fj�<XD�O��Y�e��y2�r�C1(�ޤ!��<qw$��Ģ s�j$�K�<�pvʞ)(�Ha�DB�B�0+���T|��b2�P#��]	��$�Ĕ~2���2���$��|��I��E����)C
�	@8���kZ���Od\�1@�O �a��K��f��P敝�� ��L�<��"����Ba�-3U
��	Vc#�H˥O؈,�ܖ'@���2�~�S�3z������z�b��V�,��c����I�8h�`��=�>|S����Ob�c�xGy��)ȇY}HH�֧�	j5-&h���O��=E�tB�P�� ����4�^���L��y��H
I;4���7+,
�(���?�'���� V�\$rkT	Ĺ;2V�z�b�)�� 䀊�G��5������<D��YK�|��)�(��I��R�x��f��4m����hO��lX6��{�]�A"T��Q��8mҸdl�;+>��Iܴs�~��2n;�)U��O��t���_^�NL���XjLH�'����F�>8����
N 7����'���
协�*C\��c��#�x"�'�p\q$��N'Đ���Fܻ�'hn�Y�ӹ`�k7c�$��|��'�ͩ�,S�v�)ˆ$�/o�m��'�`�Q�	��82`��M>cRX���'�ȕ����&Ĳ���&.�x��'���9B�^�Zh"��A�0%���
�'"�ئ+��P�[Q)��}m�1��'2��q�Bx`��h ��K]�q`
�'�N����D	^�Q�օ  J��	�'{T�	e(U !8Ii��o�Rlp�'⎱!�Ҫ� T8V,3}�(;	�'-4К��2t �A�ՙq"��	�'���kC!�"V�0 W U�q1<U3	�'6y"5�׮k�1w��2|ƪ2
�'.���c�A���=6�w��{	�'�n<
���5,$`��d�>y61[
�'�U�iM�m�����	r��<
�'�U�τ��|�i�%�f�&-�	�'?�p�Q��F���4	�='���
�'_^5������l��S�
�.rV	�
�'���آ��= �����Q���'�,��#%Ę8��Y!0��Ѕ 
�'�N-8wn�2�p�9׮�H��x
�'~ֵ��ɖ�G�� s��.v%��9
�'^��0���@W��+Dłr��"
�'��q�5mRO��3Cd �h��P�'��2%_�źB��'Y{,Y�'�,�u�\�-ެ�j�%N�V��'��tR�4S��b��>�LD��'$�rc�Q�.��1�L�6i2 0
�'�"l+� �!���{P�Ue���
�':�Qx�V<,6]��G,'�fp�'�8k���	F��hVL@� ��S�'5m���^"-�@2��Q#�Ṿ�'I�T�f�
[O�p�MQ)�x��'��`*�F�%�f��4���|b����'�Dp��b�z�����60*�'�	�c�#s�v=2�C����'�����ݥ{'r5H`)y�ݠ�'�"4�B�bP����Qk�F0j�'�]YY�ĝK��
XI�iar'3D�8����:+HX�vg����V�<D���6G7l�"�_�M
.m�'�<D�pED�r`!�,�" ���փ:D�D�0��$\�\�j���,�j�9��7D��d�=Y!�-2׉ѳ��s�)D���u�	���Ĳ"��<D�Bi*��"D�ĸ���	����-��+�R�sR�"D��S��:4�B@��/Tm�� D� �Γ	rJb�"a�,�挚��>D�\7�
zr$@�3`@9zv�c��'D�����N= )�qjX�]r� H�9D��:�W;f�����Ip�p�D6D�Lr�&(̢}�҂G
�ʵ���4D��`/��;�L	4�P���}�ec'D����m�'��]�`O�����'D�XP��\�@g=H�@�:�:`�VC'D��`Gg]<KCTC���C�2l{�$D�� �e��l\/3ꢁ���M�
�J�"O�<���6'��%�KoZ�Mcw"O����\fe|M:6��b���"O�)��d��ue�x�Eb�5��U"O�|�"I�G�Ԍ�tb�&=��`�D"Oh�
`��*d=�t�@ֶ1��]y�"O��	��:6D��!؝Ju�y��"O恑w ��* ��ٟl_d�"O�$�gE�iY�)�!��1�~q��"OҨ�"^�'�$�d���-�,��"O���.]4�r���-ڌ�\|0a"O�D�u�ͲA��)��-�$�#�"O��Bbo��	y�JCH���ѳ�"Oj����\W���d�2; ��"O��1w�'F�$��蜒"O�Š�KN�.48��0#��c6"O�a2�	�e�\�I��V E��[P"OT�('�ɝNm� 80gF�8ݪ�ӑ"O��	#	D���Qh��2��a�A"O���-\�pF����'�6�"O6��7���e����
��a"OH�Q�
)��X7)[3�ԩ;�"ONqb
0w����n��u���C@"O�1	��/�ĭX�/�(�^�X"O�-� �^;,kV��įZ3L�zA� "O�� r-�$� p.У.y�e�g"O���#oL}���i׮T0Zvj�Ñ"O��#ǡ%�݀ ��e���"O���a�X�!�#�SjW���"O$iBӆ�-=����E��F#��`"OR�KO�g3x���A�@�q!!"Ov���3U��A� �9`mB��"OZ̛����-��	�A)!34Pq�"O6�Ѐ�4�R��f F�\RV��"O�E����Dd����[�v.�Ӧ"Or��EFlC�-�����zr�B�"O��AD�Q�k��h�#�	}nD@�"O���̪��u�"!˽KZJ�"O��
��	J�D-^�F��"O���a��
��Q�l��_?̐�"O��kem�Scj�;�ː�zZS"O
|{򣑛'���g�°��U�t"O�+ ��f=�� !�g�l��r"O�L���f��`Q`Z�7��0Q"O,�Q!�?�U�rD�ir���"ON�k��.B��� �S�xg<tȢ"O�h@�bW2��M߷H^8:q"O�M�bŮH�b�c�!\�4�Zm�#"Oz�;$ĕi!0#�1w�a�G"O�	��j�v�Q�"ț��L�D"O�4�B��oj�	%���,d��"O�cJ�.$y��~^�xz�"O�$��� 	Nfj؃�@�:��3�"O�u��]� �����1:�a��"O6���FiQ��1��f�̤�u"O.�*�ڪM�T�6��=���8�"O>U��(�0�>|�%�*w�� "O̹H��A?_F���O-l�x�"O~�b��=	����.'�P���"O&���Ɨ?.�z�& �O�PՊ�"O�Ī�C�k���Ё�R �"O��-u����� Hrr�6IĄ�yr \p;����5`�C���yB��"gj��a�$.Hz���^��y
� �!��ɍ�;�@H�d��bmfe&"O:��CB;w��)��I�8J��Rs"O$��A&B�f��y�o�8у�"O���1B�+4"�pm'3v�I#�"O��Ѷ��L�̥0V�/v8�Mڗ"O��8cAPbqJ�w34�""O��WO's4AZG*=w(�\;p"O�d��fÅ'�����Q
Pw:�)�"Of� ��Y|~��4gS�&`�9��"O�(�Ҩ`I#*J<0�BT���B��y��Ǭ |��Ƣ�1-}>�)C�.�y�L��[���a0$�S�a��γ�yR��>M�:���6R���y���3�y���;QJ��)@焉M���M�9�yb��S�z��`a��F������y�AVkEt}��I�<!9S$�y���2�^A@s�^3��iZb���yR`O�p�h˰G�|��1�*W��y��XUQ��O	
���R6�]�y��E
Q�$�0�!K�~�$ E��3�y��<~u:A�2��5y���:"	?�y��Ɗ,��a+i��Iΐ�4IL��y��N8[8|�sgA=	�^�P�D�,�y�i�C#6�����-|\4rC�,�ybh�y_��2c떄b�0Jf���y��)?��a�DޮTOF�bei��yR��2��x�f"O��	r��V�yB�	_�	1Í�H��K�"���yblJ>:Hˆ�K�?�A�D��yr�B�2�0��ȁ@�l�v����y��?�x���$C�o���%��y�o�,!�Z�!�L<:�"����"�y"�4?��d�򬎾H�u"��]��y���>Z���ҧ kZ�T�	U��y�?	�t���Q0fnpU��*�y�CK�3���b*B�[Ь�y�ח�y��ݺ9��I�_h�bEg�&��p��'�t��ai��_dɣT�X��A�'�e��ɘ+U�جq�o�xU�}��'B�͒3�,b~�I�*�g�h��'�RQ��F�,�>�#&�K�d����'�@l�V6�BY�����U��	P�'�0���1HK~�`��_Q����'R�K�D�%j{�`j���$F02h��'9�^+H���@�Q9>��b�'-��L�<L�e:p&ϧJ����'��$� �߮D�b@�W�
�P�<݋�'�T�ѭB���+'�
�V�z���'[����	��"�x���G�D��ȓF�Y�� <
ڵc�$O�
��h�ȓQY���������$V�"U�؆�pnr�صf��H�i���T�B��ȓ6��Q����y�8��Z
-�,=�ȓ����ȟu�r�c"��2�����m\:Q�Ā�/]��CRD�_�����u�	Q�#� %F��d�Ӧ;g&1�ȓo{��A �A8.�2���;S�0��ȓV4�5�(�&crM��(��A��X��R�t� A�)#
V�X��."4@I�ȓ{ I���V�&��R��A`.u�ȓ�I7�V�5fpP`�,ˀQ��ՇȓH=V)�C	x�v��aEϱM8�p��G t�8rk��"W& �6��,D�l4�ȓ)�>�"�mZ�p���'i����S�? �@�FdGYqa��H1�9� "O`[��E�+��ɣ7���:oD�s3"O�)I��|Ip��!��~^ !�"O\P����9=��\�� 2/S\Uq""O*a	�'�S�
����^��"O���7�
�}-��Zvd]�cg��"O�pkŌ;�~��ը�y p�"O��A��������6�2�B"O23� 
  �X     D  F#  g.  �9  E  2P  �Y  �_  f  fl  �r  �x  B  ��  ˋ  �  P�  Ş  n�  T�   `� u�	����Zv)C�'ll\�0"Kz+��D��h���b�&�ی�y����yb�҅w+��`�\�;®�"f�YY������$&>=�0jQ6U|lq�UE�-��NÖ�����A�d�)Z)F6�(�M����;w�
1AGM
69|"��v��&vK��V�C^Y���Lk�'�?�5��
Wi�07��!5���kcL�CC�Pi�a�:���Iw*|£��*	�d6�Ͷ<����O��O��D��#�d�Bnـz�p�K��>{���d�O�l� �Ms.O^�O�� �I�O��$Qt�ɀ�͆?��̓7��@*����OD�o�۟x�'��-@<�u�O�$�\���8o��l�U�R�SdRl!,���F���X���'�T���	a�Phs��,B �	�)��?�lIy �@}�7O��Ob���  ��,ed��2�����I21f��3E#v���'>��'��x�����Olʧ�y����l�F�"�l���?�f�i<�7��즁��O�~�����䦍�#�ͬ]0�/�(>#��eΐ�6x�vE��HO~���HTو�:w�	�>7m�Ϧם�O^8�x0o��{��V���[$�2��i���XэPh�Il��M#��i��Dן*�/�N�Ib�$J���+�	�;��QТ�iL���1	��}�4���#�
��M���ɳ�8�WksӮn�*�MC�O�'���
w�Jd#,�e�nLbT�G-[�f�#�iڠ6M���"U���S����`�(��h��c�������)A��I6i@��^���˙!
�xtO3�MkðiH�7�S	�"�K20z5��ƿc��{��O, o����:���0�o�����HL�B� �үЕ�}	gd���T�?��F��J�9�� �^���ܷ�?���'��'�7M�O�DU,fj��$�~[�AZP�
t74���O�I����O��d�O�9`"��n9��� tPQ3�߉,x��s�戄Z�V9�U�R�	�����PQ�#�f�m�ucR�Y�R�����F�{-��ǎ2S�(�bt��z &>�d\DyRƅ��Osyrg��0�
�!�O-4��	y��X��?����?yJ>y��?�+OP�$*#��xѵF�m}ʅj�R�n���O�*!�LY,�O��9O�	�՟��懘�S;xs��H�p���%��O�˓R�0�jT�i*�'sb�O��x��'�,i5��B?Z�K�Ūa|rۦ�'���ϧ#�X'��N��h-�xY�`B���V}�Ӡ6.-���1����0�*��' �,��)Y"��EM��[CQ0kЭxe����|;=;4�ɾ}��p��
I3���|�ɭ�M���|�T�B3^"|�p+	m)�%)�B�ȟ<��ß,��v�O���"d�¥<Q��[�Ce}C���Q�A�ڴ�y�i��	�4w��P�	A��X�`�@��B6M�O˓������?I���?�(O���A�D6C�
�4XmBBD���I�Y�"�	˛+��!�S>i�S�l��tB����$E��'��@R�ۢ4	f�t��3~ �ca�AET�rc �8@��c>ep���w���ǟY�������4��Aǚ�|6M�Qy����?Q�����|"k�$C]PD�TJ����ղ1��'#�)�禭�Ĝ�lWl��Ԫ\�}p؜�6�'F�*t��o�^�i>���yy��CS�������}�l�$�<�^9���+!��'��'���̟|�I۟�s7b��NڶQ�l�C��JA6"���f�2a'm�(X����"'�|���<�5��=��|cF���cc�R�Gj�i,e�����F"��y�F=���<�ЯH�Q��@�p�A1q�i����-��	8�M{q�IM�'֬A���9u>UZce��&d�.O ���ʚz<e�̃�f��$Z�k
�e��'
�6Mݦ��'TN�YGk�P�$�O<��5��$�҅3���p�P��7��O���	!~0����O���͍�T�Z%�Q��7m��Cތi�D'<E~�;�Rb��@��G{ a#�Wp�drs^C�6��s�C�O}��#��J9��1'K�jG|�EAr��P
I�Fp�M>���ן0��4P՛��'��Y&ڬv��rĠ�.0C��#gU�Xo#�?I>�cܧUB��@u�Dr����,��:"�y�?�I>�����qナ��ABYa�ϒzn�{��M��M�����A���}y�ЕEC��?U{ߴ�2�0D�h��q㐄'r*��u��+�?I��cЕQ��)j�BS0O8P��l�<�:O�Q��m��^/9�b�S!Np�|�'��;�G�u�F��ύ*:�|�QMI�;t�+�뀀����Tw8���1��p� �[Eߏ��D��-e����K|����Y�'�d(G�П!'�`B� �䓸?�J>��?�+O�����%�TWMw�Vհc�y�'��Dj�����ɦ����a�^)��'��:�:�E������4�?���?KW=lN2�2��?q��?�w�`�SlZ�<���%��n���{����~� M��lL�7mTn���?���M*ezd��#_<>��p�[�hA^}*7*�dF��r�=&���╭D��6��/}Ъě*��%b6Cʩ��.�C��!��1�
h
cM W�6Hyb S�?y�����?!��H����9�(�y���1cޑ�L>	�\�|��	�,��f|�I֟4	ߴlC�&�|r�O��P�L,x�K�P�c�E�B�Hj�h���ʎ*�ڟ���̟���=�uG�'�25��4#�i�3u�������g����d�K�|0#�B6k}���U�D�;\U���(�(O �(ۻGĂ��2�����Y(AƝ.ָ�������CMЛ��!�֠�(Odz�
�#9�>�A��t$*�:'EȂu�b�'�"�'"�V|��ʟ~��hcgF���"{�	�D���U���Z�%��ڴ�?q)Oִ��VЦi��՟���DG�w��8dG�oW�1� iğ���� �lt�I����	�^�ȴ@+»~��0o�O�H� x��2���#k.�`��c�2�(VEJ��Z�I��D��"n�)�	>Q��a�U�D6,�̌�'�݅{E��"D��##h��m�O����T�D�v�&�O��ɔ�' 7m�FyrE�? P�l�6fX䑫��������d �SB ��;K��\��lL/I�`Q�ԩ�M��hO��~Ӯ@�2���D�t��%!�p@�֦�'�����`�����O�ʧ{� ����0,ل��c�x͉�c�!�����?��kڇz8�a*���I��P��I(�N���	�;;�k �O� �v�85
�@��I-���r��(ǎ�d��IxmX ���/��'v�m�D��4�@j�B�$	��'3�	��ɧ��і�J��Ѡ@���R�uC�"O���΃A�>�B�L���
���I8�h�xJ�%�uB�x�7�PS�����`Ӭ�O0E�"(����d�O��$�<�"aR��iS��
 A�ǂ�4tfe�2&��=OD�I[�}W�=��i�`I��(���Ŷ=Tx�T%���8�ʊ=����@g��\!R�10�ɏkp��qJK-	:�˧^J���e��+5��3��T�6��RLXQw��#�M�Y�ЈbB�O���:&�8CB)Z#Cj ��B��� ��l�ӟ�	ry��'G��	��P�BS���!�A慍P���Iɟ��44�V�'�b6M�|J�����"5��{�K�~H�i�@'m*j%
 [��e����	iyBU>�̧mhx����]�=�0`�#��n����C�W�Tڡx`G��`P�U�ӂJ�Ձ�c0�R�=)�LG.�:]� ��	/��pB6Z��v�C1�S%i� �Ɉ�U�)+�K&.���K> �K%(ޠ�1��?���aI��W�@!����M���	b�'d�=hE�0|{���0�N1i[䀳���<وy�!�-9�MIӼ������6ƛ�jӨʓ4�F��s�imB�'iL1�l��5Le���:]s�4�t�'��B�"f��'��,܃OT}��#k����?�:H��GI�_���2���w�8����'hy�TA��5�� �ũ�ex�A��V�4�ri��o�����˄GQ�!ш�$�.mSb�x�LI�'�,P`]y���8���K)��K>�	�;�f̈@ �D������D!�'��{",q�t�!E���&G����\!16��Ϧ��'���)i�l���O:˧<t����]j=�`�|�@� '��;���?A�# �?��y*���r�j�gC1u�����he�'���"��ᓎ�d��s��(U�ű3�4g��R��9�ɯ��S�O��%�E	4EJ��S���S���'rzQ�KѴGv�XN�r����$�>��I�Uyص6!�"W8� ���Ӷt��(Pݴ�?����?�W,�9�R�ϓ�?A���?��w�m�b.ѓo�!�M�E����T�ԃ�νq�"�90��������Jt&� ��	D�Ł-V�)��H�n��H�ㅤp�lRe��y��c>��vn]Yy��|`PuD�5ή,s����;-�&��<AFe����D�L>Q�$�8W,�a��T|� <KV���'��	V�'��ѱG+���n���r��[y�p�Ԙo󟸒�4��i����'}�B�rk��}� f�F�`&��"o'��I���Qyb_>ϧY�ڈP�H�#"��%�DmD�]��%/T�%1�ݫ�<��Gm�&o��Z��V���<q2�ް|x�A�U(E�7�p�Ӕ�͍f�ū7�үk���R	
�}od�%�]!N�<�� �$!�,\�џE<iA��N�T��E���M����K��4[`��V��LHVU�"e@�j���`���?���hO�b���sꀔhE.�胭�)(Zl�0�D劣�4���_1�����O^��ȸ���Vh@*f@P\뒢�3-S���O~u��d�On�dl>��n[7am���C�Z�0�\z��C Ptڴ���W<k�h����V�sZ�qF'�_�Q���i[<R���b��*Zh0E�|�V%� >�� w��$�rp���N�W;Q�H[���O�$�,�$a�p~р#��E�T9D���ELӄ;�������LH���"�M���i]���2&�c(��kr�ԤzV�h�<���2 �lZ{��i���'8ؠ�@䁡�:�J3��<xB�`��'%��I������Eޖt� ��aG;E��hCp�Ѭ����-5��i$�R���H;���*](�Or�A��,ӓo����񂊩��CU�ـ]�"�ON�E�C� ����q��>1�$0��Ohy3�'��7-�I�O��	���Kf�.�qk"�R�|��'���'�2�S)iQ��ʱ#�~�6��j��C���=������c�(�O�)���п�>E��(�*@���K�Ҧ�	ϟh���l04�["E��\�I��(��ּ;V)'׸��ċ"@ԴXq���P�����ψM!V�U�ɲ���|����/&���� ?�T��󡎸;5��`���,趕���˵
?N� DǇV����b��=��p�Oz��c��2�y'I }����2����ȏ�`�&��<�e/��<�Sz�L>�7��'1�`�۱��aʬ��ژo!�DM�XA�c7q~�;A��m_r�'�"=�'�?�-OĬsq�����+D����I�w��|����`�O~�$�O����Ѻ���?ɝO�,a����-Uj�qt	�d�z�RBB�jl�+���}�Ȝ�D�3�� �2 �e�'Sl�c� "��#�9K��a�w���`3Rx���=^F��5�-ouPѣU��WI�����1h�t�O� ��ǜ�)�F9U\��a"2)^�B�/t���Gz���&U:1[Tb�$�(xz ��Lʒ��D"�	9nec�h�/.�A���Z5*��Oh�o���,�'v�s�ý~�d�t��4⏜C��EY��
n�������?��,�?a����4�-�.���	�\�` Y�	�s�,=z��M�R5b�0œ.0[ڥ�V��c�Ey2��fZ�LH`��
7%IҦ&`8��#h��>��a�"�Ӳ#`X�1U@���`Dy���?! �i��
rb)IAS�!��iw�2k<)&���	 �f�q%	/ӾSd�B K��@D{�Own�䐂E@��B�O����+���;+U"Q����M�ty��'�4��d�I�/ؾ��a�en���"�Cw�"=��蟜I$`ƣ���q�h���R���΃R ���|��0�@�QfL�d+�ɱG"���� ����R���$	p���[�qB h��Im�ӇLh\J�IռR���E#I���y�d��"�M���i5b�~⩟���DA�a�޽���N5M	��s�'9���J�3�'��|��EW�J9S�cșa��?R�iz�6m�O�mß�1#Iߡa���C��.+=�(b@���Mk���?����
��'��=�?1��?I��y����X��Yɕ+��(���aBe��'�v@	ӓ1�� ���"m��بe'�6o�D�<����o��D�6aɩvXmi��ђ@iA�z&��O��* �'�1�1O�ІE6��,�EΈ�Z�� ;�"O�UI�E�����Q�b��d��>�q�i>='�h1F,�)�̌aÂ����p�a�CR�(�M�؟,��ğl�	��u��'�27���ō�#E����	7���c�;*��Ur�bi�hD�PK҃KY�⎖>�(O�Ub⤍s7����P�p�qB��e��@��(l� �ɂ*Z1Pv���(O�1�EWi�����V�
�Ps��� �RA)�O�`(�n�P&�����w���R"O b�Un�z�h�]�+�U�1�|�nb���O&��5��Ħ��	��0�ařVrj8P�E#�A������,�B������'u�X�1( :;��Ҁ	��w�D�s&��nG�lr@��j�J�J�	�ؠ��#ʓyG��s�
ú1��};�LG�>cj ��NЀ�E,	�UG�9!5%WS�B1���5ʓy�\��	3��8F�<C`��<m����Txt��ȓ$$$`��H9��!��$b�<��4�O�>�?�ď�52��8tj�o�����H�S�I,����ݴ�?����i3t����ۥly��(�(Q�_=H���FJ�$Oh�$�O2Y��O�b��g�D˖@:��1
R�ʃ�S	K��O����)�'4w�}0Vj�j*"9k��ߜJ�'�\DB��}�ɧ��5����k�0�C6P	@rbP��"O>́�L/S�����*�
:U�UA��I��h��phR(�|mV �A	��j`�i��D�O���ƾ+%� $�O����ON��{�Q��,�����@+̊��l��V��,��4��B��tRe#�|Z�'0h��@�V?Q�jΗ?T�,c�wF *̡y��� ��1fLhm|00O�4��(�l!��c�,p�ڱ��A�mC�,Js��]�7���u�I�;����IA�gy��'���.�_�(��RE��5��"��'�ў"~
Ǩ�{`��F^vf�34���?����"j��O�Q��c��7�`��h�1�\ K�Z��,��K�%�1��?Q��?y����$�O�����%��
�F�0�'�6��� �,G0*��3ύ�'�8�3�*o�l��I"J<���Hֱ&>����Fgvh��  �%�v3r%˙+�(x��:b�p!n�,>n $�|!�H'QrA8�gY�	����#��^.���[¦قM<q���?a�ҍʦ8���
��ڂV��a'T���O���<Ac��"5�`��ú�&2W&�o�I.�M{ �i��	% *�ˮO ���<�0���!�\)�P��7���$�O��1���O��dq>�`s"T�1D� ò���䞺F�PTq�.�-z�2��M��8 <�k�Fy��]<d�4Ų�$��:��.Q1�l�t.�84���I5����2sɆ.r�0Fy�� ��?��i@��d����) F�|�sֻ6��'�0��ɏSb~yQ4JN<9���@Q8IG��0F{�O+���Z�!AI�D@ۼkw���'�(�2Q��	��M#���?!*��u1ҥ�O�8c��YF���!N�r!��C���O\��]�vt*T��B%D����gٙ52ua�� EO��v1Rz�(
�sրp� �P�'�r����_����
p;��pty�����毃nk�Ȱ5k\�1l>��ב���a��O�1$�"|p����8 ��!
K䀉��G�<�(Z�ye� ]���VeE�'��ɗ�HO@9C����O��(b�
6�������̟����_��e�UG����͟��I��# �цp�:�hѦZ��i��&1��ѱ4�U4D���S�F�� �0��|2O>�U�F@�u�.�Kyfx�)o����_#}���C�!H�j��,�|"N>� f�1�ʋ�^p �ʳA �H�~�� �'a�I�E���D�Ox��.�I*�����d�U�"\��
�4 �|X��TLv �fM�2	�|��pK�&'�H�'5�#=�'�?a(O&z`�޶X�J��sa�I8PP�j�!�H�b��O����O�����#��?9�O;@��Ф�}��"F@�F�蹀gMҍ9!� ��&��d�V̐�H�џ�Q�g�1xM��ᑀ:A`��K��M�l��B\�[I�����'϶�G��S�q�l����,|�ѱ�� =`�P����?!����'�>y�!@�'%9TQ�e�\�Y�$��n5D�86��Kq�Є���T��i&�d_����	Jy�)�}�맄?��B�$��P�G=kU�ek�'Ï�?��+����?i�O��ɑf]6Z3�5z��·F)I�Y���ˇGc�����甁i!�Nc�R	Fy�I<K� ����:(�H���@�SŢ�!Q�X�{�$��P�X�Г*J(LP�Ey�d��?����О0��!0����N6japڜ
�'#�'�T]�@ЪU<�M�C%M�xd|K�?���#O@��`d�>Ipu9�����?),O�ݻ�����S韄�O[H���'��y���Ņd�z�`��߭��$Q�'\��_3&m��)G."��� H�^���h���.��Ӎ.�l�Kc( �!��D"P�׼��C �U臦��Jv�2��@��]w"��Q�PC�����E2*����>2wT��Q@֒P����|d����O֢}λ�\@��fȤ���8#��� ��#�'�5���@�������E� �)��d�O:�Gz"&�6c.P<��BЋ<B~�	RGϐ$�`6��O���O�c%�S�D�$�OD�$�O
�D�$�ZAoT�95��p��@�@E��"��	dV514�]�@�)�S.1U�ڣ�O��3�Z�]b�l��b�7��`D5)N}�$�G�6O��*1 �/hz�|�ċ�\A��̻NgBpz�&�W��<��Zt��	U~BIЃ�?q���?���醿3bK2-F kXp=��d�f�!�Ā!Vr&�`ƋX�?��4I��zB�'Cv"=ͧ�?.O�-��
�&C�,�#�L6Nീq�<j��PJV!�O���O���������?��O�p=���C�4�x��2�� *�ᑫ ��@�IGU����(@�b{�=ے�T�',��D(�9q&T䠢���Db�9�u��#��jDA�r�l۷@֝[�Ĺs�n�q�'��K5�=Pp ��S��c��MsՌ���?A1�i��#=����;k(����W%�H��5M!򄐯*F�p�,74��1���D6�'��7M�O�ʓ0M�e WZ?���F���p舷WV���4�k������ ��
��`�I�|*�΅�Dk��7o]W�M)w��-R �BǊ��g`�0���D��$�Z�f��@�Ģ<!�j�S��@�"��U�A��N��@ь�)���H'����I�� ���<1J����iٴZ]�	� �`���D��iA�T˶�\@�O���$ͯTl2���X�]�h6�E	I�����O�Uo���4�8Ǥ��5����'��Ɋ��Xڴ�?A����)9r^�$ܺcҚ�8D�?2�t�
�A�a�����Oh�B@OH�	?��֤Y��,�ׁV&��$sg<�%j �p�Dɘ!C#<�$ ��r~b��zN�x���V̬�1���6���A`��S�$�6H�F�ϻV;�0��'��D���t�v�I��Mk'�S�|2ׇN�:o����f�� �lH��V�<!G#��H�<���^�ɒ�q�w�'�̣}�G��(Vr.���T�l�P�G�M���?���q�Rm��kC0�?����?����y��5���!$#IU�m�*ڇ%�pUPp�BU�T�(�,\�F� ��d�=�$�1r!��b��ń�ȩ���K��KĂ�G�L�"�*��R"�*�)�*�\�[A2�Fl0�a�z��qT'V�P����	f�&!�'�T�����ȟ�'����`K�<�����G�)����"O��##LĻ
���b��ͭ?�P�C_�����4���ĺ<Y���z>��Ʉ5}U��#⮘�o��t�VJ��?���?y��:�N�O���l>Q;@c�9+J���,�9$�<T��gùe�����'���G/�8B���2bdIKZ�De�@m�3.�h9��J��~��Y���X3��Ba�����	�H��y����!5cb`������0		4��O�QnZ��HOr#<��,m�Y�p��E~�l���W�<Y!��X����J4��!�n�w�ɫ�MK���dº!�@]�O�ₒ�:�vAY�O�8���4!M%��'<d(��'�=���Ad�*���f&B����bnI�,�\�T/�a�JPk����\<á��(O�(����^�G�h!udW}�XhãHO]ޖ�;vJ}ļ��N�.�*�EyB���?yB�ir��b� ]YpȎVQ��*��x�T&����	�6���V)�,^�Fm�6+��$����d�ܟt[c�ѢP(Rm;v�W�m�n��S��O�˓P���i�b�'���7>"t�ɧ >]����~_������B���͟��5�1)\��8'L�P����I�a�� 6>�'���@AJ�r8�@��
�#:�d�'���@c��pl4�� A�s���2V������ƪ� ਴��O�?��+���LqG��O�m��H���3� �� tϾ/VqtDڝy��"O�t��>_*`���/j�i�U����h��,`_f\�yR�$v����f� ��O
�$Jg�� ��O2���O���b�ňt	[�h��c��^�=p(��ϕX�zՋ�`�$L��JP���p�&b>;C�(G��$�3w|(��a[��nu���5�C#��Kldu3��ҧ}�<%!��I^<M��P�'f�����؆�t,�$.��KX�P�i��ʓr4��I�?����;Br��J�tq�/ĺd/u��O]�<���O�BhrX���
�P�*�+L�dy�f0��|j�����b��@�Z�h�]���	�Q�P�ӁBЍ����O��O��;�?������Jd��r���g��R�M�2�6�(F�B=�؉R��U6,�\ ���X�lFy��<$A$p]�~��5y���$/�� �� ���$/��0��kA8(��Dy�O�2�b��`�V \��uq�+�D����K���c7��O�]�g.�.R����7_B��"OR\���W��ͣ�b��z9B��|�p�p���<�eY+o��&�'��!X	0��dK��ηa�(d�4ᛮ{B�'E @:��'�1�R�*�i�@�ɷ�O�gM��"B��c��	��&F!g,hE0� ��$@��КXQ���J!wC��H��;.��$H��݂pwh�TLV�Q$��*Z��ytX�v�Q�(I���OLQ'����mO$�,��Acн��YB�>D�Z�腾�`� b�I�,�"�c?��w���D �O�@����u&Ti
dC���D��|��='�6��O��Ġ|:r�C�?�3�W<��x�hޒ��Z8X��	Ɵ�J�I�;��m����]�H�	�/�/q��L��.M�dg��4��ɀ�6����Чك���Q�X`�%�&gC�%J�Q�a�*
L���'Oy���L�n�Wmm�yC�߻Q �-�6l�	�MCT��|2�'�H.�@��4|j�!J!�I�<� �� ?�)�U��.S����w�'���}�A�$���#��9�� s�ˀ��M���?��~�N$ �����?���?a��ywn����a�Ie��KW���V�hcfU.���*w��|�RB��$R�F�����9����0n͡2䤑	�/�� �"?��S#�)���:��P��.�+�j�#��A�uU��ݓzV	Q���>&�r�2��ć���O|�2��'H1�1O�H:��֩�D��ܐ�z�"OZe�aO g�Kt��&ή](b�'�b�0��|2M>aW�ϳ6K�̱B�[?E�����
#0��4�4kO#+&��#t.A(+.P!���1m��jugY8F���#��#���$_��h ��A�<_6 !QE̴�?�����?���?�R4�"���Ń 3 ��z$.����3���`�hNe�����X���Gy�'�0I�nʍ_�JaZC��4��%���Z�^4XF�\��,)��$��d�2�2Ol��'?q8b팣%쀒ӆV�OjT��J�<)���4�S�W9D6]�DdI�B>�O���'�1�0�%P��b�X�J�![,O���7��ަQ�����O0���'��G�!D<0�!�re�����$T�B�Ɉdr�d!���F�Cd��"����Ed1���x�!�:�\���ě �=b9Or� 0*�7:"p�1pf�(1�qѢ�Q�
��|��d7�邻oRE��e�;zA\�x0�׳;|�ĕ$Zy��u������'��	W*O�D)�N�r7\p"&c�'c�!�L���m8�mD&nPj&�DH�ў�،���nc���P��%
�����&��
74��O��A'UP*M��C�Op���O0�$�Ժ��턀xG��R)>At�� 8;j�K��^�H����SO��5�ХR/��)<ꐉM�X�u/]�B�p��c LY�qb�A��j�v�zǦC�h.��t��>6Z�'f��zg//}��ߠy_��p��S���26ңi�	 &"��SԦa����y҄�(4b�=�@ـ)�8�Ȥ�ΰ�y�%ǁ(M@[7���2p�f��?q%�i>���\yRB�%=AD}IW.�0�$XP3�8Hb�m�o�6r���'w"�'D����d���|�D]�F1�)ʆ֊W{��Y���qX�4MK�_��yv�	75D�3d�,|�h�<A5h�����7l�<���+m��9��.Ǌ=�p�����-�h�o��,���<�b��s��/PYL�ZG�Q�CӸ�	b��M�'��y�'z80����V J��۷)���'�����`�!&�n�BU�X�S�f�!/OfElZ�ԗ'k���T�~������ń:O#�X) ��wծ���L��?Q!��?����?�� ��!L��e5E�vhZ�@�P:�,�0D
�yuFV�r�aJd�1�.�Fy���0+�\@�>H����6J�
��=�sɟ�%9� #!�M� ���  O�W�"�Ey�O�?��iYB���Ze�N�$	#8����Z�t��	2`M.�؄k-#S����LH'G]�����Xy2F�nb�5�v��=8.P�˶���D�T�m����g��(����'�<1����`�>��aE�X����'�ʄ��18�`rH�
����	
P���r�)͐BG��[�����:q5��
F�(J@#�#B�`v�A
x1ҩ��Ȣ#[f[Ui�|�7b��WB�᠗��Ϧ����<A�[Ɵ���4U��)�)<� ��IN�[s���CÄ.j�E�t"O�$ u#��E�4p��k��K��Aр��O.PFz�O6x�04��Fv\8��I�*������'FB�'?<�B�c��+��'�����'q��{Dƚ�X�E0��ʭy�����W6fQ!��9T����m��S-?@��6�>�"��S����A��1h�ȝ�|M"@���@��)T�ט�P�O�,M��N�t��I<Y����-�J(v؃��[j���O�*%�	��MΟ�'��䞰-� �B��YN����E��!�'CgHŋ���T~�LJ$!SM��i+��|����dV>�����C�l�`aGغ zX����.;>&�d�Op���O����?q���dL�M��h�3��<]@�� ��Y���$ �xպ�	!Pdf�)����qk<dEy�#N�.j�U�@	�<	��-a�HǤh��U�1��:#��|��b��"6��1 ��ɂ!�z���!w�!r�*Ȱ#���qCY"�$nZ,�HOD#>)��]�Nq�񂉧)_Z5�7� V�<)w��`&(-�wC]�<���
e�TyBOa� ��<�4�_:v���'��1�N�����y�*�	 �Q"$�����'��@��'hB�'���$(�o��x9�a\24,�N�J�8l��D������JѸdA&��F�=�(Odl��B��^m3��ܣt�(%��l?Q��a�4-��I#A� :!�ܾ�(O��ˁ�'��?x��%Bmй:�R�V�L���++D����,�-p��pP��[�@<���(?Y��T>}�-O
�Q�߿B�P9	�[�(K���D�O���Ol���I5j�M�:�0a�ʑ9@§��q}�5O��ĵ<a7R��>��6�1O+�u���ܙJ�0�a��2�I�U%���B��d�M%L�(�ySlD��H�t	�6eg7��O��@��`�$Ҧ�O0�����dr�4��I*x�r�$:g��@a���> �m���PA�L� ��1W������
A�dm޽1��,���x�|i"$���CA��'?XpH�6Oם�8���?����<���[.���'�L��41���	ʸ��ܟ@K1n���@���� ���]Y��dg���TSR �P��sޘ-��A�O�@��'X��
$�'�?�����vؠ���';�-:�A��$���u�'i�p���?��lO,�?���'>�!���M�u���ZhFۧ��f��8��@�+�:���i�V��T�&�2�'>��/�OX��ݟ��I�?�[Uj�+l�9B�S���m���N O���Γ%o8i��ǟ��\w�2D�OLPʦ՟��*�6�0X9C	o9P�X���D(,)h#Lc� 牪(�oZ�Mk�a�y����	��i�$* �7�t0��N�ųs�æ9����<�4�_��M��i3��'�<��U"����\ k�Ąp��i8�r�i�W�:6m��R�lZ��?��4b'���i&h�)�~"�'cgt��u*vrf��Q��0nY
��"O��R���������ʆ6#Q�i,�R���	���I�O�$�Ot�d�&c��	S�W<���al*3��'������'�2�'���O+���"���+��j���Yֿi$r�'���'���'V���ɚ%�v 9��@��,��.ܡ0��*޴�?i����<���4/n|<q�(K�H$D9$e�/^��^�IX���d��;t ��KX�`J]�d͏s���o�Fy��'6��~�/O��佟�R�*�)�N�wA��Q��P�Ba���$�O��d�Of�Ŀ<�'��~:�$�ac�o��4�����A�B�	>b/�U�W���x����Ɔ�A��C�	8:��[T鉎J���	�/K��B�	m,^�����/���h��J��B䉜
�l�ѵ0�RtXg(BvB�;����+�,xؠ2d�͎��㟌p �/BV��s ܑ0v�� �ꐆ6����۰wx�HR ��'^�j���z�(���,y`sƯH�a�ڽig	�3P	���� �d�h�	��]�����	�=-�K�ǎ d6�@f�D�l ���>y�lۀ-����3n�6��Y�C[ܞ]8�/��7��D�ä2z�qb���2��gC�~z�T[�cׄE������Y~H��@70ha�2&Ѡ��d��lE�\�7kN��bs��Y���J1E�4x���k�οQt
=�eѲ,"��"HB�*���`o�ݰ��]x�$�%��l���!Yh���(�?A��h�"�ۆG�'=�b|у��?����ʟ;np뮢~��� UC���Wa�)FF �׈���20&^0q�M�o��x3�E	X�*�{�Q�����ֹ�f�#&&M�'�͒��?��ibӲ�J��ѓr{��Q$[FL]�"O>�#eC�\m���MP�^Œ2�'���<�l�I[.�t��6IMBu�W�!,�T7-�O����O���`��7�����OZ���O*��� �d��*]>ܡ��J�`��0�s��M�:9���k�Tx�*��\ļ�x�'��@ã-(�a� Ȕ�`���S�)
)�bM�fת���	"U�q�*��G#\�ӂB�.�T1HՄ�e�*a2�n�*-���O$q2�����ēA&���W��e�S�	�����ȓ\����E	RLf��2F�Oܒ���?���i>�%�0[�\�&]j"혟`���Xf�
�n4��u�&�?���?	�� ���O��Dp>��Wa�;��Z�-�.c*$U3�/,�m��i�1��y{��_��H�璜�Q�԰� �}���8Q��1��̜ �l,#6��}/+����+���N�+b-|�d<�JD�9q3��BK�ը!V�rļ�(�aҟ���b�`V��d�}c���1Z*6�ȓ*Rʝh%N��l��#��۫8&X��=� �i'�'���� d�Z�dmӄ�"Ѝ�h[���`)m�B4�TM�⟐�I�Pw̽��៬�'K4<e��X0^���˗KL�0��(�#OZ"Re��?}CD1�f��f�k��7�Ee���a�$Nc�婥�:�DL��Ƌu0&��AOۙ#��]1��J�h~���?�B[����;��	'0Bdm�0�P�of�� Q�K�4C�	�M%{V�	 G"�#��rC�	z�������$X��"��6m�0;2��J�I(�Pp�i>E�Ii��3:��y�̈��灀%�n��C뉵|�P���O>H!1΋�B�ʆ��O�����Ù%��(�;���E�4T��A���C&����rB�'[X��F)
�}�Ĕ!� �$�Zd �f��l��'�"� ��V�a���J1\N�$������O��$>�'�M��8.�$\�'�Dk�&LA��N\�<!!��83�K}D�Rg��8������[�|� �i�[�F�[��!�Z̹�4�?����?9tj\�i�*����?y���?�]�s�6�y��bY�#ׇ��Z�::�o�	S�u�ܢFU�+�H�+�O:�ɋ�G�0�t��-t�l��HM�i1@u���
;|���Aѡ¶�2�e'T�3���4��d�Y�=Zf�ݯ̰3'I)�0!"�.Q9X�*��|R.�?�}&��� �7Ef��j�5kZ4KA@(D���QE��C�n�0g@�(�H,:6E$}1��|�J<q�([#@Ժ����:W>|\p0��G^v�ae&U�M(��'y��'ں��ȟ�I�|��˘ ry0�/���Lys	��y�`����^ �h�$LĔ�|�d
ƁR2�<��cڀDk���`)M� �(�ȓ�X�~M g��?�H 3��[�<����יD��<q��ܭ�f���C�ZT�JҢ٘f����	;�p?A&�(qx�ʶL�48���pKA_�<a4�L��R�Q��	<)2��Y�k�Ƒ|B��3��6��O�7��)$���c��\
��D��:�< �����jf�
��	�|Z��f��G)^�/����h�+
�4@G�2������6��C�A�@[�<1F�2��@��(EfP{���PM���GLZ�'���)���u�>xy6ɦN�x�<������K����	^!7l�����a���@%M;D��Q��*	�րhr� r��zf 5����E(cu��9uB�1��h�Ƥʛ8P�&�\��'D؟��	ӟ��OӒ)��i�*�[��L�+���\������O���ee ��]���U��@�;+ `� �,� �'=	<����	?��8%Ŏ*}��'�����
�$u$�vM��p� c�
�(����S>%ӓ3ol��U	S+% 6 aw�<�D�VL��'����7�z�C5��.��"�iz	��'����mϫSe�Ӡ ǹpʅ�BPQ�p1��k��̢�����f�	d���'N��'�<�⢇�:���'�����+V��,x�U��/\�`����aջr�@Р���]�*����>+��[E�IY%+zVu*�y�P�!a1�@�2�I?!n@m���ɨ>s�����2�d�s�'�θO]&�P *m�)�S���q���J��S7C�,��O�2x��'�$���S�g�ɲ�f���@�"O�X�&Зx��B䉷Bw����c�F@��W#4���'�r#=ͧ��hX��ScO+_�z3�"*R�E��ʉ;�E��'���':�c�-�I��ḩH)��,r�4 ��M�"��
���S,�!�3Tċ!�N6g�ʹ��/ʓSڑ؆�ӿ?��ZE	c�]�a,Ye�A�P�G1V9R���fzM�
d���(O�9ز��o`��C���YPFIq���-��+�O����&R/{��r�@F i/��!�dױ>��4Ca*�d��K^�a�qOL�lc�	]F��
ٴ�?��4C6��uƘ�6"�頍S�X�F�3��'w������'Nb&Ҕ':�ɉK_�y���3���%>����ʔ�w��kce�0	�ڹ���� ?ٞ����'t�� `ҭ9����"ʠW;h-:�*�8��	 �m�� bD�P�D�;BؠL�@��&���O�H���'m�7MG�mZKFUX��Q�:���"3�D�D�va)O��'�i>�%� ��A�:��!f�H�f� x����'�ў�S�qjd��S@@"RSL@�`$ .�0rA@0�M�(O�-Hf��˦�	�X�O����iʾ��f �2nW�v)f\Р��O����������K�Lm��!�"�@�h!�;AGd���t���(^���H�0G6��'�4Q�mގX����v�~Re�ƫL$���`^>�b#��4��G״��Q{#J)�O�i*r.v��ED���P��qm��F��kRK��[�����"O�$����6��{��� w�ܴc��c����K2�������HQ젊�N,��@H��j�x�d�O���H6	֭�'�O�$�O���w,���Khv�C��d[hY�O�_窱�e%�'}*�LQ��դr.b>�P�b�>6"j^1� �Qlֿ���jWE܊�8m�Q&�?.��Ajc��#GD� �l^9X��O��htdi�� �`zVg��o+N����D"jz�����ԟ��'����|z���'��(�c	*eήQ�H8F�Z���'�ڤX��(,T���eR=7p�z�'��(��|������ݱJ�*��+p�B ��H¯*�y�d�u�D���ɟx��ӟH�������|J�Z��p�ro��GxVPjdH�\�i8�Ӥ��pGA�>u�
��v��hO`@[�ۇn��������0*U9+����WK��m��0P���3����a�6�Xr� J��������R�'`�1E��ȟ@��t�'бO��`cͽcP 0Oà;O��b"O�(�"��7r�y�"��3=��������TyI��06-�O�6M�C�p�5�֘d�8�`����I��|��Mʟ��I�|:�ۮ^��	���$/hrD��N�'��<�S�N�:�B	a$��$�t-H̞�4�<�R�N�:��P'HY5��-����$�(��Q�~�H���Hs�8!�[OĢ<����D�F���9a���@m �p�	c(�RU���	��b�YD(�l�x�#Ċ�9�Px�Í,�9&	#��+�m[���"�|�ϳTU�7�O��d�|:�	��M���C�<��� ��߱{�z�p�hZ�B�'�t�ڄ���j��s-&�!fIR�{��H�X?��1Ì:i2)U.���V���M �D�5osFe)�!�^\�<H$�C�#�]�5F��� J�B�H#�X�;Rу$��'#�'p����Uɧ�O���*��Z='l\X��"�(R�ЭS�'�J��R�S>?A�;�g�%CB��
�1Q�����J�H��� O x�4�����?���?���r�����?��?�����tH�����j���j�K
����y�úi��\��H�(%�x����N�2��D��\��㋖�Q�^���V1q_�:��\�Һ#�
+2Z	S�i�b��I�5�R,��A�Er^��6&��\d������l�Oё�<��oB�����9�R\Q�` D�`#�4����N&<X�R�.*}��7��|�������j��(1A��}Z̕��/U��T�Ц
8���I͟ �I�9Yw�R�'��J uB��b��8�脰����r�d���0F�"�1� mc4-��IW��A*����!���r^����U�;y)q�o��b��-�
�tq��BjgN�B�%P�v�r�������T:޴[����>�g�ʻZ����M�ez�i���D�<6��jC��bE�+2 Ʉ��j�u曖�'�	�2a@�;��&6R�)�2���##a���c� 1�I��`Pa�Ph�	�|�D'�!�L��ȑZ��-;qm�;-6� ���-�3�0�e���͖f�|�<A��!�Z��0�-<cJ�[�3�=�c�кDV-v�ܽ(���e%���Fy�o]��?IB�i�|��3=�0T��K'Z(��ņ�8K\L�܆��h��� E 54��y���*�>�<���4�^D�gǝ^�TA��D�;�9��A4v��$�<���LIћV�'��V>� f����sn uV\�%n��F�S ��?Q��R�������@�"��lk���v�J�5��9����[�֖"�r�*A�_!f���q��x"fϤp���J��Eg�@J �3e@�x�W�^C���F�U�����H�R@h
de[����� �ɀ��S�|� ��M9;��0��'� ���2�ħJ�!�H|8� Ӯ.�ɇ�� �(O�̡@ Lg�$�� δ2�,*��ܦ��<Q�t���D>$��r�/T�z�� v�S~�'��'`��bG��A@��cKK%
o�T1�'��](e
[� ����DmWQ�+�'P��iV�� *h �Ȅ��/���'�(TI�4	�D�!�d�T�(�'�^���d3@�|��iV�X�(p�'��,���BW��J@�^�U&�2
�'�d�(L4 �*U	��Q���	�'t%��ڬ].d=�����d��'�Q)5��!A�1pp	�ZAP�' �a���ޗbv�h�w\�|�$��'ǼEJ�`�:p�)�	=p�°p�'�X)��0^���D�(n�r���'���H�1�V i�e�V��t�'v~�A�o�_7��;%@�F����'f*,�/ܔ(�@�d�]/<m�5��'B�1
E�,n��{4�X f�tI8�'�d�S�)�`��K��a�r��'��٣A^s��-�&�V�O�����' �\Җ���
!+*b�s!+��	�!�� z9��/m��	;� J8E��y"O��A�ɷ:�P	�웅+��8�t"O�-!�چ=J����,��`�N���"O(0@M��/�P1�K&�vq�S"O�<i�*ն@xV�9g� �ڐ!�"O��� ���-�N�y�͜'�t�%"O��@�~��5���l�04"OHt��*��8�����*+3�ag"O�X �OL�#v��f<(k�"O����WL�ܩ�(�'�D�q"O��P��4��H*)�&I��'���B˩i;h�)t$>i*9��'�������%96h#e`�l��'%rQ ��1tX��7.h�
��'����#�����l�OԢx*
�'w�Ъ�㏞/����H|~Q�
�'��l���V������PgR�S	�'��@��j2J�*ur�k��B��d;�'�X���Ή?n�:c&W;�����'Ѽ��C� ޶IXr(�/?8�*�'�<B�ƒu�|��Qd�6^�(Ѳ�'�:-bR�ظe
2�q��<R�k�'�)�(�>q,4��p�����'d�1���
�
ӫ�#A-�� 	�'1��≜\d�,�fQ,Z\�	�'��D"�E�/_4���w��?,;&��	�'��`"s"�+9����͂�RW��'� �7�C�2��+��GB"�	�'��-����X��b�όh<���'�KgJÌo$<��)�@ʔ+	�'�f��%H�#b%�O��~Aڍ��'cu1f�.[z:�2�	��w&OX�<�i���Ucc�[�{�z$��W�<�Aψ18J4bS�[
$��%񂌅\�<q���SQ�	ׅ��5�xs��]�<!&�V�n�Z��"��u���p(N�<��$:ʨp�s%X�n���X��Hu�<�ˋFs���:yX�
n�<��W�7�
L�vF˙�hГ��LN�<��`e�HE��y.Z�#c�R^�<`�{�40[�␙?������W�<	��A���!�>8LH3��G�<YE��aqh쒤�\.\U�\��@�<A�X;
T�%�p��94�|�<y�k^\�����Y�{*"�3j�v�<�g(|f�,Ч��	n��8��E]�<1��Z0T�Hzs�F,+��r���V�<��ƹ8�i9 ˔�E$B�YV�<Y�EQ8���`�k�>|�P@�d��V�<Y�F��^��r'��>vX$+fC�Q�<��,OGiT�e�4a�Dy�g�T�<�P*�$O̤�rdV����h`��e�<i���"[��'Q��Y�5I�c�<��Q{�Y��+\�WYԸ�v]�<�ƬνC+Ȁ���&�||�'.�Z�<ف��s���֖G�,i*�\�<���Q�FO�{%�ʙS���fJ�Z�<�e��x��[��k�>D�e��Y�<	vn�/�����c�%oD�e
���j�<Y����0����% �%[�l
$�K_�<Qc���	t�p�+��tЈ�+�D�<�c%�f��#uJK�$ۘ)�	I�<�2\+sѦ��e"�9{(%J �G�<i"$+����v��91�^r1�G�<� �`i�Ί��00n�:jș��"OP�+ȟO�B �B-��^MX@ba"O�C�O�b�"��G+�0�YT"OL�fĊ=r8��r�I�T���qq"O� �ԇ��zܱ��ܑLѾ��"O�,�FbłJ�@ e�а8�d`"Ov�*Q/��"+�Y�K��7���
�"O�ͨvC͋	(�T��� A8��"O:�����C��]���
2,P1�C"OPS�	-h
"��b���R���"Otey�o�#,���+����EE����"O|�F�� ��h����U�t5�"O*@�F�]�+��s��ŵg�ryG"O�]C�c��W�|m�7LPf.���"O"�
B3�L����S:X~��j`"O�u82jJ�8���۶�	7:����"O�X�%��C��`YS��:7  ��S"O�!�j�-.����d0L��p�"On���($"x�8u��9'�r�)w"O� �┷"np��������Q"O�@���Tg��P�+�;l޴�"O��A�i�_0-рJ.f��I�"ON�sjǹ]Z��3UG�5Jz�T"O���D.p
ԥ�2S/`j�"O��8�)^$7��I�Ɣ�v�V)QU"Ob�pFI��
������\�����"Op�!����lErk��y�5#3"Oȹ�p�C�,{n���?Pn�$H�"O�U���;x,i{U#�'R��"O`�K�o@8"]�����ۿL��2f"O^M3Tl�8x�`��d;1l����"O��)��
O2uHd�FS��yQ"O�d�5��4����@/VJ�Qq�"ON	�h�E�dD�w�zFeZg"O��y�@'1�,���,1�)4"Ovը'oV2�f�ǭԟ/���1�"OPP�#�1~  ah�
�Z�/X!�d!d��h�`$X�
�0�D.k!�$M"j�ź�'Ȥ^]�up��C�LT!��4�d)C��DT:��2BWDE!�$��,�ʰR!ʕI���;!�D�&H�@�Q���4�씁��25!򄇿<w����£M�.T�f%ۄE�!��'*5���!�la�EEV%}�!��.,`Ѕ���E�*��� j�(S�!�$�@��H�th��P}���H|!�$���qw��6n��Yu��Yb!򤜢n���5�7m��-�CHY�U!�$Y�F�VM�u�]��dp���+X�!���k�NM�%��
Z`��M�{�!�T�sI|�jb,%:�v4��fW�J�!�dݐ�>H�vi�H���w�L.l!���K(���wE�$h���!�>U!�A��i� �L�0��A�q?!�d�57.���
%9��P6���s�!�$
'�NIP�ӀT��P0`�>�!�$4qbƨÔB�F�p���V!��[������ƽb����o��!�d�3,��4���V�F��r/�2H�!�D�[M�R��(�PX��'�
�!�ĉC����@�P?}H�xňF!�D֡��[��:�ՠ�).!�$�3J� �@p��t8�}p2jN?s!�
�{��S�e��]#���ꆄ6!�� n�S��
e�l���&ƥy<(�y�"OHA�g��!->���qe�#��@��"O �[��	?��u�H�q�R�q�"O
p�pe��s;�r��&v�2��"O�Y�s�h]Y1�]9BY�@"ON�
w�ƓsV~ȱ���:�� �"O 5��߯l��xKbD߭57�8%"O*�8n�q��%�!Q1�41�"OT�ô��[[Jg�
L����"O:{�	Y�Tt��.�(
��]+�"O>(2���^�RD�Q�/y�D	�"O�4D�!"=&�Sa�Ӌ;����"ODd� �лsSzQ7��W���k�"Ot51VJњw��U�V��+�N��"O6�8�'�>j�v)I)L�%��EpG"O�t�EXN�-�F]����"O���&eB-3�T1`#&Ӹ%j�\�7"O�)U���P{|�zT�
�L`9R�"Oc��b�t}JS�F�S<��"OZ�^�8���2;/6�p��I�!�ʝZ�I��+B�7}�0�A���!򄚩o�0�{��Tf°�T�I!�E�4����X�/ ��8�dO�5�!����
Ēŉ�T��	�@�*>�!�ño�X9#�+X�g�ĸ�"�Y�!�˜H�$��ҡٲ��p@�F�5�!�df2���G�K8Ja&�XT��n�!�T�d2lٓ�+Į>��EY�L�#z!���Ej8��^��8ZGEީ`!��I�W#)��P1 i���CP#W!�d��R���狃PLJ���cR!��1�p��s��1=�K�횧p8!��Ҫ.\�C(��q�ש�w,!��ȁ
ϊ� �"y�1�p�N�1#!�ӹFb�{%I7b�}����
.!��Ͱ8^H� �J�Q���K��ٱT!�d\'*�z�S���2?���� J�7'�!�d�Zy��ycF���(�H�K�!�O�x�����$J3D�2��E9&A!�2�43��	� @T`!!:!򄘰��Z @�[@0���G%;'!��=�����##D��CS�ۂ:=!����~���AB+�]��>-!�$�%S�o�[�ÂL��&)!���7֑�W����R��8�!�`�!@cĬ^8�5� 12!򄗉z���$�C,+��rG�=2!�N��`�s-N=]k����	�v!�dK0ٺy#��q�R�Z���d�!�$L0:e��0�f��| ��D.G5wB�Q��s(�y�e
�o����$��n�6���GK�!���	�ɑ�(u!��%{"����پ	���i7I�2-	!�!LR
�F�4��Ȁu(A;^!�]�g|���B@RJ:Zy���S�#q!�$і�N�QÃ�B¬yV���xY!�ė#k�P%��A[�'`��
Y!��S,�б�M�[Ѐ�O��w_!���2J�衳�՝:��Ј�E�'Fd!�C[~~9�E��5
��i1�JG$!�d��h�Pu�G�8��I��jL�Lv!򄐎߶q�ǮJ�I�&eC���,|!��-� aڥkT�;��ato	7Af!�A's��AoNQb��F�[�!��;~�	�V�D�,`�kYr�!�� d�Q���$Hv����Ҕ��%�p"Ot�`�-�"�(��+�Y���s"Ora���c�IR�6<�Frd"O����oփ*0�#��׃�ʱ�U"O�G���X�8$޳3weQq"O�|����8��dp&
����"O$�kr.̫�	�N�"a3�"O��EcJ)-��-H����)("O(��͋� ��R5l��	��E��"O���bC�;��E ���S"O��p��X>_�)��N���<��"O����F�� �ek�C�"O�0B&#~��i��ԼUTK5"O��HP�Z�cW�LJ���YR���F"O\T8qIK@jh��kԘV�T|[�"O~���ʰ��Es�/L�_-�=`�"O���E�O������>`�(4"OBј���yAD�
���d�B�	�"O�E2���t��x��$��@h>�h�"O�mj��2.�YPn��tIvT�"OT�pf��f������3<���"O ʳI�
@-�l���ݧqVD8�"O�-p��J/Yj�-aV��MN(1Z�"Ol�H�N�-�}q��kNpd�2"O֌{f-ޡ\��t*�l�(fO��*"O��sP�4P�죷�IE�)��"OܰKdd�T4����ȔO�v� �"O|Dcq�N%H�`"Tb$5��Pؗ"O@��kЀ�@�WB[}�t�P"O�� �
BsD���!w��t"O�|˗�O���e�~����"O�hç`L�cw�)*p���I�TT{u"O�E�#�ľ+O�M@�͸_�6�*U"O8�� �/Ji\CBK
R1z�
�"O\E��M"�q���p���b5"OR�r�ڪ��p�B*"���[0"O�����+A���KA��u�p=�"Od@��%D?���§ƣe%XY��"O
m�PB&<��-��%�R����"O�0��ҥx8��q�� :xA�"O�M��-�j���p��у{�ʨ{r"O�L��靆-�b��\�q���I�"O\�۲#��Bc�*�Z�N�,��"O������z$b]`��B:�]�R"O,�x�N4B��t0�(i ���P"O��)�[�l��B���/	a��k�"O��ڑ�C'�԰c(��n�	��"O��V�0�n�:sR|*�A"O�yF��/���xF/!�p=B�"OJus  M�(��D�[�2���"O�]	�9$�I��[�)�T"O*��U�K�L%�UH@*Ex@�S�"O�H��Y�$���t���Cj��Sr"O^��� ��1��CGT�-��"O&|"!�\���'e���ж"O����Ӧ0zm�E�N�r.ͱ�"O�يe�J+6�.����B�@���ȓ"ON��å�pDy��FJ��\KW"Op=S'��!��yA2��Z��)�d"Op�����!_RF,��CY&3�Tq��"O(��nE��U"����ȑ��p�<	��]4��5�?D)����I�<�������(Ҳ�8c�vMi���C�<Yࡍ�*rH��K����DI!��B�)� r����(��,�%��)��=��"O��!F�@<4	m��É�\��"O�|��&[�\��$5:�h*�"O��g��L�d���PvĜȗ"O�I����]�����R06;� $"O�|�BX$E�m+�L�0W8�*�"O��W䪵+C�B�w<���P"O���o�	1�U�v �?J�Qcc"O\�)ab�R\3种xf�"O�H�B�W�b��,ʴ�r0��w"O�"3���F))���-P_� B�"O�u�e�����	>&�6�k�J��y"�E�z̪Ys$��0"�I8�G���y"n$|��EU`�,:�å��1�y�NV>	�B �kJ�y>2��DA ��y��e�mz���$)e`����]$�y�MŲ�P�1�
.l���ɑ�\
�y�F��f�!!J�c^qZ�,��y����.:��� ���Ќ����0�y��P1�D=�#B��W(i[V�I��y��Z#t��9 R$�ر�%S��yiЦ6���i�8~ހhƎ�7�y�l[+�&�C���fl` qA!L.�y�Ƒ7g����b�_�Lg�YR`7�y�KZ/�j�RP
H�|���{�%ѽ�y傒v�Ll�3��)����G���yW3*x��0�!��!jv���y�C�V,�ˡhL7Zx����E��y2-�;�Z@p1D�9Q �)B�y#C���娈&1�(s�]��y��J8n��r4G�* T�-�4m���y��>Db��Ƃ��-~򕚔��y�]�(Up��Ã��,�D�	$�M��y�Oԁ#	�!� ��%&U~�3���;�yb��Z:6	:��'lǪ�!V���y�I�D���0��0s.��q���y�*�0�x�#,�D!E��y/�9���p���"8��� �A��y�`	 ۈ�c��6��t��h�>�y �	vQRm�B��� ���*w�+�y� �gB���������k@�y�F:�]b"�޻k�(�r��	�y��W��b��u�O�d��,M��y�N�?�2�#�D��`��-���y2
I)Q���5Ý�|��,"5�-�y)�:a�MY�4&\�qQ�N�yra'	�%
��'x@=����yb��|��iӃ��Q�Ԩ6 5�yR�	,Z���"$\�W�t;ƍF��y��{$x�Z!�Y"KQ9�R�K��yB�E�R�Q���G r��@��@"�yb�Zl�̰���m�U���F"�y�K	�D٪Iw_4k���0+ �y�OZP\Y��h�$m8�}!#��Py��K�^y���,�
lRLa i�e�<�d�$�����  і��T���<y� �f䱕,�>}~����z�<�wg�X�\`�&W�\�Q�6��s�<�S-
+$�p�y�C�s��
p�t�<I���>9a��ZĂ]mH�]j�)�M�<Q����o"�r���m��Q�2^c�<�Ũhj���V�*��H�[b�<)#I��f`"!�+j��d�'�{�<9�G1)���vȆX0�[4��y�<� ��*ĠĤf�*�qV@�0�<��"O��B(�k��5&U�I?,��"O���,�hZf��6o�136���"O>	���� x�XfΖ�v�*���"O���4�^�
����bY�X�Z���"O�+PF7VB�J�@�d��I�U"Ob���Y�nL� z������C�"O,��nA�$a�b% E�3���"O�ȫF�iE� ��ٿ�mQ�"O����P	G8TX{�F˟`m���"O�L��!5-��l<I B"OҭpQ���9<�t� nD�|L�a�"O�z��R?2Y���%��1�"OF��0�%I�~�T�ޒ2�T¡"O �BK�9= �A��jY]�^��"O�� ˏA6Pl��F�p,>䫰"O��"�M�6�P��	�W�L�s"O�P�Q��4@��px��Mf�DpV"O֬�D ��<Ed��R� =�\ɰd"ONЂŧ��"UٳiI�L5���g"Of�{��G
LGj�ch����r"OTM`�"�(�̫�n ���c"O��)B��*Ԝ�UnϟKЁ�"O�Ű�΅�8���t�\8z��<��"O�!�p$� ~ܼA���e�,�0S"Oh��#�G�~Y@��] G�� �"O$��v��,
r�`�H	"6 .�"�"O��"�$@+�q�v	޼#�����"Oڍ���"�th8	ȧ �^��"O�
�MM�#`$��	i�vAa"O~u��/�_��U��M2k���l6D�t[a�W�&���CW�D$Q��ф(D���N��B� A����!��IƬ6D�d�EJ�<|�9�fm@�d^�x!��3D�t���۪��Y4��w��k�o<D��@QC��d�&廄-�x�Ջ�:D��
��S���
rI��%���a��9D��R�O'Y��I��˜0�4����'D�h	E�'
A<U�V��KT0��!!D���*Ƶ>s�a��4]�.\XSF2D�,�P�T:A��Q��"Ue�$���J?D�Xbq$�p;��I� �u�x[p� D��B��_�E��S
�q��ద� D�@&۶ �0��@1,��]�b.D��Z�e�VͰ�'LϜk�Bl+D�Th3
1I8�98m�Ml@��">D���F�e���3�hՑm[���Bc(D��bU��v��ěNU�AǸ�ۓ�"D�`�B[7A �����:x*�%D�@�cO�/OB�Rgӏt�$4;�g$D���EIӏ���Q��R�EP�p�-#D�LK�k*z��l9�L��^X�a��!D��(T	0B�ι��H�T\b0�-D���3J���p #�:RqP�ę�������'r"���%Wx�0;�6w�]�P�7�UK$�"D�$GLԡ7�$DY�B��O�zG;D���F��A���a�>͊���.D��r+^=Q���	�-�\�б�*D���d��̺�5�;'�@���)D���������5���/����#D�4�򭒙wꀴZT_���6�%D��{B���
�"�K��:ϴ塷c"D���o�a���Iw��_W�Ց�" D����N�8���w���t����3D�� J��V"§.<B�I�hMc�r5{�"OF4�0�P*'X�J�ڈ�Hщ�"O��i�#�V�>}��0nA��$"O����ˎ{f�`m��y��%��"O���FhN�4w�Pڕ��8����"O6e)5BN p8n��fH����Ԑ"O�0Ht�8�ba;�fL�<�
�%"O���GK�:m�`�Ȃ�>684��"O�%v6�ؔR�a�&;ӆ���"OVlKc��5PH����+�B��"Ouqf��%'��ʒI�t�h9:�"O���`׷�v����Z<W�T堥"Ojt�%���5�H)��"Oj >!!�(Sxl)�Ԅ_E*����DF60!�]�!�$�(s,[����Ã�-!�DS�Z�ih�Őe0�@	)x!�$� �d�A���1��E��!�D+#���`�Ju���&�g�!򤞾;\�b�:Ď=���  |!��ۻ	>,P��1��9��f@ac!���l�bE����0kI� �Ä#x2!�ē�k�d�q�ɑuC��㥃�!�d&	F�BE
�2�BC�q	!�DǘYbBE�	�%M�(�ՁU�s!�$Z<R��������P�X󦇂\!�ӡf~��{Ɍlա�唳b�!��ׂwt��&���)�*��.�!�Dذ?�Ѣ�@,[��\����$
!�-3��B��/W�����F!�wr�H�e�t�f���@EIU!��F���U���- x��MJIt!�Њ-3�)$"�m��d`a��bh!�H(W��񋜴 �(x�#�M!���5MXLu)�����y���ŕ1 !��_A$̸��!Jq�AK��7)!�dH�,��G�Z�^}2%�P(�G�!�G,����*��0��� On�!���#0�NQ�@�ǿ oHݠ7�$Bm!�d �"$��l�� �� ����_!��A%Wɞ�*E��e��;��
|V!�ǜX֜Աa��,vن$SC��� �!���g��s��G���%$�!���a�aa�RN��D��m�!�:0,|�Ve��m�@=����f�!�D���� ��1V�4ҷ��h!��X�>��Ԋ�0$�8`��$�!�D�4C-��|��
�!F�;!�A1\�^�in
2���'�<�!������ҞK�B�`5G�e>!�dƪ_�0�b��;hwZ �E#0R=!�";�9����4�6�I,�7 !�$ślx4��EQN�\r��  !��|ѡ1 �v7�q��Y�p	!�ĉ��T ���Y�/4d�k�Y1
�!�Ȯ8)T4��"r��dqgE߾c�!��I",\(� -��qb���!��6%Wx�a׃� }nT9Q��Z�!�!��?>��G�Y�m_ �ԈF?q!��xkBFٺ^p��e��=}Q!�*CW!��!�#|�V�9 X5�!�Dɥr{z쒥 ���`P��f�*P4!�d�79���w,��k��p�	�P�!�D�O�=�DC].R��:�č� 5J��W"O
�4V�C�%)���"O� ���p%^�h��G�ӱ�Ta��"O�����V�<�1eJ�b���"O24�Μ"C��I!D�
Q2�83"O�a�!G}�n�l�x;|\xa"O���" GؘS"�0)�L�'"O�X	 7'_X���AG �ah$"O��f�M}b�B%;> J�Q0"O� K^�)7�X���/Y��a"O�D�v�Ƈ8�Hq|=&��d"OZ�#���^����.YhT:�"OH��0_��Cî�-b~�""O��07�ݫ�D-���0|2d�"O��P�-��%⋔5J|��"O�ɧv�t��Q�DLU���"O&�@���%6��<�F�h4Y�B"O��h���Cd8urA/�w\p2"Oʵ���X�`'��CwkS�B|T�C"O�|4�+xᎅ���M>]&x��"O��:" ��v�
�R��*�칸&"O�� ,����q�T�'�V�1�"O��ڦ�K>�}"���' ���"Oαs��EhHHQ�a��H���@�"O��� @e�xd��JS#t���"O����,�9F�"��-˨	�"O�!�3p����2�ǀ�1"O<�Z� 6lZl�"�+պ8V����"O� �B̢�,HkVAk�]B�"O}
�'�k���c�*�ڈK�"O�����K�`Mz�H[�b��"O��!��k �`QH	q�(��u"O��""[�MX�q�T&�p�Ӂ"O�-�C���4t��Jۜ-�Z��d"O4��' �FƄ$@�DX`�t�j�"OQ�C��&��`r�E+H>���"O(�n�,R�����P�R��c"O�t�����qI��u�����Y�""O2��#hߩq/��Xv�z�� ��"O�Ͳ@� �'֐i�Ë�$�L�1"OJ�b��;��A��ڱ+�x�b"O�2Ƙ���8䊈	����p"O,�� g����Q#Jғ	�V��1"OB������g�n��ע\�4�b1)�"O|�Åo_1� W��YCT��"Ota�v�Mo'B�!�	�.7����"OͲA�/N��U� ���FL�-�"O�"@� >H*�t�!h�^�	� "O����/��<^`!#�1u�m�C"O��
������)BR���k�D��"O��£_�9�&�0'�&"S�lj�"Ot�z�)��l���ݯ2��@�"O ЃuO��:�&��ŉ�q�t���"O��Zsj�W4։v�U�<$�"O�����D�p����!\�G����f"O���Gb��TS�	�
��i�"Oh�bƃG*t�F��'�ؠ w�!��"O.X	�[����EڏdB`ڱ"O��@��Bs�H҂I�Va|���"O@x�F�KmLA�FBe��hk�"O����6�4�a��G����"O)9R�,(�#S��$A��Q�"OH��5LͩD�ff��(p���
�"O���:f����m��=�|Щ "O��� "����1��L�2����"O<1P�� �n�	�U�~u�@t"O� t��,U?;Z���Ǥ!j���"OR8{��\.^M�7��}+���"O��B� FR0�SgN,b�@y�"O��j�;E*�a�C�H���S"O1�&��8@G�I<�3P�L s!�dI�0�J�`�Z;k[tP��d��{�!�ĈJ���'B�B�@�QC>�!��Z�P�|��Wm�\喑��=^�!�D�!�d�j�L��Zh�ac�)]!�D�g��0�4)C*=�#�Z?R!�L�EV  r��
5<���n>!�J�/���Gl�[����+!�D#93H�􌇼y�`�����2H!��Tm���O�cԐd�c� ?X2!��9M��[�,E�v-�Bѣu(!�ܨyD蕆����<�/N$�!�Ąv��=)��3J�j!��"<�!���"c�m���%�D,��ˀ�)!�¹9�@��IU�X� ��Ą\�j�!�䄠+�>�1D�g�谤��%�!�D[ B���(��&T�³h�PyB��3���ڐm� $�j�1����y�m�z��Eaʫ#!�L�JK�y2)C-�R%����� �R8�I��yb�חh_�4㷇�$ �`�b��À�yn�7c�8ro�@����y���#�>T)�G�'��d��Y��y��37��!��&4�"���yRa^�c��iE �)��2A����y���3lI�fė)�����C]%�y2��.
�~��H�#p�H��ƕ�y�IL�X+��J󢗪hZ�У��&�y��K�y�πIp�
4h���y����oҴ���2<w�!#S ՝�ybm"�i���'�����J�*�yR���n�����/��N���@��y�@��4�L���sOj������y��.��5���Y>G ��ᘼ�y*��I�t`9G؝2�=�!�ǲ�yBg�rfܳ�$��u�^T�tȓ�y�5�L��#B�n ��9$�B�y��U�xܞ�YB	ѽa���Sj���y��#-'���K�\&�\�P�R��yb��Mv�@B�[�z �Sk�*�y��-~��� �
��b���L��y"�B�nKJ�%�C4&Z5�aĻ�y�JF8g]�uA�L��M�Ib�:�y���G�p�+kAz��P�H��yBM�i��E�����Fgڰ�d��yR�C�
8� �F�m�dtZ���y"B8M%4}�`H�7_�zh�Ak\��y��Q*��1³��7)��Z�����y��A�4!��c΅��̲����y��ҫ�|�җfJXx��d��y)�y)j��B�X�
��80e(��y�´u� �E	W\���%���y�fѸj@-Z��J%2��!�E��y��� u��k���f���JH��y���(�F�������r���y��2J��I�� � ��a5']�y�D�5S] ��#E�-�*�IS'�9�y��#��l�"j��HE+�/ ��yb��?O"���g�ʘb� 	�yRΌ&��!�g��%��8�f�-�y
�  I:�.4R�X�
P3ֈ�"O�Ļ�*K�?��I)�`Ą%��|Q�"O䅘W��0(�z(i���5:FDq��"O��S�L��+L�\��E��M2�-IG"O�@�2Ϟk���Qr�I$;8�C�"O�<��N	jlz9"A�V��P"O����Ka�Dh�`M�ox�9�"Or$���=D`�ٱ�B?8\��0�"O̴)��͂�`�Y3/��RL:�{f"O�m���	�]yv훕� �%HA��"O𥻔c:Hޖ��3JԴM1��;�"O$�3H�-�d�J"�ɺD^1*�"OL��H�VB��JR눆>�>��"O�Ey�#��l6��l��JQ"O��!��?*�չ�m�"R�� �"O8U�!FY?S�7 �9&"HH��/D�<zG��T��I�D��8����(D�H���ST���		��C�B\��9D�\إ��7'�I�S�8d��`֯7D���V
�'�&욥kK?^ �02F�?D� @J�[Z��cF?x4��?D�z�f�]��=���;t�ґ&/D�y�O-g�d5ڔ�H  P�*q9D� M7q�0�
%�X��p��8D��"��ψ(
`Ta�N�Z(0ql5D���� 	S��D"&H-!7��C2D��
��3'�(:�2o֬Mk�>D���=gfy����Y�v��R�:D��Rf��j�XM�ģ�,7�i
C�3D�0���_�Z��`
�B�)��3(/D��k/0��49�L/���E�.D�8:6D�8q4܍�ʌ�E��L�gj1D���m��y�����ʉ!���)D�hSS�Ń''�}�5,��?����(,D�@4+ߢTwT��̆)XvM��6D��0�.C,nU`�x�������3D�L�V���n��;���R'Qʁ�2D�x�� &0�8�@�R1J���BŃ2D�Ԩg��NV#�N&H���6�2D�D��ȴU("؛�i�"J��8c k4D���E%�j���C�M�1&(���3D� h���Cq�L�!��K��H��n,D���C�\yJ�N/g� G�,D�� �Q/p<�(�JǔV��R'D�T1�c�7y|��
�́�~1��2"$D���£Ӫ9�XH��A]D�<�(á6D�4��//,6d(�,���Xm��*O�]+�m�/X������-�2��"Of���/OU����?B�k2"O��e��;�h�K��Z���0&"Od�Z2�� R�iR'��5�e�"O���tM߿6���pe��Pf"O���Ԏݚ)rU��T�&��YiW"O��`E؇U#b��
��lj��zD"O
�arn(��9�hJt�EP�"O��Kv��*H�j!�xx��"O>�V�����rG�3m�Z4"O�̳T�V�<Q�l�%�	2v]�u��"Od�� �Ӈ_�v�3b�E0d;�"O��Q���'���`��2#�]�"O����C�v�x ���?L9��"O.��������ͱЯ�?��4�"O���f�q�����n �s�^Abp"OH��J,b򔼚l�A����"O� �;�gH/}\�4��� {u�D!q"OPhX�H˵]d�g��n���"O��$�6W.��<U.U�p"OT�0�
�,>, ����#*\��"O�I;�ϰ#,��y�d��t"\XA"OV���'Ӏ>h�٪�/"a�H�"O� �b냝���3�[�iKR�"O��l��H�j�:��БgD8�!"Of�Pk��+*,�(f�؁?|;�"O Pj�K�2n:H��� ��2"O�)w	^�TJ���MQ(p��1���'*��Pq�$F(�ҨZdn�b�|�xrd7D�d5��PH�$���X:�2D�hY���Ja8d� O�;sVd[Ҧ2D�<��h�J���Ff&r%�-D��R�3K�n F�TUg��Q4`-D�hqIP�=�8��d��=zȑ )&D�sEC��\ �Q�-��0�'%D�8���O�J�"�x��S�����T�/D��Yw(B�0n���v�T�� �?D����Y�2>�<(�
<H@T	��
;D�8B��K?���S�%��Q�5D�$�B�1u��(RM
L���n2D��y�^�Xp#@�?C���P��0D���d�*l���A�kG�!����&�#D�|�A#_=*��2��F�Qn]S�%,D��B��f��%e`ʬ�Thi(D������ ���<IF�� +D��G��Z��� "Q;&/ޅ��m(D�ИC�W���{���jD���J%D���fJ�.?�Uӗe�w�x�!��/D�L���έh2��bk0�����#-D�tP���J�ٺ�n<g'\�)D�d^���-�Sb�����b*B�I;���X���̺�`�B	$B�I2��p����T�n� g���g��C�I��"X� ԫ?8@�KB�C�	�:|��Y���y4Ј'��y�LB䉲gR�ǝ�jT�X�4/ �3<B�I���)HFI<zΌp3l]�	cB�ɢ\��191H��b������aB�I�92M��ěZ��\�`#��C�I�e�y����7!�H|���R,&%�C�		�<{�O9~����@*D��C�ZN���߸z�*$��>��ÁO�E�O�#h*y�$ �h� �+��'ױO"M�^J\�@'.P҆5c"O&dR��oD����3�"A[T�x�-ȡ�O��,<h���,bn���O�@1ʲ"O�2"	�t���(�f��M��"O����D�+6h8�p	�:'q�T#"O�)C�4@閍e"A�GU�ѫ /_UH<A��ͥQڌ}J����}Yg��'��G�'^* �Ja,E�H��'պo����=� �H�x�W�5e���'�#=E�4��0����JU�`<��Y��ۖ�yrLL�nˀ��CF	Oْ݀���,��>�"�'��H�&ؐck:�X��9��T���Q��$ƗW��Q�c׾@j��A#�p�!�8�� x��ڪ7V0�SaE둟ti�Ӧz|H|
eKI�A�@	qwȀ:��C�ɎD�ʌ*�GD8�F��`DK�B�8?Y����	) hA�U�݊oP�(�U�G�h�FB�ɶKjV<��� p����rh B�)� 8@�,�;�|d+�AĊ�"O�|�R�ڒ=�tE�0��1�rP��"O��r � *�0�"�&X����6"O���3�jLV�����A���D"O& P&,��[�Z�

Xw���"O2ę��іi�X\c����Ѕ��"Oʔ��J�u\� �3��+j� ��"OXee���R�c��<F�7"OV[�)�i�zx�0�Y	&�(�"Ota"*�*o��E]�Y��d�2"O����]7=�l�� (�ux�@)�"O�V�9o��!#'ѽ0���"O�5#�KA�%�ڵ��F�P��:r"O�9�A.??���"����U���  "O�q � ܙ�&���-����s"O�\�`�U�P�z�z�	���H�"OZh�6��%T��2��#J���T"OlxHq��)F�
�+���\3�P�g"O.�
e�F�̥!�@#B�9�"O����(O�L0b�U6�e["O�ȩg��^0@suΝ:O���8�"O�Hq���R����N��@�	�"Ox�hBɀ6*i D��n K�0��C"O>d�W��7/�,����E�l���"O���e#W�2��9+��8Q$�0��"O�r�FT(4����k�w��"Ohy�`� !-lqF���Vp�Zf"O��)R�����@B�
��Y�c"O�G��md��p�J%k�x���"O�D����9R�
E�_8){��"O��zPER�������kr��V"O`�b1 �'�rp�r��0ʪ��"O"̡$eG��i��K�A����1"Op���	C
W��l��B�I�C�"O��w�*��XKu�P1"G��4"O�@��[/���TcO�86�d+�"O>�fN�*�� .c��I�'"OrQ�V��
� �7d�AȚa��"OHZ� ��I�R�
$��.��yE"O8 �F�~���7ǀҦ5*�"OH��� Ѕs]�T[3�=1S����"O��;I� K��4��#�^H��t"O�|҄M͡#VH�"I�NJ䭱�"On@���0p���J�H]�!F؉z�"O$�S���9Q2ԫ�AX'7�r�{�"O���+}��a@>f,5�"O�Ie���0LA4(�k-bx�"O`�jB / ��8ɑf�73t��"O����ީ�a�@�"�u�"O�:�o]�3�~�I%�3g<|��"O�\iP�@%���˱MW ���"OP���h��2�L��V>���A"O:X(�ǔlRqb�U�g1YB"O����虝Y�t�
�-V�*oj�p�"O�����2vq�Rկnfp���"O��s��.c��9���bQ���"OT��3J��c��PaT/ �)´`�"O����	 ����E?;�=I%"ON�@�U�j/�XpU��9M�|��"O�Y ���'\��da��|�&�3b"Or�aVLT)'�E�`��+�\�zP"O��EH�`�*My�	/<�hI���O�y��L[��M����M[�R>�s�l�T��æ�a� X,_�����V'?f~9��*	�nK\�&	�0F0���`f��1�FtP��4e�(1�.�b��{�E�Gѻv����k	z�t�$@g��s�g¾>>����]���3��;E~����\� ֜��!�!c�8���C�~K
Y���i�2$��>|��b�<�Sm��M[E�%~�lJ��"��'LWm?a����>9�oד��ÊFNs��b��mܓ�?	"�i�r7-3�Ľ~���4����2@$���!
���'1�%b�hF5^��'T�':��ş�oZ4��xq'� 9#Xqs�#�0`8^�;��,U�]r3��V`�b��U��rÖ=J��'�¶��s=�|�`O�6��y�iݠE(�Z�a�&	�a�P&u��?+��)��&���"pxd��%�O�L���if����I,p|&��Q��QK<���?�OP�j�n!��� E
�6��Q�O����u�@��n�w�|D������f�Y�D��M�þiZ�'��SGy���P�c%LN!~��]�7X�rIVuZE
�P���'���'H^	�'�?��$��+sn��S�m�vfǸO�,a��GZލ���@�D*�dŏ3�A�7Ps�'`�V�	s0l��$�|���㳊I6k0�R`�v��`���&.�Z�  ��j�' ڬ���r���J����eh��q��:P�¼�թo��6m�OH��?�*� =*��ߒ.B&5�s��"'V���"Op3�ǁ�\]L]��W=DP^E�`����4;5�&X��!�$�=��D�O�'}��۲�97E>=B!m��D�E��˔ +���'��hوOܤ�*L�%H���r�ؖ~�����`�8 �5C
���9)�(A�.�H��2�"sd|���]�i�z�z� �ZP�T�O�^0P�c .+e�$aC�J�d`(��D�Y��k�Of7��OL�J[P���� 7�*��D+F�k��|���+��O�,�矌1�E�<��]Bw��:v{�*��'�O&mZ9�M�ߴK��,���;J���-��k����: ���P�i��'��S-f��9�����o��B-�GÖJ���9U��Wa�	�Y)3Z���,i����G��;����3�N����� ֘QI(�0��D�rqJ���)7+6��F�CS*j��%�@�cN4;A`Ee0$�>�X�Y�j�c��Qn�/�)>16׭y��Ij�b������i��Iv�L�G݀�7�%K��9��'W"�'k�	� �ةए%Gݞy�HN7z���$�ɂ�M#��i��'������K�*m�FmBvN(AL����d@ȟ��I�{0���#���������/�u��'
�v㉮���#6[ N
���F�E����5X&xI(����"m��r��Ĕ�I]�~���f /G�0��aOA�?k$yT�@&^i��cDK	��+���L����8ijh��Ey"`J�y�Nݡ���"$BHr��X����-4��	r��h$�X�	�8�'��K$/`��`1��-p�H$9I�h��ɐV��0C ]��!�f��u�L�V�i�~6�7���*��0�dc�r�� �  �(   �  t  �  �"  >)  �/  �5  F<  �<   Ĵ���	����Zv�
�<@�h8�	gz0Xj�J�=r��	�O�{�`�@-7��!:7�� 2d01G]G(!�#��Rb5x�͒� �b�P��j{r�a��܃;�ޅ�S/����9Ge��p_����8��ָETP!0fB)�բ�NPP�x�����4q�i�d'[(@�<%�U?Jt�(RĘ�QJ��U�Xs���Z�@K�XaQ�����y�KX�-�T��eb�&n:pa/�!��ep2���q=�E��N��T��bH-�(`8��ȿO�)J���d�v��u,\�pHd$"p#�F�X���<!�:1���?���?q�'�?!r��Pƪu����i���ʚ	+8|x��>yO�ة��Ė�칙!V>�P�a�^�_��A�l_tPeX�1<��!�c�$��18��U�BA��¢MSz��搜`v1O��8i��n�Ѐ�D�]�J�Re�\��Z��ON�D>ړ�~�o�4��1J���i���RV�W:�y���&�a;�s�t41�ʱ�MA�i>e�	\y�ȝ�l�t�w�`�	e}��3f�G:�f��g�'�B�'���x���I���'<z089�j�/����_��A�g�SV�\Q�.�	|���lT�6$�r�'ʓDV��Pu�F
nDZ�i[�D�����+�P�Hm	&FJ,,�t�ї�đ^� �IVH9�g��u�I�%>�� ƕ��䵊����_lؕ�'Iڴ��� ���ɓH��"޲-���(O������\��`��R'T�`�4��tb��i���'���",�0EZ�b��Oh"%	���M+�F�9N@R�'a��r�(-�ƍ�]��C�@�>�VdH��bޔⲩ�9n�E��%�#@�P�ъ���(ӱKP+	�F#�:v�P|�a� !�^��E&�����sS'�;tg��a������N1�'ª�Э�2J�a9�&\�����Pܞ�)"	�YYdHp�&^p�̇�	����
�� �'gC�v'����-�( ��	�ei�3ٴ�?����)ʔ"8�D�O�h���,'qHM)�/ήj�|��NǦ����)K�}�V�K�y�6���]�j  @ӡ�\�'XX���ޥL9*��%�U��(*���2��t��ol|0fj6 f�8*P��8xV��>�!�˒7(�F�:�	*D�-��N�ğd���OP�&�"~�flÜ}�*D��Z�M�Z�Y�/���y�($˪��/04T(�%�HO>�G�
I0]E���dm��)^�PQ�S�S��7M�O*��ĕDrDK���O����Oh����N���L�Qo���}kq���3�H �I�+��][qn�0�)@�酖p�哠I����<AX $:��*�ׄf�z�Ca�5T�C���#�vm�L�$�D�O��/1O��h���+l(��8�_=y�
���U�����O���<ړ�~�A�s`�A�̜!}� �3����y�)�(�рE�^�n<;����M���i>��Iby�c���Pكh�/&�^5�e�3w�<i��O
;���'B�'B�֝����	�|�Vϖ	#tp�� ǂ'=�Z`;��;z�&ܳ��@2Rr���kK��fڴk Of֢<���@+R�P3�č7���(۸r��ɹ�أO��1`
^�9�`A*���T=Z��o���?aV�΅B�����Mqm��S�A�S�!�@�K�^$�wLE� Z�B�OR� �!�D�3'~���^���bu(C)q�^1��OR nl�I&N�� �4�?������N4)���@+S�����*"�MkcB��?1���?�4��&`�@V�X�c���xP�X�x������0|˴��O�>|p	�ȉ&�Fy���0N�P}��IU���D
�	!a��b$
��u��AUiS�Xq>���̗.w�Eyb`��?Ya��	K����#Y��Ѝ� M�C��Ycx<�Ңٷ_�:�)�hS�R���Y~�Dǔ9&�i���
I��D9���Ď�<JHl�֟�	E�t�=0Z�'3�@��f׆oע�Ѫ
J�S�Lb���3kV4N ��CЧ�0@I����E�:�F�
�5��.[�p2�N߶�~����lhx�ɶt�<mk�J=�N탵��o���C�Α,H�q�89h�)�#G2���+;l���l�O|(rD�'���O?�@g��vׂ0CRc;e�0�XQJ�s�<���!�$��4�����n�p�'�x"2��Z�h�����X�����?a���?!f�C�rxi���?���?��'�~G��-=ІL �e�6
[0�H�)��Y��r�k�[^)�cĚ�G��]�.���x�B
�ēu_(��6M�Li��-]?@�c�u;��ۄ��,�"I�$�m���2aڞ$&�,su� -����G�X���aͳ<�ߟx3ӓ�>p!�Zg�Z9S��Y`�e�ȓ=' ���Ο�@Y�dk�M�{�|nڻ�HO��?���:AK<�B�C�K�zl�@D�4 �B$��
S2���Oz�$�O`��;�?9�����L�4jp4��k����tA�Q^佊�a�4_n&����1LC��P�ӫRtX�Fy2cH4mn��Ĵ��ԛ�@�kw|E�g�D>tD xċ�Y�D��ZC_�\Fy���%�?QW͝�&"���V%؅�&�铎�0bJ!�d��b|�L����k��p��f�!�d/ �� �
Ҏ �ڥ1
Y�l��ɶ�MH>a����jӛ��'\ٟxl�t ���]���
�t��f�i*��"�'WR�'�L��dα1|n��`�ëu�I9�*��-^4d`U��!U��ʷ��>{R��ŋ�(O2dp���1:P��(��J���W#a�� �("G�Τ7��1�ҧ��J8���y�'N4���s�>1���M�I�t�H4���FO��0�g%D�"c�m[� a����`|ȭ��j(�Om�'yfp�@�G�?��C0h�j��i[�OJE�u�]¦��	��P�O�:�s��'�8�6�J2B<�a�#W�x6M�n���UnK$lѼ�b�WEq:��&�PS�z�'�Z�!J+=i�7���M�Y��,Ȱ�b�$G��I��-|����'
2�d���i)r��O�|J�(�,{'C�#�B<;�Y��?���ퟤڴKܛ��'b�O���?'�n���'5�^�)�fF-E<��'�B�|��i�AQ���	m�ę�o
�B�Z�qd�=�I��x�ش
���|��O�
�Jb���j%�MR���L� ��hӞ�d�O�Xs/��q?���O����O:E�;�?�Sd��v�H�,X�o� #���'Q���H��O��8�Ə�5�i3QR>1je���'���Q��ؠ
����L�:�x�K$m���ի�ʛ�q�H=� Iݥ��	
�_R�RN<i��0+�X*�,Z�)j�c1Η}y�@2�?�U�i;�#=��'Ͳ	����~%2Yj���/!\I1�'�6 ᣅЦN�ޕ!C	,x�b@qf6��^���4�'g�	�GJ�H)�
�@E���2�2�Υ1 +Ѫ���ğ�I�pAYwy��'"�	i3� �s��*|�(]�z��ړ�B�aIL,_�6Hs*���|�X��ݐ��`�@7@	����+m�;t*۠<��L������`1r�`���F??r��On����'����-˲|��в���n��8J�c���0��D��Ms��M�C�Ls�GC���m\�<����A�y&���5��w�|}X&�GNi���Ms���D�
�p�O��ݟ�Mˡ�́�@�A0����r�iՊmP`�'��'P��:�KUHB��G��x3E5]�DZ�oC�i<�J�k &>*0B�#ړ&��@�3b���hC��?H��H�%>I���#U�k#l��W��4X<���$�f]r�'�q�BL3�� uQ~P㐮I~�V�%X���������j�y�`���HE�A���Nu~��7r
�ϓ~ɸ�1d�T���T�\���m�ܟ���f�$Q�(s��'��M�����8%�¦�8Q-2r(h�ViZ�D�]��F8q%��1O�,5!�3�-�S7l\N���h���a�J=�u�I�7e�ScR���^
X\��p� M0?{q���(��ҜAl�h�-̨�J4!V��O&���'P�O?Q�5���>���A�	\o��(Y�<�D��aP����FJ(aa��^�'�#Z���n�R0�g[tn�IZW���eG�V�'�2'ƛpYB�X��'�b�'cR�j��i�2q�C#<��#i�	0�^4��,��"�D1R�
�D�p�*I;�|ʧ_A(�[R(��/d�2�a�c��s𙓢���8(RuCv/N�B)�G��,J���T>�a�hPEƉ'y��WC��6�zX��E�	K��j)O���U�'] ��đ61�:�r$I �2XFl�QnV�N!���� �$Z&^��sN-r�F.+��|*L>�'Ǣ��0����p1��P���i�
�?)��?��� ����O���m>	
4 �#u����>̮u�5(���n�(��^��jl�R*�\����)�V�'T<�$j�$-��!�2	D�[��*�(��*Δ����P��,��2�r<���2ef�d���b ��^�sG4EKI��^]n`�'�Q���f�����IgBU�|$�v$0D�@9��ѹc'�h�!�T�f�����>��i�[��SRe�5��)�Oz�ӯJ�Fu0W��.3g�
6c�Y��7�=L�H���O��DԨi��uR�L�>M0<���Jǿ�M�'N$�(B7`G�+b��|�|�S�	 xMB��4����T"��򉃇1��8����M�n,Jd`C O�ў\����O��n��O�!�5+_�`�����+$�K�O����A`
X S���:c5�Pq��a}R!?1���y��a��ߌk�Z�����[}�''_�d6��O���|��E
0�?��8���A�-�H��G��Ԉ�Ǽi�T��7b�Y�`�2D�&�p��cIx/F��c��M�z�P�D�%RN�y�X�}����(9v�#��lQˢAB�l��Rc>�OS̴K&/\v8�p�U�T	r����'�����K�B�<%?��O�V����ܶ�9���PXXs�"O�u��.��a��@'Q7-�j�9���O��Ez�O��)v��')or���� +j���+a����OмѲ��/�v���O��O�,�;�?�Ql�S�V� n�=���B
�����l-<����'K�Ѣ녢���@ K릐�I<	�N�$,�\�* ��X�,1���æv��ݓ�
[!?謈/��~H�ܗO��x ��g� I|V]B�Ʌ�nh0� c'�$�nʓ溹����0=�A��! L�b��?j�$��ȒP�<�E٤j�܄��E;`��b1�H̦�`��4�ޒO
��A�4db�0"�&��U��H[�7��ȓW��p�̒�&�c�n����'��a`�X���H�/�7l$ڔ9��� �zd��9}R��A�^=r\���"O��:2��4f���jŃBI����"O��{a�;h~��q��q�F���"O�0��[V�YRP�H c���°"O2""(=�����`P��"O��"T#F��T}녢�#W��<��"OZ�a�StC�`��B�z�&���"Oj� ��ְQ����h�$s��k�"Ob	�j��f�Z�ZA��0���%"O�4�q�ɄF=JD�3�Ît��
5"O��7'�^Q�5�%
0L�Y&"O��ahT&v�v���
n	T"O��@U�30�%
���0H�I2U"O"�{��A�b�v����Bz�$"�"OVR-��U�����X�nf�<s�"OɃa��-����L�`�P("O�=`�-EO���Y�'ބ'�t��F"O����� �rp��S3G6r��"O Ց��O>^�$A�bQB�Q�"O�`)���<O�,ae�ܐrt����"O��@(�5Ve`U�Ŭ���	""O�00�L$�1�����r�2() "O��`lM"����h�y��Y�"Oj5�7�+<Ʃ�sZ 27,�&"O�i(A!�<aof�ͣT��ȡ"O~a(��7WO��3�_��flKP"Oz�:�eą^��,M�ޠ��"O��#�Θ/Hg��`&���~$�<�"OR�r�Ά�؂�`"æY!T�b"Oj Sf�241k�Fʽ/�8+a"O(9��PL�q񃏕(G��i�"O.��F@<LC���%�$yL�:!��K�z��y�wM�S�,�Y��G�y!��$6��]Be舷[�SR*S	2{!�d_>{�p�Y��	�
�:\�W�D>;t!���
]E,e���`�v���F��U]!�$Q��l�V�L;e�	a#@܌8"!�D��Bφ.mW }Z�- o�y1"O6T�3$�H㴤z m��}[|�3"O��RӁJ�n���#�TE8}�"O��8A �>T�d�N<���E"O ){�,Ѣ9^6(�7�@�3v"O��`aK�<���1AI�0�P�@p"O��'n��wi�ygY�':r�2C"O���ƖQ\<��
���ȝx�"O|�*�+��L�l����˱|5ҵP�"O$��m��[����%�¨$`@"O�}X�BՕB$�1#�ĕ�77��H�"O�@ F]1w�ąA���i��y�"O��86��5:� ,����E�V"O�!hQ��A�l����ӵT��Ź�"OpI�t�v�Z��E�}��"O�M�`L�;%�H�S��F��{�"O\-�5��(G{�9��HΖ/�a "O��Z4n>~��P �
9j�}i�"O������d��$�T�e�"O��c�.� �|�4���P3"O����֖ �kFOZ#88���"O�Au�VV�YYa�R���=R�"O�����(:l���.��H*.Q�V"Oz�Ӈ��%`� $�	pD8��"O�*��T+ �N�{S��8
b3�"OV��wF֒¸-(� \
2��1S�"O:)#sa�$�G������"�"O� ��!���	p�<1Iaף�V���"Ot�X|x��a߆|����c"Or}����(0�l�de��zl�b"O���4�Ĵ_D$�%DD��脘"O�2�h02��r�ـ�Zh:5"O~�2���k����FGߒ�3"O<8�E�6�rd�7%� ?��x�"O���p"�Sx���1:��a"O$8[b$�cD*�2�$Lh*��9t"O@LK���@�H	�Rv"�p'"O�<{��m֠�@4Lr�D"Of$����M��ԣAGә/a.5��"O>x&/��Lg��A3�[{G>I��"O�����WAvM�'�K��⥲$"O��D�B�����.�c�D��s"O��$�-|�l��q'�5��	�"O��d*�=!��ؔFZO�L���"O���j�&{��bCQ ,6$ �"O����7,�p��ᯞ�
���i�"O�r�*]9}av���H�/K�RUr�"O���F���)���K���P�"O��v�J> nzTɷ��Ix-�"O�y�G,�oy��a�rr� �q"O��i�`�5RI�m�8�I2"OR�y��!}S^��r'	�QF,D�"Od5�v�<i�X�*�%B�KL��"Ov�`e�X9�Ш�f��Z1�"O�a ��(_
Q"��G���"O�����>L�:��e Q��f�AG"O�I�50��\�����" "O* 1a� ��f�k!�H�"O��hM!�8) ը�	}�DU"Oޭ��ڜ;���0eQ�6>%��"O�K��I�;6��*6n�"u�T��"Oz�� ���HӤB7hkڅ�d"O��z�Z��>%9'��$�\Qp�"O�ł�cS��d�H�M�)�>�k�"O*��$,�I�$�1�,�HYn�:�"O��3�M�kp��QLS+*Hp4��"O�a�@˞S��0��HJ(��"O�}Ȑ�݈\�^�Y��J8 �z5"ONt�EBXx 6�Xb�p'"O���g^1#˂<Zq�Y���"O�8��֙zi��s�L�<b�����"O��k���?ȼP�sc�P�cA"Ot��`��S�����ި#w�(CW"O}��fC� ���2�Ս�H�U"O@\�c��K,�%�''�4X5��"O:Txg�N�R[x���H�J�X�"Oԑcr�Ύz:2h{��ģFz���"O�MS���.@��h��*�ZpZ�,�y҄�4!]�H+@�M�W�,��
��y����v�p��$�ΩMU�e#��Ӗ�y��ݞʂu�,��h@P�Լ�ybD_��jQ���B4*����U$�yRK����vLD����R`"�y�G{6!jS��`> hR�����y���*@���h6��,w,A2D6�y�M�	?��Y&k�0
@Vx�D/��yR�Z�3�`�@5���>�l�#9�yB�	~��`C�nE n�.�2����y"�B4G
�gK�U.�
���y�!S��^{C��G{�� N�y��
�v(X�OC7uʜ�6�Q�y
� .�&n��5&d���c�|�p}�"O��#Ē�k��0���Юq��Ụ"O���3h��/YtĐ�C��g#ڐ�"O����1u�6�r� 4#�(�"O���M�;� ���R�(��"O6�*��ύd%h�C"V	z*y�4"O s"W5a� 1�a�[.L��"O�1'i7���f���W2r�:"O°�«0?y$Y�iK
LJy�"O���׃�"D@a�ϸ�!Z�"ONE
rc� h��y��í-�HE��"O���ׯP�0�YAo?,��a)�"O�TStJ�-+����톗 ��р"O��Z�K��!U��1�D����"O�äX�U��Y�Eǂ�jU��"O��j�f��|p乐��*�ܸ"O\i��b��Y��1�is(�
�"OhY��k��sVτb��;D"O�5���c�TI�N�
Qb���"OQz��/���aMZ�H@�S�"O�%(�"����U�/����"O�e`� T�m����a�̋~�:�[Q"O�aj�H��Z/:��̙�?��%"O�H��ҍW ��Q�CEe�DE�#"Ob��FHט 1:ܓ'`�vo���"O^X�H * ��x�t��{�V�b�"O�	��$P�&�%��`�+	��"O����(fމP򁃁�pmJ2"O�Hs�	
�0+N,�$���
�@�"O�q�gç\�ji�d�K�y4p� "O�l���8L`���%��!�"O|�s���7v�Ns!�R"f:��a"OhU��ɜ@<
@�5-\�ge@��"Ox����H�_mRI v��=�;E"OJa���_�#q&�����.�Ts�"O�`��Q/hA$��M+CQ*�j�"O�ţ���2S<�ȁd�K�ީ�"O�4���$�����_�4<"O��	�0!�ErJ_&(��p��"O�Yc�  D.@��jȉ7����G"OR	cT�7��EJ*�L��Ib"O<d�� �	�u� I"#��T9�"O �ӗ��v�������ؘj�"O�0-F!��KT
o�� ��"OP8��瘌q�peۂ��5@��Ԑ"O��ÔD>j>܄A���_ŢR"O��A%o�Vb�e�m҈,&�V"OQ٥eH�k2�(�LR�O"8��"O�	���6c��tY�CT��J��f"O�U)�FTOu��
!�M�t&z�"OJ�Q��-	T������P�����"O��.ՁH��4`$�d`і"O~�	"�_v[�=����T>�%8#"O`�5�/1#��%Du@v��"O���6�	O�$���E�79��m�c"O4�q ���{� Myc�SA�n�I�"O*t�9�b��*����`��jB�]˒E�C�	��<е"�WI(B�I	d>(�9��#Zg~�å%�u��B䉦"ƞ��HX�r��@+E'$�.C�ɂ�Vh��H
�)��B�A�C�-����aS/�슷 ,]��C�ɴ(����ݎhI��c���+��C�I�o� D����t��,c�G�:�tB�)� ��I��Q�Pא� ��ŗ.�Y�'������A�T��r%��~�P�cDH%8�B�ɼ%�̔��
'�B�����#}vC��w\��4�U�n�SE��GhC�ɖ,���a#�(���s!�!%��B�ɳx�H�#��,'���4خ/�B䉾�`YP�e�����LזKH�C�I,|�n����)�	�&���%�C�<��F@�8V��B&�U�
�'��:q���$� �2�FɁ4V.4�	�'κXI!$<!���,(���'� ��1K'�. ��';b��'�;���Z�\(G�ٿq��
�'Ŝ�0��a��`��܅n��� �'������hH�9��B���'�N��)r�ԝ����$��:�'E*�Q)˓b�HS!�'��	�'h��ë�0J~��A���0��'K�\rUN�.O0EB�ͱ>�����'ՈX:�bJ�0HN};�$�:6lX��'<,��C0N�X��R�'�Ze��'En�Մ�t� d)q��l}�
�'7��AW�	$r
�� �ܚ ���
�'s��3�W�{p^�ᇋ �gZ�H�'�������&Z:�xTh�.X�8��'�&�{�K�?Ib,�J'F/P�ٚ�'y��頉&#����6�A"'�8�'��ۦ�$n�x��ei o�����'����#p������,@�'�f� ��2"`z��c�YT���'svu��b޵�����	����
�'Zv�"�G�A+�ȶF,Q
�'�B���+�;|u<�6OB�l��
�'��Xs&jҠIy|�#%�L37|�	�'�((��	�s��L��l�� N��	�']��/D�z�z��q�]|��I��'�8�q�~���R�w�*x�'������:\��ED�-fy���'��T���-1��̋5��'&�-�ʓY=Dl��ɧ�|��M�p���gǫUj���r6�҈N'4�ȓE>x�v�B��dHoO�94.A�ȓot@JQBj1��2̯a��ȇ�H\�#�`�!K7��)�K^"6R}�ȓ+Gj�K�m�#Bp���	`�:���y�� �p��`����Wm�8l,�ȓ�ʜ�2F;[��<c��]�L�>���=Y���2�E~9�9[�bÞ9*Ή��GUTԢ34ۜɪ -B��|U�� �軧�7l�HP�4M�]��ȓ7��"���FTh�WZb����u �14ćc�8�5G����ȓc����g�?e#
��&� ;.j��E��-S5B]����$��:�ćȓ?�V���9���R���9���2��xD%�D��*�'ùm0����4(�D�m��}P�jT��W�)��8f�����$-c>@�V�Z!t�<��ȓw�Asg�I-2�UɆ��;��Y��&�<�R�AF�Ft.�� �Qq��ȓXת���i��g�%A��(ܵ��^ʒɨ���Z�A� F���фȓcLx�C�e�<�(��'͞)\<��3��5��,��:"!{"i�W����S�? ���cR�x:��y�DƏWrn�$"O  zAIבJ�����a�w���ˡ"O,u)�N+>8`����yz��U"O,�S󀁐ET�M�լ�pE��"O h�P
96��%Iͽ/�HB"O.QQ)E�?�z��q�ܑ#ĸ�;�"O�	��Cs�I�Ы�y�L���"O
IQ6g[�`��C*�2�����"O"1���L0k�L����=up��"O`:�h
N6L�r.�a\�j�"OA"� ��U-z��m�)R+��A"O��Y���c��ȳT.]24;�4"O}td@6DR��p�&~�r�y�"O�c�1T�VM"A����I�"O\��ڜ*�X�q�@�U��ْ"O�	DN�)8�tQ��	���p0"O 9�1��&Yh,����-n��)r"O0�æ� �?���kӤ��ql�y��"O�����?l`퉕�)l�=
��i�ў"~nZ�Fl��!E���"r��IF�OڌB�I�d�
���@� ��a6h����B�	�l��0���?�AK�A~�B�I�e�����Quv���C=9vC䉜^d��PFM �c>6I˖��.<�PC��"	~��էf�Eŀ�|�NC䉗Yς$aT�G���tL�~p�C��uP�HE"@?��ء���{�
B�	�:��qbA�0�j���G�+	� B�	>�2w�B�Bj5X����>D���`�N�<l}�  �*	���>D��`�L/"��$a&�+� �U <D�lP�-*��b���@n��;D�l���W��lі�8<�ީ1�;D��q���1?��� ��Ar�r4J"7D��Q��	��L�	�r	���3D���mE�.�d�y��Nx�8i[�1D�h��K��~O~h��@>XQC@�-D�HW��2!��ۖ��#��
5�*D��B�l�$ �>I!q.�¶9�T�;D��j�!Ԏ�t� Ŕ>2פ��:D���6)K�"ݞ�3̐�B��i��L8D�@�`	����E&Y�yҮ�׈4D���"	�,��'��#6ll�b�<D��P(�1Y��q��EҪ%�^�G�,D�����^���`�"��]�^�P'�7D�����k�M*�N�}�H�`�6D�PAAϖ6[ʐ��eX�j�hh���?D��I֏�-��\�[�;L*�XtF=D�\��#�O��ݻU酬Zu�A��;D�H�W��=:S��*UaF�;��s�8D��Z��� �#�9���s��;D��{�> ����bf�K�A	B
$�b/��~B#m�s�=@B�Rae{���C�<)��JR�+#()�8�:���V}�)�'PoBأ��^)���	���$^�Q��-*��1Q�#�&ĸ%�A�'�,��'���
�+���iuҍ8�jq�6��7�P��ȓM�`�I��v&Y�� �_ۨl��k��<��Z�$r�#R��,FQ�aF~���nl�����e�<�*f�;n��B�ɢ�x;e�]�(e�� )b���	|�Y|�>��vX8Tl��/{�8��N�F�P!��7B)�׫N`��k��ڲI��d�	���?�POP�1k����P�y�4�:b�|���A����� ���jFk��`
���;��Zu"O��S@�օP�(lɁA�z���3��o���S�?K����:�$d9��͌;��C�I�[��`�M̺p�\+@M	��Qˏ�9�g?AQ��/�h<�0̓�Y�晹'�t�<1FJÏxr���a
`�X��Xs?!��F���
�KW��(PB^�V�P��ȓ5�fMPWL6�j�#�ǎ.�Ն�ǅ��ylj�s���������~�<q@�3�pع�&W	`�&T��jBa�<�V��	���`��T��R�d�c�<� j��j8a�H�@)�Ū�Kt�<�!#�L�m:���5�D��z�<C �1x���u"J�2;�M�r/Ov�<ᥦ�5�.�	��K?,j�(h�Oj�<��
:
�"����6�}Q���e�<�ע��\s,�㬕	5ٰ0�!	Y�<�VC,�^ �V�ф�U�<q��O>*��t�4�B�l�>$ 6��i�<eL�m����K_ @��䫆n�<�F�/��%�_j��H�c�Ne�<�r%��\!&�t��K\k!���RUB��	�W�P #'��7N!���swh-a`ID>��EӅ̃�&3!���uXJ6�XdT�,��DE5�!�dI� ]��p��_�$4�'d�7~!�D	�	���`@l�m��|�ECG�v�!򄑵}���T��1Q�2�Q�H�O!���jp��sͥ>� ��3�M.;^!��(t�-����}�B�T��$Y!�dU�<��|�����yI�I�8W!��4K@�ҤC�!d�u97hT	`K!�!y~PT��g��i�cgϩ[/!�D��8�@����Ŭ�8d�?T!���Kф�S�.�s�����& >8!�Ę2M���;�L R>iKD��N!�D�f���Z"P$g7Z鸕J�+e�!�D!q�&��2Լ I�1K ��!�d@�i����@�Cl���L�+o!�Ą��f1X�Ä�3�1�b�1�!��եZ�ش�C�Ɏ[ FY#V�A�!�B"I�2 )bbٮ v�ҡ��z�!���	p��x�'��4Ϊ�yG���!�$SY� di5έ#���!EF�z�!��>R
Bt��6�c���p'!�$/0�x�b��Y�v�1e�*�!��8w8*M�A�4=��ӓą`�!�TM.N|�%�tK���1Ζ.�!�D�.k��Xc��8V%(�S'�H��!�ĕ�>lt {�/L�9�T1��C��g�!�d�9h6�dc G�d�-@AK!���Abl1�����a�(��၈k�!���\�����)��|J�@8@�!��s�i§&4���ƥ���!�ă28�ڴc��ó}#@��B%җL!�D:Ji���#�^����1���P�!�$�Pbr��t�\I�D�0a��4�!򤍅S���
��%q���Xp@<T�!�$�?�Ь$'O)@ ��H�!��U3h�j��nF(fP�"��Q$r�!��ɏk�I�E�!3S��a�LB�!�$�LY~A�2ER �ʡA�Z�!��>_�ԊUg�8N���G�>�!�$[�u9 Y��ޭLA�ؙƪC9!�� 60���\�<���A�s.8)�"O�ka �? �tS�Z/��PP�"O8��aX	��J֭]'6i##"OhA���7���A��Ê�T�P�"O|X"�C%�(p��(�&=H���"O��р	�  ��6h���'@  P�:"Ot-����7`�8��6I�����"O2�s�[�w���f[,.��+�"OPٱ�3\
��r
�[g���b"O.��%�!V��`�B�0H��E"Op��cJ^�?lZٱċ�t��HI�"O��bn�o�@%I�A�7��X��"O�AvgC48Tf�;��ʮ-��D��"O6!!sH2h�P ����	{���"O$�xP��6 y!�b��w�3�"Ol�"��O3��up�C�t�4��"O�sgb���b�$�8Dm�"O.�����2z^Ո�ꈩZNB���"On�JgA_-W?N ��Iځ4i^(�"O�	¢�F�A���"%�ޓ"Yvu�"Oj��c�B2H��(C�J��$�8�y�"O�i�Ѭɿth�q䂜�u�$�)$"O��Y�CF�ư:��ՙe���@�"OH@� _�1�bB���X)<�'"O��G(��8, p� 1�"OD��Dm��$0��_j P�ҥ"OHywE�;i����c��s����"Ox�w.Z����Ad��xi����"O����Λ�O�>�2#�L^jm��"O�� Я��3s ���@$(��XY�"O�)�t��� �b]��� !eR�8�"O�y����hDHr�f�
MI>d�S"O*h0�͡N5V�pc�pԲP0c"O��p�d'mH2m�MN
#��"O��4��k&�U�4i��aR"Ot��c&�����J��O�N(�;""O�h��N3��i O�'eBXp"O�M�7-� i��*��2@W�<k�"O 2F�R�,g�!�%]�	D����"O���"�T�!2�	Ɏv�b�r�"O�5I�(�f� qF�Z
 �j18�"O��[G��=�.Q������H�"O<]��P�\&Tam��n1'"O�L���G�]� �p����� ��"O��Kqh�U�����)B��H��"OLU�7m�1w�@'L�ʦ4*"Od�Qs��8%�� {�ɛ�9����F"O�z�*5.��[�F���xT��"O�@��8��[��M1bPP�"Orx�"�5%���#6BA�1N���"Ob���FY��(�aC�gb�a"O);Wό"� P�JE ε��"ORa VLL]��	a*ף6m@Qs"O�4+����G
\D��	�)��11�"O��b��%S�k�.�,�420"O�h�r��<%�f]��J5-qP=z�"O����2y���Ή4�ʙ�U"O��@��}?�ekg�'T9���"OP�1���(���UT $�D"O8}Z���6:x� �?�,i��"O�I賋T�N#ԑ9d!&�PUQ�"O0����؂v�U��^��"O�1r+���V�ʶċ�1��0"O�Za��+E�(��Ǹ�||�P"O�Q�7O�.C��0���.�-E"Ox����ȎT��p�P$�w8�8�"O� !` hW�/�9�E$C�|��U)�"O��(@@[.X$�jț�0h�"OfAiVO߼ a��Ã�(Վ� �"O`�24�%���D1���"O�0���Z�1�V�qqm��N6r"O �3F�2e �+T��m,�ɱ"OРQ�ǆU�r�8�m�"Gx8� �"O�)z�
XP@BDK�ad��"O�%{�Q�*�&-P�҄g��]��"OF��ǮD:#Ȅ��LC�����T"O^���EL����R�B��B�,�5"O<�@hN/j4ND��l׉u��`�q��b3�Q�s&�'E�άJg �k^6M���<劒-Jz���e`���!�DU��]A%�L�\�e�C�B4+�!�d�&n4)�A��88*�(�]<E�!��]�m-I�<E[�ŀ2���[�'8�B�A�<��o��`��ix�'�j�h�%�	�h��p@�&`juR�'�h}ل�ě$�x�K�!��	�X��'�`m�b�Y�z*$�cDI�r0���'#����JY�j�01兹!l �'��h�V�W29v���0@��$���X�'�P���٘S������*"	.ђ�'U�H��=����c �FH(��'O��e��$%Y ����Z��	�'�n���K"+P��֪Q�?�|b	�'����'�ܰZ8J����+~��H*�'�$��V� ;�ec��BxƸb�'�)ȧ$���$���;h+����'R�!�C �:'l@�v�	�wE���'��˵mX,��aV��f��T��'�Ѹ'BUmZ����ޞ]�@��'b�|�rF��&@���Z�	B|��'wu�T�� ���ƑV���
�'D�I�
a�:h0AEN��9k
�'�T�s'%_�f�"��)n�^t
�'�~�ƌ}!ȵq�jG��0�'1��RW��+(<PfB�^Dx��'����DF�.��if&�)i=���'>\`���ȣMĄ0+V��9Z`���'>Na3�C��Y�jH�O��	�'/��	s��-e�q(�ȬF/�TX�'�<!�±[�uQ��Œ>�8H�'k�iXRL��h�D8B1e��6(F��	��U�$M�$���I$��F�`�<��/_0	p '��i�y4CEb�<	1IN��"��X����ɗ[�<�S�͕i#��A�`I
���nN[�<���ǉ$nN����=��!(1,X�<A� �?%L�� �A;D�|�K�!U�<Y�fT�
[NI���0~YH�K�}�<�P�F��Jq��)F̼t��Lw�<�CkʟM�!z��٦9�ܨ``�M�<Y�f�9<�n1r��P=�4���H�<��Ş�F|�q�ƑPB����|�<E�T�2���-�yU�0��%�B�<�u�΀<�X�,�@�X]���x�<��j�L�|�봇
�$�� a)]u�<�#̞a��쳂�»t�j��$%T��A��W�[�f�B�{h��B� D�8�$�SM�M1d�+Tq�98A� D�HA ��,���," ���6�:D�H�c�2s}��t��z�����+D�@����1���t�
1���I�(D�� ,�
��@�8����5����"O�����+����d�3nE�d��"O���͔*X�Bɪ�9F�7"Ods���u9SD�<'�8i�"O`XYr�D� =��$Ҍ�6`�"O~pz�'�'t�f����ۙX�@a�V"OH�������);�BK�Q�9jP"O�-J-rQ�)p!��|��YW"Olx��X+�y���>G����"Ont�@���k�����ؗO�Ι�"O�0b$A�$`��D%MšUX�Sr"O��H��R��C��O�X��}Ra"Op�ط ���2�{T�ʷ?�P��"O~���c��f�"0d�0;B�(�"Oz�j��H?� U�06��"O]@RhF�2H4)KcÐ�%��"O��3옝C�\�ǉl�2D�a"OxHх��k�UҴ`�e�6e�f"O^���f
P$)��l��Ϫn�����b� ����}�$|`4%\&&/��ȓo�>��qn_�t26�Pc��z�&���rf���R����8�����Є�Į��H�f��ܲ��4";�Y�ȓe ��sgS�'y�4�e#4NT�H��"x�PܓQz^��7ƀ�c����E�}�w�)\��ˠ"ݧU>�%Dx��)�,΂F�R��E#Ӯ7F�iڱȝ{�<�Wꍱ8�X��L�*N�|�!���.}�6"=E���xqj`m�-`��񇪍 �M��1���F�M�?l���?e����'�~bܘc��]���,�،A�톛��=1��|�&��T�t�hF.O2<\"ș�y����.|�P�}�><Q�Β���'_ў�O��p8�-M� 0&��dX�p���	�'�4Y�ړm*����](&���C	�'�^�`nћ~`d�fNK(R(�R�'�b��!
ZY�e�eL/s�t�'U,��փ0-�8cG��n�����'l(p�r�̡.vl��d���l�h�'��v)�jtc��C�
@��'-�D7'h$�!3G3?����'��4���=J@H�.��1��|s�'�H��e�Ӱ4���i�!X2W�B�	�',�HP�b��E~��h\::�0��'�I��8b�49����/�J�p�'��
ĉӳa���P�V�!O����'���x �H	u&t�Q*�/d�a��'�$�IѨI4c�&e��ޒpX����'&�p��,خ���Bp/Q-g��u��'Ю�pt(
&,c��G:-z��i�'���%G�vG�2�O�+ɬ��'b9&��!:ȬA!���:e�m �'4D�����4��4���3"w�z�'(uF�^���X��P2d�l!�
�'� %�%����x�
�#a�� ��'�R4	�G�37��t���ƯW���B�'FȜ�EG�w:PQClC�~ZPQ��'U�)���8�qB��x��4�Px̀"�P��w�V5;"��ا��/�yr��7�� �7��;<#�*WE���yr͉<o�1i6�ߖ6�$Ij׎�6�y�jӃmx���W�I83����*٦�y�@Q�\|)DW�v��K��ǨG	��I[�S��?	�-��l��͸�l�76 �h�!%T�� �3��ٖd���Y㬅�:��ҏA%<�!��K"LS���ЊP�B�|}94��=R��z�߳Cg�'��c�h� g�V%k-��x��b�'��%��EF�I�
o�4���{"�A��O�O����&�
	B9ص�Gj�b���'6|����!�(	�k���]��O�=E��KM?6}��C�@�Q��� �yH�>@! �X�n:�]8���M�a�O&ea�F�,`�U����rx�DGVF�݅�	,��2c(�@@+Қ>P0�;�+�W�@��l�q9wMV$N��D��/Pg����?P�}�آ�$�ζԺ��K
C����u��T�<ɱG�)��i� ��l����eC�ў"~��#�(X����9O�b��#�;A��C�	I��� 0�Ɲ;���V�Ƴ{�pC�Tt�p d�!��,��ޛ->C�ɖt8�1k-<]���fX.,C�ɓa8 MP�. j�<�b��<[�B�	�j��(��"�1tMz`BA�N��B�I��}���Ҕq��{p�_8x�B䉫c�S�A��(l��@� :Y��C�	af�qtBV+X��@1��+ZöC�	���}�ƀȱU~$i0�_�)�C�ɘW�Nq���G2jrp8�GAP:B�I�B��x�V��.m ��]� ?B�I4W��P�v%�/u����`J�,=�C䉜Q>Q(��H�l��8_tB�	=
�v�Q���E�(�Y�)b=DB��_�,`I�!e�9��Bn�,B䉤?ar4f�=N�D�R�3,kB�6 ��5�'d�wx���P�;�C�I�p�lzc-��W5�y�WG8O�C��9����Y�4ؘ�Z�$Cu<B�I ^֊)q�@*UkZ�Ɇ��'B�	�M�&� #��#�IB�$��C��8deV���A( ��B`�Ր
ʴC䉡F@�dȖ�S�^���c���i��C��+e|���,�3\y�\�j��@JC��'K�.�
�G't����_��C�I<�ک�v�@�1+*���ٱ,qrB�ɛ��hH��P��z�a�BK�B�	'_��M�V�X�Cܰi�)G6CStB��.a�!�O�"{=ʠi��5qJB��13��W�<*�r�c�[ �`C�Ʉ"�.遃��@n xc�#@�<C�ɅEw|P
V�$o��z5�W�j�ZB�	n���>��r,֌o`C䉭gQ����);x ���8l�B�Q, �@P0~=�<����%��B�I'0CV�`�`Rm����Fףj�B�	s4�yڡ�3u�����>U��C�I����b�#�G�3�
����C�	�^�N����E�w(� 䊼P�C��.-��ab��20�h����G�BC�Ti ��P�8n���r �) C�IIpm�RaV=$*Qj0e�=_�$B�ɧTkD��!E;OTV�ࡏ�\<
B�IP����N�720�6�ϒ5h B��/|�L���x�x"�+�\�C�ɀC{�u��j,Y �5�N
�j�C�<�>�"�̃|<�wC�B�C��(*����R�ӭ|�)�k�k^C�	�B���`�B�9�P�0�-Q�s<>C��~�E.H�;BH!
!��m(C�)� (=y�	�&��CHȶWOX�"O 3fk��?t!�I�!Q ���"O����Ոy�jٓUEC��)�"OH���R�&�P�� �0���"Or�آ���aP�reHJ���i�"O��X4F$c�Q��J�gw�V"O��d-�%X�����\!{m��"O�z�`@�{��� ����;^5��"O�2���KI��pjM�E�TEx�"O|�a�$�3���x'�ե:���
�"O�}#t�^j�(↪�!1����"O���iY� �h A���0c�,͋f"ON�+D[�7&��`rfT�x��ዷ"O�D*P+�����S7�2�"O�2U�+Z,�����R�gd�h�"Ors�i�wd�����
�,���)�"OJ���
�
  ���l�@m)�M+�o�뎓i�\�I�a���I�$�Ucul^' ���.T-R�U�Uā���)�FP�+m��VZݛO��qp������ߴUC�� �P��! �\�H�4*���9�n�l��x��Dx��ʓ*�$����O�	��G�ޱ"�9aH��k��Ƀ �>����,�D��7�>q*��N �:%c��'�\�D���t���A!1���#��*Ӕ|�k�8#����4O�� d,�%T������]ؐ�O�i��R)wV�'>�MQdI���\�F� �爖+�\�a�C�>f!����ze*�O�(҆�v8�'Z�|��	z����m]0\e�qZ�D83�%!O<�-Y)3�T&�$���1"d�`�ȭ��ۏr���fL��<�z���J^1�󏧟�c�'�@��o�jy�O��lpP���q��8��]�?�bСS�<��� O<��C.du��??Q�O�gS��&��|���W�.$vRЀ ��=�� Tqָ �$.���q@����>�@�Ҹ|%j%� ��E�l��A��
ov��dW��~fj����i����?ݬ13�8;��%{Ƽ���ɺR���`�K�HT��'l(���;���u@�G��<�֪�H:"�� 	^���6�n}M�.4RB���'��I�1�@���T���&�����"X�@:���@\�KMH��v,Z�#��	g≄#,�'��6��,tA��}�fpa6
хdP<���Ö�^�:�&E�l�"�9��ʽY&2|��'{H��&�} �Q��'��Q�b�G�8@��f׈cV6�;-O���!�U�Q;�'���W��ēX��(���I�/q������8����/&T�%��X�>����dE,53x��ƳA�`���,n
bI�$D�<0��   ��(V��^�D��9p8�b�U��EPw�|����:u��U�L~�@�&R܂0;�^�0G˨X+L���E� 2��u"$�w�젴NC����#�'��X3:�H�3�՟$]Γ0���W䙺����S� 9L�����ҽrˬ��Й�|!�
|܈H��?�×�ϱy��*�Ɉ��� �� + ^�Y %�!���s�'�,�� Z}� s>��4c�/ �$�O)6�!`��!R�&8B�NE�E���       �  �   _+  �6  �>  �I  �U  \  fb  �h  �n  0u  r{  ��  ��  9�  {�  ��  �  F�  ��  ʳ  �  ��  N�  ��  ��  D�  z�  ��  ��  @�  ~�  � 	 ,  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P���G���к�ׁM;(�2�b3eR�35pY(aM�w�<a�E�8��h⎗b�h���[�<��aV�RP�����4�P����N�<!s��^��lt	�!�+���Ky��)�'4����G
-T��#EcA+$�ɇ�r���Pd,�!cx&D�C��"D~Ї�x��EcC�O6(�=�c�Q�*p!��\G.=���ݮ]�4з!�T2ȅ�N�1GɊ�� ȗ Ρj����ȓ�.�#¥P0�g��F0
����TH�	B�X�.Ⱦ5�j���ē<k���V�*�Z��U�W�`�Z� 2�}����HÃ/(U��lx��	�O����O����ъ[(����?L�* 80F��I���ǟ�'���ڦI@J��o�,1j���qp�h�$�=D��E��n�Ҽ��cQi������a�N���5Ox�O���IKVl�ТO�e1�$Ч)/}7�C�ɯ��M� E	v���v-C���B�I&׸0�@OElP`P��_�x|p���O ���gkb���l��>��*wZw9!�dT67�칣2��� �a# 6�h��ȟ� "�@1n�O�{�$�"h�D4y4"O�|i0B��l��)�b�V>~b᩶�.�Şw��0�hE&��	��*���H�ȓ*�М�V�ԙAN��[d�`�D��'��A��'g�������( �l@�
)x@	��+D�t:�A
*�������:LjР N5D�$چḽL��c@E�`l�y�"�O��=E�4F�]U�*�5s@��c!��!we�p@CĈ>t/x|jaEG	��'ʓ�hO�h���;[� �QĂ�n�� #G�3�O��'\qY���ezh���Y�7G������'�(	z�@�M ��cv�j����'̊!X�hɐ��`�@�
���F��Q��0=!w�?f��[7
��|^�1$�ȦQD{���i�h�m!+��A�r�
�x�C"O��h�O#F-���(��n,P��<����s��6x���JfԸ���8@g�=��If�I�Na��'�I�J8�\��l�-^�����:�Dθx�d|]��j�~_!��+��h)Q��@���Z'韜U!��E%1�u�7���l�l��&N�=\�F{���'�
A1*,f#�9���yh�5x� �S��?��'�T))pK0��!�H�<���S.viƐ:�L��o��[�,�?Q�m)�	�(Y�9�w�Z�l�L����C�	/{&R�(�΋k��-�%�X�5�n�=��'T�>A��&X�4��yC�/ ]J�i7N!��hO�S ��Y��-]��jRTp B�	�2y���
�19�DҒ�Ζn!�C䉋=y�ڕ�� k�T=�2,©os���p?Q��h�pK�f[ {�T�! �nX���O(T*����X0>��s�
�!��"OZ�*Uk�X���@̾O���"OB9
6#P�[<dS1OI���6"O2-���'yL�#��^�>|,���"O���5�EF�ɥ�K�:eR�"O88��߻Wp*q���7f@x���O����һ`���+��7*J�!Z�:���rx�,{pFϼ
l�Vi�J<R�m4D���U��˪Q[�ܸ=F��o%D��s�O
3sLmJ��ۘ8-��0ʓ�hO��6��� 7塀zP9[�B��+&h�� B]�*�r1�u'��M���r����O�t	P��S�"��B'tSZX�AY�0���
{1�io�� �z�`�(���du�� �7{h�bIv��9$c,D��HΔ�b�Bሆj�z���b?ʓ�hO�iy�,�Aȗ!%"�0j�i_�gR�@ F"O����H5OZy;R�H�i3ZdC!"O̍	��g^�9�B��s4��0"O���I��vT`k�#L�YyU"ObYcK��l�tx�����X ��20O������D2Dϋ�~��1��eM�uz�Y�� �$�~�'I�'p����0_�ZHrCkX� J�I��'�<U��#N�m�L@�B́یy��'e�9;g�N�gA �b#�qZ�	���y��"@ԐS���;. �� Ƣ��?9���P�q��Q%bU�D�� >^h�ONb��D�����H�@��'�77��i#3�:��'�O�uaP2�( Z��H�sO�%�P��\S����,Q++R�ŋQ��"& ��h3�O��={di�ߪy�6M��ޘZ�<���!��P�B��H�l!c�/��dς�Zd"OL	��J��T!�%p�+�׎�)��	`X�� * @��]��#V�Ʊ.Ҫ�#G�'�O�=y�U�uu����<#"he���S?��)�X�c�Ѧ)��q�.�'h&��?��4�hO��;`��y�D�8��kr�׆#B���O(P��h�K�n�� 蒜>�ԅڕ ����M��󩔼�^�1�^]r�S���5n�,�S�O��Q���I�|�dHI�,#5����
�'p�	�▚. >U��Ǝ	.0��	�'�$�*EH�oqȭb�4X���i�'4E�©[
vLP���욷a��q��'ab ��(_�}u��G����R"�yb��,�f��\�|�J0@�n��X���	;�f^�u4z%iR�jפ��W|R@�@��(����!�"m�,n�b�������A#�`A��َZW�����]�y�߸0��XP�E3*���#�����y��bV����A0�l(�7�"�yo]8#0]�b��,?�@]�@ �yR��*���/�*/;f�#�K���c�$;����$I.YS��#gň�$�p�=��=)�y�6@@H����Z�pL��y��B0\�и � �zg���yR��"G��!���߲5���1d���y�Ƴv>��6�W�z,d����'ɛF�'Z
���.�#Ĺ���G�4��$h�'/�%�ǎNݰ�z�F�	���r#�5D���ࣉ .>�@�bH��\��!D�!�Ȟ�jUv0a�_Ȁ�т�#D�آ�ŕ71�d���E,.�JA�&�	k���8y�~�fM�8S|�bE��b�VB�IsL�8�&�_!MEȠ���[�B�I@�||p�lX(_$�h;2`��B�O����Fفs�1����|��B�	6_�I�%? ��%��H�6�B�&n�h��	#nɒ�I@$v�ZB�	�bQ����F&��]�@��&?�DB�	�wК�q"U�@�(� E͝�<�B�I<O��T;"�e> {P���B�I'���S~��;�"ْ)HC�ɮ"
�M�A-[�b̙	B(C�	�2v8���
Q;�<�j���2�C�;I�Jyr�C��r.��֤U>Tk�B�	 n�ȸ�&��J)��_��B��3Kߺ����TT��bJ�KtB�	�Cg֌��Y|��K$�H�4�B�I�~jN����X����z���|��C�	90H��)]�8�vi�E&J�y�C��;M���4NE�E�p50a�[��C�~6� w�M�]��j%��@��B䉜#���xA�*]P8�2�B)�B�	�Ь ����b��X�b
�=��C�	5��Si�-kl���.	-/��C䉛o��̑0**B{l��g��	!�,C䉙Jl��ĴN�fcW�X�	��B�	�}@�����/7A�&�BlB�	�x���0p����uH�k��Hq�򄁮#��ia�8ȶD�Y�6��'�
�C䫔�kɔ��"ԥS!n���'d�ð���y�������P�DH��'����$��].��"�Z)A�M�	�'�h!K�cC�}�&�Z��Y/FDs	�'���+N$xW�e`Ek
�l�H	�'�&Q�w�ܯf����@�0mb�P�'�\�IG��	
�u g6�z9���� �cR&C���	qDG�� P�y"O�U���г����B-�t1�)�"Oi����.��5���3;9,|{�"O���l®c!�L�%%��2�"O���(Яr=v���.)��0�'�r�'�b�'l�'~B�'Z��'��u;eKP�d���S���(\`���'�B�'���'���'�b�'�'�x4�Ӷ �<$j��	6,:�iӔ�'�R�'�B�'�r�'�b�'$��'����� lD�l��]�*Z.!^B���㟔�	��	�$�	ٟh�������3}4�q�X`�򤫄��EB���	������I����	ȟ��I��H�I.y+�p`pL�^���ܿ;��q�Iɟ��蟠�	ӟ�����������D�Pf��!���i��$R���Iݟ���ߟ ���`��ٟ|�I�P�	-����dJ��r��'�X������	��(�������͟��I��I�B��<�S!��&P�����m�f]�	ܟl��ğ��	ğ��	��|�Iɟt��w��,�s@W/ Ҝ1`���e���	՟���ş����D���h��韸���I3�9y��K�fPv0�T*A����Iܟ@����@������������8��P�ͩ!�Q#�)2o�[�"�	۟�I����៤�Iҟp����,��/�Lh#,	q�`X�pj�%����	۟4�I�D�I͟������4�?��WI���p�U���"G	�U��#�T�4��\y���O�<nZ�FFp�C��%o����N��b�����4��Da��@��Z�(X���W��
bz�-�NĦ�ɝq� ZAl9?�/ЗH��A��>��m��s J���
�H4b1C Įߘ'5P�D�D-� d�Q;B��	C9�)�5T�7m�,E1O��?] �����+��~���R6_�!%Gh��iN�<%?x��N�9�r�ɔ9��D#��RG*�L�BM����22x a@��%/�G{�OR"�@;��W�)}<@��eԻ�y�X��$���ٴB�V��<��i�.<�N���:slՃ6l���'Vl��?	۴�yB[����&+3�t���=�P��v�(?1D6 �N����}̧*�BU����=�?A��V����i��^��^}A�����<I�S��y� �� �xE�w� M �B���y��~�Ѭ]~��uӶ���97ub� ���� ���L�IßlZΟ4:�F�	97l�D�q��<&w:���_[2�����tĒ`�s�G4X?��i�]7l��m��7;F4#��ϛp��cG�؋_������B>D�A���0�FEƊG#�ISk�a5�@0�\�A����B���d��èl�@#�jI�X3e�$ț�[^(��6���u��L�aR�F���[�@/c��;���K#^ŋ�ʞ�OfXDR�M� w����8 j��7ↂ<���2�ǭ�d!�@#�w?VX(�@�:%/"l�Q��:@�����( �3�#�ҮɪVU+w_�aXAF�_=�T����W9�M���҅qg���'\r�'����O��J�'>,��'��<�N�2��,�J��?)���?a���4�.�υ�k/�]�R�V3X��݂�Fݟ8���ۗ�Mk���?���:�'�?I��?Yc�׈G����!�B�XΆY!���R�ơ¥9r�'��i>�$?q��+O�A�!��aS4�a䁢��A�ߴ�?����?q�@[=T���'b�'o���u�����M�NY��鈇�Ԭ�MSM>�Qa��<�O ��'��*��p�9ц�!p�r(�K�3�6�O�=��Φ��I���I�<ѩ�t��O�r�(t��'F�3�?j�6��ezl�v<OV�d�OF�)�On�D�O����b��J�����B���$K7�@��������՟@�I�غ��P��?����I܄�	a �M��m�g��*�� ����O4���OF�d�O$U�����I��(�-g&���/�(5�13&��M��?��?����D�O����<�����;�4E���3��*�� ����O����O�$�OR���N٦��I七i��4���1%�~��6!I2�M����?)����O���6�ʓS-N�!���[6`Y	4�]���{���?���?��	�|LbԹi���'�b�Ot<�t3\-��jf&N�fE:toj��D�<��I��;,O���|n��1
&X��D�;44|��PDV=W��6m�O��DL�C��n��� ��П����?y�I�	3B}��c�Qc����cE2X�UX�O"��ǵn(����O���|BN?�*Q�R&�.��r�S)fuPm���hӰX����9�Iߟ��	�?���,������i��X�R�˱k���v 9��M��e[�?QO>�'���?	+��J�.@��"��6

�� :����'���'�<���>�-O �䳟x��C�8P~(A��	�cb��1Mr�r��<i`��<�OD"�'��C�OHV�*&"E�;b�zC� �7�OL�؇g�̦U�I͟$��񟬓�����3�,�b��5B�xr��-w-<�G�(5��?y���?�����O�|�"��Z����^+VT>��Vb̤M�Tnߟ�I��	���I�<�p�R�[��WI�M��oͅB�(�X�g��<����?Bb���?������S�F��m��W(�9� �¤@�����+�2�{�4�?����?����?9*O��D�)r�i�L%ڵLK|/���
L{��o韌�I�(�������/
�@�۴�?���V�����Z)aP���D�,��[g�i��'bZ�\�I�6�Sh��7���󉈄&I�)�د�&�'0��'�"���w�`7m�O����O���Ϭ>xX-�� ��v�&�@���poZ�ܖ'�H����'��i>7� ppA cߤ8��ɐL�8T}���i	�'Đ1�D�b���$�O���X�	�O��`��ݻLP	�A*�h���rb]l}��'O���'��^���v�鉲�Fh���$#�N���:��fo]�J9�6��OT���O��)�����O��d��Ek:��%`	�K�V�� #�`�mZ�{,8(��� ��Dt(�R���?Ś�o�ÊD`�AJ�;޲�WI��M+��?i�PS�5��x��' �OD1)4�ߏKy����eԅ?dp�D�b&1Ox���Op���(i �+�	y*p�� '��l���T�D����ē�?�������+�$h�W+2Y&6�åeKd}RҾ֘'���'�Y����Ґ�@1
��bbv!Hs�G��<KI<Q��?yO>Y(O���V��h�� �)��y��_�b1ON���OJ���<��-��
��t�Y����؝Q��ŗz
�	Ο4��b�INy�I�����d��!���4V偲Eԥ
����<�	ӟP�'xv�*�/�Iٰz�eB(�\��pq��'`jpo�ӟd$�Д'�4,j�}"�S�H�T�/�#���"I�}��4�?���Ĝ�
I&>!���?5�$�.N�5�S��4��2������{��'�H|+��V�s���B/D�(R�lZIy���6-PK�$�'���")?�BѲ6�3�#��Uc�A�i��%�'ӖTa�����A�Ь���L�7�1)%MP�]����2=�7��OH��OJ���r�����n�0u�e�>wS@y����M�Â�b���@��]�b�Nd�1i�K�`+%+G�V�2�oZş��I֟���MR���'��O��s��*rc`Y{���Bi�����$%!�1O����O�����w7@�#�S���l�#/��GcJ�mZɟ��/�ē�?!�����p-�C���H�����R�13'�\}��ј'!��'B�Z�T��n^)FsZ|(��i��JR(�A���yL<)��?iJ>!-Ox�Pf	��̖�
Á�	�v����:�1O8���O�D�<9u��|�A="�^�c�3"��'�S�yn�I��	u�	Byr���Ď Cw��q���� ����.$P�	��	ǟ$�'����>��1��(k�� ��fb�����lZ�$��'w �@�}��,?�| �fM�GF4��R���M3��?	+O4ݹ�dK_����$?�&8��_B�j�8ìR��<��M<1)O���~�U�W��[�
V2f����X���'�i�ad�,e�O���O�@�$|�lR!���YʙаD�gU"�l�]y�䀽�O��d�)2ͤh%Fh��K2K���#U�i�y�T�d�����OJ������>�2I�D4x@
��ۏc�lH�&�q���a�O>���'Rt<��ɀ�x.��6N\�'�v�3�4�?����?)��%�OJ���O�d�n�5%���Tj�%��Uqql�p�`�D�<���?��I�ڙ(�PbblR�bN�bYHk��i����J�^b�������5��&(6�C�.5}J���������s*1O��D�O����<A��8I�EA�,:��}���c��L˥�x2�'F��'��Ty� ǻ{<X	;ҩT\�Ĺ���:U.�:�y2�'m��'��I�F�~���O'�0����1R��2	���9A�O^��O0��<q-ORM)�Z?9��ɔ�l�X]"�ʜ7`6�x�F�>���?����dO�p��'>a2զŵ���P+R�j�B�3�J��M������DM�H��O������6Ҕ� w���<g�i��i�2�'�剓?�fP�L|����i���,�UL���@��0@ˉ'"剀	r#<�OeLyQ� {BT�yD��6F:^m�ܴ��$�	�R<n���i�O��)c~R�Pxd)Ǉ��P�؇�Mk*O  Af�)�S�_PaQ�E�(q�R�sS�k͞6�_�%o��P��� �����?�j��h�m�D��)�jL�+�6cߛv���O>e�I&\j��g�F($�1%iG�	uh���4�?i��?�bh�.=މ'h��'Z���2�h�`�
���2%��-��OP �#��O����Oj��O���848"qB"�W�\tgAH�g���nZ�b�dJ1���?�������"���� xf
��v7��h}�*��t;�'r�'p�S�4��Oȫ��[��	�4eC�ϛ�B���aI<���?9J>�.OL$:����Z���!�,� �$8�aZ��1Of�$�O��$�<1�������<�^���K�Z�|Ȓ���_��'4"�|W�h ��>�FA��8"��g2f��q���V}�'���'��I1;�ҡXN|Za�~���	ц�=6�4�q�	����'�'��8Ahc�����͑A�j��!(��}�~�)U�oӆ��O˓y)��Ֆ���''����eHԬ'V|Ui���v�K<�*O����i>mH��ǒw%<	�u�D��~=��
;�M����?��,$��v�'��'���??�"��J��`%��')��{�DAئ9�'ޝ;���)3�LH�Ή.��q�Q�XP��fе��7m�O�D�Or�iz�	��6�#���q��*s,����F3�M[��\�����D�Q�? ��H��
Ҳ�كC�#!Y�kw�i���'xb��e%hO����O
�	j�.�Pv��
Z[�DJP:b�ܙd@8�Iޟ$��ԟ$����3����R�IJX$;�M���M��B~a��x2�'�R�|Zc���;�n̻Q1���.��b��؋�O� ��d�O����O>�R��Ҥ!��Hn��kvF�$i����@H))�'���'r�'���@|�Qdʕ&�p�؅md��e�&��۟��	ß̕'>5��n>m��~R<���L],� ĭ>���?�K>�+Oy��Q��pŃE=9��#�ѭt��Ycg�>����?a������J˦,&>�`!�5G�쀙hg�u��O��M���?	*O`���Or�h�?�r0�q��	T/��0�	������'װP�qN-��OV��CSsJ(ɂ�ÛS�t����0HnIy��'�R�ö�����s����	+�X��3ǃ��.L�"�i5�ɈEn�y�ݴ=b�ԟ|����D� o����3Wy�=��@��	Q��'3���j�O�xϙ	^�肷EH�-Z<Q��W*�M�����'N��'�$>��^����!�5����q��73���ٴKۦ�Fxr���O�ш ��5���X%���\�P��#�Zզ�������	'0����}��'>�DITdl,�D��m������pF�OhQ�t���O4���OR���Ě�R��3·1��	aw�DӦA���{�KH<����?�N>��J�<9y#G��Xh��F)�
����'�*���'����	�t�'�P�P�̲�� �rK܀n���4�	-�O��D�Oz�O��d�O�:��,u�z݋Q�R���E`�N�>;�1O����ON���<��E�8y��)N�.���Bf�um�t��D!^�T��ȟ�'�P��ȟ�Ƀ|�d��ě(s_PU0t�_�s�&�b�T����O
�$�O�˓ʂ��F��ʜ�WJ�٨B'hr|0p��)m2X7m�O`�Of�D�Oܤ�6 �O�'�(C�]˛������I립��Ο �'W�Չ��,��OV�)B0㬽	F��3{v�:o�>|�%������(�������'��V���`��*tɀ�e*�0���i��ɳhB�Hٴq�S����3����(�|!Y�e�w�a�'�ۭH�6�'�B�Ї�2�|��$*ӝeU�;�a�dx�`p͐��M�d����'��'��� �d�O�,�u�R5V��C -2eȮ�s�,���a�n@֟%�"|:�`�ly�c��.�И0���N ����?���?I@�#d։'��'��ÙX0l�Ɂ���G���5ύA�v�|Bl׼�yʟ�D�O~��$$ԍ��F�+2�ށ��� �[H� lZ��X*��؅�ē�?�������ҥ�%[:*��d	�7�!"%�{}�`�~
RX����ʟ��	ay�_�żq�f�+	���C�#���EPУ;��O���%�$�O����������E5:��%���Ǉ	�����OX��?���?i)O6�9� F�|JcbZ6�-H�,�C���
4�@z�	���%�\�I��|�I|�T˂c�2��`�ԓ*�� %	�����O���O�ʓN��:e��t�L/͔���S�5�ؐ��(Ӣ��7��O��O8���O81٦#�O�'k0T`�
\�i3r�Sf�u����!�M�[�,�J�$W���$ZP�����w��)�lW� P����mZ�_D!�F8� ���I��l�X����>+4f�p�y��i�Fn/!��I�D���17��=|�!���+?64[�H¸(�"��Z�/{�	U�&��\*a����R�Y�@Ϋ]���"M͢��Yp�W�#�lz�^�2��j�(�2�m��/˭O81�)��#Dզ'�(,D���nh��IM�MB��O���O<��LvȌ8���VlP� �(y�`���y�����<Ѱ�S%m���g�Ԫ{
2|b�HGܓ$x�%��#l�(0@r��XK~]����A���A~�#��?�}�	�$�	:"QY�mF��	�U�V�0Bڐ�Ɠ':�q�E�YId��A�F��-�'Ll#=�O��ɀ
��Aw���=ۤ���e���
��7F��a���h����I_w��'�rK�T����&8Ar�BwCC�\��i6*R�
�����)|O��S'��<����7Qм<ҧÈd!3l%SN�./0}B�Ȫ*�xDy��1Vh�b;u�@s"H@9{��;�Nc��igӔ�Ŀ<����'b�;�,��L��+i���O��ZY���	���\pB�l�/V���O�-r�l���'�����Lq�)�������3�V�x#��-but�	��ʟ`�ɸ]&6��	ޟ(�'��E�fbW5QU�u ���M3��Q/ԙ�@g[g�!�'̅y8��YD�M�mG�Ub�Z,-���oZ�	�\T���_������N"P���~n�'#��'��Q+�<j�x�sB��Bpp�E[���I^�S�O�BE���Q;j�N�1R�6�l�'f�6mȖe�Z�Ң�R0U1�� F��PK��D�<1FDM;�v�'�[>]ST̈ӟ,�CLޡg,$���>׸���g�ៜ�I3����k� D���i�|z�I�	Ś���	(�2�`�f�J��N1>�ݙ�FǕ%]05�C�i`�}Y1��9;Z��D���'k�hͺ���`�,�'јu��g��	q��-�3� �풵��V�d�+��Hr���A���O������ٖ�R&)�8H�S[�z�ax�2�D�7J׀�RI���W�`c�i���'`��bf|����'�"�':"�w)�գ��ՙ@L�QQDI��Ơ Zu�U5~J�-@'�u�*E�dt��$?c�؉w˒B-(-�5�9\���G�h���ע^��?i�#�+��>�Oh���S�mԜ�;�X�l��c���O���'.�}@�S�矰�I�\�Ec�M��E���"r=Π�d�f�	���	a�O��`˂7&<��7Dȗu:��C�OZ�mڠ�M�I>�'�b(Oh�t���)x֝Э�=<̀���3O�ŲQ��O"�d�Ox�d��S��?Y�O!
���Fۮ��≒k�nɻ%k�mlm�^�PG\�!$�ۥm�џD���.6�}��|)�� a޶BVP�b!Wyaɔ�V�9w>�F2-�u�����R�ID��`�߄.�|Dx��h�f�i�4�j���&��|>�a`����~�Q�f�U�y2ɉ�>�Z 1�͜�t�Z����'�
�����(8nӟ�I ]}�u2����L���@4�	���-�I�Z5lɟ����|*�eF�b��(q7+ �&��d�pj%0iJ�J@4a��.��x�?{*���C�<Ԏ�I�xd�d�6G�8�$��-;����%�b�'�I,V�d����Hq]�9���#���	�$��i�S�O}�X�;V,�\Y��r�Z�[�'�r7�Ħ_`���A��Ӛ��P�B��<�j,H��	ʟ��O���s��'Xn���odl���FşZ�HW�'�B��7b�L��MX(R9�����|
a�.��s�Ҩ!��т��q��D�h,���a�@M��؉����-Z���X%28��s�`(��Igpp�ɻ�M�3��?� �)
��t��cnE��@��U3����![n�æ�K�9��S���@�ax�D ғ���CcF4mL�a�iǲ��@�itb�' 2O�1pۢ����'�2�'�r�p�		"ǀ.	�� �,ĥ2�:�:R��	� ��
0x���K��]1w��|:��>���%��� řr����*L�6�C�ܩ*7^�Y�K6!����}���>A���/,vYH$�$<h�4C��]>@	��n���N0�"��Y���	���3��L=[�@P�j"����ln.m��J�nb�a��IʣF�2)�'":#=y�'�?�/Or18�o�H����a�>��u"O����.p��q������"O���3��	G��h��L%��!�"O@�Ba T ��D�J:���"O8��/B���QAję�:�S"O*@���B�I���ЀO����Q"O�j��`��C��p�8��"O|L�� �6�I��c�6��"O�Tj�\�֕A����F�`�i�"ODA���
_����:b�d���"O�!Q�������p�W$����"O�IrT���>���KM�:��)�"O�\Ð(��Vv������T�ƕz�"OL��7��*Q�`�R��˛es�l�q"OB��ïŝ<4�y3�Mf^@�"O������K�ԹvvN:�ئ"OXy��ٔb%�c�QK�@"�"Ot`
��S�i � #�[x[v���"O�
g��5�D��g��E�
�{#"OT���C�SN<3�`�1�+�"ODQ@�,ph�����T�Q�.��W"OV�0����<bD$�?H�9V"ODyv�P�u/H�J��r�`��A�!��T�*��a〳J2�*�]�t�!򤈮=P���.E�1b%F�T!�ę�aB1��g�Q֣�f�!�dڊޒm��E�#7r�y* ��z�!�d1 a����m�3��5k���!�!򄀪L�:!v��?�v��@M�< n!��	_��	ٷ錦H��������DB!��N3����M'>:��ذ	!��K_BЉ�e��'�t�Bi	�!�DH&`H��W�����P\�@�<)G�Xo?� �,��pQ�槀 ������V�l!r�㝝^��Ц�'Z�1KE-�)'8��IRI�RnVu��e.}r�r��|?q��K5n{�eQ��O�Fj���v�ңgDb� �k���{�E�ˆ>}����?���C&�:�.
�?���al��h�)���?A0�:���!L�I#��L}��.!��J�@
y?��_yJ~b�#@�Y����9o�p#�O�J8���ƅu�X=l�����(�	7�6Y��#.dwP�� 	L��'H��	r}�HU�`G��`@,��B|ŊF���O0�f遊`A�QM~�'JL$��2Z�� ��"2�@`x��T�_��D����`���
���HK5_�9+��M	2[Dm#d.`�U��/��b��ӧuO��"�'a8�S�-���GLG8}c<D�N�H0�I��,�d�6F�Y�3?Aa`=��\��GW�Q҈����F?AH����'S���OR��O:����E�
����k|Ӧ+�KA*\�$�|�'9�0�3e�����⤂?���AD�_.� Ѣ�$?���*|�		��3}Z�~r��@q�-(�\p�����
��OVX���7�YL~�'XH�Qq����b��f�%���T:Uw�s����^� 1�&�%��D8"�,�VO�{!�Ts��nJ�!��2(u��jYw~@!�=�g}��ȦK
�}(�NƄj4��T����@Y�F�Ӏ�BZ|��2�Ⴂ,�Q����+3glma��m���b �z:r�0 ����O�S�F"��b��6/xlk�+I���j0)m�h�v�	�-Mt$�7�QҼ�d��F�Q�-HV�zD��M<�l��1IS#ɐA�Ę(�gO��-�>�̓  �X��,]�d��g�\��'t�`�����n%�Sj֑^gV���:<�N��(^��z�[��*���G�J�,����|��J� ��q��,�[H����i=,OPt ��ݾ�ԩs�й)������I�z��V���0U' ���e0���*�(H8�lF���j��lP�٩�'��܋��I�r�X���q#��ߝ8�>��� ��u/Q����D�p!�w����X���0{�h�&0� ��A��t:��!&Fa��Ƌ&i�t��ap�i�L7�	< �)�A�I[���[�e��Ov4�+�.,D
a�	u��P�I�=f��l�
	c�65���TkW�<1L�)C�+'>���P*;���� �ĸrT�p��C+�
��7b_JX�lBu��$h9�r\wp�2-�&P�H��ig��rӨ'kS"m@q��6d�8�?)�)$��[ScB5* �P�)ګ"�Q��D{�O��t�A�7m]#��I�L��� GɎ�8W��R	Q���Y�;���w�viYk
I�J]����'R��<���hO�O<,�:��';����$������F����mu��(|F%���1P��&�<$���s�ڤ,Q�l�-�)lU�s��<9��$[�3�<e	eK�=@�E�ޕ++h���Y�{[\I���	�8<��᱊�i~�Ի�ͅ4Y۞ъǫ	}��?˓(Q:բ�%J:)�D�jS��"~z��'�V��Ѯ ����b-Z�4�EK���'>�ڌB�a�($��@7���y���ԧ�u�*�>��C,���3q����C��C*�D���OӨONq˕#���ʼ氱)��)d\q� �^.+��e{�S�O���)W��4�FG�x\�Q��J���T�VB�n�j�k�'��B�l-?Q�JԄ�����	W�Q\���?�\�O8��O&��禍���M-�(z!bҸ|RXũ���%vg�`Z�3I���#�E�Z̈X`s�'�8 3��:�dF�'��1	�J��@�j��*CI&x#)OP� E���$��T�"�­��剭K�	��(F�Ky{��"Nظ'!���N�=���?�N��|��=���Z�긨5ď	���#�΃;a�������@��1ﺰ0�.t+�u�b
=V+�����A����?E������Ő��8 䬫����-����"�҄�%�K9L�@�[S	y�l�'(�j���3�u�Q��q��@��@�ݚ�{���?��T�ֳb �RV�%����(5����)�t{��b�O2Lx(�PU�~b�I�������O�)`~kJ�.�UH����]��+@D�|V �f
#Jكŋ/�ZA��ǡJ��Nģ�ԓ �͓?��'�����\�)Ήg�B#x��(�M�/M q���wɬ9x�b�2_���P�0�O|�{�Ċ�W�����A_�S��+j�� 4��y�<��x�코'(�9��F�ɧu�'�@HsAf�6O����Rpj.q)����b$@IqEn�Z� ���dO�4wD+TdO�u֢1:&�^�R!�DJwo�O�%%�ֽ���+Q�c�N�P��t@��-~�2Jǝ,~�\�#�R��d��f�W�h#t���/�>�3}*�j�S,`�l��!�B>����P�~�@�ɶ(��I�T r��"�2��g��	ö�)u+��~�F<C��2���	�7���3�'���"Y0�['�Tk`oʣ�yZ0�Y#�Dc�'�a��g�C?��&܋7]�h)CLJ/	Df��@��J�H"6c'JE�䋐F;�yi�գ� ؀�E=N<Q����뛰���� D�:�3f�b�+$H�K)� y���6`O��q��1z72��e�U�A_
d2`DU� �s+S*6qO?�I�[�I���Ѧ ��a��d�1n�aĀ�_�qO?�	6㊬��-��
�� +%�D�q�ɺ^�H���'�*<ѧ��^����E?I�$۟'��I���X�'\�Z�=W*=����$�>��&@L�f������i���	A�b��/OϤ�������2S���%�)J>l�f'��A��1�)-$&f8*��[��>9s�W/L���+bOYxܨ��W�3�x����bvɧu�u��*B�nU��#��?��H�g��K�O�(C�2iB���I��y�鈘Tĉ0��O�|�OD��N�
0�@L
D��8�B� �T�^���~�d�C�R�x�C�B�3�I�-�6\ض��R>��kFo2d�ɥ��r�2f3�Ԅ��?���iT]ë�;�����hʐQx�=s!Hŵq<J �'%�M�'�����y�[`����Av�e��(��Y� кA	&�)ҧQ�艣 "d�ZF�:\r��N�O���
�3�D�@��4������D��(�0KV��"�����1f/��X��pܓ$B�I� t�g�N��$���NX C���Jk@\j����6HEP��I��z��z�S�'�4���a�0����2���-O���4��"7dn�js��cͦ}A��	\�pq"eÊ3,�̪��W�Ph�@�1�?��G�P���=�I�?����Rn>��Dl����`�����F�=�7��0�\�N�8V���$�9�	���3|f�a��ߞ��',�tA�E����;EU$������Z�p�f�� Hp��Fx޳
�I������h�
���d�|��u��!�	=��3�oD�)-���M��M�M>`֟�6D��=�zMk5��|��G�6}(�,,ic��q���)���N�T�2�@+wk��1�i��@*f2��<jE p��~p*
�+�����6`����` ̏P�"�-̨���	U���*�@�4I��ԓVcG�|���S�a��"HTH���'u�$ʡ�q�u�O|�I.mN�lڵ"1��#�^�Y��ީ"7�]I%�1zj�3���{��9Q����аx^X��@�0^d���5[N��Q�:L� �A
��$V���'E�
A���҂Ę�)��屳��9Pfc�l;rF���B"�&�h��֦'�A��N�^�� =U̴;��pc��ǋ3,p˓�(O��kw,��@M�W�X�@Y�@���x����4E�/�`�C��Nt�ȊC�	���!��&]Tء�F���qT��0M�Rla�GQ?�Ҥ�P,S�N�c�MY!�˅�z��F\��u�\���a�}b��s�,�	�+�.��TCE/m�����m6����t�-nu���ԭQ�=�f�`a��ħ��q��xuϟk��q%�� @�h�`�^�w���n�?b�|Fy�'`��i�d�N�w�|ux��F����C�D1.���	��K�G��[b�R(��� (�M�<xS��7;��h0� A�O�xli�o5z�OZ�YDL�>N_�1���#D�>|�7��a�T����~PL���Q�j������!=�>�
Ó2Ty�N�_V���6�&<@��[\!�0�40��9���#t�z`K��2iӚA 5���wӸC��d�� �4�p���;��Ҥk挭3*�R1)E�35~p2��>Q�jB��j��` U�4m��iVE��d��J���1j�y3��Ti	�!G�p���!��7Ә�J#E��$P�O/�'�d3r*�F������%�Yc'r��Ei@�Q���>S%��!�A&�2Ax��*�
+M�>��lа/��>��Se��p�R��	Ǔ,�I��B�5mz�(���$P�t�zB�2��8��� !Hֵ�w�wS�lЃ�)R��&����t�CwR�N5L�{�j��p<��55:�2�灊�ļ����z������VK���I�[��٢���>O
�h�ԫ!�E����O����������?��ěD� ��'�Q[3�2?��	V�_�:Y��n�~���z�a�'8bT��ut�D�!jSA��8֍K&�ܑ�'�]"F�`�`H|�	:�:ql�"y�24�R�X�R�4��h�>L�-��"Sj�D(���
- VQ�ǌlޙ�b+�3+_�`���-)��)�񎍩Kv�9��e&����8��{���45HG��!ܠy�l��8y���e�I_;�hh���=b����$��BĪQ�N� �}�K+M��*�&���L��=}��8�Z�j�O)�2Q��:;QR��c��*�$����S����-�i����y��$��|���I$`ְ1���@36��j�J?��>�b��	_�E�M~�'E�,!�BG�+U�A�͝�$i4$0�'�t�'����2�����S�A�������p��|8U@���]�5��,7}pI���9�#��sv��Lm6��E�s?��k�ny"b�^�L�ֽ�DCo�b�<���ۃ*	��P�G.WJ�ɋ��kD*�����2�D ������L�9M���(�ER?	ӕ>�{�dև'��hpR�����1��¨���2��l(����>SI*����O@��^~�mFK?������Qe�߈\TJ+��	 ���OF�O������C|1��Ɂaޠ����!%�<A@c
2Z ��/�(+�:kА��(~.�S�����S2��}\9CӮe�~B�	�^��b�e�$B{!&�!9h1�o�X̖'�r�$>�
E䕸l��ɗo��F
ٮ�E�plXVB ��D�o_p!F�@�oQ�)�mC��XMr`��?b�U��'��Ez�b�#[4�E
� �	��f�p�E��%�0�H�I<$��Hrǭiyi�M�l�(�$�wK|x����#a߶���Ɩ�"�!�C�BqqɆk�1N��ِ�c�IN!�A�)������-M�lIЕt_!�dF 85���BA�Kp�)C�&Y!�� [ʡ�W��J�K�E�sX!�$��EsL�R�nW�+{��{&'"!�	�-��Ѻ����x�v9w��7b!����L��ש0"z�uXD�!Z!��R�s(�i�6m�,R'$P�5!�M8i�����'b����դ�!���F��+6�V�GT��Q#݀9|!���9��(���_%���!����!����ݱp)��h���KDU�!��e���X3�ʛl����`	.�!�$�(딀� ��	w�&eQw��*~�!��I�V��(`GL�=��)e�ڳ{j!��V�f���IX0
��s�"{�!�D��<\Q� Y�u r@i�N�6�!��]%B$@�!Z�5��q�W)!�_4�H]���=�,e
A%ؤ(!�D�/2�Z@P��˘U�p1� �}�!�DR�_Ì��6�V-S�d�
sF�!���I"�8�L��*��G��!�/�%I�i�<x���P�8Ǝ �'�*	����7�ΨP�7[�ԣ�'��[Ṕ;�bu�f)��8�'�(16W�A�&髀BB5.�ZE��'�P�:��7p3�J��̄yJ��P�'���R6-β04n� �Cʍf�.�8	�'�4 �&��>	Z�#�-Z�u!�'cxR�_u`� �+N�b���'dQawe��M���"�Ƽ�Hl9�'�ΐB����K�$0c�a�9	��D��'��y��/F�!�8x�k� �����'3Vd�'�J'h���a�~
`�
�'�z(P��߾r�qc��H�98�

�'�	r���"� }	0�8&����	�'z((�3�V?2!�X�l�M���	�'h|	�������V�"w6�i�	�'@Ա��r�t���ߞr��̐�'�uI�Rh\�0H�"^�o�@�
�'�� 8��*`Y�hr�����}��'tX�P��EK����O?]��I�'&^��)�)8��bF���~a����'8zh*��$ >��J5v�
	��'1N�Q����j&T�J�!

ri��y�'E,I#��M
	S��a%"�
�'�@�D
c��!��RU�d�
�'�4h�F����p�%7`J�	�'�s�\ b: ��}��H	�'S�����ٳFcb����(v��h
�'�`�9x��!��f
�݃�G%D� ��C#+�P�+��K){	����)/D�p����#e�#N�]���-D��ڴB\�OޠX�@NP��PP�4�0D�� G̚�6�\���v�a�C+*D��q���]�P�{"ƍ�6��ȃ��'D� y����jln,[C���p!s��%D�H��*]y�Hq� @�v|��H.D�<:�H� e���#H��HL$)���8D��Zg#�R8�
�`L$(1�Ij�N,D�XH��6�ۧL�]Z�!0D��k%f�&I�p�Ԕ�ɰ�!D�� �h�PA/(j���h����"O�e�C�6w���T(�cҙ��"Ob<zCc��zpx� 2eѰkJ�U{�"OZY��h@�sfmrdj��@)�"O4�A'�B	p�AAX::�0�3"O8uÃ�פ�@�& ���!%"O q���4 �)�r��P���"O��Sȝ�@Y���N͵R�T9AS"Ofp�䐛l2�hV�B��!C"O^��@�~��`��R�!�Z��E"O�ٲ�Q�Z��h�b�!x�lk3"O��dʅ%P�����$�+v����"OBXy�
��OApdR�"	�$$�9e"O��s�ʍ
�`Y�
�8�[""O����H9z�x5`ql���F8#p"O���/F>;�t{��B'5����"O:���
�9�Mӳ���z�8p��"O����C�n�pEY��NT' ��"Or�p����{�&�'f(VК�"Ot�x$��B7 ���W>�B�	4"O(�z�̗�7\8�6�9D��k�"ON�[�	��'���#�b����"O��m�9����Ȩ(�~�{@"OB��2n��@�4!�'�@:���:"O8e��6G1~Q��D���>�37"OڜKb���ez�p�K &�DP�"O@�X��
t28A�ʍ-?�n�)"O���6��(5g��iH���w"O�	�� &�����h�	��"O���c��J��0��O�W�5�%"OZAI�@K9xHpC�45F��""Ozɨ�*�.,�b�!Ƨ�*%1D���"OE�ǉ6Am���̄�R����'�qO�)�!!T�(�t|y��@!�$J�OH<���ҳ
'��[Q��ti�u#��Nd�<Á�	��� �Ӽ0�Zy!U�{�<��
2E�@���ȷ@?�TA�+w�<�VO� 0cB���)6J��dx`�]�<	�ޤ=����a�;���d��N�<�5lG�/�"�b�Ċ�"���CU"KG����R�$��&��T6�8@�,A�x�pm��x@��'�'}�|DzH�<&,e��7q$c�h�U0
i��']�jH�$��#��&�-²=
�޴�4�ȓF�Z<B��(��E8V�IV�����B≍s�JЀV����+���p�nC�9+.z�R�ƛ��>(��+�B)hC��UR9�A�P�J����02TC�	�*QN�"����"��	t�P�&"O���� ��tx�ʧE��"O2i� $�wڦm�5�m��(E�>9�U��a+F�ܶ:�]A�U�ﶍ��a�\�!�7*��`E�s�)��+�����1G<	�PnS�}��ȓu��Q�FO�y����i�+k��y�ȓ j�a�씍6�����$���H��P�`F�/���iV�H�{���ȓ@Vʤ����^:��Q��M���5�ȓ�4��%� 6�a�+����I�<1�'/ʴA!J�!p�{уE�;�A��'�&Aj���Tw� p+X�-^X$��'�l�)�%D/�P�y'L* ���{
�'��hW��x�lP� O�D��K
�'��� '�. y�M
3��D�x�	��� f�j���T��M�e���R���!��̆���9��H��"�Frtdb�C޿MFC�I�$|�;7�d��@���%�,C�	�x���PeC>�rV�ݣ=s�B�`ht8�MM�(Ȫ)��C���2B�I���!{S�Q6~9��S#e!��C�	�>(�|�q�9O����S���@��B�I�'��)H�ͽ#p��D�ɵ[�B䉶.��5 ��]�C�8i �k��1pC��}���h��<<��J �B���C�ɹ@FU��j��8.�Q:a�_Z�DB�I-;�����g	F����a B�ɓ,��R��%���Y� �2<0B�	�g���8H�*:ry��+�=:�.B�ɶb��D@��d�y�HJ�F�XB�	(_�,YD��P���@�	�*�TB䉂�6�f�%HMR����% B�I!�z$�#��+8t���'C�h��B�.Z���.��O�@����%d�C�Ɋ	ʑ�R ���b	;�xB䉋@.M��fY�nͶa����;D�^B䉇&��#7�1Gf����%��C�I� ]���	{tu��˝h�B� ���J��@&J�ܼ�ECJ�<�B䉼<�DlбNN�(��
�.�/S�B�*�� [��ʹ=�~����(t�B䉛-�E�!�S'$
�1q�坕z&C�I/xrJ�w�|�p�Fڕ$/TC�ɨ;��	
3.�%Ș�g�>C�ɉv���CG�;G/�yX�g�;'�C��{n�$f��)K�q�s�� t�B�	��3s��Ok�9��.K��B�$|���C��
�]Pt���B�I3�D�R��ܞ��L�B�nB�IFwtY���,;�9��Č6�,��0?!�"����	B�A�/"�鷧Z~�<�NX�2�M8�$Ն]a0%9"u�<Iri֐x�h@ZR�V>t��Ć�[�<a�`�(|#� �Oɶt��` $��W�<���>8��鈄��m\���p��S�<Q�d�/�:-AD��z��O[[�<ѡ�+B�����C�9#lTkv*"T���$��7�P�KEN��Ȭ���7D�샷�ѽl (r�����ɚ�8D�a3�?L^���J[)kۨ-��f1D��Y�"�>W:���r �_ۂ�S��1D�T ��יE�L�#�n��T�|�!p�<D���3G�<66��)�Kf��Q�C-D�4A�gM�s<2}�P!¯L��$�r�,D���T����a�3�8f�Dʤ- D�\��m2�|x���Gm+�邒�<D���I�?p�l��AA�mP�Es�(D�芲�G�o�:�r#)X\v	"!�!D��a�(�dcle��!�-:�?D�4����\��Ǡ�n�p����;D����^�D��Y���ݠ~�Tu	#"8D��;�gF��&�(��	tXNa��4D��d��'O,�B���jvB��eh'D�ػ`́�(�d�+���-X��@u�8D��ҁ� ��a��7��T(6 1D��3��}}z�I��)/����b�;D�[7$�w�(�FxP��H�5D��B"��C�~0��_�*Ypz C7D�ty$Kӊ&�B�'�2gj�P&0D�� 6%a@��[��P�Ӭ\`�""OZ��l՟zG�|��b�;{g"O�=0eD�"G��tpĠL.7���'"O�(�2�Ƒ3bJx���-^�pekt"O4�r0���X��x�G�F��$�"O�(p��`�x���%fʐ���"On4�+I<2�����
���"O�DK �ɉ@� ��'�J&h�P"OըP�1@p}U�\4sJ���"Op��	��z}$-@,N~�m"OV����9JLX)��B�y��k"O�l+GNbXF�kdk�?`�A"O�Pd%�`Bld��	���Q�"O`D0S#R�>�re�"���;�"OD}떀"���g
�7L��Y"O�l9rb	��|�8ŪL�;��AC�"OA16@��9:H��G��9k��I{s"O�
"�X�'�"\I��L����&"O<�s�@ �.��ؐEW�pX"O�S�i�0ja��Ѧ�����"O�	�V�]�~�x��I�9��	IT"O�0����9�U�A*͓XQrt�"O�!ҖjU�X �	0�P~@J�� "O$E ��5��HJ�ÿ;=�D� "O��K�c��;�zpc�o��&7�\3�"O[�Ӈ�<�F�XƮ�S1zpY3"O�0`W���g�xA�ƙ	��,�`"Oz��C��0S�r@E��� �� "O$z��J-ePH݃C�5G��)`"OLA��%Y�b`35��~3�uCr"ON�Fl.\��u�2�ޤ��"O�� D�L�wDIB�d��m����"OvtK�nW�q�xa�☮F�<d8�"O�D�7�8OE*,��	6�|A"O�j��eTh�oѨ
*��""O�= f��Hި�³N��UBl1�"O�P���oh�\���I�eA��r�"O� !�ߋujt�3Tm�g��AE"O��憜%|I�s1@�P "O$�g�+'h�щI 0�c"O4�A�O�#u���V�U%� *b"OyZ�̚!��&i�:$� ��"O&�YS��5a���A�27x�J "O�}s�k )�dQ�G�+6ɀQ"O��#�n����cC�����"O���I��p�b�ߝ0���R"O�cF(�
9�x�	�⑫w�8Ґ"O�P��B������X��Y�c"O~A��R&�ƴ�`�ɴ&t�"O2�9S�,,�5h�N��	�gI*D��(���C���%�_37��1
�
$D����*]�hX�yڧ������C4�y�Q
*.H��7�J�A�$���)���y�>/{&첷�V9fl]ZRN��y�#�5��.ּ'� �)�AͶ�y2-
sb�0��E�!�E���y2 �I)S�d݃h)1��GX��y�P^��Hc$V�5q�d�1����y�a�"C���bf� .9ʘꑂZ��y�_{̖ݸ�� AFu�` C�ybl�/��chUUr}�,Y=�yB!��x���ce�ǋ~�~��`BX�y���i5h��b#A�>/i�׊���yB�̙h��#�Ґ������T�<� x�ʑ�M�T�XIs�f1u�e	C"O��Yp��a8�+��#pH���"O,8�h�<vr%;v��i,\�9�"O��O07��`��*��Y|6xr"O��PJ�jx��� �Z��0�"O�,�� ��Ԥcfa��m��	��"O���G톌M�hMg%�)5�BU"OZ�I� ϑ?�zlBUB�mi\��"O&��"�;4�ۓ�E!�2���"ODUp��=��ݕ{t�R�"O��
�`�_�l�����;m��DU"O�dBS�G
_g���G��w�L "O���eD"E��5Gr*]v"O�%au��7<�(�H��\t��"Oޭq׉ؤj�FuJpG�TnZ\ �"O���al[	���hW쒋vP���"Ov�������!��,V�n��"O:x�BؓX�)���Ҡ7|�ܐ$"O��bGX��+7��sD.��"O%suk��s�?k�)u	!��N!:  ��7�B?���$�>b�!�d�0�� �G" &�n�!�!�$�R���Q����~��!+�m�,8�!�dD�P'~ ���ӂP��\)�lּ�!���:V4Š�]��B�Sd��!�Ѣv�r�h'#H�t*��Y�M�!��{B��;6B:o�&4łֱ!�˶>�Ea�b�l�������q!��(�ԥ�W ��ʚ]i��I�S�!�� `[��e��s�`���s�!򄗇x�k1N�$� �pG홻.�!�D��L�^����N�@a��i�\s!���x�8&-�=;�$B�ՇM!��%�9��c�/�6�2�ҙa�!�d��|�D,,e�J9qӬT%��l��'��Q=Ū({5+Ϣ��*�'��xY����Q��rXX���b�<񂦒�?���sBdB���4�Хb�<�WŃ$Q=r����Y7y(P���^�<����"&�i��	6t�`1q+F]�<�w���ī�e�\K�lH�k	^�<95��4@l��"�P�w-Z��v�JN�<�p�+sA6�8p�2�r�*�)�F�<!f��
�V���H/+D j�WF�<��jF�v:�Y+g.��(*����AZ�<�FF|��ArO��J�q�A�Y�<�iQ�"���Y�_�%��|�<����'58�@��ԯ�\Q��!O�<!$��\� p�𮍩�
Q Sc�<م�W��"ܲ:�Vģòq&���'Oܑ�i�N�ҡ	$ބ"/ȸ�'ꂝ���o�ČJ1���'tA�
�'��E��J�CG��@��Q:6��R�'�
I`��3}6:��� SfFp��'��$A�n�"�1WiQ;4��a�'܆Pچ�݅,' h����4C�L���'�Mh��,Mfd͚�@U4@�Ȉ��'������tqJ��
�3In��'#0�Cu�د+3��ꥯ��:p���'K�{�G�GgTȴ�4{ߠ���'��L�Dc���e����Dx��S�'T�s�'�/c�å��?mX�Z�'>V�����4SOj8�'";8@ !K�'o�h@%��!Gv(j@�@����S�? v܁��Lo�d��N�_��t�P"O-�dn$���#'|�p��"O m��S5~��pP�N��)m�q#�"O�!`���]��{����Y�4���"O��b�ռ_A��P�͞�]�v�9�"O���&�B1Rm9���	������"O�%%�R�Y���遉E�<��`�"O4�rꑛ<���*Ǹ�L�����"O�;�G�n�H��צ�	l6n��"O���
?1SPl;#4Z1P�"O�5��� �C*�p��a�**1Z�"O�T����/(H���"ʮ~�("OlDA5G��|۬m��P�~��M#�"O`%j�+\w|�T��B��<=1"O�"��U�n�2L[�G�01�ZAS�"O^����;�-p�`�s���"OD	�Wm��C�XI�� o��E�"O���	5�x� 6��t����"O~ �/�Ir������3��	H5"Opu���Fl�5  Έ=���a�"O��wI���D���A�4E	��k�"O��q��+E�q�6�� $]����"ODؐ�8�z�2G�g��3c"O�r�A�-i ��E�����"Or!y���n~�p�4?������\�<A�
����}K661�HR�*@D�<i��%-s(*�"�w�����H�}�<1W��ID$�!1W�{�2�Xu�Nv�<���׋���0�(X�#�&dXe��r�<�D�p���Rŏ[�2�)�`,�p�<QC�?Gt�ywF�@���CsD�f�<�� ��AQ$��#*�t�w�Sa�<�W�]Fj �aLWd��x�(�d�<��/�Gv�M0G͚zB�����a�<�I�(WV]KQK��6A���F�<�G(ׇ�A� FT�VXe��BB�<Ic	K=�\�r�.���dd�<��	�#�l�Z2h�<ت��C�<A��F�<N��1eɒ��B��g�UZ�<y���n�`u㣉T�[��PZ�"�A�<Q҃^�����V�}�|�ADz�<qՠ�7
���5/�,K�ΜQ"cVo�<aJ��\X�(�t����h�<��I
{2�`'��Ia�����m�<т
:�E��LR�:��Q��Fm�<�Ë��R����LH��$����_e�<�FJY�S��E͊!f��L!OH�<� m0�� �%�V��a
���A�<���&?6t�����|��B7��<��b� �zX�� 9JA`�s!]v�<���P2�@1����f9l!� �t�<�s�Е1�=�fb�V,��1V�z�<�'kM4cj��3ҸQ�����Ry�<	7�K$R��k�aj>9����t�<�2��#'���	�$��3�����q�<qC ���(�e��ႈR"�x�<a��_�?�\jVK��y"�j�r�<�(��2��|HVH�,qF��%��w�<�gg�"���{�
�!i�����Yu�<��Ə�@�}ӱ�F8RgP�0#�m�<��㓜$>�eᶇL2u&�����q�<aaA_�xb�Y�¬Q�v:8�+5��q�<�3���".��r�08^ذ'�Cm�<�2#ݳI��sp% O��РvI�M�<� ��;S��9T�� ��j.�Ȱc"O�QLD�& ���ݺm'�""O���'J�;E��: �Ԛp�zaR�"O�l�4B�Ry��s�$�	Ď�q"O����Z9�"U`E�g��q�'"O��a Z �z�� J�$�rxs"O��G��=,�.��D��3��y�"OM��)�����E��t��"O��R�Ƌ�ك�!��m��"OX�2� W� ��e�J��2��{e"O ���Z�%�-a�O�$9	X�`�"O|-8�� vq����Џ���9�"Oސ�!kA�'�,���JU�H�z��p"O�I�(��^uXM	P/`֔���"O̤:U�� .-`Cw焀[(��"Oz)��		4K<�ȺDT$ ,u��"O��p��N�[�Jɸ1�P\yn��"O@���s�0�R��*
��Ɂ"OlQ�f$Ę���Ü�I����"OPe3E	��A�Z�X�&w�l�p"O�5B.�B���:���	rhNHa�"O��'�ֈ2_�J5iA�DGpB�"O�\����+PI��I2�T�h���"OjlA"���P�M낢N>W�(���"O4��U+��z�&�I����"O�l2��#\r��0 �+�$|�c"O���Rh�q���ۺo^H�`�"O��sP�T:j/>���$��	Xrm "OX�A�E[;?����$
�5>�"O6pZD+Z�  `a;��ǈ#�5��"O�C�#N0�pH��\���8�"O$�{Τuj�٤'P�_Y�z�"O�Ԓ�G2�b� b��q�bu�p"O|a�q�&m@�m�8�ԕ�"O,��'�T�u� T��U*[�Ҕ��"O��"�k���"ŨEaOP�|`RS"O���@�W�2h��Tt}����"O�@KdL;��g�	��S"O�kgl�{y9x��޳U��� a"O�4)�k�9<�I�piؚ.�nBF"Ol�qæI�uRZp�@(G�Y�°��"ON�9US3y�:�p��d/�TAs"O��q�ް.�.E`�h^u@�!"OL�(4��?Dl�U+^6�e��"O����J>IJ�	RfՏpR�"O6�{�(�_�a4E)j�J<�"O.HZ�F̋:�0r�i�) ��\Aq"O���ɁMCT��hxV� �"O�Uɗ��=��Ȓr@T!5EB�"On� ��לeM�a�V�U(@%v�[0"Oh�����\�(C�V����"O~9��+��&�Sj	�G�"�!�"O&��bϊ'�p�;So�'@���h@"O�H��-(ǰ)4d@�w����"O�"�
D�\۪=1F�R(v�8!"Or��
ʝ|�XpU![5iҖ%��"O��Ibo�*&�<�@�<3Ɏ��"O�))��|��@�`�G����"Oly�@bY#�`�	 �%�<�y����Ԡ��j`�š�c��yb�IX��%CX�
E��U�E�yR	������]�5\�T8�y2��z���aj-60�cT.C��yb��(G����@њ0�Q�� @ �y
� P�Q#Aܨ nv`(��7�v`�"O�@[DMm�:�S�g�?2�d��"Op�0�BP�"��]K�	�f�� �A"O�}�BA�w/����ӫb�dݒ4"ObjW��Z�VUiq������%"O�Hw"�,.�e*6ᑫw�|�"OR$Bp:�pp3�O�'G�tI"O~��&�B-�}I���8�P��"O��a/Y��t-�a?X���(�"O�dbj�2#N�i��ć�m$v�[3"O>�h#W�U�Hܫ�E�<r(U�b"O��P
%f����fڎMEBA�"O�(���<4�>'�lBL�2"Obi�E"��"|4��F�F���2G"O�1zR�f~PC���*?�3�"O m���.��4`֥��a*2�� "O�)�S�R1WY��뷃��o��"�"OX ����B��C�RB�a�"O��J4C����P"j�4oP4X��"O4�aA��ft�J0)�����T"O����\֐r�j"X��S!"O�M@�e��(&x��T�D�_�K�"O����ꍀ|tb�3 �\�X�t�C�"O(%���܋P������9���AD"O.@�܇<5qR���*A�]+�"O�Ё(ҝ0Xx�x	;,:��0�"Oਁ@�)e֬�k�!� i6axf"Op��p�$>Vn8��ԛC�²"O�\93��n�����W$+,�hP�"O��qADO:��Dj��N�o�v��f"OR�	S�˭uh	2��i�<� "OR`Q�ޘ��BUJ�<ߖ�@"O�rMWo��%Q��+o��|0�"O�L��㏘@����SL�i�6%X�"O�Г�շi��|�0�=r��Th'"O�P��_�~!�"̣WX̩yQ"OT��#��VMx���<A��%"OȝC���vrHT!�%����˗"O©l_�ز$�H#��ո$�*D��0E:>�p���Z8?�Av�*D�Ȕ����h�޽-xH1�r%)D� �QHŽ`N���M%\")p!�9D�䚐�ִ��yf'�%���F�8D�ly6��=D�`eȴ��T�`s��9D���ΥT6�3ֺ��@�5D��p�gS�*���8 �C������5D�`
dm�%1!�`���)��ɠv�9D���i�����R&Sf& 30�4D�ĂG�C�p��\�Q����L�0D��P�_�;���ᩐ%��ac�)D�pj�k^�0?.x�!"t� �Y)D��ˢ�M.7�0Uxv�HbN  )7M,D�DK��T�=�f�
#�  L"�Ii�*D�4 �n\4*5j	ṍ�8�"q��#(D�,�f��g�J���^�Em� 0�J&D�d�V�P6x�L�2��] Z:Pe�%D��i��z�譊������5%D�X!�LA8Z=�Y��n�>w`Z��AC!D�� ���V�Q0s%�" +�q�k D����Dcb�0g��9��%�=D��x��rat��$$��}��C.D���S��!���I"��p���1D��2����ek��ekw�IlW�R�!�D�y)�Q��M[Z�2���
Ԃ�!�� �Ly��1J遄H߇q�f�!W"O�!��eY; ~��eU?�d�9!"OpA)�H �PV�b�nl��3$"OxDC2��)�ڥ˅���4n1#"O�uم��=6�x��!A�H|P��!"O��R��s&4R�τ�Vf�ؐ"OڍAUL��4ߖ욢NiU��3w"OZu���:B�f$�%.õq>��1"O&��u$�IŞ4�tϒ�$+4-��"O�\Hp�B6X�hY��B�a*�m�7"O�cѭ�(	��y����u��X�"O��i��@>yÀJ�-M��u��"Ou���{9�slB*D�D�"OЌC�aP�
��u�S�u�p�!�"O�E�����YC�XUO@ �y���1@ED�0A�4��N��yb��2������.�ڭi)ɿ�y��Ĩ�|\Kq�)w}���0�F�y�j���<�cI�lRd��d�	�y��7~�&�Rł�j���[��<�yBiQ!:��7j�h-�����C�y�(4����Q =a���JUH���y�O"wx���ԐT	�u�O���y��-� �3	��C���Ҷ��y�@^6�)3�DϮ	� �6�7�y"��"<�]`�C��B\�&�ɼ�y"`\�/X��1�z��if&��y"ܲWr�*t+J�;~M� /^4�yB��<K�r񨱣���)s� �y���cf��b$Mt[���'���yRj�Y#�Y���T�l�&5���%�y*J�2�8k�	؀/����bT��y2��a�4���2$��X�h��yb*���d�8uhY-x�{e�V��y�KŞ(�J'&i0�X4���y"�ȟt)� qL�v܆QB����y��@�@h�\�BZ�i�dmҒ���y�OƣM�Ȝ�����L�q)�yr�ֵ^��`��B �����8�yb�����V&�5���@�� �y�口7�,�)���  :=� h���y����O��໵���@wY��L��yᇽ`E�����;j�rd*�)�=�yR�� Yk�hA %C�a8da��%�y�I�Bu	P�S��Yb����yr�@+�v�pDF��]m����b#�yr�ŷ<���r���S���q����y�T�lu���V���bԈ(�'��y�ԽD�,r�bU0$lma�$�y2�L*t�
�:҇�����.)�y�kk����"L�z�@�Y�D�y��y����'I�oZ�q!-[$�y��$RʧDq���a���y���$`��rAYPL���9D� Ƈ�g'��@��T��z���!9D�0�3�+�|���,N� �<(�"8D�Z���k�L86��)U�B�I�~D��S�L�0y�	@��`ܜB䉙\'���e;ơ�4j��B�C�I���ه��	m�Q �J#l�B䉈@:r�!Q ɴU-j)B���y�*�B��HҲ�]�Q�~����ڀ�PyboBZ"I�B�ۦ,�\���x�<��I79���*�	�d)k��u�<� ���B(4����e�b�"���"Oh��㢅.GSh�AtϜ�9�6 8p"O 	+c��
t� ��쌚)	5B�"O���wC��eg���E��wV�j�"O��u�
��cU�W1oK���"O��A��byd% �j�)-E&���"O��B�@_��!:���Q����"O�i��.նM�$��89���A"O��P*&ے�kE'�42���`�"O�@�d�*VXg6F�"i�3"O��"挝(3���3��Q
�1A$"O��c������W�S6<9z�(A"O�Ჱ`��t^����C��ƱJ%$%D��p�_,V�����CƎ�X8zB(D���ոTU&hD�-=P`�O9D� �Q̙�t��� � �b�s`�8D�8I��)g�(��-�*l�N�Y�3D��[�	!*�֠!$��	6���;��7D�X�b#[8O�Ap3�Z� ������4D��ks��4B72Ya�d�$xĈ��\�<����v��	�&�δ*��5��\�<��LR'a Ju�˰1����A��|�<�2a�)2F��u�۫H(hq�~�<)��D� ���)r��[S��y�<�`O7�*����,p%RG�s�<Ѣ "a6�+��Y�&�!;Py�ȓ���[����Y���Lq�$H��4刅k�D�D$=봈I]�x��R�̰���l�p= �i;��u��q�,��\�YƐ��oCg���ȓA���)��1GZջ� ՄP�� �ȓ7�t-ᱪH%v9���e�ʼ�ȓR�J���C�~�E�K�w�҈�ȓS������dw�!��ܖzY�`�ȓ*W�$p&� f~��FMÕ'��A��O�N�ط#�~"�� �7��`��K����q�K�^"d�8֤�1z��p��zg���T�U�8���⇃#O'R���r_�THRcÇ�<�j�O�_� ��ub��"3�UJ���I/F^��ȓBSb�*��E	�h�%I�?��Y��!ԢH��j1$�� �׽?��ȓ@0�丧F�8�B�As��o�H��ȓ*l�d���\�x������{��I��0�`�a��1K�.X ���,8�4���bWHe�%`��{D�IX���ȓu�8����\w���3G�"
�zL��f��B*�7+�HL�VH;����ے�sb�˨h��F�L+qK���ȓfl��a��JpE�ǚ*PN֙�ȓf���{vf ."������P$&�P��H<̐�	�w�l�2��A#L�K*D��IP�� }��@!-��`��؂�	9D�(�d��-��1�����1W�$D�$B�%R�OL�|W�G|��I a#D��p0��4yLL$���g�T���7D��	CL��
\F���拖w,���E0D��� �+6������Pd���-D�|K�K$~���u�ѻ[��Љ@�/D���G( o<|l!�HU�h���.D��іE�"r�Qv�J^�37:D�l)!�\$^�x�/5�l��b%D�0�f��t�X���l^��1��#D�<��Hְe9�a���
�Ekv� D�� N$�����T�fdHK,\wҝC'"O��Zq�J1pg�Dx�G�<OR"���"O�T� l�+fP� z� �r"O�q��*�fO��oX|�H-"�"O&� !Ĉ�*},)Gc@Mߪ�"ORԘ"hN=&�����@���;�"OZI�q��VR�R�/S>9�H<{�"O����OJ�LH��B�{�����"O ���ɯU�^�ˇ�[-E�~m�"O�BAM^��p�t��<l�$��@"O��H��P:��pp*�?N�m��"OL1B�K%z ӅɈ	��c"O�h���/ ����I]!�"OX������j2��)�+�E�p"O�8#�Cq6rg��1��Q�R"O�2E��u���v���j>{P"O����%\�\��`G\�,��h�"Ol4q4B�.Im;�fD:Fx�"O��T�b��aA�FX&-����"OL���j�&)��	8��U�ݸ��b"ON��(E��Ƀ�$הe�� 1"OnC �,��2�d�$m�Y"Q"OȈ���:I4���UM��ײ�p�"O�9P��(8a���ˊ5��y�"Ob��	 `��A bҾ	,=�t"OX��i�Z�I�T���j�Q��"O��2D��� ԭ*�m�$W0QQ"O�� &E(Z�l��͖_VXy��"Oֵjs��ELaQ�F>3�H���"O�M��Q��aQO ~>f��"OtQV�ۘ+�R����IU�l#�"O�͛�녛k�
E��lS�Qz�8�"O�8J�"�6m:�9�eƷ}����g"O�,�|�UIV
~9���UB�!�d�4`�b��W#�9�S'��h!��J$j(H��2O$� h���f!�B(#L����-@���b��6!�$�|��E8Ƅ�+��@����}�!򤁤K89�&d]'	N���a�<e!�$�\p ̉&k�	c�Hq���*a�!����b��?"�T�*����!�$��d1��'R�Z>����V�!�$!?6(��٘N,����ǔ�
�!��1���q�1 {*�[�$�]�!���FX��C���`�J�EJ�<�!�ڔkQ����$l�(ye%��95!�sE��teӛzÜl���'PD!�$�2�-�h\�|��m�MP!��܌;lN9*!�J��~�񉘧?!�d�(�dlrCW
 �4HR�)��D3!򤆄R�ʴOM��(x8V�Z�I!�Dܸ2��H�%�=m���h��K�g?!�$��Ne��g���tі���V'!�$7�v�؀;Ӛh�Q~�!�D�o1.J�`�;;�\M	��*�!��:+���+�DԤ4�8]
��~c!�DRE1�� ��4*����w]!�$�$AңU�h� ��� @!��<���C��<��%���%WF!�M%c�`�R5���p�$b& W2!�d�B�X[�&��b�`ȸ1F��I2!�d�4k�Z����ۯu{d}�Ѥ�)!�䆚�JY��b��OdJP�qcſC!!��Q��Q	D��\W�� "���r!�� � S��T�D��$@ue]l��ڣ"O���7#��=��) aOOV�����"O����#Ċ���xpV�tn��"O�tK�
���3�)�`�kE"O���4Dڪ?����q��x���K�"Oh٫�i�|Yv2���I�4"O\�C�͜2)s4��(E�
�2"O��f �,	�,)1M�{T���"O4����I�����4�F�DT0칣"O���PP�>xH9�f�PK6ܘ�"O��C.�>�EsP�<IH�a"O�����ޣd��,���ؿN�Ѻ"O~!�1A��O'��*����1�"O�%��ՃY�DCpX�E�8���"O���.���s�c�7�d��0"O�<���D	�d�1�!�o|�ԁe"OX��G�.w���W��%v�,�"Oda���QrH9�7W.aj�R�"O��c B�f6a����L[R��&"O�5�� Z7ky�-�QeČw�:�@�"O�\#�#�s}j��&~v�e�G"O刓n̪f)���"h>��F"Oȉа��t8�3�Le꘥�7"O|I��J�� 	"�ҵc�"Olc���?flm腎M���]��"O��3wfEF�D���
LRdP�0"O8�r�J��5p�(S���߂T��"O$1�ۤ!��u�'�ϊ`И��"OhM�"KQ�Dq��ܠ ��"OJq�RA��|��1ڮ~�HzW"Ore����+�Đ�b�|lP"O�L�@+�g�z=��W�fEZ7�1D��`��)x�D̙���fhq�r�0D�"�#
�`8�P����K.D����"W@P�p���4)���6�+D�DX�c��<PD�.Y�j�P̹��.D����Ǚ& m��QPeC�1���+:D��)p,�(�"����[�wF�:�-7D�����0R}�}�-�c]0$r��3D�XH��ݔ@/D-�c�"��=�e0D��{���9�`�'�?V��i�T�/D��1g� t�D%K3-X!u,ƥ�/D�|y��-.x����"y��[M"D���琎	�����yj���>D����ϝ�+~��jE�ɫ!�P��a	;D����);v܀��F�{��x
��=D��פԪ@����F36��[W�:D������
��\��H['d�u�-D��bSOZ��X��F�w�P�w�'D�lq�$T�:��ZB�¡?!�LpQ�0D����*�&� �m�4y�=GH+D�����͙L�H�9� Uo���zqO;D���t��33�d�+Q%��b+9D�T1�!D�[���v-]P���4*2D�۠�#tV���E߳
p����#D��tȓ�KJ���sMZ�	�$$D�����.��đ�C�ZIP�I-D�h��Ŕ�S.]i�)M,Tɳ֨*D�@�)fVB���j -�<��+(D�� ��uW
��H)��H�!D�tSɏ�$�T�aҲR�����
+D�`�' ��	ؘ�$b�@�H�U�#D�H+@�ՙQ)l��7a�#��}�c' D��)��R� �eE!`9�i��<D�� ��sU#U�7e��v�� S>��3"O�12Ģ |S<�[�c�J���d"O,%���M"�t�"���KN*��"O0D�eIɊPR�0J���\�>��V"O�A��ـO��x���%SzHuBw"O6c$�@�U��U�d�N�u:n��b"O�耶��oF�)f��_3j��R"ONtk�$�r+�� �ʘ +��E"O�c@�S4#w���"��@�A"OޑQd'�� ��E��#�<D���"Op�G��;&�tw��fX��&"O���bJݺR�4��W�J����"O�UѲ(��7��֎� ���IB"O��q7f_.� �$n�1��� "OZ���ͯ5�!ٷ�=8�~<�T"OjH1"�	� �)5���&��y�"O� �"��%S�A�H�)'҈�a"O`9g����%�֬&%����"O�pBQ"G9D*�9���P;�m�A"Ox�'�$# �8ċ��.���"O\�8D��U~6U��(=o��p&"Oh� ,�6�
$�PLl�ct"O*x۳�E�A�v�#$1MHe#`"Ov�Z$�
�e
5m��43�C�"O|5R6cs�T�@��Ηe���B"O
	qb��9�4���W���	�'򚸒�_,f)�4�1� O��p	�'�@��7s�  pGO�N�,� 	�'��Q�r�\�������v�콛�'�� ���!l��EHd���{
>�A�'��8�f�`+:Irf�JN��'1*5#���$]��t��h�X�
��'AD���Ʈ7>� S�1<���'?,�$&�꜂�G
@_V�#�'7P�0��{d�5I��4���'0�)1IPk�e�F$Z�`r�'�0$�M#_� E���&���0�'��}�r/K�$dn!Q��P���9�'>=wО)��Y�`c8}� ��'#*��Ũ	�Č�U!F(r�`�J�'����
�re�ċϭ;��x��'U��f,Ҝ~FH�K��F�/��Q�'�@�Q�M�`?@����&�L��')��y�F�s
&i�0������'��\��`�U%v@`���l�- �'9� ��f�&M���������
�'�`js���cd��q&�%��=��'�t�%���[N�11L��:�`�'���k��j�.H��!ކ*��I�'���A�̩nc���/Z1"�,[�'ޘ�c���)�bp��K�: ����'���7���$]C��;re�p��'�z(�c���Ќ�p���0��'�0�y����ƥ�k�,�X�j�'V ��c`R+c�4i�F'�>q����'fd�b+I��sF�Ҧ>�8���'w�t��f�Qu�����.t�|X�'WЩr�kV�I����֠Z'���	�'�,��*�Um���$T���b	�'c 5�l���=X�-�
\�H��	�'�"�
�������c�Ҝc�8C�'zB���,M��5�r_%NpM`�'�re��!F�.�R�ۡ�gV����'`����A�bVpɖ�Rn�Q��� �0�2���d�F-U����"OJ����4v�j8�4mO:1׮%��"ONq*��5����푂OӞ�Z"O������?v�ty򡦑�(�^�8!"O<-�$��Z V��G�W����4"O�<�aC��O3��HGaO���R�"O6X3�T��vjȺWT���1Cɥ�y��]�tc���o�"u������y2��<gU��`�
	4��IC��2�yb�rtV�S���j�԰�C��y�`����0�+[�ZM���I��yB!�3�(a+�DֺfuB��C�y"/A=d���a ��t���Ae�)�y⎈<s������ep,Q�NR��yHל!�Ƹp��ߌe�hp�-�+�yBȂ_�@��	��]0�͚�dO�yBĀsV�[��0���
�t�!�D	�jV��s׃H��.\y�F)#�!�D��#�p�k����$�@KԒM!�č�d�x܃r��"pi� @��ԟ,.!�$�75h��*S�o}����I�!򤕬S��9�7�FcuH$3��!�d-D���r0�Z�d\��;�	� �!�d�-f�$b�Q*R\|���g!���.F� ���A�I���0�"�!�d�!z���[D�H]����t�Fx�!�dÐ0�l�t$C�8xм�Ԫl�!�ǎbj��K�!ɤuT�!q��k!�DP*
ʄ�22mܙWL�书�9!���kU+��#��2+ʵ�!�Ė,:���A��jb�Pc&�	%�!��_�Ga6�#C�xU���3�&/<!�$�6��3!M�6P��$X=�!��O�
�|�uiK�2�h�B��0[�!�d�>�zIQ�fQ<aT=!4+��M!�d3l����(	�%"�!�P�X�b�!��#s������j�,j4��N^!��2~j�k�,��Q1�]I��(I!�ĝ7�Xm�Ëњ�a����!�䖕<�<9�?T��|IU��72�!�Ď
[;�e��ѳF�By�4�I�5�!�Ď�1�u ��>� �Is䓫Q�!��Ƅ1�c��U�h/ Q��lU:\�!�$ܼ91v��#�h��웰%��*�!�ތl}$\XGe�	q�|����!�dY
4� )���ψ"w"�s�D�Q�!��DӓDZ�;}ޭ��h�)u!� �D��%f��;�ș�]�!�� �{���x��be���F�Q!��z�x�hen4pcjE���]�::!�D�?"��:o�k����T!D !�d�=[{H���lB�4���ʷa��!�O�I����
� ��� �I4!��LP���)J6��� OOD1!�ݙ8j&<��E(���.M2"!�D��d��kC  �Y�t=H���!�T����S�DlښR�bQ�!�$6R?2���G�5� ���(Lf�!�d���<!;���'����P%?�!�#w 	��M��^��]��ͰR�!�dT�a�<j��M=t
��Bg�8L�!�$\�yK���fQG�$�8���&f�!��Ζ��@	���Hjw�P�!��*�ځ�E�M%"p����C�%�!�� }�wNL?L}p'��o8PՃ�"OF"�bQ6$B���CY&J3�@�V"OZ�hG 4J��t`'(H'dfl`!"OLx�@���P$�"���#ꜱ3q"O�AAt�@�I&��B��ρe��A�R"Ozy�R�}��AQ���ʲ��	v�<�S� %g
�=�7HS�`m��[��LV�<�5˔�O>�KN�����O�<�uiU�Dp���/��1��fA�<15+�u���K���Ar��`D. H�<�sc�C�<a�tB�;����B�<	�G�r�*�pf�D�I}j����@�<�2��4TP��G'L�x���;6��`�<���I�4ʸ��5,՘.�|�IH`�<yQ%E0AcL͉�	`�u#�q�<a�
*t���q5JϗY��<C&c[t�<	��O�y������;����Kq�<)������h.�T��I\C�<)��G�*Bhj��7|{��� �@�<��#YL��K�
G��Nx�B�[v�<I���nT��Q��F)o��;� �u�<� ��%jt��H�J�zLY��H�<� �
@���.
%IQ�y��lF�<	s�՛,nc��$:�X��f�w�<�U�h�JTI�U&�$@��jZ�<I���54LC��v֌=��MT�<A1E@�Mf P���N��0*rg S�<i08K��R+^�[mXY�����{�8	R�*/p=��H�>Y��ȓp��Pc����
TI�>Qm�\��f��C�Ý>V�,�(�dF�sZR�ȓa�������uG~<� (|2����Z�9�3YjHĸb%�$��Ѕ�p��)���x�&����ȓrv�2�CP��:���}�q�ȓ-�� ; �9)9Q�8e&�T�ȓ{}܌�&UM�F���:\�ȓo�<�"`N�RL�$A���T���Ki��c �	IZl�07
�)) -��v0 ���x�ܤX�d�$k%܇�E�ɚv�DV�A���-v(-�ȓ<�Ơ�!��		�Lx� V�FA@9�ȓ_|������7T�h��NT�n�橇�%|�;E+ǀq���S����k�J���i&�h�R�W�l� �[Ǩ�6~��م�_gx���h��((r��ͅ�gn�)���ߟ���`Ė+YU� ��3�2U)P�άv�����ʰ*L��#n\ k�X$��{��ȓp1Ԝ�c� �2�Q M�>�P�ȓC�8�2�[���I��=�f��ȓa.ļ�A��X]����Ϟ�z"�ȓ�:�k���BL���c�&Jq�ȓ{���c�'��\0����Ϡu/6B剶If���!�� Ɉ�Q�Y�+��C�	cu��IP럏l�с�nX�B�0D�s��2n�К0 Q�	k.7�PZ�<q��F���ݙ"� &����W�<����>�LL�3�P1��V�<!���K���Ye
֑$�)⤋�K�<���N'��
�kL.a�R$�E�<��cL�u����!G(U���Q�<�cN�	�h-�0d	mx�7d�o�<a�NU R)��: ���2 �Sa�<� <!eG۔m�����j�G��u�"Ox�I�E10~�ij�+�38Ĩ��"O"���-WS�`��F��l#`�
D"O�KDg��=� �Y�]�a�7"O�}h���Zְ�L-0�B�R4�yr�Z,�0H�a�˅o�J����y2��Z�D��d b�����Z%�y�HITH�Ȁi�p+�+˃�y�J��oN�b#�U�K:61�v�+�yr�܎B9���'AȜ[6@j�D �yr�8v°�F�%[F�P��"�y*�ru�U���Wv��R����y"�RL��8c�W9���Q]$�y!�M�x�6m^P0�n
��y2 
?IӤ# �ߚ9
�� V�M5�y�]�!kf��<5�N�a�*��y���z2ሓk�.�,�d���yrc�$_�&0��EʏԜQ����y"D�+�T`�ę�ed옡f	��yRe9�1Sԉ�+}z�ñ�H.�y+/��|p#�0p5�T���ލ�y�'xll
%f�S#���^6�yb�,:?&�!§�c��Q���)�y���V�Us
֙Y44tc�A���y2j�<��1�a��zA��r�o
��y�GU!芀�����w��\7�Z6�y�(��eQ$�)}�*d��@��yR�	"��53S喻*�ʐ���I�y�j
,R��¢�t>�y��,���yBL��E!TN�(���r����y"�
[ܮ\� ��&EbL�#gۻ�yB��Mmy*��l4d`:ăE��y��ϭ4���'�B�;�����y"��(��8� �S; �z\z�͖�y��&b:���^t�C��^��yҢ��j���|�а�D��yB��d��l��(C�IR m�s�æ�y���+�|y��=<�ޑ��E4�yb&L�1#f�q!�8n����Ԃ�yri�6@̺�
Ο7�Ҭ��G��yk�]���i7&D7{|3����ybH�w���V�Z�;!��t���y҇;�IH�]*�:�����yrN�r�0K+y��|Y@�:�y�l	�9��]8�i��<�(�*�yL��l�V=��/	m�lҷ)Ȗ�y2�C�` ��c��6�:`���5�y��ul05!ֹ&bJ��ς�yb�"�0�b�"S�P��Ty4���y�F[�q���+���H�����;�y�t�ĉ�e��;c~�зm���yꊷ'f�����և:Q>�Z���y��/@N���=9��t3Bo��yr
�9>��<aF*��0@�zQ�H�y�jF/;:�{G�G�Zh�x��yR�" ���FU�K�`�c�^�[�@B��!u�J壢�Ixj����2�B�	��&��F�~�촂��\�C�	�8A)�#���xA��M�ou�C�ɕڶA��(hG�!�˻;��C�ɓx:�A�D/6ut�갃� !�@B�
�t�:%i֟�RA0�B�!��C䉞R :Đ'D��Hy@1&Uf;�C�	+s2j<6��"�<�X�i�0W�nC�)� ؠ�����V��	��1j�
D�"O��AFI�$�Aף�1�l�hp"OP��$.������"O^�(��E-~�x�t��R�����"O���RiX��	2%*L$^x�\�a"O�1'���6IP� ��L8��"O�P�7�Y�� 8æ��uX�"O��`��[�G�(,g��$ 8IkW"O��K ��7��uA���Qp���"O.�9��,0�����kVl�B�"On��$A�/'Z�5j�̂�,^0��"O�i�#�H(��{�j֐9Vx���"O~l�ѩ�0������Ƅ=P}��"O,2���� ���N�U�<� "OM2%�\�8�����%7&\!�'�41�'M�+Bp��=�ʤ��'����C%N�cSr4����:Ťu	�'�D����_��vI��N 7m��Q	�'���"�ؾq�}���$B����'�Y��*ś,fB9趋�c�Z��'�P *�NQ��Es�֍X�����'�+!M�Z\<�2���NČ� �'�ؙZ!.ݻ����̙0P?�,��'�ri�@�<[�x��c�,B��|�yr�'��e�党rX���E�8�,#
�'�:���h�u����J�+���
�'*��TO� ˬ�*� �r>�`�	�'Ep�s��0:�D��h�J��i	�'
���
�!a�����ԉux�9�'̖�8u�8�cDL�{�5��'���VkQ��i�e#n��%c�l���'�Q���'�hy(t�D;Z^��"\���	�'H�4�k�7���f�K[�`��	�'3]:�kâY)JD�U��~�ֈp����?�u!ˀ=t޽3�NB(b3�s�k�d�'�ay��N�f.$���n�;B��X�f���yb+(SX耠B<#f�+E����>)�O഻d(ƅ3'�ᨔ�X����Y�"O�T`ذ+<<��W�Qc*�3"O�6LڡL�}�4�� ���2�"O�р����֬���N��A���IF����A�Z%������q얡�d�G�]�!��W�@@U�܊]�6`g���!�� �W�&T�
΋"�a�gm	J�"Q!�"O��:r�0#��x&.��"���q��I�<��)^4}�DE�$DU//��芳虌5�a{2��C3e��Q����~�{S��b���hO��lJv��Tu��R�� $@���!�S�n��)(�oB�i�v	����"�����	[����O�rB)��n\�����&p�u&��Aj��G�'�PJ� $>�@�6��yV���	ߓ٘'��Z�ǁ=A��q6�T�xh��!�i7Bb���S�O��Y*�m�b*9Ye![�rrbı	�'ΌaIg$@-"G�% u䜷~���	�'�:!2F_���(*#A�9���'��O��b�G�s����F�7�*h��"O,�JV��>�θ���ƨn{N�b"O4����D/s�h��W.4\��9&O�����	��$`�,[c��吓�X"	��xǖl�'�:�@�L7����`D+`6D�
�'���lS�
�:�Y�R �XM>���iA)d��-��=eB���(G*��IW�'�?!�f�1o�XH�$�JP!"��*�<�O�����E�6������r�Q9E�=U�!�� ���c�]+V��� �F16��"f"Oh��"m��1ᤚ�3��� 0On��dJ!/���3^%�v����ZF�!��T�-h<�� mZ��1�a���Q��F{*��Ԁ�T6�`�kW��8J&*p
�"O���陣B*��-�7���3O�=E�DM-z΄X�J��d�\�:��/�yI�#ژJFd\�\
���j��yBaݑ4\����K
��H��I�0>�O>�7"�2��4x�$G�J4�4�G~�<As'W"B�Ĉ7���r���a�r�<����L�,���c�
�*��Kn�<I���1��؂������BԂt��eE��j�ß� �z؂��>b�<��ȓL��ܘ��̙N2�J�F9=bʕ�Ɠ5���mn6JM�1���j�$�+Ot�䘧(��8:&�,R�Q������ "Ox]��ƾ�6%�֌��:�܈��"O�=(c��ȤC�k˷~D �z�"�Z����r �~Z����o������ڧ�y��^����wFP�i�>(�/Q"�y"�:=�Uೇ��KPt��� 	"�!�(D	@�k�˚������w�ɠ>
�me��-��r�%^�eM(B��$,+���KAf���RB�I�"��lr�];4�d��*Β)�B䉋�|�W�"K�J�r���E�B�	
:�����.m�P�`�kdB�ɟ$E$*sd0U^��4fE.�<B�	�(Flycw �'w-Ҭ�Í��`
0��Ɠcf��!���U62H����.����38�x��->�.X��.�"|���A��@�aΘ-?�.MRǋH�Ҹ�ȓv- ]�a+W�e�@�v唜d.����O�8E��	,�B\:!���OqD{��T"De���'��=��¢R�yr��0a� A�'D��WR���o����D.�O�5��c�t�V6.A�0V�8���:ړ�0|�t���р�ᆌO ��`��K]�<y���$z��[s��s��H�2��A�<��]��i�%fF<V XEM@�<A�h�F�lؓ��3@�J)C�[}�<�%��<���gA�S�2�
&��v�<Y����0L8ȳ�U�iji��q�<ٗ@��/�p�J ��9���� i�<��ȗ�9�fl��� =��;��a�<��B	 w��Jfc�>SR�s��hH<9 `_V����G�jP���'�� �!�dؠ)ܦAk�56��9ku�B�b��'�a|«K�D�R#M��1��5���y2j��JP��I�->a&Y����y��\�� %�ĩ�~���(PCO$�yr��~�(��qh*r�U�W�C��yR�d�X���+Y�.p3����?�f�h���G$��'�?��H���ũ�D(Yu�I��I?D�h:�#�wv��G�S�d]x��ǭ>�d'���~R�j��U	�
L���Px""2��ٱ"O�-eR%�@��(fv\�ӓ�'�ܢ<ikZGsHBb5:ЪX�t'�\�'3ў�0jj��@͎N\���앪l�pA+�'�&a��	osp ���Zx�n0��'l�x07튘St%��C[�oh�	��'_�Ɂ!�����2�N��}�x�K<я��)P P#�Сc��Ex�!����*I!�� ���2ڀ7��������*�JE�)�S�S+8�\s��� 3�&���ډP�B䉪lk(�+��U�*���e�>5ʮB�*$	�t�*�1"���A���B�	,G@l�w%ڪbǒ��d�)h~hB�	�Z�ĈUa(>�>,'W��,B䉐qB ��I��q�� A#��,�B�	$[L��A��
��pp��&XT�C�I�����a+�=�Đ�ɒ�e��C�ək4�H��G��Y�K��Rϒ#=y�$q��j�ς�7/&	�Woߣ/�u�ȓq����k�NB.p�3h���E��/�]$�>�H
r"ӛL	��i0.ec���벰)��[�HK�ć��K���D��)Dsv4�R�E7zxC�	*Fh
A+�S�xyZl)�HE1C�� q9�(T&יL@�
aꝌe�:B�I*V� ���'G�P�QҎW�7�C䉎H��� @O�hc�˓�f󂼅ƓD�A��6��@@�n�V�t��	I�p��Y�r
ݮ|������ $�͇�l!��aW���=P�#�d�Ň�R��̰�F�~�YÅ�J�9K����&``��_�1(8`c�?�8�ȓ5�����Y1xl
t
�d�ȓ/�,{�h^~�H�z�*T�I�`5�ȓq�N��'Ό%���Z0L]9%���Qj�K�
1������	�Z���DZ�[6犹E������ap6���=*l�:�LF��mX�H\�z�*��ȓ#!�LI�ǻEZ���ԏ�@��ȓ|��z��9T<�� ���9�~)�ȓI>i
1�[�2�X �Շ��g/\!�ȓ$xAa�ύ9��Y���Xޕ�ȓh�|ǆ�J��hqt��_�ІȓI	��8T���n��f�))����f>�h��GP�p0�ߧ��k�'� �J�r5^�@����B�xi�':�	ɲ��S��$�G價d���
�'�,���A+6����,.D�-�
�'�Ȕ⤧GA��������'�H��fʘ#G���S@K>~�0C�'�|��K�*|4�+�͏z<uB�'<�����ۻq�8��D��q�|��'�1�!BoT��D�Q�oVR��'�ވ3�Ѱ"&���f�(X�����'��X�- !Q�i�Ư�IҘ�'���!�vkbp���DF5j�'���1ä�U���1�9a�D��'����fH�7���� e��	V��
�';���F��;
�����ŗeLЃ
�'#d���
�Y���F�O�v��4��'�6�8�i�>^�*٩V��z0@�'����C �3s���pE�%�1��'"2!�c>^'@iX���
�q��'7~`I'I
w��y��N1~-����'�@Q�Rf^9�V�_:{h��`�'�2L����{��H梁�z&u��'��YXR��`δt�̣rnYx�'�ؼ�cL�� ��ق��(�i#�'�Și��ܹ�T�Q,���|3�'s��aJ�cC8��q-V�H�@�'bB5j'�ތI��#a̎9i�x��'8&�J��K-o��2tG�+i�
�`��� "�s c���  �S��ξ�zv"O�MC��Z�mk~@ ��(�ԙ�T"Oਲ਼�W9\.l���Q~� �2�"O��挄�H���!ড়n� d�F"Oh�Y��ބA����B��Rz`��G"O�L���G�u�z�xtO��qX�Y��"O�=�Q��xΒ<+��ْ<kl%��"O�̝����!^��@"O��gdУqD8���
7R�,��"O~}a`̑���x�gO�4@Ѐ�a"O��c�%v�U�VF�%?��IB"O���>?"ޡ� �U|�V"O�P�A��XD�a���U��r�"Op��p�=9x4!�+�6:�J)�"O@�å�'U������K���"O�-y��( �1hg�Rʦ�U�<	 f�bMJ����&Y.�a���M�<�-�y��˓%�,j
QA�˄]�<хf�$��h;נީ[Sh��D�WX�<��ǅ#5�9B�3x1�q1V 
O�<	wmK����g�. ��YRD�<��S&~zȲ�O�0H�m�T'��<Qp�2U�j��%�,q2�����v�<A�E2u6����2�4i ���j�<y�cc.a����&b���%�g�<���Z�c�1x�~5��R��c�<������$��M\02�p
�Y�<A�j� h0<�qG#�
z_ptCLOT�<�&�^O�i�֧�������T~<���M�p��V�
��~Ř���<[�(��[�N�SCG
C9�� ��)M��YG~b�S??�n80Ą΅2FԸ��T�F��C�g}�]��*fe���$A�,B䉎�И+�m�8,$�	{�iΈq3�C�'X_��ж�EOL�U�Ek��,50C�IR#�m�B�q����!� �C��/�\r௚��X�q�B�ɳbd �n��{���*�4\"�C䉼F]�]S3�I3<�8��'��96�C�	I���h��h���Y�R�DC�ɷ,B���e�
�P�ؼ�u��B�	Md�QC���5��\�R���C�	R3�m�$
$<���2�"5m�6C�	�R���Z�'߶H̞�01oQh� C��,o�� �(O��h�8F
�P�B䉑e����~׆ K���>>�TC䉳Q�ihP��5J�p��	��qv�B�	{�ܵZuk0�R<�%l^�<�B�*]2 Ar/."���QCQv{�B�!�<(I4�h��ag�PQ�'D��B��Œ+������ͮ��q3c#D��(pM���(��p��A�e� D�`(�z��ԋ��I6Sf��u�%D�P3o�<|���n�4eF���'D���4�&U���G�_AB�!�'c7D���b�νd�pᣠ]b1`��qm5D�(�c*k ���tO�X\H��5D�x�'�In��R�ͬ&(�0!a�g�<1#�	�q���cq�֫x��c��y�<�ɕ�"\����äl0���c�z�<a�`N/-�X�ؕ�A8@�������r�<��AF���q4.^7;g�t�cu�<a�����l�ʓ�ۻ^q�ł���d�<17�׹8BI��G�� f� A��Yi�<� ��t�]�M�b�@C��5l����"OTY��O���]<Poޘؗ"O�A��gL'���	ϦX����w"O����A	
B��P��h٭o��xh "O�L��#iRX��@S���1c"Ob h���h����-���Q"O���l�)��b-�C��U9w"OL}˴��fp�-E&��a�"O�TB�C;[0ƩY6k�'3s.��7�	�KʖmH��	^M!�0�A�T���W�A�*�!�Ą�]\Pi�GK���%���D*q��ʻ?X$⟢}��^]rj�F�33�@���"�`�<a�LW7�&����[�F�@�c#�X��7.������0Z�&!JR
�)v4NtkWŀwd!𤙰Z�Z<``�e�����@��#y�q��E�R�Rfk)�O�1�T
(<� �bD��VS�{�"O���R(E�%"��9LtZ�"O�1�Ń�%�\���>�� �"O&���CD!j�U[��?D��"O�Z�[$3p�2�l͏#hi�"O���@��':
t���;*`��"O>�3�OQ(r^��`��$b���"OFh�wCJ�(��[��Ĺ;P!"O�$(!�!�*��k�T�8;�"O�T�ש�U�Œ�H�POb\�B"Ofi:CE�BVt��*�!P��)�"O���"�(_H���[�i�SK��`&!��W9L2	�&K-<=hz��$�!��N/{�"e�5/	�z?��� I�\!��Y�7-�)����@����$�Y�.R!��̈N��[&%ˢ�L�R��&�!���]E�hJ0�� &�d�1�
�`�!���w�b`c�.�;g�]�d�!��C!�҄��6^V�"1h׌E�!�D^�b�Fq+E!�l!A��
!�D��"q�����a��(���!�D������X��&�@v晇h�!��׿y��@�ݼO��=�p�Yr�!�DK:]�&�q�)t/�D�d/D��!�0���a��[,t�*x�C���F�!��7���c6,�}�n�q�M�.t!�D͠x�^D�rJ�Vu���+R���'K��˅XVF	0���UL"��'��Qb �{\j0���R�%z����'�����Z�(�8�1��� 2ڡ)�'���k�J(~};���_G/�9V�➄G��'Sʜ�1ȑ���hQ��b��E��'�&x�4B�/sv�q!�'_#jD$O�N ��*�!W��0>�(T�%g��` �R�^��D���ux��h 撀\��T���x���A #^a����U���HpD���y��:Q7b:���r�|�X�(N��ēQ�P���$�Z�q���(�4�AA���%�R)`4"ܕt��\Cu"O����-?~���*s>=�xb�9,޾��G�.�?�s
ǡF���'��k H�@Y~��fy�VI�'��9B�̤E� 	ɱNJ�MT��6��#��P����p�����6�E�Hq�M���˿F��m��e*O&�yg���+��'��*s��i���u��ʕ�����hʬ�y�dL�"����$�$������V����ɤ	LjUa���/3���i!Dߒ U��?Ѩ �R�e%=,�� ��dN:D�0��f��I�����&T�8�e�a�ّc��Ȅ(Y�kDU���ߗ�c>Q$�в��T:Xk�ARĥ��!e�5��*�Ԫ�A705V���Bϫs�&�+b패R�lC��+\&�b7j�; �Ȍ�OH�9�.4�IQ�ec3%X��R��A#V�8��ۛ+��d�'��m� �ZDA�)�ʸRT���y��p� �@�N��8�0�,?�$� s�.��?� @u{7�U4XQ+1�7K=��KR�����<k�lLYw+k�����Fk��p�����Z}IB��`� ��u�=) F��@Ӽ��O�D`n� bM*Z;,-���9F��4+ĆW�$�������	�+��t��s�&��
6�`w�?vjM"�`�F���� �'WNE���]�Y1�`x�aO=5p#@KC	�uҵC���kc'1��I
.2����d�� �I�M�v ,,�6b��x�F�֡��Z�\�r��-CHF��d�-��S�؁�
h�O�1�'G�����O����ǩN8E��\�v$	0p�Z(J���mc���x�d�9\�0����,r&
�y��yL�h�ƚ��bb���&E�j8��JgN��̸{����l9H�)w!��ZpN�:F���V�Q�xb?OИz��Q��������Pq�O�HY��K�]�D"�'SDSN1�Q!�1$�����픡`x:yY�4\O ��G"���:��
�~����'���"�g��v���,�̦�Y%�B��P���b�>,�Di � 8D�$ڄ��p�h�AV�ԁyM�}�7'ȸ��KQ&_?��[3T�8h(���.a�1Ƨ&D�s��p�脑�if�}H�� 0��T�{��(��F����W���`��5�5D�����=s&u�VEݰ�dIA��2D����-'����]=�%&]��!��[��u�"�D@ؒ�!�>�!��
���E�5ve�� �N��!��M�z�:rI�- ��E,L�{�!�䚳&���K2�8��x��D8!�ٖWdtMs"�ޚEcF��5)B=h$!�$�}��n�GP�\QG�9w!�$�y����g���BÉ�!򄜽~�T Qo��s�D�G��V!�$(`'��r%J�}�>i�猯=�!��œ-vlB��G"0��Dr@F�I�!�䐤7����H5<_Dsu�P�g�!��!z�,̀#�X�|�t���lN�!�J�\&�MX��3zuJq�V����!��[�Ș��Z�Bf����2j�!��
ps0��E�S��sM��B�!���@m"�Ӧ.�$~&�˳Mٴ^!�Ą�Lն|�QJ< ���(��5LF!�����|��.QC���kԻI!���I�������*�6ĩj�}!�$�y��)�q,�.�ֵQ2I!�dM aZE�	Y|^��ʇK�!�dȉ@��,c�,O�R�d�q�)�!u�!� �7
���m�!NL��c��6�!�$�(^��W"Ժx+g��_'!�d�.<�&,Ҁ�ׁ���Y�GU. !�dX�{,��0��
3�X�kw�I�\!�R�^Ԡ)�b��Q�� ���q�!��-&t#%�[2XVԣ0&F�5�!�d��3�j�ѶeC)Y��10�D�!��%L"P�2��&@ y��d�^!�Dٗj*Ȉ���| 1� !��x�����b޵�̆�2�T��?�.���H^�X�)���:����2!�Ց$ǀ�װ+�Z2tVt͇�dh"p �h���Y��D�dPZ���b
5��V&b13h��WrF���O2�$HOϣe�|�ja$��2hR���SC��H!��AP\#�g\20�I�ȓzֲ0(��5���.YmJ���ȓXz>�Aց
8p�^t#0&��%HR5��o�(�7kD1��ZP�@�`vpC�Ʉҕm�P�m�호L���h�'\p�zBǎE�T�Z��D�@e
���'�B|�aO8~
���`��3m楛��� ��x��M�kH�{� �T��H��"OlUr�>�HX 3@�Oy��e"O䍐�G5-�l�`,Cb�ȳ�"O�(�5�;�f\+g�Ӆ$l6�+�"O�q�+�r�3KC�`#���p"O�̉��־T*�H�1�9��"O�!��I(J�p���S{.�C6"O�9���g���W��(���"Od��
�*��� 83��A"O�a�����Hj�Ǚqj@5��"O�q*1e��ƈ]V���W"O�X����N�FD����L���r"O�3��ֲim$��F�U�Q�ș�"O�m	r���`עY��#q��V"OQ���Ś6��Qv�mb����"OP�qAI��6�S���3xBX1i�"O��c@���-��Ż%�):ʠi�"O�]b��P��R��E�i;�h�g"Oᘇˎ�D��Q��� '$P�"O�e���P�v@a�㍬2X��#"OVt�!!��,h+/����M#"O�h�r�B*^'����OE,wV�z&"O��R�N�]b���I����c"O ��ìH� 7�ih�G��~vP0k�"O�͸2a�����S$�G�wO2�p�"O�|��JWWj�l�#,�5998�"Oʀ[oK
 �N�Z�N�/%Z@ZC"O��ۆK��a鈐J[�Hv��j�"O@�äVfƒA�≞�]�@s"O�dy���\3��֧h��mzc"Oٲ�lS�	uj�ٲeM�i�q�"O����#����ń��y�A"O6��o:H�~��B��F��Y("O$H����%� 8�T�U�%���P�"O���ᒍi`�1 �X�Z��i��"O�8��$�9X˶�0���#Q�N`C�"O�c�N���C��"\�P��p"OL�P��?'����@��h��pp"O����a �lPE�:r:Hk�"O�x��՘D�T@-чqƘ�9�"O��"`KB�D���3i̙+�R-��"Od1��dA5�𝩷.������"O
���K�T��9��BF}3�"O�)����L� 2,۳c��MkR"O4|�beӐ0FDM`ҬJ�D�f���"O�@��K[tX]���G0=tΥX�"ODـ6��
:8�/qݦ���Β�ybMO�y�&��-ߔ]�~s�,�y2���I]|�k�i�,x'DDڲ���y�gنdJ��؅��s���3.��y�˄� ���mߗn д4=�yB�	/s���$nE�bt�x[sDO��y2���p9B2M�K�(��Gė��y �����)6}��ڧ��:#t��'c��DǛ�y0��BPa�8)y|�'�x���
� ܚDa�\�az�'�x�*��#�2L��nZR�z���'�>U�� ��uify�c��6U%� [�'�ڄ�H3s�����G3�	A�'��q12n�8�-0p3��3I�
�''�Tj&��@#R�*��J �ū�'�&\q���58Kr�W"a�^�	�'�T��C��%���?[y�i��'��(���#إ�ԧQǞ�
��� ��5�֥B�t��"/�2>���"OR��1fO�4�|e�l�ˢ�)a"O�!(%��j� �Kc�'|��mX�"O���&C��x��ƢH�9��(P"O±�����B z���&8�J|h"O" i��z��B� S�:��ESP"O�u	�(͞{)�,;���w(���"O S�K��T�Aa�	�7X�e"O��4G~� ���ޫr�p�@"O�dBcXN@AI^��p��"O��xe�g���0�P4����s"O0Ls������`�P<;��Z�"O��Ssl��zX��?Ez��a"Oe��	�Y6|�z�XBC�!�%"O0|�ԍ���hUI�	k��/�y�j�,jd�(D�j��.@%�y�␋D��sF1ad�Y3	ַ�y���*�(
�m��`SƝ��y�-6g:��� $s
[��M��y��$ΜAK'��`��Ĩg*��yr�V�o�����#i6X`w��y��8y�t�
��Ȏnۈa��_4�y� J% z I�c�΀S!��UkJ��yA�s`-j���22A�d�K��y���1b�����3�\8A�[��ym�|��u�И"�i���yR���"�\�g�J3#h.��Ү���y��1A �ВE5 �pظ���y�����R�ot}��@��yb��81�̕%k
�{L��g!�y�,�/0�$Q�����T*E(�y�!�\\��(ڔ��EF��y���-*��c�j$�L���k@��yRc�h�p�n��-���`�aB��y��@-J�ҩ{�H��@���3�K1�y���#���m+N.FX��0w��;�y�bH�B��6E�8!��:7A�y"��2�����"FqK&��\��y2��2��Eg\6v <�E.L��yr������dP_���ڒ�˼�y�'��t͒����X�y�A ���y2/�(fR��.��{#($��]4�yR�	X�B���#{]N��2ň��y�'G*�x�z���w�bĠdd^�y�T8nת�ٰnP�t��9�#V:�y�M�
r�"��o�~��Jޮ�yr-�b�P�
`$�:^�(x�bR�yR�RE(h���C�Phq"n�*�yZ%�h�03Nŉn�<E�;9��C��&�d���Y#�,Yk�D%E�C�'j8���$ׄ��z��$BX@C�.e����Lǻ���#��M\�B䉐3A�0�5��t$>���g�B�I[a�Ճ��U�B��*Q eC�2x�3c�/q��9Ye
�^�XC�ɀM�\Z��3��mpԩD�P
C�	�Wj�ؘ����zt�ÑHy\�B�>^��t�@�\�3��mC� n�B��E�$p����>T��"A�~�xC�I��V� ��
�8��ܽRGC䉊t�jT���2F������\�&�C�fD���2���0Ԉ�c�g�hB�	���d�<X�$`�@mY�I��C�I�L��	#�W&4�Z@��D  Z�NC�)� 2cP͝HV�����F�	�r� �"O��:5
W�#�m�>zs"OV+!�ڲy�pU���S��X�U"O��9$�Ŀ"�2����.b�����"O�8�q�9���X���%��� !"O0-`g! ;<�i$�M��y�"O����n)�(�\1M>l��t"O��8�lʔ8��S׃�+<yx�"O�1x,�r��D��I��c>�x`"O��"���n������w
z��"O�p���Ӭ�L@ig��	b��"OR��� �8R��M0��X����q"Oެѓ�M��9�EJ�qվ�#�"O6 RC��{����eܐZ�N�q"O��A 	V�H��#FBU:2�l��"O�i���U&b�N4S�!�i��5s�"OиIg�D�mf���d�&6�e#"O�8�d�%~`�kO� U�t"OT�˒� NH\a0eo�>^Ұ<a"O�ԣ偈�-�,q0�F���"Ox�0��ϑX��䫡�W�p2"O�L�%K՘,� �[VCT�A��A��"O�)� ݾ[��Tڦ)"���"O�� JTv��h��{�l� u"Ora��C"0�$��q&�9!�j�s�"O��hs����q�[lM�U��"OL� �)]fv Cr�V��켚�"O��BJl�hT��DP��Q��"O��j��U�-.�4# �hؔ"O.|���fA��B�MT?}c�ұ"O|d�m�ʜ�#�AOh���s"Op�"�A�'����F@/)��[�"O��PbN]�t ��eX�Ux�(z"OJi�/OG�.A��	P"5d!*V"Ob�+�2#j�� R
�}n6	H�"O8̸��*i۔��h^�dC���"Oj�ɐ�'����Q� "��9�"O��r�";ztXd��!��"O���i�-�Ƅc�O�>Z�x�d"O�ig��yqV,���[. �t���"O��9���,H�k�(X�R�S�"O�T�-B���9s�^#7�����"O�X"����D��6�S��ea�"O��G22~���E@�[/j�X"Or��)���P����9����"O�M)�fͼo:Ա����2�,�y�"Ot��wC��	�� E*C&��e�"O~�pweS]Zh	�/Λ ��p��"OU3��E	���C�Eh���I"O�-	�#ÜjT��N�a1BL��"O~��&I�5@�"<,��"Ox�H5��A�@	!ļY�tH�"O�M��L�5�4@�k�pT�"OHr�G�v��)�A��m����"OF���A��x�t�:� �9M'r�y�"O�ݐ5�H4>d���� J��y�K�U u�ǌĵo�q��]��y"M-,���q��]H��t���y�@ݭ?�0�(�H]Y�"�#�b��y@!?h���	�Y�B��Z��y���_���I`�V, _Ftbb�.�yrjW�3� ]s���wx����O��ybk��e}p)# )3g|���/=�y��-2D�+�mY	7��j����y
� �@�W�B���aD�I�h'"O�� �,Q�$����C�e���b"Oj����Ɏi5F̹��C<�ܕZ"O�%�.�&=�����o��������� l�'�v��}ӑ>�����ܠR��\�rn�)oz��'�0Ŝ.S߉'s���dE�qx� ۉ^�L2�Ƽ �BT��r7U�����<pa�B�Y?W���`e�%���b���<!��U<}��y�P&�"�H�4D[�)㛶O5�S�O�T����"}p0�`XDN��c9��0|� �1"a�0�k]�p���2f�@m���hO�'X�j�����Ga��2G!+X�Z�$��:���I�0�����g{0������E�'�Q>=�������N�f����5�v�4x����/$���8��β.�T@��G�]�@�Fy�	4���]�'M�]��N2�I��6{� ����L�� [�'��i��F���
�(���Ql�*l���m�Y���	b�T���l"��2$'�O�˓�~�'(��$�q�A2iʐ��
��k�.�p�L�>AS��>�p�	��H���(T���q�ٽ���Ni�@7͓��(O�?��beQ�tx��B�\Ĥ���Sk�'�8���/V� �%��
�Z�Ҏ:q��O��GzJ|��L�"I8�I�bQ>Np��{�	~���OY���Y,e*���:à=/O��=E�4�Ӷd�h��l1K:Ț�)��?A����x܌�2L�c|Xt�A��5{B�Dz��|Z��>0�zS�@ެL�F$�$��<	���p}""	e}���(���4(aK:	K +C�I�e���'��	X���[�O��]��!_��y���õea�С�U��X���=�)��srp�����n��r&�����FԼEGJ����ƻ�M뢁��6�|�"�YJ����R,_\����.���y��Ƈ@���!��@�q$*�!�y��&#���#��2y�F|@d�ê�y�Q4p�`j���>#�Djs�^��yҫ�"�uHE	6�Y{Uj���y�% �'L�*�
F�YxT�Ç�y�ˋa��9 $��L�s/���yR�52|1pm
�n�k�����yB�Y23zf�bw�@o62�M��y"$�*	�YY�[�0��Qb���y�E�'QT��b�]�#�tx�!ɚ��y���0�Q
V�ۨN�n9��j��y¨ζ"�m�tJ�/1q�������y��B/!w�B� �90v�y�����y"�W�f9�&K�U3��*��T��yr�	�R⼳,ƩQ�x��� ��y"��`�f����@EX������y���Q�FѠ��)>�l��d�=�y��j���s'��;r���dP�y�(��B�`������4�����y��z�x�b"�ƾ %�!�A\��yB�(IOɹ��;�a���Ѓ�y��ܧoFTQ˗)B��HA�0�yR!P9���B�ԏ{�p� ���yRcT'���bh�x�ؐ�w��y2gŪ?�Xѷ�E�вg$ɢ�yB#�!G�cp�
�"�!kƛ0�y�ޅ�ґG�>S��h ����y"�K�Yd,p��+AJ���q�)�yN�@��%@Z��Ĺ�����yb���T��ʥ]���x���ߗ�y��/a#b`����r����E��y"+,N����!�[�����b�'�ֵ됈P�,�p'h�1j��(�'�  *���a;�Xw!G�Lj�!�'^�t3fK�9~���#8N������� l� �7��� �G�p�ؕ�W"OD`f*@Pa8�A�:6W�H3"O�xӦ�!#����� &}=�5""O*8Po�\J6/�9~�-�w"O�q��zBbT�u�ȝ_��"Oz��uL+j/*l���	v�jp�2"O4=���Y�0���S�P�v�V��P"O�`)c�ֹU�2h��ʍ+�ĤYg"O�H` �Mxp=D��!�����"O� �WC��J5�䰧��><`"O
���şu�}X��7$,�C"O ��rmM�f������BZ��"ONX�$��x�2�Ӯ'��y��"O����O7�	��
�[��9�"O��r�O�%zD�qwig��yQ�"O�{���=�P0hU�O%����"O"��,��55 B�5�a"O �`�*�R�[r�+z���ر"O��qa�?7�r��tK�;Ǟ��"O��'� �P�	���@�:"Ov��ǆ�w���r�N8���"OJ@����m �*q�^xL�{�"O���ƎC	?�xl���\�,YV!!V"O��p��0P�`��h�@(%c�"O��	!I���	s�G�2O�p��*O�]Z'�����f��K�&C�'i>,H�mL(uwX�s&i��J��I	�'�Z���Hdkd5�&+�P�	�'7z�+��0��e1�B+{�ɳ	�'����l�/%f��4"69\8�'~��2�˰%�p��/[��L�'�L1�	q�0 ����bTU��'�h{�"�\�}���".X�S�'���:�`�4;`ab�K��,(� �',h�)��i���O@~�h�'��iȦπnvhb��A�]
H�`�'���0��3�V�ڶ��j�h���'��Xp�����80�K0!�4��'6l�����FH���u�5�h`K�'OH<�H�;�4C���u�R�'��������5���8��A	�'��Ǐ�|��<Q��X�D<��'�d�ӳ�D�w�1b0߶i̙�
�'X0���%y �������'6��ʍ0m ��e%��e`	�'�:̙f�e�0�x�蔥}~<x�'������\4c���?~N�H��'� �:V�?SV)90n�#�� �
�'ߖ��I]�g��� P��.!�"	"
�'��Dҡʕp6��0�2z�ջ�'��0I񣟅ZC��v�&�v��'Q
�6�%4ز�aG��-
HH���'�� ���@�f�#7�[�~3 C�'��D����%h�mɅY ulB�h�'���Ʀ���vA �A-n��#�' .�Iv�	P�0�Ýd���'H� 8Ed��%Q��@&�W[j���'�*�R����9�CG\\���'K4��0I��BO׋��4��y�a̍� pȶU=	`.8�����y����Z�z���N�3rf$P���˶�y���t�~���H��4��+Ņ�y�/ש7�+�A�=w��haS��y��|��[p�
5�����P��y
� Jx�G���l5�CӁ$GrP��"O����ݑ;<� J`��ڌ�aQ"Od��6d'3�����W-e�B�"O�pK1��$A� m��F��O�ȺV"O�`{��VF6��h�dM�JjlP��"OV�����1�����R�g?@db"OJy	���^T�-K�.Q�:,�<p�"O&�a���n�
�kF��:4.���"O$�I��Q�.l3��QT ���R"O0pJ��L�fx 4��8E#�@�e+D�t� �Z-|ۜ����*#���*O��ZE�%D��!I�<M�2���"Oh�KW����$��N�4�8Ԩ�"O��0@&��0�����&�x���"OR��	^�TA����v�p�"O����),��`�0������"O��e@I%06����Q2 "Oh�����MU���%z�,�Z�"O�,��E��(���뇣�4�:#"O�܊eGC���4�s���*#"O.���dة!;bD�!(�\����6"O5g$�^�Rax �_��5��"O`�`GG43��27�X=�V��"O���&L8R#�A*@�t�"��"Oj�X� ̜"T��f�\�dBX��"O�]� �<�x Q�̊8�HjE"O� �֯K!3eF��������|�<馫�b�d��E틢�%��{�C�IgbPOU:� �bB��W�PC�I��2X��+��<��<�E�_�~fB�	47����A1�\ї���dB�	8�QT/� ,".�ȑ'Z�A�C��*hA��A!{�4=S �6CH�B���!��I	��t� $�9t�B�	�Q2��j$I�7�XtJC�H6Z�0C�:Q�j� U�P"	T�ق�X�C�	�36���r��1
6H��I-5~,B�	�[e�@:�Nҋ�Q�s	|�C�ɟ /�ش푯2	܁3g/�7��C��({ǎg�W�����B���B�	&�f��4Aʜk����S�3t^C�Io������	��2�]�d��B�I.,BL�d
�4�ɱm��tB䉨� i!"+�4�
9�si�38�B�I\ڼ��k�3T8��3cǵ0��B�I�Ѵ��1�1�T��L�o�JC�əi��-b��i�ܐ#D���!&C�	�����4���9�I_�DC�	�W���q�N�]F�����z]8C��/p�<yҰ�r�T,8te[�U�C�	������ B�6�+���	��B�ɉ\'b�K����{?D�`�E50B�I��8�ц�1`� )jt
7 ��C�6p�r�'�[52L3e��0<̐C�	�ic�5)��һTs"�@%#�7h�C�/�܌xA�n�� ��& �XB�	>lB�(�U	=ĽqC��*WD4B�I&&���nT�WND��̌iB�I�t�f���E�8b�6HS�1 &�B��',���n��![Z��u�ԇsJB�I3<�����2Zi@�� >EXC�ɘK���[T�(H�ք�0'D���B䉎{�D�3��W�����?J�B�Iy%r� 1�H )ش�p5��B�)� P�{�c�He�<�k�Y`���"O�]�͐!���K�>C���W"O\!�3��&b��2�-��"O��"&#�&��c�/| �� "O��(H�me�$H$�Ȕvo�!�"O��5��?]�乃��+b��y#"O,���۝�t|K¡uH.�J�"O��U��<
ݮ�q�ڰ�(B�<�s+@�K����2��7KX|X��]A�<a0�M��N�Fe�HPW��e�<A�!�]|�8C[�,�pU�Wa�<�W�\:BKŻ�k�D�� ��c�<)E�E4d�����:��A�fI�w�<i�?�(]��-�9j-V)ȁ	�q�<�%O�,t�<�cO�̡dhOj�<�W�Q+M*>4[cJ�#�v�v�A_�<AG\����y1�pb���$X�<�m��AY.��*
}~�� "��k�<��'Ξ+%"YKь�<E�v��s�<1��^�%��^�J�r��1ACl�<�A�� ��Sύ.k�ju��MGi�<� GV�/x0l:��_�?"�X��|�<�D�G%Q�6��#�+|���`��b�<q5��n����3�uRU�L_[�<!���;����E���%H����<AP)ЉM���"��V+^��JPp܇�J����ùA��)�숬X��B�'8�A�¤�U��i1��_H�;�'�6�Q��>>z����vP&U��'Sh�����;H�Ƶ+)_�t��'~�87�u}:����Ӌ �:J
�'��m�1��7Z ��c,݆ ��!��'��  ���   �     �  (   v+  7  rB  tK  ;V  �a  Eh  �n  u  C{  ��  ɇ  �  O�  ��  Ԡ  �  V�  ��  ڹ  �  _�  ��  ��  �  ��  ��  ��  � , �! �( �. 25 �8  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�O&��<i��iW�5��Q�4J���v��5Q�!�Ċ�<�t[�^�B,x����"b,*B�I����`j��BE�y�n�{ː���$��F��}@�"�i�zY!�B�q\C��,o�.y`'f�5� ��M#,��'�?EҶ���k��ͱB�M;"j|���#D�|2�EW�fǺ��p������=�dڀ=�b��>�
s��y�����$1Lq��(D���tB��9P% ����j�eKr�%D��2Ȉ36����' pp��b�&D�� ��aDA��7�ezf'G�&$`��OԢ=E�Ĉ�"qh��4-R*Ɍ̹���5�yB�
�1a���0���
���x�8?b�˓!L�[ۈ4�Ӧ݅0��#?9���l�:(B�EJZ�X1Pg�:��x�鉙_5�{`Ӝ)T�k6K�-��B�I�(�V)[�/2M.r�JU�� D��$%�S�'s��ٱgz[e��HiÃ�[�!�$Ézk�AJQ�З&�b�#l��h	2�͓�اr�y�i|��?x�8Qt��(+n&���m_)���Ix�Ԓ�F�Ud��Q�劁�I@fH�<�'^��m�ᦥ�J~�ϟ�I�� �2Q���#�ƞg�T�0"O.����e�Z��;b��Sd�|�)8|O�5�B �L?��aP�7X ���	��(O擈K�S2�T�q��aDE�%X�"��hO�>1��R�<lR`F-���.c�lSq�>1 �O�t&?�K�r]q���W	�0[F���tm��'�� �ɕ�P�eE_�h�>�Y#W����̺k�O�˓3��\q������"����4��R�'���,�--处����� P|��'-�d �OV!�ۻF�����WS��${'�|��~Z�.b�H��n�����6a�A�:D�{�&
�j��1��(��k+8ꓦȟ4 Xe&P
"��8���R=z*"O��
� F�G�ت$@ڍ���T\��G{��iP:��(�"L�MO��Ht�0�!�d�8dp�y�e]/��c�Bɳ]��L�hh�'=ў�)
$�Q��jsѠ�h�Ĭ/��0O�� d�˚�$�+_���H :O~h���� ts���bP0R�r��F�Ƭ$C�I�XYx-#�D�gj�{�/�
���4P�������͈�B-L�ִ��Oʉ#�!�8$t����5%��:@D��H!�U<P:;e�B�>B����ħ4!�\�9R,�`lӴ`4�X���G�e�!��RX��#u��)���x<!�d�b��|a���7�J��%j^ 银hO���b� �BA��h��>6vt �V����(mZ5BwKG���<C���?��B䉐���ABta��> �`��=D��c'� ��իeU:td؁��mh<Q���)�4\�%��+E9����rX��EyB��8Q�%��?�8���Y��yb��91���4
��:HT������8��d�Oo��j�h�?2�ՉS��(.�L�r�'�d���m��Na#s+(.��-ON�+��D.ʧ07R���֖RH	&��U����ȓE�00`ulS?����I
0 @Z�^����'�qO�T�I˗���O-��A���c�ax����1�y"Q�85�HJS�uo`�&��.��'<�z��T�&�d[w�8��"Ê ��$QI��䧀?q�쐀 ���'dʛGȞ���	V<Pc!��t"d�c�T�D�HA/��w0a{��$[���z�+˒A�N�H��UK!�Dζ^�����H%�+֢�^^�O¢=%>���K�j}������Q1T�+D���W`I�p|[r�_�qx�I�v	(D�@��=.D��4�	A�p=�F+D�<b�f�rR$+�BT+.�j=�c�*D� �U"R�U�X1�3	T0Y8!��.�>����Ss��ʏ��z�D� G��B��ԐT� ��E ���c'y��'/a}"ɋ�%UH�'d
; � ,ð��?9S=O��J�雈%�T '���3E�,R�"O� H�)p��J��Z�揌g8��ɶ"Ov9;�n1{��$��� RE!'"Oh���ʞ7�B -D=H��A�xr�&�O���7	@�&��eҳ����Aq"O����e:� `S>�ցJ`�	Q��򉍀t�t�28I&�l��4t?Q�DG{*��t8f,͜K��|�&^�8<t� d�J��O�}����E�ͪyǎ��N�u���S���g������<]�L��fȎS�8!�& D�'���U؟lR��P�js^��@oY�D6�eAu�z�\��'N2}q�&6U`�	eߐI�n�'X.�(�|�.����G�E"@c�'�4�`��k
Na��N�(G���'��P �U� ��0���Ja����'����I�F&tĺEU�mM�	��������!Y���1���h��}�62��O�6� nX�,��n[�Y���vI)+Cx��.r��E{ʟ��Oc�$To�X�U+�u=L�H�"O�d��g��.$xpéP<"#>� 2"O:%h�iK�,�b�C�gדꅑ�"O�@�j�H}�F�� �f}�C"O��b P
��q�Z����"Oq�F@k��J�ň�&O΅K�"O�@����#0�&I��c�z�у"O�E�"��";<d�7�`���"O ������~C��P�V2q�"O�����FQ?f��g��#o�0]�d"Oj9�We_�d�X�3��
bVڄX!"O.�r�I�8\����.TL�,1
�'�`h"2/�Y����1n8
�'�X �c.Ƽ<� �@�J�v\��	�'��)R�
<�.iE	�5q6� 
�'{2(Oƒ�A�P��-r	�'��`�V�G�/�<�� ��]��d��'�d�c�ɀ"^�!� Gэ]r��'D�⒋�	�r	 ��T]���	�'r�������#&�%�1�G�<��ܞQ����Ŏ�X\�Y���_C�<�a�"d��t�&H�i���� if�<95@ς/�T���&���� �\x�<ّ �#:�pP��D�w�>Q3K�u�<� M�fIⱦJ�
���D�F�<���$Q�>!J�h�1\��`Ҷ	^�<�0�CB`��IT�Z���z���T�<�	?�L䐒D�%;�z��3`�Q�<9F ʻh�x��`�<d�$�Q��O�<IB��� :�a#�*P^B�YGK�H�<��CG�TԉV�$W�� @�C�<AHJ7^k�١�#�n�jp��
I�<a�BV�A�Xe��ꈗt��A&��M�<�&��d�Hx��) $�1S�M�<QV+̤RK��&M�A�(���d�<!�P1خ  qNӘcDI'SI�<ل�Q⢝ziՈ{]��ceDH�<q�'m=X!�X�����B�<��,�=�z��$gS ��ǣ�}�<1�蔽5gP�!e�9�䘅��w�<ѷ+ӄn��$ �ʉ�>� �  oY�<Q�f�eΆ\��璄#���HeL�z�<���K��цA� *08�`K�M�<QamT*W�����G?���ˉq�<�W��;�8��s@C��!ʆ��U�<q�-'i�jp��$O0.PࡑF�[S�<٥��)-鮁 "�t���C�Sg�<� ̅ A�W/!�l�����1#G���&"O�4�F��w�m����vh�`"O �Et\���բH��q*�"O.�W/B� ��T8"�F�0%"Ope(�ӕk����C����l1t�'%��'q��'��'��'���'*ԨR��	3(�U� ��f�jKA�'���'IR�'Or�'52�'���'�|Mk�HM7h�ڑ��A<q�a#�O��d�O �d�Or��O���O����O8�h3"�$�u��i�F9fr�#�O����OZ�D�Or���O��D�O
�D�Oh�C��PCM)C٬2>���*�O<�d�O��d�O���O8���O"���O�;R��l��D0��8$m��7 �O����Ob�d�O��$�O��d�OF���O �+@͏�a�|�%L��B�H�O����Ov���Oz���O��D�O���O��1�oV>\x!cEHz�i���O:�$�ON���Oz���O��$�O"��O9���{H��6�Tr���&��O&���O<���OT���O����O����OQ�!Jd�-h0�4~�ĹI���Ov���O��$�O����O����O����O��am�=�V|0jԜy`��Ѭ�OJ���O����O �D�O��$�O`�D�O�(ԂG5C�$�r�ʈD�Y���Oz�D�Ob�d�O���O���O����O���FC�`[04����%-j�lq��O����O|���O&��OL�D�妥�I՟���W֬�ш�:At$N���d�Or�S�g~��e�H�cf.-рI�3��E�^� ��)d�I��Ms���yB�t���*���n剠H�m�X�E���1���M��-&?1�*�gq6�#�a1����*����Ê09�&��@��Ř'��P�G�t�]3F����`Kܒ,?�=1��)m]�7���1O��?�;���f���l�Zs.�����튴����q���j}��t��$7�]ə'�z���&ثx�*�P��S���'@�=�w�	�4!��i>��	h�h-! `�'�`���+ǃj�(�RyB�|%g��8�$��*lIV��gB�Yv"��d⊗Z���8˩Oցl�4�M#�';�I�:d�����1n���@X'�:�v�R*󌀱x���|�Ṕ�{٣�1���A�,ݢH4�yfi�(�P!+O ��?E��'��Y��/�.RD[�� ���� �yB�{��<�����ݴ�����
I36R-h�M�q��G�]��ybu�:�oٟ�2���$9�'���cE�ևVNИ���E:�����!�8
Τ�IFk�hO�<�H~T��gz�t�NZ G,P��DM~��z�|I���$$��XA:Y�PGB
B��A���mFz���O�Ulگ�M��'ՉOM���'�N���M��kx�p��	�U����۞{��6U�8X�+�L3��yk�� ��ɞp�<P�0�EP`�{�%Ѫ��IEy�^��%�ēٴM+�0�Z���@��d�|��D�	���͓}m���4��^ҦM�ݴ�?F�X�"���%!fH�����M���XU��I�N`� *�..�	h�ݟ2�� ʆY�1=�vy��B��\��D1 o�eϓ�?1(O��S�O*����Ù ��X�n�-�� �y��w�8 k"����4�?�(O�x��K�P��%*PM��yi�Ao��'��6��צ��	,Z.eBT�a�h�b�C/����GPFk��P�͘�% �B��L(u��P���M�IY~�O��	ҟ$�2�J���G��+d���{2�e��%���۴W���<��'�ʷ���t2$�� cA�*�DxC���J~b��>A��i947��\%>5�S4&�����H�U��(�D�W�O�Z�cb*["F��0b��7?A��x�v���б~� ��^�S"��g$ �<�~X��	��iB�P�G�B2gzz�i�m��,���;f%v�T��&���8k��]*��ĩI�L,А ���T|H��� 8HZ<I�͜�P�џ�[�A�@� !QDH�u,\鋂�@7.����f�>r]Y�slڒX�#��w�PC�� 1ӎ]i%�8:���� (^����j׈lf�1 	��k�T�@�/O�C�����_: ��Z��� Κ�Y勜)J�����S�쮼��Cm�I��S���E$)F�bA@���`���Q2n�a�Xt���{�	柴��򟔖'���'�<=s�T b�� KF┤ҔY!fܢn�'>��'C"Z�`����"�M�1L�.X�e�A�N��"B.�-�'b�'�\�<����l�Pǽ~�%"�k��4��aIZລl}b�'=2�'��I�nz��KH|*�!�M4&�S"l,K��Cca����'HrY�����컱�<�S6�M�������WEZ�ZSupٴ�?q���D��vQ%>����?�أR��2R�G1)�Q�5k�#/�F6m�<���?��O�Q�O��ܴ	D�t	�%D�REc��G�?��mZRy�lQ�\6M\���'����%?q��>��"�/(���v-XӦ�����q���uyʟl��x2Jŀ�����,E1Vِ�+���M+���q;���'�2�'i�� '�4�P���._7r�V�Z�ԋ/3.�cs,	����jyb�'H��Ϙ'cҪ['r�$� � �9;��ACpJĞ?9�6M�O���OV�'�X�i>���������<��uiV)c��+�h���d�ON�$�YE1O�$�O��I3�\P���1��Q���&U~7m�OH�XƆ�<����?)�¸'͢8���'>1���2�P�&24��OP5`"@+6z�I؟��	Gy�'z�4BT�c�R�X#B�,b�&��" A=F2��ʟ���؟��?���� p�c1ю7�y�0h��*��'&�i,��'B�'��	ǟtx���} ��!t��8O5��1J����ޟ��S��?Q$��I�=n��Eh�H��#8߀p�IԹI.:듏?)����$�O��ǻ|:�7dR�2�*tD�`/.}�i=B���O���ϯR/�'�:̐S�Q�"-����d�x��ߴ�?�*O���-d�'�?A���!�W.^�^-y3 ȮKY P+�	.бO��d���B�T?�sσ�/�(ٲVB�}O���0k�>����hՃ���?����?Y������	�(��;설�7�C+N�n}�GQ���	7W���,�)��6@�bѪ��M�>I��%���6�C#$#�d�O��d�O��i�<�'�?� �Yr��;"A-f&&dSs����֣٧g��UZ�y����O��J�[�Kx�qaċ*���V�D���I͟d�	J;4ܔ����'ir�O��%GϩM"���Q��.ʒ�2��g�v�Y�2��T�'&�O��aR�D��@��q镵(�D�C�[�l���Jy�'M��':qO����O�X����5��*UfȗU�����F1��?������O�H�S� ))H0��G��#��;��&Q
(ʓ�?1���?!��'Ϣ��7 �u}`�ì��Nu����H�^����O����O�˓�?	R����#��+���j�)C0X�&�b�ܗ�M���?���'����_�ds�4��d�c F.�J����2��'�'��	ޟpQ�I��'{����m��C�(��D��<�05��u�v�D;����9ŋ٢s=O�� "B%��@a'ǲf���aP�iJ�Z�0��	\�ՕO!��'B�D��4b��Lj���.r��q;0b�����~,L�!�F2�~���U�.DP�q@JZ~&�a�@YM}2�'C�T�c�'�r�''��O'�i�uk�7"^������pǖX qΰ>�`��P�A+�v�S�'r�����ぺq��#��T}f�m�~Af@���\��͟P�S@y�O2RO8�m�#��'Qz��4@�!C5�6AM1�����Ɵt��
��К2���'�s3�<m���	�D�Ǭ
|y�O��'���6h����<=h�J5h�$�v��<���̐[8�OT��'���w?�Q���KX�P�C��P���'֌�BpX���������e�&6�%�r���`���:�$x:"�'7��`�+.����O�İ<��o��)�J�c��g㌶SP��u�F!����OD���O�\��"Ep���u�Y?����@/�8hڰ��Ǔ!�f��?�������O�}�$��?)0�镌*�J!��BY��U}�*�$�O|�d?��ϟ�:������7M�%n��pI�i� ��;WDV�S���ɟP��iy��'f��T>����M�E跩ޠ<:<̓����hpE��4�?���'�@��à)��l�B��g��p�� ��mօPZ�oZƟ$�'�r�وH �ܟ����?�(�O�$%r �H�Z~x��f@���'s���!�ni3�y���������t0���R)���q\����#�2e��ܟ��I��(�byZwwP��G�}��yAbD;$�2�O��	��DxJ|"D�Tb�f��Pȏ�)6� �
�æ�������	�@���?������'���ؓȜ4VH�Z���#L�6�yV��>I��]���O{R�\�Q�<`�c�3^����N�"uCF7-�Of�G'���*O��O��D����TB"!�r/�"4�x�����OD&>e�I�(��%���@���e��P�k׫t~uo⟤;cBUyb�'���'EqO�!���Y*o"(��'�
C9LU�e\� ��"@���?�����O����*��9%R9"���8B��d��C����?���?����'�������E$I�SM�	>}h�8�혵r�t�0�O����O(��?ɓ!���D��!K��F��$XRdŊфA��Ms��?�����'��L��|��4[�4,"fÔ"� t%�Y�%�P�'4��'���Ɵ�y��P@��O�yZ�#�Æ�K�	ӀuX��ӵi���d�O��(R�N�3��'�X�D�>>�e��LbΩhڴ�?�-O>� �	U�'�?�������V���3��_J��sbľ)�O��DS.�e" Ř���T??���P$��C\�[�k

,���Ɵ�pS͟�� ��]y��O�i�!�"��*Bx�`�GC�p��Qx;��'C�F\]r���y���(��p�ɂ6����u ҭ�M��$� �?Q���?����)O���O��H&J ��k��'x��Ex�#O�����2�c�"|���Z�h�B�f�a�#7�U�A�i=2�'���m/�i>���ʟ��m�z�H�Erp4��L]�6�(����-}[�4'>U�	ʟ��SJ����s\����K��@\Io�,"e`
uyr�'���'�qOnh�CCݜmNX�QgM�La�U�0a� 3E����?i���?q)O�d�Ee�R���Sa��j���-�-[�!%���	��@'���I���b5�ϊ/���C�dT�Q�
D�Ei��Op�D�O���O���<i��
�R�6�˜SR�P"�ɿ8M��I6$��^6��O����O����O�ʓ�?q����|�"$đ �8Y�c�Z�����.�i��'���P��'`"��~%�^�g՛��'�����z���*����,�����斗� 6��OR��O.��?Y�mD�|�L�� ��K��ǢOE��!΄#���:��iw��'r�'R��Hs�<���O�����d�a&�*P�0t�^0���B�'�ͦ��	my��'I&�O�R_��s�ș�@�گ{>V��� �?;�|�!�ib�'�D��ga�&�$�O���ퟜ�I�O�Q�$#J�>�F�;�C(MQ$H;�#c}"�'�d92�'�']<�z�O�'I<���%�5y��E���7�n�&���޴�?1���?!�'�����?����>�Qu �)3��P��Jګ �d�ķib��t�'2T���Y��:�˂?���a��fdLM�d�ު�M���?1��o���b�i��'���'CZw�<�Q���9��r���/�.���}R�2ݘ'���'����;W25��n�׌U�a� o��7��OJ���E�]��ƟX�	��(�����1O,`	��⛄�L�тNI�N�7mړN~hP�5O��$�O*���O�$�|�
�����J���as�T#5�ĂN�K�i��۴�?��|���ry2�'[RT��`ҧ��%P�L�r@dܛ�L]1��'��'���'��	%N��Hߴ�Py��B@=n&����;̸��i$�'9��'w�]���I�V�v�s�$���ߐP�ܘT�?0��:�\�`����ɟt�I#�p�1�4�?q��jhnɓ��,K��|�Pe�-��}��ib�'RZ�H�	
!�x��韌�w���A�����S�N1֘o���(��`y���x;��4��ំ�7��F�M�1`
�i�v��@�u�ԟ��	���	c�~B�͔�7�8%��'V��T
֭�򦝖'v�e�t�r��(�O"�O*�_��οn��J�F%_$rpo���	?n����	O�)��(9V�)��B��u��պ�-��7��_��l��t��Ɵ��S�ē�?�`�T/8|�
p�H�\��p��
4ӛ�A%z �[����W��[���IܤaZ��A	 s�� 2��M��P��4�?!��?�́��'(2�'<��3��3 �I�6� a[��[7u��&�|rHķ�yʟ����O���L3fs������0�Ӂ�V�ތn���@sE��	�ē�?��������aX�M3pT@r/)2� Qx��b}�	�yRX��	��p�	ayroѓ����mW:Q
-k��� \���!D*�D�Oz�D*�d�Ox��X�m�mM��=pqH�fR�{i�S4O���?a��?�*ON���E�|���(�r$:����1�L58d�Vy}��'b�|��'�dD�v�"�F,t�����}���!D�z't듭?���?1)O��(DO�B�� ���1�����K��}�{�	��q��I�I�t��w&�I_��E�v����,ϼ�@=��C� ��6�'��Q��(��Q��'�?!��~���re���z�xv�_v�l�x��'�Rf��y�|2֟�����}� %���٧�H�#�iy�ɗ/ �*ش.b�S����S���	�!6f=�f�O����H�dT�&�'�b�݉9��O���hzP� R$�h��#ִ���u�i�"�{d�d�*��O@�$�ܑ$���	�2 68�@å,���:e��ٴq x�Ex���O 񙣫��|���&�T��$�Jɦ��Iӟ����
x:�2I<9���?��'s�E��i��@���j�(Rs�jI�ݴ��_������'��'~ ��A�!0=���	Ğ�8&�v�P��w�p�&���	韠&��+|��M�Q�Yy�T���D�aC�Cx������D�O��d�O�ʓl�f���C��T�AiL�)z��@��d��'&B�'��''R�'��<�r�ղ,V���S��tig�34�Q��	ɟ0�IGy"LU,q���ӂ!�0�"%�1�M2�T|��O`�D4�d�Ob�d�%/�����/�|@�v�	��N���@#k~| �'x��'�S���A,ڳ��'�E0���,̡ؒn��]��q3f�i�ў��q�&�����'Y�:�Sv�޻LX��6�V/8p�l���IKyY�Mu��j����kl^Y�΄�O�%0ltD!+E7H�O�����I����O�b?u3�lȈM���cV�"��ֹi���'��XY@�'�"�'���O��i��:Ph�6�(��w� DD���$u����O���`WA�1O��d���#���I�Ń;H8��0U�i�:L�Q+u�V�D�OX������I�O"���O|����FdH�r��D#RB�,/�Ĝ;4�O�i&���O��Y) �
���	��=qR�ݦ��	��x��!����ȟ�O�R�Od����O��6��s�I�5��L���g̓
p)�u����'!��'yx��,�`�6Q6�̶X/�hfuӒ�<h�"���Oؠ�Oy�|�,_4��%���R%@��t9�D��n=N�Z�Z��M>!���?���?���?ԘZ$�)"@8�ueI=\!�ݓ �_��?)���?����?QL>���?�'D��
��J��N�	���A�S��'���'���'���.����Z5.�H��ͅ��EK2G�\7-�O��D�OƒO��d�O(� �e�NJ����
�(��jO�6����կ�����O����OR˓w�x�	�V?����
��E�a�Ѽ���a�=T���"ߴ�?�����'yzuz�}�m�xg�)��fA�%J�0�M{��?����?�v	 	���O��d����KE�>V�ܵ��N��k�f1C�n�j���������!�B�)L1O���X/v�c�Z�D��=�֬�D7ͥ<&�6���K�~����"��l�ŀ��k��
�\#b,���@s��$�OVP�7��<ͧ�?A�g�)� ⸓e�ͪ=�����B��"=�Q�iԸ]"խt�x���Ol���j�&��S&C�i�r%ܽHWX�;� Y0^ɮ�jܴ�ny�/O��$�O����ۼ?�@�PC�O%�b�"C��'m�ز2��t��3(�1P�5�'W>ЋD
Z%S��Y�fa�1T�V=���nN�Q���R{\�RAߔd(��R��7j�䭁�F�-S<����A�-5ir����NC,m��Bؚp ���ӧ�=F�T�@wC\��f�Q��~��	#%

5��5�!�-0�J�͘=L�h��h��l�QA�oĶ�c�T�k��iP�)O>$�Y�͔"����h��Z�R��	ß@�i�7�=8���$�O��S#w�zуR�P�l�bh�5qp�Z��O�50��>[M �B��	����剜<�0₀��Z�)�TŘ����O>MU��h��&�Q G�2[t x��C�F�pSI>��C�d�	�k�"���f�s��}����L�'�h�I؟�?�Oh�d���C&k�ŢM��i�`m2Ó�hOJ�©�D�������20O�@o��`�'b=���~������V3w,��ܞ|��)���B"�O ���O2��hF;�9���5����@ώ��\�;�rg�y ���4�\�S�.Z*{XQ���Ă^EG\�0#�,I��@R��1{;�-Y�����3�3��\X�m ��n���W��6�.���O��?i!%� 6l��r���<�Z��ig����0����	 9�a���"T#V��hO���H�I�#N~(�P�S�	Ǩр��T=1���I�a�"��ܴ�?�����	� �J���OZ�D��|?�@��v������>ay��$3�r avM�0p���|^�(9�*���L��!H�":G�4�e	��)���j�͔�,�6��p��*N�*l�Al�F��!�1�и)����Cw��;|�����n�C��5��N��h\nd�gk��?��������|�.	G�>�Xe)֩=5fyF,���y��wxJl��Φf��mxP�����'��O9��|��,�̐(�""��Lj���=pl�\h���?a�蟪/�&�k���?���?������OHX`4�ʧ/J9�u�\�B���@Iܟ0�1F�8iG�)F�ci��Iy3�{�ջY�&�v�̎1j<��n���n
_'nL�a�?�=Aa�ĆBh��
p��^�~pp�,EQ?ye�����ğ��?1(�b��g��k>¸��--<� E"O^����J�Y���
am�K��A
Jp�'�N���2�H�lD��Y���Ms��T���T�C�:���P�I��d��Rӟ�	�|�Eڎ9��8w
�d��!P'Η�~��(z����_�����9p~��,�F�&lX@��Nm�lS2���/�rX��lB�uw�]��I�%_��d�O� I�#`X�@'M
2`\"$���OB��<�������)B"2�cƋ&�]�G�=1!��A>0��|b񪇺M���a&�:(�X}"_�4s�n[��M����?�)�B��e�{�|�! IT�2:I[t���V~�d�O����'uU�+Q�ZIخ�QK��6F��Zd$�358:�{G�T��uhCmR2%|�����.>n�qzv W0f�u@o�Q�m��'$@:н�r�G�h�ͥz
Zta�	G����O\������/!�zP
ˣ#�p��.O�%Ҭ��+�)��<�a�Rp��+�n0
~�9 Ƅl��kO<A@JրT`(�Z"τ+R�ܔ�1n��<�qG97�V�'@bQ>�`j���	ڟ��퓁|g&!)��F'/ftXVgH�a�ڥ��`��aO������QHT�G˟H�%�|��fZ�ЃKD=A�$\�ⅰ5�V��T����{^|i��u+Lf���$ȄkLq��eՙeߨ9�À+�(�Q�����@f������W~J~������8?Ny�K��؂���n�H�!�$/q�i�f.E�;�xFoT�+�p���4���T9����c�ֈ�nP��o�,�����O$�\�
�����O6�D�OxT�O�r��&�d5[&�K�`��tbv��6���SN�fq�0{��A/L�����O�X�*�cTp̓D
���H�:�ݚ�S�O����Vf϶�V�{��S6.�~%�G+�vj���R�nc��C"i�E�޼є���j�� k�����<Y4�ן8�	����<A�����?T�(�[�'�rR�!�L�I�!�O���]��-r�� aCT.c}�Fz�O��Y��B����M��$-f~A�%T�2�di VĆ��?I��?���`��'�?A�O���)��[�I"A�C	��-��Z��"nP�4�΁
���[0�<5�>�cs �^�'Dl�C8��rt�}-L���K�7t�����J�G��9Q%�J�.ћ���0V��@>���02"~�x�r���1����@�"t�@ձB������ZyB�'Z�O�j�x�h�%J�z�٠fҫs����#�4E��#b6B'���g��%ΓVݛV�'6剣</��޴�?������F���s����$�� �-���[���O2�D�O>�A�"<�lr��Cy*�:����}�>�#,�
*�����I8�ڽ3eP�m��p"jG*�(Ac�O��<Yc�\Y֩Z�m�DS,�򤀂`�|��o��T�O�y+�M�!sκ%hd	�%�eJ��'��O?�I�t�������1��p�VF_p���dJ�;Nԃ@�/]��K$�ۈ9���	 "o
��R���H��Q�$Lżj�B�'

� �馁�q�.q%'
�R3N		�,�Yvp�`��֣kh�*5�މe��5��EF�,c>�N�)���1���UU���P"�t�[��4�NqrvBLKnҙS���0%� uHs��wc�,S$�n�� ˡ����f=!6��3EE����OQcϊ�rV|lP�C8� k�"O��ѯT
r�\pA���!ϙ��'D�0��|:�X�h�BF�%�����ź�0!Y��?iCj�O{R�+���?����?���R�4�Zi�En�*#����e�6�ެ�dfX^��	:��/@^�{�Ú{��\�d�����y��հ\��Y� -H"��uP�'��`�c����Y2�ؗb	2�C�O�r���EI̓lKd��fF���Qj_͒���j�����y���My��Y����xyBD5[lX!
�*\�y&b�+�y҂�x����x8����]�@���6�	 ~�5�	Xybl[� �ם3(J�[ ��C���@��S6y@������Iȟ�qV�E�|�I�|R�N] Q�4B��Q%��A��p:"���4,��`XQ���FV�x#D�4i�ܣ<��L�)�d��4����� 
�q�a�5+B�8q��� Ojp����.��������e�	?�MKc[,V�XY��K����BF(P�Z�f�'��	��$�?��Q� !^X E_%8^:Q�2M��0<9��$�[���!D �lA2�y��K��D�զ�	Fy�%͡>7�6��OD�D�|��M3#���`����5~.=87V�Uj8S���?Y�{�� _8�0m�'��S�,�|aZ5A�zUh�xt��B��<1��Ԝ<������L0�H9w� "pr`��:��3���}(�)H�d��lO��<��$��p�	/�MK����16�J@��	��5��a(҉77�pmZL��D�>�I�8/�����VS�\��勣nJ��]��	�4�?�f���e��a�PD0�%���<�m�w���'�^>u%N�����t�UDU
(�b4�"䌨x<n�B��3p1�=�1ʋ:<@��L2R�J��VdY��0&?5�]���Ҧ=��\H%���t!�Ǔ�?>��ါ�g¦${��1y8Ͱ!`��q.��ߠ;�HP�w�Ĝv�~@������	���'�L6�Ȧ��	m�S�?������L��Z�v��@�Ю8�Ą�0��ݟ�����P�	jx�p�O���@�r(��! d�Fc%�	ȟt{�4~e��|�myӺ�i��4;`�q!��F�hIC�ʯRx���O�,)��іw�����O����Ol���?��P��|�C�� d<y��V��Р��C܄����<�"��Dѡ~������jr�-ڷ`ïX���wHQ }�@��H�$�����ZZ1剒q4�\�W�_�7�f�RW%�<Z����c���ā��A�K<����?�.O��bT+Ƽ�B(�'O�ufD|"E"O-�b Vl蔝`Q�ߧdI ɳ�e}�'���'�ɧy��S6v���R�*u@� �ޔ�y���6w�PQ�L�&��s�����y�잪U�8Pp6h˖q���Bd��yb�c���Kv'�p�� `sK�5�yR恄'�b����@Ak�-��y���XS��V�D�Fl� �y�J��gSLd`T�.�MQ�ƙ��yrh�C�N�c�*��1kB��y"뇗MXv "�	ds@���y�}�	!ƅ=V���oCB$�yB�Ot�J�i���Ov2M��P��y2D��F�CcsV#�gݝ�y2�4������w��z�_��yR�3^ ����d�@�`
��y��ǉRTZ���,1f�(����y
�g�6�a��.K�"�c�-�y�,�+ eH���l 
WА���[�yM�npj��N�$X<Y1�G	�yb��4r�B �Dg���G��y�#{�6X�5(M*1RVe;�瞹�y��7e��(qE�7cj�f�1�y���i[&i�E�7xA@�� �y���6d�|"enH�_�&%z�I�5�y�kZ)nx�3s�W�� �刚�y�Ӓ^}|�1�[�J-ĥ��,� �y�͟;5ن��IŻ9d�=PDD��y��&M�ȸA��5`xR��P�ݫ�y�� I�L���d�(VkdQIg�䍆�DW2� �-�!T`��V�F�; p���s���{�P�'�����a��~|��S�? ���"B�7��P��	-�B�F"O��cH�70x��s��Y�"���"O��2DG#De��+0$E,z�:��3"OЬ��K�V- � eb���1P�"O�#�� 44P� $��A��Kq"O��#�O;�*�
̜�)�.1Q�"O��qd̅@��-����z�պ3"O���%c.dt@�T��� u"OJ|� �Q�4�V��Q��-o�l�[7"O��&�)1i�Q cd�l���P"O�I�D���f(�"�A�{Ľ��"O��T
4a��;t�ֶ"��ZB"O	X�+V�%d^I�aI��r��"Or�!��d��摟���"O�����I ��(�UC�?����"O��
@��gu
����Y�=X���"O��0j�'c;l�򫖅1J��b�"OV�b���1c�H֊��5>�P�"O�P��a[$0��7&Z�Pb�"O����l7tW�1�+O㤨�a�'?��0F�
[�������P�,��1�(>�kAkԾ'h�hQ��]�����M�V4F�y��'�d*s�
s��Q�Ɔ0b�q�}"D�88����ܕk��,(BmX;�ē��`��6=P�4�v ն0��4:�����O���ھ&^���J��yGNA%��5���U&l��:B���p>�S����QT�R)^��$1b(ƒ6�]���� ���e�.U�"��(�h�+��ĳd��Fx��\O'n���F��#u.p@�l֞�(Of���L=�n���N��c�.qB�T��H�%({���'��`���Z�T��#���=����R���逢¦L����j��py�pR���
�:M�Ш?j'fJ�J#gE=������0�
0���r�1��m�n��e�I�}|<M�ӌ�|��H��c�.g�D7�®U��M�w>�9#t�~�(�$�*ړk��}&ό-$F|����3k�(c�J�	�BJ�RYKpB�&,��I2��(���rƯU٦uH��V(/�^)����F�D�M��g^8�o_�d�j�(!?qdϞ~�l��Q�@�
�H3v���<�ʇl~�k�0jp���i�-?r�Xb�#�MS�B�qq.o��)�H�b� �uB@�õ&߇%>���D^y�Ě[d�uJ�_�hLV�!��W)3�\���NJ�`	�ԋ�'pK�[���I�! m�x��nѡx�h�3���-T�=@T.�%=b<�C��WV H�FM(�a���`�8S��\0s(�D�nx���ӑ%&�Gz����J�r����'iP �q>đ�2�X(��<s�p�'@`��� 5l�-h�s:b��^<+ƬA
t)����P�X�Y��	��ē]�NkF�@٦�b�dܯ�1�7cʫ'E�x;6��D��<�FIO)>��zP
'?y������Kq�,+O�a���<)��|~��(jr�� �
�/$�(uK���
�MS�M��DanZ9N��*!J�p"��ӷ�
7���*aʓ1\:�&/�%��D��!�8*rTP[G��.z�A�b\�<�Gw����ͳ�@ �I� �$��J����#�&VT(P�A=U$��e�<�2��I`�hE����17�&7`*z3D	/R�FtFz����љ%Bh�'?����SjղAA���`�,04p�ׅ�Z�'��X1dA2A�.��$I���خ�4Q��NM��!0�+�g��r~�'��:aI��M�"�5 �`��f�ʂ�<h���@A&���N��zhl�藍�{~b�3}��U'
�3{R��� �$�yR�-���:'��i۬E.�ڶ�ۑ[E����f8,M�ݴ��M���G3<�"T��-35��cʄ��DJ�a����taލt���ɓ@#��X��
�
���JC4O�I��~��b!�ꖼs.&��̉q��;�	��6���{cjCIޝ�b�^�'�Nl�s�E�`�F8yht�+3b_x�L�;���]����;#nd�R�T�_�F��nI`�u1�N�hOT)�������K�*��Rh����c���fߎ��$H�����?l����&E
���)	6C\r6ݟ@L H�++�Aq0͛4�
X	��#�6�1�������<h��l�g�mŦx��I!k!�0��̟%I�dD���ӻ8eV�� �?��yҔLG��M;��ͨS��`d/��ȊV-΅3�ڍ8)Os�'�uP��[p�W#d:��IgJQ7���[-˛E'ayΕ�$f�!!dcA�T��IEI��ĸ����mM� ل���X�{� G{����98��Z�(h4b�ɍ$�Ҩ�����ߪd���!Jf4��FܺI����z�X����TE��K�Ś�Uj9���	�~�ּc���1)�Y1�2ﺄy�.K^�@�60f-ٳ_�x��|�А��kȜyUҜ2��j��	;X3����-�7�]�',D�z\t�	�,ǒS�
 �
�')�]0����j��@+�l�sJ�d �� ���v�oӂM{�NȿHHRu�dQU~���$Ȕwn�˓zjR�����q��}�@PH���b>�@C��`�4��:΀�饊�)%` Zf�d���e��"����q��I X�'ͺ����΂W�٪�I�R	����y�A�����Ԥ��^��:�f��nd�iȞ�KE�6� �pJ/>4b8y����)Q����B��Tq�">��Nox�Y;!��8����ԶQ��۪=>Rа`��|e��ORѲd��x��S��3AT��耧Z�AS�K6`"[�q�ǜ�t	�`�6��`�A7Z��I�$����&����rE��
���3��T��e��(O�LC��2������3s#�U��]�QĢV�ib�xrܤm�$b��0%���"���g��L��E��(`U#��8�4�ېu�"-`!Lb�J�)�ǈs�[�&�"V��E"ҧ��r��9G{��ڬN���H7Ȉ6@��<�w�D�J�$�A�'�hv.݃�(O�T�"D����C�*��A�Q5i���=��	�#AF-��ȓj?fϻp�Љ@�A�h(��>�6y�=�G�5��Wg��04Ј"n�6��)�i �d�q@VEs~R�0�X����6�@�B�N�"}�0���NH�ibB�O�l���6lld��rf��\$�re��K�l�I�m�v�A�'W��H^}N�X�EƫZ%��oͧ^�D���E�d���Y i�F\�w+I�?�$���oJU�Ӏ[H ���a���b�d���D�z��ԃ �'ޠ����i�L9�R'	2�ԍ��ř3(ѴȜ�5A"/Ox͢(O@��?!��_=SD���q芗2e���ګg�ax��#�,�jUT�<Xѧ�	b["q3���o~bM�фQ�z9��C�\�Z�D��?M��/�4[��D���N�"p1���:��Q6�ÃNΠ 5����d��g]`h�fQ/An1cS9yJfxz��	�B$���b������%$�� "d  5��Q�l�H����Ј��b¼D(b����8*��Ćj��ƀ�):�j<�$O��B(�m��$�*�(����Γl��9(����?˓zϲ��0�u��� �Y&��9c.�6:� @�	

��aJɸsfB���`�vX�MP�Ɣ��0��!19R��1d�O��KcHALs�ɰ}�<`���O��y��ףJ�1�e:.����'O�):2ʐ�(8頰nX�f���KiF+p��G�5qp�m�j���� s��0=D�Qo�Vy��yB5���7(I�Y-�@�B�?s��B%W�$�8�i���o�]�''�5���C7J���@MD7,<�u�Lß@2p�$��$]Q>�A%�:�d�ЀM�3�ƙC�>�!�ŠF���ֽ��I�|�ƍ�"���ψ�� �)vi<?Y��1?�.���L�s�d(�_;@�D��-�8;ʉ' 0����'"D���%�b�9w��~�A@a����b��)��>f��	��)5��p�~4*cJ f	�pp�L�?	�W��~R�cy�bM�O7ȕ�5��04��y,Z�N[�mV�4p��@��$
Z]�=
%Q�m^6��
����D�xk¡�C�K&��l���V�"�	�o٘����^Y�u: κ0(�����G�qL 
� � �`AJG%�;6��6�)e@
i�e{��o�,O�sӌ�a\� �%Mu�����E�z���cX�"�-]95������U��p<	c�m�TD��j� }���f��pv�hӢKU$9,F�'�s�>u�L�f"�8�FGč?�R�x��S�)A�{"��'w*TۖL ����+��D �(���� ML�$θ,<�yI�b��IP����Oh����_�f� ����Xk���e3U�D9���޽[���ܸa��q]��ȶ���?"���W�n��X�%bnX�Bg%��%��z�(�HV2�if��(0��X�'��'r!��-ҿ"�X����I&F\Q�0	,`y� ���3��6͘*�6 $�3�`�p����d"@���|��/W��k2��1���!)�*:O�8�v�N�bk�0Z��ΎX����l8O٘5 �^�j�5� 1�4�����P�ΓT��-RS�' ��y�O��iAU�w���C��>��ͫp`�1&�����C�}��{��ΝL� ՚�C['H���
KQ=z�(]CH����Ɏ 0ԡ��b����P%L���J�O.�# ��/:@���r9��1eέ-�����Og푞8iLN�Xdp��6�F�V��Y��/s���e�V2_2a�6�׹���y��A$@�x��!)�j�	����GYE `�F�2`�����Q��:k",4H��#a,�7��s���E��F���s �ՙ_����5VDY��|��9�N���R7n���l�7��d�g�D�.tᲩ��@�}�%=Oܢ1'�61)v�C�(Ŷ/�D�Ӂ��Z��l��BL���'������S���@�A%F �e#MaT���`B�i���$�.�&��]�q�2�PhX99k�@ G�z\�5�ɚA����D�)� �"ot�%i0�A�5u$q1�b'J=�L�5~.�eЎ�$��z������S%�]	�Wt��6z�^h��
�t�p�;ƨ�d���k������r��p������즟�	>D-
�C�׮Em\��+66Af7�U�u��ر��+|��<1O�s�1K�B}+�(Zo� ǉ 3!0tH�%,��2	�����<1�T�mB��(�dC3���{�� �?�"�>������[��651d�>}��Y �hV�+̼H�N����>I�F��8q�ћ��̅u�`!�
IY�����	�l�]��'�1��M-}>�a�㉰Hi�H�A40&QQ҄�#^���[�Q/�DHGχ;�d�P��X%j�ڜ�`�� ��}��'X0��v��;B�ey���.x�C���Vny#H���O��X�DV?Xq�Po�D�`��'��ݑpBM� �\r�( HM�웟'��e���WQ�O?�Їę?d��B�Aѩ�?D�� n���*�v4>-��B�)��Z��>Y�Z��RE��Ɇ?��(0,
M��y�pM�"l��C�	� �hq����k"��+���C�	� ZT��!�KM����$�/+�C�	�k�`9�Ao8���'hǲK�B�	��D����q�H�!��}FB�Ɍ��H!gm�2u�������k��B�+vpY0���B}l�P3�� ��C�I[�������wA`!衈\\o C�ɨ2CN�KG��6����$@�B��:cSlmᄏ� ��`�V Q�,�B�ək|��Ӆd������O�BB�ɨ6z�1`� �Q��ˀ.K�B�LB�	H]P�ʖ%'^0CgȲ+�DB�I'i\����i�$�ԍD(i�B�I�Hb��1&K;4�<c�-�[~C�ɻkl���ʛn���b�B�,�FC�	"��ER��N���3K#3K�B䉵5G&�����VT�ԐqFɜh��B�I���*�@	[O4�Z�H+J�C�ɀ��ibIP33�(yإ$2,^C��	yR�Y�3�@k$a��%yi"C��,�p��4*��U��%g�C�I|5�X ��Г��@�J��C�i��]����\�vQY�BޏU�B�If�"�f
/9����?>�NC�I�^ybՒ ���	�G',kC��9h����s�H�A���k���,!�B�Ɋ ��XQU@�}��T�s��+�B�IF7pW���
�p$I``�&_S�C䉳	%)�>7�8��%#H01��C�)<t�}Xf@)�*�83�Ä�|C��4`���:G �"@��9��b��'lC�I�I�$��ΚC�2d�֩_*{�FC�ɕr����w�
U"PA��@�.�BC�I�i��`b�>64�2�+T�9�BC�I.y�PN�E� �(� ^�X��C�	��tۆ�Y:^������?X��C�	v�EI /
hLpH�1�@�^�~B�IV� �ԅՐ[�D`ۀ ݭ)��C䉣I���A$��1*�\�Y$˝	t��B�I�{Rj0���A�$�!���"	JdB�ɵ|�T`��
�a� ;���\|C䉾�
��r���{ĎG�NC�	fL�1��k?����n�x�0C�ɂ?"將��4*fZ���4T��C�	�%��i��N4y&m���,Z~C�ɡe�<`s2�ؕ?B�2֖jADC�ɝb0�E`�훩6����t��s�.C�	&Oz��3� �<Nۼ�(^�)ٸB��"esr��C�v�L��"�^�;#�B��,����%�vذ��~��B䉐*l���G,�n��(M�yjB�	��rl�6�
<8V��4��9z�^B�ɤY�h��Ƥ^.<�z7�~�C��b���k�Ǖ�ɖ��A.	l��B��+�.4��臵<ƈ�`��ϖB�	�%�R��t��@PbS BXB�	F�`�2��9wi"��vʓ
?��C�� ʼ��` $��`˱�N<W�dC�?	��W?&ܱ�%�LRLC�ɄI��,q�ʌ5�$�U�	peC䉦QȢ�p����*���"�E�!k,C䉫~6rej���!��LS��D-"�B�)� �i����2��4�A��!
ZE� "Oh�薂&(�]��
�MvY�#"O��Y��*\�Tq�
�0��"O�CO�I0�yS�I^�����d"OZ<pA)9T5�nQ��v�)"O
�h��S6L�3�M�<ڈ��"O��Q��jR�<
��B�9+ε�@"O:��k�;V�R��^�1���[�"OL���  \L0��E�X!bas�"OPihak^*_�6�p�Ǵ+;�UR"O��@�Ė�36��A�ŁU*NB�"O�!s�&�{�&�����&p �1"Ot�ڠ�H[>�$��o��2��=K�"O:	a�`	
�:y�h�7e���"OQz���#�n-P&h�']���X�"O�� �٤B�:%]A��ၢ"On��VI$O~�l��!����\D"O����	��-����Y�g�L�br"O`Q	ѭ�,l��Ux�kL;h�ة�"O�0��I�L&�pY�+U�Ew%��"O
t[P ���8Y��dVj�D�V"O:�Yd�U��|�S�ET�R$��"O�r����d\�=C�ٔ�(h�"O�p���J+nȫ7��w���"OL�ٷ�"7�I��Ƃ~�:t��"O<��V�M�e�&��%Tsɤ��4"O��fD��\�́��˼	�@+"OVd����Yn�"0�O+����j��#<E��',�$���U5����~l�Q:�'l��s�Nےn���Z�SZ��
�'U���UC�//��`�3��
˰�#
�'�X{����1Q u�4�/_�t 
�'�Z�0a��T(�"��@/Fވ��'�$96���JP�`J@�(İP+�'j21�D��/���é/ �lL�
�'6yK��1z�� rӮĦɲ,)
瓤ēvj��1b�x�5ƙ|l=��7��a�o�0����و&��ȓ{$�E�IX#bx��+�7����ȓ9�Ɛ�t�N?
R�m��k�?%�B�ȓp xJA��(h�|���M�-p΅��DK�i���]7~�*��"�
5V���ȓ!��� ��7;t81`w�6(r���ȓR���ذ�.niP�$B� ���ȓ�p��V8/l;wCS17�Z���W���'��h�J�R�.�����mR��Y�j̀Fs�0�#H�b�؅ȓ3~�H�E� �{TK�/��0��B��|+�	�3L��1�G^�]A�%���qÂŌ
x��I���?F#r��!��h���_�g'$;�dՒ���]<Y���/�E)�* �g�
H�w��N��&��9tb�C�@L����4����L*D����FM�+hn$�aLX�Gl,���M5D����j�.�44���*7�\)��e3D���s&л"��4�<��T�A(�(O��}�ze<���	q^Դs�� �-l��ȓ_<X|S�I�4A�X�Ig߭XD4���k<�2���T��ʭ�p� G�æy���)��a#2�l*��/��	`�LX�!D�$�Pᙿa� �B`��"���R35D�И� &��hJ$
�7Q��ѩT�>D���q�R0=w���LȪ;��bb:lOh�d˃R&!��Ha�@�;u�@��v�:D�� h1���Z�tt2xr��͈Z��a��"O��&My�>Eh��[/z�=�r"O�P@�ŕL!�Xe�B�<�*q�"OP��W��7v�Ms��ND���G"OdY�5��8�8�Q�٩� �""OxP�u$Y�N�b��΅�RcָK��'����rN̵YEj%��!\�&=�}��*D��vb�	5���˖!ي���eDHԐx��Ì�Q�v˗]3��:�@�yBnC�z����Ċ
W~��M�8�hO���$?[�ΕYb�	����$;�!�$^;���TK�Rc�Ab��Q�!��21��˕ :ap��Ft�!�[Xj ��O�y[� ��挩[�!�dH*Il�8��ðSp��P�
�!���i'|�2�%�RF���S�ŶW�!�D��!!U��<2Z��&)�{�!�d�$(�:tx%ɩ+)�9{�g/m�ƝG{���'�ȉ FZ~Ѹ����Ҵ4R����'S�����ە �B�U�*l&T�'^��
��1a�hD:�H�O>}y�'B.U(DȟO* sf�F�Hp��'��r� 8"�v����
9P�'�f�Qr��+��#�i!�fɛ�'^�m�`�љO��l[��I�R;�A�'n�q9��Q�}	Z�`�H��4y��8�'���uc�DtE��Q-'���'C^�C�,��^ ��Z�GF,)���C�'Ԥ 5OB0t�y�ć
�8�I�'�*��$�Y�nD
aB��:�T
�'u"�h�<Q�ڤ�վ{L|<�
�'�b0����%���@u��n߀�
�'����]}�:`���e%P�	�'���y�(~���Sw��(jɮ�1	�'����%6Ӥ���+�)o��$Q�'�,䱷��zc^���B��4͢0{�'8@	�C�`��'�"\��Z�'�:��+�-b�	�f	�%��Y��'rx�pD��*�4�c�J�j��
�';bP*f��J@i����
	�'��P�3��qɢ`�lN��'���$��0jg*�O e3�'Q��+��V%S��Ag��6y�YP�'rn9���ϱ
6��@4¤*���'=�p
w��,��q�͒#*�H��'u6�00eJR��$I�%�p�s
�'���[�5�q��?ƼԳ1O�0�y���28j��  B�<[�`��D֚�yR�ϡHf�P�*���ʅ�W$�y�#϶(��%�*�����B��0�yӚqIR��"Y]�!��"�yB����T(�p{ ��9�y҂�,s@m��h>�BX@���y",ǈ7��C$�Ҥ��`I���y��k��]24�,�B�@�eH�y�����3��I�_
U�V49
�'+�9���+����H�Y�`��'�LԂ4!Ęo���iF,D�t��X��'��{�&�'wM���B���V���'�H S����y��^�����'t����8Y���8 �\�Rj�%q�'< �AbJ�#�L���X2"��Z�'��-p���6�<
E�����S�'�pUB��e||D���ƈ#��I���� 6���ٕڦ��ѧC���"OY�a�Ĕ'��P�B�-�RH�$"O$�s1�� *e"�s.�J�"Orax�,�o��H�g�{\��"OP�����;c�8T� ������K8�yR%T2
~����@�&Ƽ��%@��yB�X��2����^�.C8xH�M�)�yr�KO���*W�u����u�0�yRg�d��JD�h�x�F��yBZ�zN��h�ɇ14\�(�jϰ�y,ا<²䁷�I�Z���
3���y�-&V�LX��̚d����!+̽�y� �	M�
���#ϊ��AX`B���y�Eޢ�<j�H�sx�:��H;�y��Z1E���)Z�.�����H��yBi	7U�[V�%��qy�^�y��,:�����3���6�X�yb�N�N(�f��^W ��v����y"� t`UB��ף`�h-�1�2�y��������_��𢇊���y�.�&w����dGY�rrE�9�yb��+i�,8Ug)Cb��s�N�
�ybۈf�b�r��A֐�c[��y�M��A��Pi�ND5��%�J��yR��d-rҨ_(���)�yR��?(Va+�%�j��̇&�yb�T�
�| ��Q�������y� �+#J���EU�l���ybc[�k��!GA�� ���XP	
�y�h�6wz0T��Ӄr��ip���y�LBd��pi�k��p�N��w���y2) ��M��U:j�lwIP�yҁ
�V:΁1��0p`=�vC@��y�h���"����")�D��qg_�yRLZ1�� ��-�j����Պ^��y��
�HE����%J�t��L��	�y��P׎�@��sI�������y҈t�T��d�33�`;V�\��y�P	��-!	�ׇK#X�༑�'&�h�S�0p�:���+��H�DTH�'���ug��%2D�Y��=��HB�'��`8c�Щ"@��g `��=��'\��dV�%��	�M]C��q��'�\���X#:4Z�ٝ8{ ؐ�'��Ն�(A��m���hF(-��'D���3Ȍ��$rfO֭g߶�`�'�hq�Ñ8mڊ�`v/�e�p%�
�'߶,��L�;l�~�ʦ�b����	�'�\��C��.<����[�o��mr�'���B��qXk�n��6�x�'�p�x���X ��h��7�iP
�'���	Oޏf�%3��k&13	�'�lYb��"Xs�RvM�+����'	2�3�c�V��G%��3씂
�'xިӐ*��F.�)�/� FXA
�'����c�� �m��b`��'�.)b'���I+n)������8Q�'Z����4��*G�� sc)��'j%�PjY3i��0��M-p[��(
�'��� �!8EF���,"df���'���6/?�[:�Bd���'�a���,~W�-���`?Py�'����O�٨�ۇ�X�_��I�',���t#'�P!���?,��}��� D����ń$-��R�����lz�"OʅaW�C�T)�dJ�n��}�(�R"Ob�s4+M�Q�
�����?U�"O�!���	 :�z6LM,C���"O��s��E)`�̓��IA"O�E�!�[L���pv�1�Ԙ��"O֑�`��7�� ِ��PP��7"O��p�9&"d����>"�"O�X`���a�N�z�/�`7���"O�� �K�/NxT�o!\�䠁"O�Въ��jk>���C� ���%"O^�#�,ЏD��@���U"a��2#"O��*P�ZwÒ�8!*E�86$)z�"O
�	��7��z 
Н-��ٔ"OH0c�M�P \E��j�23����"O���� �0%��8��U�@�$"O����F�7 E�6��>�v�E"Oaq�-�9�~�y0�ݗ;�`��"O���RII9��zT��:>2ԫ4"OB�˓A�!U�Zh	u�]�H��"OR�8D��vǞ�	b则"�J}��"O:̱�n�w.���%�çxP Iv"O�ű�,ْ?%`�
6�
5� �"Op�@a��|��c��ӽR)Z��D"O��k�#E�IY��X��-x&����"O���"����<�Q � �W"O�q��hO=/FQ���0D�0�"Oj	cseP��ј�I�'o�<�I�"O.|� ǃbl�%Q'��`�fرP"O�hW�3]<���ƅ*i$�X�"O�=0&!ӯZ��W�,B�-S�"O�Y��.�/P"����ާ�.E�!"Op��	�T��eq�[?v-��"O�p��(�-}����m�N1�T"O %`����y�V9K-b��P�"OT�� 5bM���/���[�"O��*�
:���ID*�d"O��BBL�gt����� #���T"OlU"���5���𧉆�Ĥ��"O^q��Ωݮة!�S}�8,�D"O�L���ڪ-�Z��% ր�"O��� 1h�:U�1N��s(�0��"O��BT���H�<u�U,��!�-�"O��3�⑏vT$
�ͅ;Tl�"O`�O+yodIK7�L"V�:�$"O�p�.�1?�y�v��Ja=3g"O
���OlV*S��EPU;�"O�}��l�:|�\93�.�K7�m��"O��aW��T~~e�w*U����"O��c�.:����AP�a�����"O4Ԑ��v$�����>"�<���"O�5�d ҆"Yƴ�����{w�u�"O
��W��;`�8�j�թy�J�3"O4(	Չ�	���,�/c�*\��"O��HsڒB�ޙ�-��jڜ���"Or5��d��ڈS�+�k�X�ȗ"O�4�1��t�P�X+�z���"O$��En[���Q��ߙikR���"O�U;��
{nV-�a)I�E["hZW"O<���=D�����ۋ�bti"O، ��G�����7���@2�"O,�R�a�G�2���g�EhF�;�"O�Ta��&�bp��$-b�\"T"O��"W�6���ȌB$a�"O� <��cZP���JJ8z��"Ot9P'@��\S@%�@"��Ѐ"O�g#/9?������Y��"O�X��悬3ܜD��:���P"OԈc�,��p��U��Y+3I�L{�"O��U ���b�����e:\d�B"O�ma��./�����ʬ'"���"Op)Q@n]�]��=I�DO-k:���"OƤ���Z-S��l�G!�Zn���"O`<��|��Փ�mӱ,�e"O�9�Eu� �k��3�0��"O6<�3�Z�p�Z�sk,-� ̪t"O�-�흘 D$`���@��0��"O��nQ�B?��HD6���r�"O.T�0���-��A3���D�"O0�# ��	+�cӅ֢-��d""On�#!$ٝ&P��'�y�YQ"O��1�-� �PxZ�e@�(�f�"O�1f��5��jU$��epR$(�"O4�'�[�e'ɨ�>X��"O�H���Ҿ%P�lk����9`�8D��s���f���"� CCn�YP�)D��v,�`_��%��	P�Eqd�+D��  ّT�^Ur"'Z5�-(��6D�k�̦gBR,bahW�I�0�9�8D�ԑ0 �v�FE ��a���U#:D����@JF�
5����V���@��6D� � i<��g	C=Z�C B0D��+%��p��a�A��I�X�IRK!D�@�u�٥^\^dQ�^�G
~!3D�0�`LO;?���'��B�� .D��1gIA#A֌����}�v���&D��@�'��h�X�sFؕ�<c��#D����G�:X]t�xb�U�zz:�K(.D���W��j����Ҙ8�ޭ3G.D����)ڡ3P&8	�*Қ����D�(D�p�୏��l ���051r� �(D�h�k�|�楐���x�P���;D�<YO��n�0A�"#I:'8Y#b
9D���f/]�� �a��nʬ��5D��)$hSg�ڰ21L�O�ryP��(D�����ȟR�ntR�J^��X�ȕE(D�r��V(a�ڜ���' ��a�	2D�p�,��ⴀ�'[8/
0�:��.D���@�Y�Pa2��;A@�i�g"D��9��G�v�rE����ZZcS�?D��p�I�@�&�H�	��f!���!�=D�B�)_#Ur�!��+ӐV��8�C
6D��q�JѾa':�ӕ��7N�ؚ�6D��A2�f�������w��Ǭ?D�����*}6E���֋k����&9D��"�FC���P+GD�?"!0���L6D��b�!э�ze g�Ȋ�&�8�5D�@�d�d����KImް�k��2D�d��EU�M�<DB��Jg�9Y&j;D�D��c	��l��c)��}��=D�@�s�I�I����CN*�U[!�(D�ȣ�͹�ޠ�!�˰o����Ri%D�􈱎	j�v��3���8! D��#����e� I�mX�	Ȕ!��B��6Q�A�u�Φ.Q̅H�*oNC�	�n���{���k����C�� ��C���®X&�ҹ��bڇ	� ��"o&D����>B�̡��".����%D�� @xEQ�Tƈ��n�<v��0�"Ov��F�8/��ٰG�.\o�X�G"O����@�_��#��I>3oĄ�"O��j6�o-ph��l�MQ�4RT"Of̲G�)4���J��Z�d�i��"O��s4��<�b��5��O�Ɛx�"O4���;X�|�V��:#w@h!"OX�Z��_	=PTu�$M�\r&��S"O�D6FS�	��붦iUܡ��"O�D���Z0.l�]�Co�5T��rf"O|��B��-�&,!��ISh03"O�%3F��m|���p$	�%Lx��7"O�e�C�I�]���7m�3Yc3"O����L/#��c4�D�N'�dY#"OƤK�o�/)9�բӋ[���"O����&<4�Ҡ#Pm��8�"O���eh�n tL:���<�>� E"OB��'g�~�(�ɍk��9��"O>��F��P��eD�f�`�'"O��%�9/�)`�
�Pa�)Ȁ"O����D
�5���7b��b:F9j�"O�8�5C�q��葑��0K��j�"O���פS#�ɉ%��#F�2��'%28b���lM�1cQ:G��'���;�M�|B<x�@�&��'�4�a+
�v��Ea�S�38�B�'{��H�Ƃ��c�HB=0��1	�'}@�K��\0oT2��0ux�#�'W��Ո�%+D�YC���"p���'� �P¦ �f�2��!�J�Q�' ����5��/��_�`{
�'���J%�j���A��|E̂	�'|�����'[�jl����*t��	�'֜�E�&m�"�x�$�K```�'e���f��c��$�Uǎ,Du�p��'4D��Mvq<\{%�N$x��y��,;�>Agϗ'�B���'���y�O�2Ϙ�8�h�,N��ô��+�y�\�<���ip(�9;�T�����y���a�(�hA�١9���УD%�yBL�|R�s�IN!	�M�`�J?�yB�!&�zӉW0*�d�׋���yrI�DڜR%�H�q�2EC��%�yb�P&�!�5%E�A�R�a&�E��y�+�r��$�Cf	<M �y���y��&S-����� #��̹Ġ���y!�(clX�3様���5��.˝�yR-��*5�hT�	r�Y{����y�_1 R�����U�b�9��ҽ�yJޝbBXa���C�O�И���׽�y�dP�\�.-�֢ێF5ҵ�D���y�n�&6p-�'i��C4nM)����yR��"��\�:�r��@��y҅٨@0�	�3U�`2C�Л�y��.�n0�WǇ;�����;�y�d�5#/�Fd"3R��0L���yb���
��ᑴ�� V`�po�&�yD+�Z��O�E�M�@��"�y2�R.W�(+���1.`�.�=�yk��P8�h��,h2�yg��?�yrHf'���N:/G�5x���'�y�i�iЂ�q�C�o��}kG쐡�y��*B� :�Rg�|5kGn΃�y�
S�>�J�f����cB��y
� و��.}�^ �����wb�1�r"O�|��P�w��i���)�4-PC"O.�Y�oQn[���7��+��f"O�(2���et`�bTK�&ܸ���"O�LZ��1��H�CԖ��)z#"O�H���� _��)��ƭx�V���"Of��gR-l���'e�6(��u�*O����}z^� �cC�?��� �'�DI@�
&���N�5�x�h�'�Th��)��I"f�{�⒎���	�'� @!�O�������#��p�
�'��-��Mܻ
 ��$ ɀUr�'�`(�V10�8Q��7��u��'�Req�iՋ`l����7T&}��'&�ZB�� <���5ܽ4�&�'�Rm�r�8\�z�;���%���R�')��UmǯU��!R���IO�A��'ˠb�X�=*���`ʞXвDy	�'a�%X�/eh-��IcA�
	�'g.����Ь��pB��/W
>��'ϸl�7(է8A�B2��_�<���'غ�����;2���퇄Hv����'
�z�ΨZ���q-|l9�'���YY�5 ���W3���š
$�y���){���hW�[�\�$�s�i�*�yR̅�@��1�M\�Zn@�g-�yBM��l
iԖY^5��
���y�@��^a^�õL�D(ʉ�h(�y�л��a�tN@;D]�%�CH^4�y�F,9G�u*l��1�����E�*�yj��DЂ�i2噫,Ů@�ԥ�yf�b,��Ѷ�XЛ�I�'�y��Q"�8j��-@� \�7�8�y�'�=9���+�ɏoLH1�bۅ�y"g̦p~h��K��܄�3�ɍ�y�@�!��X(Î'`�H��P$�ybJ� �ʰ��͐#>`���N��y"h�2�p�೭�?��%Bb�5�yR�G �B}8������@���)�yb�� ��p����B�1q�y"N�xŖQ�W��1
�`:sd���yb�1B4L����;������yK
!W��5��P�w���x���y��܍C�H�� cF�TDkƠ��yr��.�L�%J�p�~Q��HJ��yB�U<5,\�U�B4e/���J��y­F��bDVAW�U��=�pN�%�y��8K��-��M)S���KŋJ)�y�I�H��*�} ��@�P(�y�GM�n�*x��ɪtJ��J�",�yr�ߖ\6�ؙLQ�e���$���y�ۣU�Sr̍�_�����y�Yۺ}�! �!0L�G�(�y��P�`"�L�&�x��c!]��ydV_�2M�!*�<GbB��B瑂�y�	Z�dU�u��A�b����0�y��
���R���6�d:����y��Bz�2x�lL1($����.��y�n	#���b��
 ̈́=k��0�y�7H�xk%�EG���ꚹ�y�.Hk��BnH���*�
�yR�Ӛ+Z�uc�K=A*�T���y�(��ytE�0)��4
Aq���yf�;������(y�8yCO�:�y
� f)CLן;yF�uʛ�?�|��"O�(��N�0!�l��6)Rj$��e"O���(��*3Fd�VH0F�Z�Rp"Ob���oA������G��*�9��"O�䫢�R�0��ՈЇA19�>�H�"Ov��嚍`d&5�ǆ�%�H|�5"OL	�p���&Y��v�+D"O��0"�D9F`0��/YY���s"O>i��l��Ek��y�"R�]D���"O������Nx���H�	��ęe"O�Ț�.�cn�����: ��(s�"OtP��P�%Qnhi J�&�3d"O�=A�:x���A�ˇ�<{""O�)�#ׂQeBdx!�F��.<["O��5����yZ�@9H՞q��"O�ͳ�"�7�p��2d\��"O����
�2yxV؋���":"��U"O�0[A��,xR1�qb��|��8�"OL\��fEͬ��F��� ��c"On؈��ǻT}���R��F�XJC"O #�\�ƚ��a �"�
��"O��#'R�BH��A�� �n=�"O&���e��?�ɲO�bU��8`"O�A�"-�+z�XG��0n;^�q"O�u��b'c1"I��럓B)� �Q"O���B�ԫ�h�d��o#���"O"�!ꌓo{��V)��,�L�Z�"O�\���_�5��5��-]<�H��"O����#K�W�=p7Ǌ�iHp���"O��)��u�� h���k*V��A"O�|Ӓ<U$\�$G�(�j��"O�tk5b	<����Q��$�@d;D�:1�B�b\)�v�RQ�`�8D��:�n�	Mw�)7�.`�P-�!6D���Q�H�A�0�1#/�V�i���2D�X@�I�v�jܢ�S$c��(��6D�����=e��	kQ�Q�M��ˀ�*D�� �8G��A�F
O�(��$&�-D���Q�lH�ȥnAi�D��E�,D���V�œ���C0]�|�U�*D�0+�F³-S0��!!�2,�|��b%D�l:W��=K�(ձ�e,WR)��#D���Ȧrd�
��Z@�ѧ<D�hӁ�̼�#P&�BU� d9D��3rœ#BX��Sn�'[Z1��"D�ct@�'1l	��+ M9rH[�H+D��u�ͥ�l���c��XЀ� �*D�4IFo�}g�8&�8$|���j(D�4��ʞl�<�i���0��(D��cG�:�~%Yu��2> ـ�)D���Ĉ�2採 v�B�/����m&D���h�@�̢5�T.E0zh/^6!��!YYUL���ukTE�*`!�dH���5� :�����W�8!�DN8P���1#�%~� @ipf
�
!���a$��pK:o��h�A@��r	!���n^k������n��!�$��X�@b�e��4*H}$ �!�dn3*������ 5C0ႡV�C�ɠa�r@/Y8F�9GGR�-	���"O����MJ�Yzץ2�a�"O�-���J�&iV�QѤV)�P�	"O�Y���{��D=e�|�(&"O�,��n��^M��hg�J>y�~�13"O� $]
5H"i�B@��%�3H���v"OxH8U�[�]���cEJ���B"OvK�H�7J�z�iJ�(��xс"OX�I��FhD��Dj���e�q"OVx���!f��p0
�2k����"O����gʬp�R�օZ,� �w"O�lq���qEn8RI#
A��"Oڍ�#Q�	s#m��`�"O�xIu�K�e�r9M��(Xt�a�"Oᩁ��.)�<1��6�@��"O*ثS�8	�h1���v��"O� ��	
J�b�c���,cSh�ʕ"O�\�⌨t����|P��+�"Of��w*� n�b!�C(0B!��"O��BV�{(�RRL�l8���"O{�ҍ�����C-k���x1"O����R�]n���	:9�u"OJ�Z� �f\}����( E� "O8�0�ϲu`6]Jħ��M#���"O꽋e�G"�mZ���W�8H�"O���ġڂr^���q�0���
F"O��SwLN�$�R��`掜Cβ�)�"OΔ�C�͏; ĐSqÅ]a8P�b"O����^;VExK�K�YmrxA"O(�zg��*lB�bB��tXtyD"O٩�!٫N�Z�p��I� Rf�0U"O�ձcI@�-x�+%ۖH��q�Q"O6P�ti��Lۣg�>��e��"O���s�Q�A�X8Y%@]��"O �9�	%���s1�I"`���d"O����;�p�!c��,����"O�M�`��w>$��� ��1јr"O�A���Ws�@`pީ("O@�$kB��x���.ڶ,�T��5"Oz�BE�+ϪtJ2�K!��R"O��;p�W5I�P����`�٢�"O.���N�����.)g�*Q"O��z�-�;r�(�r'MVl��X'"O��3�oB!3�D�P�R 0�ܘ��"O\z�Á� ��ժ'�T��T"O<��� Klz*b���F�h��"O�(×�M[A�es���\xۗ"O����φ�R'������Cx\�PB"O�u��iH�H��+d�n��P�"O�TI��~� P�^.N|A�"O�Ug�H�D��h��ٚvP��6"O�JǍ��z6��	�Y�K��� �"O��"tK@�A�d���ۭ �J\J�"O�� �䔊�\B7�ߛ	�D@ �"O8dJ����Y�h�c����5ܖ��"O�,�2��mfrEhv����q�"O�}��b�����ѥǊL����!"Ox!Z&!@gj�p3��[���w"O�xZf6BΥ��P��0�"OL)���Yxx�;5��8`� ���"O�`����t���ݰt�$��"O��nz�X�d��f�α�B"O�ew.�:,Rz�X5H�*�:(��"O���fL�X�h�Ŧ�!O���F"O�TZ�ۡS�l�W��/	wΝ��"O��B�%P0xGL˄��=XB��b"O��z�FQ�OO�3b�Юc����@"O�͉d>b�(S�+�.�:���"O2���,N�l���)w�������"O� @����N0*1(%�g+_Y���ۗ"O�`�D�ŀX��m�H/>��!�"O�LAoߧc�J@jb,���`��"O�ɛL� TB2A*7��+�0��"OD�" �=l��cD�줊�"Onh���%t⬳��A�8��"O�U�F��yЊ�jZ:b�T �F"O�(d.J�Y�DHC����Z�N�p�"O\�7��-Z�8آgB�y�tPS#"O��$M�aS(���o.� \B�"O"a���S�@,"ς� �b�"O$��R]
bz(�6`�A�v�+�"O�`��lL"B�`���(�)p�"O���.[1<%"�Ч"���ц"O��KU�V�0����(1\��(c"O̝{C�١ZW$!�&O��6I"�q�"OJ�XGE�Wvځ�@LȭL:ֽ�"O41�@�x�Bꑕ!:V"O��E�*]eZ���zA�"O���TgM�7%��A�&�FJj;!��t�l!��ř�hc��2��ʟ"!���FRBSv�oe�� ��4y!��Ҵ&��E��G�2b����Y�%\!���k��ű�M�I�dbU�f�!�$ľ-_����ʝ���t:6��P�!���������o���bB�_$�!�Dģ)��hq�$�(���C.ʝO�!�d�'W��C��O�~��(c��8u!�-q�!���^o3X�z�k92�!�D������I*�D��5 m!�U\ָ<��n,#`�S�뎫}E!�̋��F/(9�c`Fc7!��.8|5�U�JL�u;&Yd!��V)a��6a��+�\�c�G�!�$�{��@���_	[��c�-E8l�!�$�Wɚp�f@�
~"��to�1x�!�$�Zְh2�uc�i�d�#4[!�D������hM"&MXň�+���!�$�l��lb�G	�G��c��>X�!�d(C���t��1l.���r�8i!��ډ$zq����0(n�k$ X#]!�\(��:���,�����%�!�~�t�2�_�Zq:I�a�!�dD/�x�H$+�<ފU��?c!�F�Q"�l�� �E�
G 6pz!�D��K�0�C��B/s֠�� "Is!�R����r@W�
.��D/ c!�d� ������9Jy�![o!���3"lL��֢	(�����~�!�,�����J���t���6�!�/�09Y�u	�b��1�½��"OڝZ���O���lX��yc�"ObL���O�*�9�lV0���r"OPe
㋖[�6�
a��� 
�"O�Xd �/G����� x��i�"O��7JK�\��h�@/Ȫ,�"O�����ʧB�4�p�P�P���i�"O�EHRmA�+���PU�U�!��	�"Oj�)�)0�(�Ұͅ/`&9H�"O���lH�G&��`FmB&P���"Oz�Ԅ�9F��� �C�a��u��"O�i�
mj9�T�� x�|X9"O"tؐ�_f���	Z)0�.�qU"O�	Cp���e$���ߛB����"O�  �q��&��G��75�� "OR�Jf��n*Z�[��Z4wA��"O����լn�,��#����["OF�i�HJ�������i�:E�"Oh��%F��Iaш��/���r7"O ɡb�Ȋbդ����K1T��0-F��m��q��)�&3D���'GC!�@��_�!�P�H/D�쪒m�5u�*��7��e��0��:D���� ^�VC�p�TFŇwX�`�W�:D��b,D�a�|���GC�w��${�"8D�|���?[�X��� >6b��ea)D��k����*.�m�c��!V��bK(D���T�څ,�ұ���{&F�BeJ*D���Ʈǖ/V$IE�_8��.'D��#V����$�j�I�YB�ိ2D��C�;^�|g��;S�© ��%D�8�T��h��D�1Ǌ�J,�a@Um$D��Є�8�{��͆eU��!�#D��V�υ�x�Pjѡf���� C�ɿ	N�A	F
r���%A��/&hB䉃\x��h��)��`B��߂<�TB�o��<�'C:��0�`�I11�DB�	 �|���̙�y����$m�@�~B�I�Z��t����+Ϣ9�D�1=�hB䉈,�Hj�N��3�(T� ��?.�C�	d��x�$��l�SD?G��C�I�T�T��5���Yt�M<��B�ɝ=�4�f��RR��Z5�W?	��B�I�7=�m���R���c-�]�B�ɫJ�"��d��4&B��� ̿>�B䉰2�����ַ$��M�˛]'�B�I%w7ZY3�k�S���K�b�"C�'o�B߷;�.�9%�۽|G>C�I�9�pps��	!2YQ����g�B�I.x<��Cci�	����FC�B�I�"�M��G�WD�5��»W�$C�I��T�)SM��쑒��?UPC䉻x Seh�&��h�r�Aq�B�	:L�|S�iJ6or�WDG5�JB�I%W�x�y0l�7!��s�	eTB�	�b�D�
Sc��V��\�d�?dRC䉕|�4m��m� ;b2t�U�ʶoDJC� ?
R���I��re,�5��C䉧i��� ̌�$! 0k�j�<B��C䉺gǬ�pCk�*RGĹx�a+8,6B�	?jժ\��� _����U�I�R�C�I
T²q�w�֥&��$/4UZ��:D�<����:�	XA��f��p���8D���W=}d��BWe��i^\�d�)D��qf�H�y�|p��I������"k(D�xB�k � z��K���$\vf��G'D��ڂ�B�^�2�P�{j��S�g#D�0.�Z�Bs�-}�43��	O4B�əWG�y)cW�jǲ���m2J��C�I)?�0�V�c;�!�v&6$��C�I+\�A��04����C�Y+u�C�I#F��Y�e�gAP��d"�)��C�	4_��W�R�g�Ը5վ��C�	<���r�nSK{H0Y��W�a�xC䉭tRzX��Mƃ�@h&�N�B�� p�ĺ6*�5nnL8���C�hB�I�TW�;"@O-x�l�����h� B�	w �$3)PzH<xr��/��C�)� ص97	ZvY>�
v��H8�A�"OP��sBb�T�
�l����pJ�"Ofȡ _�
�rI��̔8�|��c"O�0��
�s�`!)^8��5��"O.�k���gh���R�\ �x%"O�*c��og�t�C�D	mJ�s�"Ob,�dbY5�<T�1FN$X`f���"O6D��E%/Ӏ(+㥋�4�z�"ORh�.X~g � ��J�g��,a"O^�Bs��`����!G�@)�(�%"O���T��!�f�@Rk�i��Tp�"OF�[��� :-P�#��8{����"O0�W&J/
⊴��*��Z��Q�"Oz� fD��T�ahǺ����D!�$�<��u ' �*
3伳�lߑ%!�ߘ/��Ւ�A�3.���T� d�!�Ӄ3��HKn�I
H�QPkM�.�!��5O\��Q�]
U���B��	~:!��5q��dsW)Fz�B٘��=3�!�d� ��9�*C?<�Flhd��@R!��ZոR��y���%EAL!�*�v\ �GilJܻ��� :!�D�ƚE�d�_�T�:İB$�yK!�DDy�n̙���gV|��_d�!���6���*a�ڈ�|,(a��k�!�ƻ1'�(O����0!V��%�!��L�E@�IW�F6����G�@!�آLF�	b[lEZ	�JӖp!�d�7JKt�c ��J� )��
�6!�ĝ�o�[T��8Bu�}�4�Iu�!�T�H����m6���\�7!�$��),i�t@޻hPp\�2�8u!�$Q���8����P ���46^!���%���A-F87����M�wU!�DN�i�4Y��U�,`]qЃNw#!�7�+i�JN���LX�C�:r�4��
��<!��$z|�C�I�"`5�@C_�.i�F^��C�I*	��������T���Kb�'��B�	�G>�;ք�3r�ʄ���1P܌C�Ɂi_����F <U�΅���A6?XlC�ɖ)n����m��n`x��@wvC䉻9��� $��Y J�cB��_�*C�	:J.܍������hw/Y�C/C�ɷ$y��:5J� �:�	�,�z�B�	�>��)R ߬bH^|S�Ҁ#��B�I�?��X!��/q�������M�B�ɛ7�0Z��C��ܼ��OA,r�LC�I%2�"G�,4Ƽ��Oz4�B�I�Q�6�Z�	_�NT�x�$�C��B�I
�t���cӓ��ز��*)��B����pB�Ú8��:���8D�d��
*C�V+4B��W�0�y�ʕ#/V��CǤƎQ�l�'c��y��b�Ze�sb��	���/�yҁ�j�R���5$ m�eO�y����h��B�\�d��E��=�y���G�nd	Ҥ�*Qզ��ä�y�/�����H̠;{�@ie-<�y2� �!�LLaՌ�$ѺРW����yr(����(P@̡�7'�;�y�)���U�"��K�m��Ϩ�y�Z{�����ڈD���K�y��	�g�Ҭ��	�6T�����y
� ��"�j��D����!�r�;�"O(�jpCЃ_yVcT�1Ъ	�V"O�Q��	.<o\�pl��#"O��a",@&0��-0�
 1xP��Z"O��ᓨ�>��doʔz�:�B"O.i�ᝦCf�%�ΉD�"���"O� �k
�D�p\�-Z�� ٰ�"OD�j�F��5K�2�k�/9/\P�p"O,$Z� �:D�d��B�%Y�H�#V"O�̻�F�+q���a��&<iP4��"O�TK���A�441��%j���(�"O�j��ccXX�Qh�C�1��"O���ꋜ>�n�H�-وq��T`R"Oҁ��L��{���8,I�����"O�Q�Ŧ�Z^h��wJ"�
�1�"O:�₏[�(*���u��l�����"OИ1v�^�H���#���R���P�"Ot%�r	�V�
�A5�I=��e3�"Ox�� �W�>�d��c-�4�� 2"O�����ǀ{�T�W�{b�rw"OL�r�K �Lܫ���4���G"OX4�®ۍ͸y㠌���M;6"Oڝ��Ƿ��
ḃN��3�"O���L�7~�	w!�_��D@�"OX���K+
�.�y�m�.� �Q"Ol���J�;
[ �c��(٨�i�"O��*�I *Bz���W��<Y����"O,�	�aԁ���JQ�׿t�<���"O��3���3�z�b��.0�~]9�"O>}�l�=h�2�1,H�s�x�U"O8��B��v�=�t%B�/V�
!��Q m;
��&M�$�x��4(�1 �!��2V-�����\
������!�.J1���TN�5�5�B��$*!�/wNͣCA=����dB' !�S$݌�iB��6?p|g��`�!�$!B� z�
�E~�J&A�,�!��!�m�ra ,2Ӑ�a2��~�!�$ݠg�q���.&��e����>�!�d� z��X%�ʡ�t�з�׎f�!�ԑ"^x�"���� �;􁉷V�!�D׿v���)$֡T��0	%�D�0�!�dؠ-f|��K��f�������&�!�dh� ��G��A��� ��C�!�Ͱ `�D�Ͻ@�1K���:8�!�D�&�u�lF�t����c��V�!��l�(�I ��$%�G��dL��M�v��ҮL�`~��3,��
a��6!pT!IZ�e f(Q!ǋO,X�ȓ'�,`���/syB@�7��,�ȓXLݹ�M<`����&B@:���q��T�I�G��
���q�����&1X��d
hv&�"G�� R���ȓ1�M��=�\zp�Z� �؅�V�t"�~��hS$�A�JB��ȓ`�UxЩ�'N�Rƍ�2Q����t��t���Wmv���%��#�>��ȓo��떨|E@�jv���<���>��-R l��t8�`��f�X��Q��]S�O'V��3h�6Q��)��ws���p�O&sP���D�P�5��?�tӴ���|��0Ss,��D�ZŇ�s�
��ъL���
�_	�4��^LL�2�`��G>ASꑢ/�I��S�? ����W�n(`��E�Gm��"O���ՖR���jT+L��"O��1�H�*X��� G�Z�L�ٱ"Of�3��UN�2�A"cp��`�"Oҕ�W�� ��*��&gLbIr�"O4��&�Se����X#���#"O�lӲ�E��H5Z�n�J�R�P�"O<�S�I�=2Z�8-,1�||�w"O���-��k� V@���"OZ!�'��6���Ó�^F]qb"O��������N)���?jF�4H�"OX��v�V=E��x���^8@���c�"O�p���ƑQ�@������A"OnL���
�����E�$k���"O�dGI�s�,Y��T	*_�%H�"OF5�d�C1
��ـ�ƞO�fMh�"O��"�M
.����5Έda�"O��pR=F��1��`��m��"O2ቔh�	no��"'){��h{1"O�Lb�F�A��1�eѼ iB9�3"O��G��%<Ov0�Dӹ{C�%"OĀb�U�4 �	8&æu8\�S"OԱ9��	)&22�Ң��3'@�T"O�$y�N��DY(��¾n�"-�%"O
ٓh�h��5������K�"O�p1�^�;x�Ya��$y� Uku"O�mA�?c�������1��(q"O�Q;e�*P5��h�ʉ(qu���"Op܊g�2'.�a $��}���qp"O�x�E���ݢg	�]I��I_!��W*H�K���XT�TC捏�T[!��.v�T�1!�u4H)1�^�XW!�D�;��`�E���A ��-NQ0!��պ~H�1)�ċb6��g�3o!�$��1��	��-�@�Bb@�e#!�V���E1�嘠d��¡ͳ�!�3?�ضE����4:7���wn!�[�Da�N���q�!el!�D��2���4�K>�|`Ʌ�3E!�D�#����&
A%�xB��7!�Ѥ1 μ����.K"̐ꄼ-%!�d�&�)��on�p`	�
��S/!򄔳D�����kJ)ziDO�#!�D� 6����4�4�#�49!�D�
E�\�S��VP`)b��!���JK蕱 K�Ekl�`�Q�!�DҔ"v�;�c�X�r���U6!�$�B2�l��BbE򂁎<5!�dӫ�0	0�X�_5D�a��9]!�O�2�D)��^�t*�	��٧'!���Ȣ���:�Y�LĚ@�!�ƮY��ua�J���!�kA-N�!�P�]´25�]���q;��M�1q!�T�#����F!�iY�$2R!�$Ĉ�Х�`�[6��)�d��>�!�d��|�@P�b׀P|��Xgn��|�!�$uHhyڱd'gs�I ���B�!���P���A�)Y��0@!�	԰ �w&J�z�)�ه6(!� �!@��я�;^���#�'P,!���'D5�=ipb[?E��o�?^�!��YI��.�6(���BhH�u<!� 7&t0�%LSz&4��3� �0=!�҂bd���տuo��5&ؿ�!�� �%jH:b�$;eVT(H�&"O�"�"�5��8Um��0�A�"O�Q� `I4^�lc���{	�p"OF���K�w�l@@+C�D���"On�ʡ�^#

h�A����E��Y�"O*P�хX�Qw�:$� N�M�"OX��)n��x5I"[34T� "Ov���	(֜�1�g�-(hE"Oް�5B��HJ�K5�
vx�2"O��;��ڧ{��4���#=��T"O<��G�ӿI�.e���Vh�M"�"O($��1k��r�W]M�e�!"O~\����8\c�ٹP1�H`�"O��yE��8)^�Zb�wBȐp�"O��Pj�3�X=3EB��01�q"O@P�舂C�b�pƠ3S���BP"Of����P�; ��4�4 [�"O�HЖ��I�j���  2b�̵�"Oֱ��B�,�p �D/�5s>�ܩ�"O2 ˛�$tDH�-��Lǔ-��"O;�/բ/&�Q��Ƞ����v"OZ	�%B� 6����fR!;�D�"O����i�?�p|�ǧ�Evj�0�"Oԩ�g�m���bf	=s
a�!"O�+�%J�	�\�32�mV�I�"O.z�b¨:�"�a6g�H��A"O��b�aY� ����س}C�x"�"OR}BR��0'k�L��D�Q-v��s"O�ԪB��$?���r�V����"O,��T����Q'`P�h�A7"Ov����%E�`�:A�@�qM�F*O<8z"	�hLP�N��s
�'����[�A�� u��T8p�K�'��XJS�ȁP�,5�$`H8!@~@�'|��PU��b~�]��җ�6�1
�'��Ke�ߟ�~��cIp{h�5�	�'C�!�Vo�q|�<;k�}b�H	�'��8�!Åq�$�#�4(	�'ߠ4�#˸bF
1�
f�X��'��,�3c@� �z,��	����'�.��Sn��Hx��"��mS�'`�|��K[�~ 0QG�0�tL��'���'�Ob�Y�S'ge�JK6D�`Q��:���Q��
b3��0�5D���@�T�1���Ґ��;X��+!�%D����_��8�`O*?B�����/D�`w˞�g�N$ɤjG$S)h�h�9D�X!��vQXd#�-�B	rF�x�<�����%[�m�����&�Ĺ����u�<Y�d�,C�v�i��A�d
$���k�<��ʋ{�������g|U����i�<Ѡ�54�����
L�ݛ�HKi�<q`ܹUT08j#`��	9H jF�b�<i��1Tp�F [;w(H@R�N�a�<icfz;�X�)޳Ub�8ڗNR_�<��lг#l>4�c��8Am�4Zrc_e�<y�C��;t���	5Wy�P���a�<	�D��XE�����31Jv�p�[�<�C��c�*4q�ɐ�*cƈ�� A�<�Ć�S(��t�M�t���m{�<��F��dvt5�Wh&�X�i��C|�<�5��A�����@�0Oؙ��w�<�[�!X񨘆|���ȳ�Op�<�VF���d��\MtH��/Gn�<� PH�-_�F,��P��>+,ҡ"O��А��%�6e{�ƚ)0B$�"O�Ai&$_�*�x�@�T<�� �"O��!��]0z�x�@�ǉ�l�����"O�$+DK43l�t��&X��f"O*d�a�P�v޺��G ��OOH���"O\��bD�%�l@/��y�Щ#a"O�<�6f�9<�R
�(�� �;"O�l�ޔ,T`s���$o�����"O�٩c0U���k&m���ha�"O8�	t�P��4��"���xE�7"O��`2�V���R��ҋ.���0"O�q{"LV0-IJ��"�C�`�Y@"O�<�'KMO!Lؙ��� eΌ��"O"=;F�'ȕ(�Ѻ&f�t�6"O�p�צ��0p����9OZ���"O��Pv�̪�@�+���	7�	�"O����h ^�XF�P!0��%�"O���f�_��]p�*�-�$�a"O��K�c��$��)"u�V�k�"O	i���3n-Pe�3G(;
T��"O
��5F�:� ڵ�V,w#P9h�"On��'�7�0v�!($bP"O.Q��Jf�&.$p�hG�P�uh!�$ϼ
[�)���Quިs� �6 D!�$A�<���Ƀʜt�����؉\F!�D��0�����esd}�s�ԙRk�B�a����5,@m�r)�"�JB�I,x�m g��$B�VM���0B�	lM&���� �(kԬ�V�M��C�	72n0���͎�Omj��ʗ��C䉤4���eDS '7`t��NI��B�ɂ ���ـ�d6��B�3Z��`H�d�54�D���¶$��C䉐*m�h���	�Ղ�B䉢!���(�?24��fJŋ0C�	$84�@��/�Z$�tIǉ_��B�6vnZA��#Q!f�Lt�n�%=��B�	� �K����(P"X�w��r%�B�	�'�xAڴ�?1��Q`�^�dI�B��
7�z�A�m�%9����B��wx�B�I�o�����;3�>��b]8��C�-�z%��� Qzv�Ҥ��8�bC�I0U��k�a�I�� �K���J��d�<���*��XZ"�6~��йUCV<��qyB�'*����ԗg���N�3#��	�'��iX�ռA�~���ʅ0�x3���I�6P]�D�1e�H�s�6���(Ol�>)1�J!D�ta��??0�8di�<�"L���4����W7b�ܤ��J�~~B�'`|���:6�`Hvn߼<�!�{��ɾ��}�!��4'@L9�@��:bC�ɜV��qp�xcR�
R�"<S�i7ў�2#DPZ�����L��*&Of�C�IM�9�#Ŏ�$�L�g��;V�����p<)�{Bd�u�"e����{�Hb�̉��'�.�GyJ|�g�)cX���5��?]N��Ks��b�<�Gh�C���b'UJ�j�\]�	T���O�`�B�h ���=���M��9�'�-q��R)e����rH�Kw����O�˓��S��O~�2�"�� ��
!̄{�����"OJu���=y �r��(x\�������O���O���գ 76`a'��9ް�!"O���E��(� �	ҲL8���1"O� �����#0��8 �ȃ�C2�@�$�'�b�>��Ȟ.V,��eI�p�L��R��I�<�p*��C��T &K T���QP�<)'�ʳj�D ���=�ʰЀ��M�<Y��Ơd�� y�S���5�`��J}"�'0�q2���[1�:3k��o����	�'s��xQ�_��j�q��G�.�#�'W�dq%�V�=�<��՟y�a�'��(`�ϧL>�p�O�:�\�Í�9ODI)���(F���I���?��<�0�=�S��yB"\�Ɛ��a	�WK[�E��;�0?Qq���`g@3A��J ժr�0UI�jh�8�'��$�P̧��sӸ�;���x�Y�R/C�d1��'qO�Lj�o�4VV|��`�Oz���!"O�Ic��"O��J��� *t��V"O��Fƙ�1Ħ	�MI�J��p"Oā�p
@V��l���S*K���z�d>|O�A�DmH*�vP�	6 }:��"O<��
��h$Pj��4a�I2�"O�	�sK1w�,i���n�5���G�<�RL@�0N��sv[��lv��B�<��� �C�i��o�O�Z�v��B�<auŒ=mG2�P���^R`y��|�<��!Z����e!�-*Ue�s�<�񈂰 �X��Ka��c�B��d4}�!X�mC��w"�z2f\�t+��y����Xm��;bKG�������0�HO*�=�O_�q�E���*l!C���>6��4�?�����s��5╍�`-4h�Q/�$o6m�<9J>�|���~r�%����U;�J	z�L��y�	��h�E8�O�^Pƹ��ݸ�~��'lTDyq��l����������A��'� uo�1�i{V�A>?!~�)�Ox�=E��C�LD@�����X��P��Ĵ�yB�\����Sl�T��H���yB̜0���8����w^�%�@����=ړS�O��Ó�ï��$;ǍO�EB�yr"O 5�MJ�����lA�k�^���>��a��d� 21d�E*u��>�p���I^�'�4���������#�M./X6�1�'� *�� ����/��u�Ó�hO(y���بi��V �8���"O���Y�1f��c�c���AP�$�p=ѱ��1�hm:��/�T*���s�<��N�(�Pa��Ν57Ȁ��� W-y�#=E��� �����[�	��-��,�8؇���?����{���RoN�w�܁�Q!�70l�O��)�3?�����m�5`B�ya�I�&Jv�<Y6g�!P���A�H
[eRa�F��t�<᠀'�ѫ����gv*���A�l�<A�O�J#\	�wK�`'�H�I]�<����ݎ�yv��:RF6�{���<1��m���@ J��.N3K�!�dVsr�b��̥"�����+c摞�F{��t�0D.�0D\�� ��%�n5��"O�L:uMP*�^��R&A\C�X�"O��r���5���FK�f_�����	o����ca�k@,a�N��e(U�SEH��C�/4���4�d�Hr��*l����+lO`�\KSe DH�+UlL�@�@x��+D��2[8GE.!�wNƄH�v�9l�h�',ў�%��.3�C��ٛ~�0(��.7r!�D2(Vԋ0b�[Z�ѫ�̞x���33�)��P9�B�>v���86�:�4�x�L0D�� ��;��z��
�O��H����l�~���&h�:��'L�&x���A./n	qO�"<��{⃌!��q*�	(a[�BƎ���yҦ��V���!���6Zv��T?�y��'�T����!$��|�5&)N$d��'BVl*�e��b���ZE���L�J���'���qS���wkY�N?LR�@����!��'R��5��!�Rt��_�m���&�D��	�|�<�۲D3辜����C�ɠW��8�JbT%si޼\A(B䉁FX�s�Q�1�h<�q��3��B�=G@�}"E��d�b��B��qu�B�	�y���z�a�,e�D|����_6C�I�(8(�����U��JV" 
��C��:�4��W╈4���Z%\�8�C�Ƀ2�$T��	)�<���n lB�ɹmp�I���?C�'�+s�hB�I�d�@�Ì��#<�M��c�^�\B�	`�0YS���(&Q�9��TD"B�K���jߒm���M��a$�C�I�����T�� w�����v�C�	%�DA�掏}"������3��C��=�I��; �T�ힵs�O�=�~�`$�Y��d2���
�8�S�a�t�<1UÊ�pˊ��PC���h3��u�<���M]ܐ���NE�d����w�<��'��"�R�a��^p�o�<)EP\n���$X?�%j�il�<�3����|�t�/6$u�֥�k�<i��l����V��|xf�A%��g�<!E��hC�HBcK�'�j٪"Ta�<a�px�Aλc�\�2�Ȗ(	_��Vx����nA�/�tM:U_�/��P��2O���CrJD�!`+ d̈́�M�8�a!�у��Lه��l�؄ȓfB�hJp��\&��IR�.nq��=�$(0 �mC�����U92M��ȓ �Y��Z=*�&y��n,,�x]�ȓB8y�ŌI�Y;�I���+MDP��luB� R��O��yʅa)T�|̈́ȓT���!D�@�` ��N���*�
�HdAIIO�x�!�D"K�݇�z �y��8�<���� ~�Ň�y�>}��h�> HȸRa�P x{��ȓ1�(��S�m3���$%;n�Ԭ��$z�`@�ƍ�Z�L��ڱ88�E�ȓ{u�LٖA�54�E�5M¬/Tl�ȓ:��薢� .�x���B*'lQ�ȓ�B8A1��v�\ix��|�.a��@��U@�k�z�����Q������	"f���kOI��q�ȓ �����G�$/ς%{'���&*ل�d����Q�Хz��cF��ȓ.4�	�k� ʒ�"�i��|�$D�� $������Q��Ύ;l9p�ȓM���'�Y�pn=�$� :���ȓ�q@&kD�wh�P�uHț��ԆȓYg�iQM���B��փ��|y±�ȓ3"���zJ��q�H#�T�ȓ/�]��ힰ1�����_9^��ȓk4&A�T@ڻ!Ԯ�f�9@�`P��<�Y9�H'&�((����~��IH0�śa-˚pѼ��WfQJ(���ˤ�B䉊n�^�k!�kH�e١�nB�)� �`@B�$J�E��m�+.gZ�)�"O�� y
�	1k�Q@���"On�XU���(E�3�Yj=lY�'z(25���Y�P�� ��:�l�'k%�pX�pt@��!�|��dQ�'Y�	/T��~� @'ޙs��Z�'�f�����	y�)Z ���q#|�#�'�LX Lj��sWG%XƵ�
�'�h�a��?~���%ي�<
�'��H"aȜZdL@Ru�L.��=
�'>���`H�u�����	�'�@��ۖ- �����%	��]��'$.4p��jb��u{� ���'3XR�L��I�l�H���3 ڪek	�';`����ʂ5����ǁ>h\^���'ƌ99Q�ܺ�pD�@��\�5�}�<���ЁH~H�{Ѓѭe��Pѫ�c�<���.%v�� �٩FAI0��Y�<� c��I��Dđ<
�$0��T�<qfÍ,z��}pqk	$$�5 ��Y�<�BJ	k�`�ˈ9]4h�b�<�A无��hT�2Wd ��\A�<�ǇD��ͻ��	�s�h$�uT|�<I�$ݒt'��+�"Z�)�|efq�<��'�0�A�ɜ"IဝCF*�n�<1f��#�JŁ5�#����Bd�<��H�Drpı��&oD풕H�]�<��_)eV��R�ЧIp@Bfh�]�<ن�!N�r�3�D�i��aAT�<���ұ>��h�Iϴ��8��	�j�<)a�52�|Z�FW5HD&yXV�c�<)�%^�IR���SLޯV��;S�Z�<A/̺{�숛���\���'�W�<������T��Ygw��k1�R8��q��E�K�!�A	\�^$����+O��Ӗ��9��<�5�'�~�B�D�8m�h��A	�S�'P���@����P,Pbc歸�R,L<�.� %���Hk���9������P�0�{�� >���$���?�~�wgS:6]��#�ɴ*<���%W��bD��>2u���$l�:����/Dab��
�r��]�+S ���J�0v��#�n�>���j���q�߱/���CGIߊTt��1��*�	�Z/|RYс�R�Oq�ІɣzL�i��_�VＭ8S�nz�8�g��F��k�[�0s��ƧI"y B�A�n�0U貵�p�B\�����H�Ɯ� �mE$$u�]TԀa,O���C�~�� �d>A�g�	HPpa��"��R�ыA���L��k&,'��0�E����{��A��A�(OԊ�@ �5oh��D��<�M ��-Y�b�f�H�\��4�D��%�A+2ar�ڔ�T�;�iPCH�/]G��\�<8�mӋZ����׃un�ċ�Aʂ��@A���6E.��H0�	$�ʀO������
L������D*�$����ST��T(�
:�A���J�������yg�0�d�&��.�!`RK��ē-^�q{@��*z~]�S ��c��:VE���M�V�R�h�:T<��K`�%[0l�TmŨV��ceC�8Lq�1E�H�L�:E(��W4�Ș��;.dbp���\�V�>D�$�Uܙ���FI���c��%O*�ʧ*���ԥ�&�p�#Ct�R|:H�&Ԓ��f�& �i��&5]�\;��ȯi:�A��P�HLj��Hu��Hn�9R� �d�~�  ��/a�|��S�ۑ'oT#��F�Ǽ�2Ə��:��)!R���g�r��Lʮd�l����Z�c�Q�OV�lS�bH,@��+7�ƼSE
a��e�g)�⟄���E�]�La�.�z�� �P�ӌ#fJ�K��V�Wc4 ��+��m�"�p��8`q~�#�&�"_��IV��镎T�	�b�"uF<M0��C�(])�1�%FGZ��rk&�dˠH���Z�E�s��� "���X>%[���R�̤��,�"@�N-HrI�V4�YE��;��%rd.U%�R��㐟V�ڐ� L]�D�@ �	�<R<�aůC(Q��2p��4<c��u&�S%.�r��/pZl����]fX�x�2��*058i葓�fD�S+6�R5�дE	&)	]�9���k�&��b�
q+��32������uirIk��ѶA*9�?�v�<�����Z �!Dg
Z�NQ�c�
�^�6M�U�Q�Dv�ȉ��Ֆ<���E��]�i��˟]�JY�3`ʌP���ȍ����M%�\�0qe[�Bx�԰�r���Ź�N����b4Z8�;�� rn�l椠��2j�a�g���#�@���]4�;qF��}�rΊ�h����J�6�pȶeR�v�k[�B[�|e�>�Fr��x��*�C,H��	��n�tSw�O���!��E��us��� R�)��L0��4�ڵ3��Zb���?�㜝@��Q#M��$X�96��M3��ɜ`�l��Do�.�����پJ��i�,V�H�����L�����z���?e�r�Z�f�a�<�g�1Z�hI�l�s\�ժ�4V>��Xs閴�?9W�A�[�Hk�#�4�lMGzB�ZNZbcԂ�F���C ՠQ#�p�4%�3C'|%����	�e�J� ����dy�r�*Ś-���b� �h���(T�Sky}6��0CI6z��l!�b5�-^�����7��x�Ai��UI���
k �Jʬ=N�X� Ɣ���@ ��  ����cD^Sz|!	� h	2��ʬ<B�-8�O4���P�Q�����1��Y���x�oFf�!����'b0�0ڗ
W�(Q$&�3j�8|2�C��'pH-�xL����4պ(г"��>�����6/u`#M�?/T��'7��X�h�Z�I-x�� CįjN�� �,�y<`�*0 ��	5T��f�QͰ1��#�r���lE��XE��|9n�"p@ �����5KR<4D��7���0�Ш��~"�P�
Z�� ���y"��u'���g
�7�Hꠤ�f�
)J�\.(|�&ǒO�4*4,�#@�@��ue�[:b���	 Dπj�NƟs�����Цs"]��`�|�t�i�߼u}� �	I�-؄#�4q�� i̼\e��)��ʙv�ث�c�:�����	3���)��O�n0���@	�]b��Qc��w���V������+ک�e+�a����C�;���A �j�>P���C���s�P��)�v��Ì��jV�)8�X�F�X�Y������Y�l�rA�R#�hٖ��5����bJW*=�P�N?���!d�v�p��ǆ��ut�� ?�X4�֍SCpx�pIAc�<�C�Ţa�d�@5�F��]@���=�J@�P�1v���6�8��A�)G'���,�?ѵ�-nڢT�I~�=��-�-�7�^�(h��h	~K`�:�{L��Վ�5;�Z��'��,��硅�[�8t��~Md��G+,8�xe�Ą���DÓB��e�Wj�"lJr�,ғ
g�b���.#���W����$�rlJ2X�D���$u6�r���+ǼQS��<�Qw�® ��<˂LJ�1Y�X��NQ�pi�iA���䏽SZP��əc�qOB����3U .|cr�-!w��ʢb�>n@�0ke�B�%�n�q�n�	8���a"��MΠ)�
����#@K�+&�D,��_�h�)��> ���1B|��<q$����N ѣuƓ�e���S�#}�U�$ѼXd:�kV�^>t/�9�����J��ŦR:`���G����$S�&�<b#Z+���-�Z��J�2�~�X�?�|IȌ�L>A�I�4�"*Ri ��+n� �f7͛�EG,��Σyg��i�R�h:�QԄS�(��&�C;<ͪ��ڃ
����58��5%TZ�%� ��.-�,X����\iw ��jK�%�,x#���a�t�y��G&?�q�gL�E� c*�~p:q��$r�\`4��0b�r�a��&0�Ecb�L����I�K�z�ApmA�6�и��
-�'lıYg��P����P�4���f��wc�L����	�I��σ��p�ǧ۩aҴ���L�"TA ��~{��J��1~<�]�O�x+%���(L6qۼ`��,qӮ���>h��TK�J�<'��R��.2V���ƨ�s޶t��⟮tپ�BӅ�n����#@H`� �ĥy��]r�I<Fzp2�|R��Mtb?�!':�Ye���`��t)V��%W�kD5��� !T������	B�Jp��T=��
r�Y�o�v�h��i@- �e��[�ha��K�{w@5(��U S�%���D
�����pŗ$U����b�)�5�L �r�.A�`�_�%j�y$�S�H��;JӇ
o��I��V�E�0!��Λ<v�"U�P&��&d�%�,��.��V�Dq�n�@dP��0�\6
�W�Bi��ӃClD��� ]嶔��"�8=d��>D���:+�p��G���`� �pkw� Yu����
4s	��A�BN���s���v�Z��#֨"%�`H�1���m]2U�<f��BR���Z���R�_�
�[F�� !�zH���8h\ܰ��]m̉E˖C
02�[
] �(Ђ1"���
Eg�PX�/�#O ��қo�@�1����E�"���0=x4����D�c�tdo�%B-�S�n�@L�áG:r"���R��"��<"�7�,xU�C�F8v*�����R�&��q"V�>lȰX�K9 P�CS��lA�An_�Ϛi���>P<5@1����-�0�J8 T��D8�zT�p��"'�%F(�?O�Y��KG�=�:�� f��ٳ$�Z�;�h|���Ϡ$�-
Fh�M�y�3�p�|�;ƅ���h8��T���Y�놼fV�i��3�p=�!$*+#�mKc��I�e�ڢH2��B"��4�J��P��e���ҫ/*�As#)�J�ma��@k�E�'���RGo�-"nph�f N�ea|�#K� yf �0�H�������Q���c(K�{���Б�^;v�8|5��?����7�O��{˃R���ȋ*x���ȱ�~�E2�˗�Ms����v�̘V@.� ��Ī֬,�����&H�]��%�̀J�x�J�:�kd�~����HP"N���1G5K�;�Z�(�HI�/���c}�!DH�(l�!7
�
�\�'q���'M
c#2�"C@�u��Q���?}Čx��C/ 5��n��&s��
b'8�Z��A�>��=�p��.M_����%?s2`�#/���ꤥ�?9�aÆ;����!@���d��W��j�-Ȉ_T���RM�3�nK�1И� p%?C��He���U��J��h�u1��Bo;�]�ԋ�2R���֩K��f:T�Y�L��<5H��k���=��C��!�I�,)�0�h��Pd�i�,&Bn�,�iB�ZX�&���HZ��0(�.�0�� Pe�Y�̌'@i�,�"	���Ezt%L(�h���L����Fx"C��[*&}�4��*X<ͪ�eSW1���I/��3,�77��p�
C>�nEK���;��rs
	6�.�C`MV�F$��S�O�54��HJB��tu+�b��=�N����*!��;Ң�u	`��P�ĜC�B��'* �yǀ
���� ���BP�wf�����G	h8ua�m��dQ���7�����`�#Q,���ʗ7\�@I��rB����h��x�=�Vh�?� ��B=����!��l�"-�l�
<���ٮi���;�2����½���� n�6	��e)%���ꗯPk`ҥ��]��
�{/�����C�"U
A�;�B�*A:1�Z�b 2퀢�0ؓ�J1{��=H4�W�'�8��S9��4�h]E�zB-� �$-l�e��k�����M[���1J�cM�t� "OB�v޲�a0iZc�	�wݺ�I`��F9E���i��`�2~}�%*W�Tu%,�d��Y׆)��G}��Wj:Q"�l-iǐ���.к|���C� ��<���L�=;qT遡Xz�la)��N A���ٸ��֖�\�'=4�1o�)��(��l�� �R#�x��L�Fc24G��@��-U*yӇ
�7o5bD�~u���Ӵ{��P�&��6@��`AW�(_<��ݶ}|�%
2�̉)D�D�<���W�$���/	 l���>AK��qez����b�h��*�^=�~�B���"�"�3���+7���s�V��Dh�*97 .��z���=Q!�$]�ʥS��_�88�����?d�E�����Ã�	e��a� e~�'�4�>��gBBMIܘhKitq��dBZͤ�k7�AM��P�va7lO�8��� �i�a�6��+�� 9��5�Ƣ��<A����3b��l30p����{8d9�Gֿ%�R �F���G���0e�����#�ΎE����$)i}�0��C}fZt� L����n��y��ɻAgc��9�Ɖ�/�0��狞?x|&�ݒn�����B:z��ٓ1g��f���f	�����Q��a��m�u�@�QI3?�Ro[�;���r��$X�J'��!(�͹#�ϟ+: q�R�� 0DZC?�8�C�2r	�q�H�M��-bJ���X:��2��HO�I�6ᖾ`V�J3m�.&��T��7h~�CƥQ(0��
"���Aa�U�f�< kH쟈��-�<,�,�C�-%�����"_���
 >�"��r�'vD@9T���1� �T����Y�O�4Y�̑�8��	`d8�c�DE�G����4@�.�>�1ƦR�#FB<�r�+\��ԈG{�)�3O\�r�H�&C1������8��U��A��j#|�	��@����RLN:�0T�&g�vx/C;T��I��Ӈi�P̰���R� <��EXw>2u��4SA(��c�)flΑ���/A�0��'�ވ�-Y��Q`��H�qƔ��L;T�H����ڇ��6��Yx�K��šU�ze�`A��l�2�eG� B@("5*�$ZԨ�,F-]r�=��E�� ��E���I�q1�qs�)Z<S��KBk�M��3���5��]�c��>!���?r5�Ek۴~�H��B�T�����ӿv5��c蓘z*�]z�h��*���
w�RU�f�Y6P�eAŤ�o��a!�%l�q[����WH�)�v�L�\���7R�QY�do�� Q�aI'j�QQǪݬ~|hx��,%o�<�uM3Od��#K�a�<10#Q�i���K��51n D9�0�4�IO<L)�Yk�f`��@#ƟGC6ᙇiE�ij�(�҄�3h�a�O��d	J ԩ�G���:�, �����T��Bv�A8�oT_�D� � �V��)$'��M����
��ϘQߦ`ԇW*)]���%�Mj[����
�EK<S#�ܪ�	�2z`���T>6ܫSg�~����[�@��c��9q̷�M�0~d�O�ݙSNa��� ���VN[�L�b��58�f׼oX�h�'WJ]٣'Gr29c��ݬJD 4��N�M�!'e����ɉ�b�>�͓�2|Z.O���P�ʟ?<2$S��	��h�9TG[���D�'�l�!dm��Z����k�0$:m�#@�hOr<�!���T��Ҵ:H��3c�iw��3�Ɏf0��?���ɶd�:e�0aF�%�r̓R�IV���ʡ&Z.�*MX*H�4d���ɵ��'8�(���)��1צƶ{W6��'�����,[؞Lc$���F:D�:c�������l�`]��H�Pj�����6?���E�ܴ��}��
�,[y^� U�P�JL^���[��j�O2������?!��	�O0,�AJ������a�c���$ô]h��Ρ>Vz���AUa}�(]��L�vkC�X�h]ےIÿ2�*h��B��5���O�4,��~2)�J%���#H�q�&SW���HOR͸��K'Y�m��ă�_��O��wdX�lO����ʓH��A	�'�<���G	�Qm<��u�3J���.|� U�+[�N%ӗd��"~򲠍:W�h�i7�֚WӲt ����y"�B�t������\-[�4:WLƱ`.��\�bͺ@�a7����(O�Ѡ�QSJ���IӪ�i�'�츣�-	����0�2kU"�+�=�@!Q�����2�
�rR�y��K$%�pLk4-���O�<Q�u������O�� ��HrL�*@`�.9�й��'3��اI����ׯ�3��'p�N�S�O�,@��8�J�J�-�5����
�'&Ĝ2�� ��5�5�-�@��'��ŋ7+\D��
�`�-pX��'�
8���=�TI�5�^���1��'�P�� n��@"Q�1�S�g�<�Rk��7��P5�'
��ɆN^�<�T�É{�)���w����'�w�<�s$O�Rd�\[GI� oh�3�m�<ɐ�BI�2� Vm�.^��C�$Ww�<9q��
1l���J�$�E�V��q�<��.Q8���z�d�U.�{�<a� C�	���'��-SB�Mt�<YAN>�0sv��)n���:��r�<1�`�,+������m�<Yū�9y�9R��Ʉ<�F���j�<���SI3 ��f�0��2�l�<��o�@��)�rfTgW��k�j�T�<��]$k�䙇Dɒm���SE��{�<�w�#}@r
�΂�xv����v�<�r�@����d �=o�A{�f�q�<�g�×3�yC�jM �	�&�Fi�<)�n��D ��k�?�5�0/�d�<�僊
@T�􃙲![�m �Hb�<� ����2x����� ��aȕ"Ox��U G4:,:��/U�(s��SC"O���g�ʉVŎ���@����"O�@@3H\�=Y&i�!��.<�v4[�"O0��У�@b6͘�%�Uy��"O��p����@4�Ά~�M��"Od`�w�ST���W�D�laq��"OrAIU1��
��]S"OdAz�@ѱ]�hTq)�3]� ZD"O|��TdoS��h�狿D�5@�"O� ���)�>E� &��ǈq�"O�]��ՃX��Hr���<���A"O���� L����S�8r�
S"On�1r-Χ<�I���"rE���"O>e�$b��\�2����>w���ID"O
M8�LZ�/�4z��GJ�0h��"O0�  FӟA ����B\��U��"OFeC�]DY����'24���&"O��(&f� 5�1E�%/l��"O$uH�O@[�v �eN��`E�p"O�Ԫ��7~��8�"�
4���8�"Oh��a-N�.�� a��<RϠhS"O��2##�,8ءc���T ��"O`}��#��C��j�"ŻAx�$"O6��!gʝY��rg�P�(��)"Or$+���*)P&�A���]b�"O�A��@�>��f��k���0"O����h�O"~$�'�'��p*"O���H�<^��8rG�G����r"OD,�(I�te�Q��� ��]�"O��a"	1o���y�ɢD���"O����l�(��k�
L�B�BU"O�YBdÒ�4 Nl�"ʊ�4��y"O��Ӡ,E&xc`)+����"O� ���s��$�2hG�5�����"O����P�\�4 2��%v!�E"O�]薆�Z��C���T2b�1"O.(����yoI��S7B���Q�'�
a�g	�$}���!`Wx}�D�
�O֩Q')�(�l���J&�c�dݚu�v�"�I�{5�Y!#k����a�s�
%R"�T�d
�$q�l@�b&�*.�Ч��K�R��n��)��WF MaS���&X>q��=F"�ͽ?Z`�'t$��P�թP�Z��s
G�$�X�t�B�V�*�(�<<�z�h��ձJq.�D�R�P����%�X��wϠ����P��RT���ߞ��T
�{�/Orv,	b&�_L�O��Ps�([�VnY�r��nEZ(����4���h�&(�~��F�?��Xk���UiA�2�mBT0���oӈ�4i[�XT�B�]����(X�C����e�<)�C�b���E��@��F��(�D�0n�&4��kׯG |9s� 6T�9�֬�f�:� 22>  å�m�.�<іG�4QX�R�%9Eu2�MO�{��hseU�v��A�cQ�1��@�g��2PF�:�KY�<@irΤr��(S��.��Pg�4�P���,K,j�@Q�Ëq2�Gx�AN�qn��`�嘗:^�n�'�t�bE/g��I3�ߞd`\zрK4)�Bd�҆X1���a��G��\��.Ć*k���)ߟdl�� ����e3|�6l�@��n�XO>e�F���i�\��P���4��"|Z���F�c�
s5�X��S��dX���10�0g��eL49������R�q�A�v=��0v���D��)Q��ؤ��4�����y뚬J��N��D�AK�>Ytf�/�2e[S�G�,�~��^:&�^�P��`�"�Ez.��ر�E@PK�/']F��7�C�<ޚ-������O6��
 !-#n�*%�V�B��d�1o"�8��B�,W|�!������Jj �,$b�U�D��@�����kLF4f��5xf�̀O^Ekw�#�rp�J܁c�� �RL����&N,N
��F�U� v��q�Ŷ e��r�9r�is�'�"1BLC�&�$�4��'j��MI�x1�x�t.\2CЊԑBၭd�<X��8!g� r�AW���qA�D��-�>���\�H��� _n��'��Q�s��}�t=ʄl�o��)�$��?�R�a�m2�CC7G��0ª?��Kv�Ф`3&\#�� �"�y�#�aNl2�BLd���LL�3��}Y���$G(�d�h��8��@z�:�Ld*��`���Ó�3��My�f;|a.�#lɺv<��T�y�v��'FR�:ņ�+��¿HZ���o9xf"��?1G�M�t�qd��6�@���&����MPTbPCϧW��e�`ςM�n4����BJO�U��Qʱ �J�j��b��=պy��A�1���#?,�~������'|�e�����ob=P�{S��R�kʷQ����>:BAi���%��Hc�m�JoTeгC�SB��)B��Q�����':HU!ě ��d󠥗5]�Ԉ�4B�JD @ ��$Xy1� � ��|����ҙ7��a��#I�?���.� ��z�_�|����3Jb�8�G��S(�q��P�/�N5�ɓ x��*��޷y��颎��Ka�4�7O2��0e���a�:~YP9�Ƭ³)�rF��"�����T�o���Ƅ��hG�B��YQUd1���:����ؑ��ɤ,�(h����s�ܵ�IY�D�2��o:>y+��=�|�V4RT�V�~u <����;f �Vc�A�~����"��1F���Q��%�������z0+�_/]��T��m'el����R�A.Xi���d��#<�lS�1��e�D�Zv��U�ۨa�vi'�[WM��24)NHe��
��V�t��1a�$�@����FY*e�z}	�[UJ��"�	���$ОH�xT:��	I�"���F/�'��Uj�L=�Z�c)S�OM zQ�[%�����!>�6�b@��P�(tH$E�?$ ��I�� �*`�,Å@Y��kR��0�l���O,��M���S>�H3p��e{J��	�#^�`�c˵�&�6�uueQ���W2T��r��N��q���!n�PE��/l `��Ӡz\��CDߤ`
���E÷Z�6�#�.k�G�l�g�bS��y�Еjn4�)�
;q�v�2&eI�gU��40�Nu
����[ϲ��"� )��t@3�եu� ��e�
�8�X���x��m����Q?����K -�� �ǈY��hOB`X���4� �*��B^>��#j��f�K��y�`@��gʢ(���I�W2D��9�'�Op� ���_�S?bt�y�|6+�O:��&E��sCK��T�V��M;�ɱT��e�V0f�5;ԏ��5#V	s�o�5h60sFk@,i�5��
+?~�B��R2Q��҆ЁM�����֫B>SE+@-�?�D
͌);z�����u����1g$_s]�A��
�>Z�,бQ�Jw@��!���4k�
г���q�d�uV�e��
��^�|���/F=F�� �T�	30���Tj_�l�{D�'7L���N��ϸ'j�E�thM=!�D�q����遄�H����q��t�yA��Oa�m�t��?*�p���Ǚ��偔&�O�����0�d�IA_���@��Y>;*(#!�F��HOΠ���Ip~"p�z�ZF�	T�*`X��� q8����Y�b�R�(EmCR� �`���y�R&�ĊT�$dx� 
s.��	!o��I:� ؕ,��S-��\~nU�=��+�<��US��˼D���k�Ģ��4e�0�0G��v h�VL�+�  ���p,NmXPL���.�hY�r.L��C4h��У~:��_�`�X5�a�D�L��E�0A*�[�0{ftTo��\({T���f�L��A�T9�`%0A/�����G2E�}J&A���B� �4r� c�� %F֓H�c>�OX���Ğ!>�j�m��K7hq��V��M;��E�]-���򉇭N�������="5N\�u���,�v����X-_U��V���PM�jumP.f�:�B��N�b��0��Y W�#<�*!_��UJ�d�\!��*\-82x,9�a
<Z�����Đ�l���ڃ#��#���5JM1���90~(�!J�\�����d�>���@��8��#�pȸp�DMl�	O��1q&�]��<!�HښC?tp�4j����-�5
��!b6a�>H!�)(I�x�@Q�$�|+�NÕB���J�D��+�4�%>٩v%� $*�U�N�8}@��o[�%(���[��p1aSf�Չ&���!"�5.N�.IHVQ��5�C�o�1� #��=B �Ő�
�8��=�r�E�����G�
��G!P0,�)�%X)B~t}pċ��{����DQ��"���A������:<�aDe٫FvziP���m��`c!	޴�<X!��#���F}2N�6��A���TW����^�h��L�g�F�?dZ\XÀ9D�$ȑ��H$|Tb ��D7H�[��K?�`����=gX�]���'�(�0è���۱��3;7�	��6�r���:��룃�8�8=�ୂ+������X$��'I�<�@gy��Y�R��X@,��%Cp����w��,��1�דN��=�񥙁[�\�WGW�jA�$�1V�9��k��{zn��W�W�N��-Ӂ�^�`��{jy��H�38���+CcM7"~�I
��  bT��k�p�!��+�B��V�U92Jx��Ch`�غ�
�lJ�S#`��@�<��v�N,�\��� ;6XXAT��nm����ԭmP���2F* S��?hx�� �	;�L��6A&ca��;`h�����^Ӽ*F�F)y��M�󧋐f��P�K�`�v��w�ٴ=y�,��Γ	�8j&.��y��AӋ{�
S2>6�a�UeǍ6�P��_��45��\$Y_b�(�AN�w�I@ઓ3:?�I��e4�P���$	�s��{��hiw��$����&jX�r:�e뷫�s^zc"*�o��Lq�TsG�J:O�a����x��YY�螨t�����h'J�<�[�&��:ׯ�;M�q���!x��AaZcے��i�?
ͼ���q�%9�Oxm�t�	�*Ĭi���7K�mI����[����99�e��ޖg�~��1���%�\��Xb/�2m����%�9.��فp{ݭ�g���  x�hҰx� �Y� '�4(��OK�T
H)@���`��IZ��W����#�$Y�dB��j5HH�a���S<�X���ʤ2�H�ƃ�&�*�O$��e�H��M;��@/�h��1���%IՙaF��"Ȱ��,^t�D���?9ҧ��.�n�����|�A��	 t�8�kѵ'$��
&N�8��Q#�u��B�{��p�t�'4��hAK��-0%Ex2�ѷW{�q��VԲsMՑ"��gY�3(���� .?�^9"���Tq�MhS3RȲc��!�ykE�ցs�܀���)�rK�C��I�ja爌
���R@�1������.\V�C�B�@Ͼ����
�A���A7��28B*��K�~�4rd�ܞs:�cD�A̸����!B���yG��29A.@#��i
"lꂫ�F��RL2�uS�Q��`�)� `��������2���YG�d
H]��]zjT��q뚀H�`�AN(�� W�D���Q'��	f	NI9$A[`%
�m�w@�S��`L]B�I��I+ �s@�3��Y���'P�������O���"��T����q����AQVј�M�)��9���P!2kZ�9dEU�ݐ!�I�Z	�F�G\@��P�Y,��㞐a�4¢��d`�.$I��Y����8V���_jI���XAD���ہe�@m"%���5DD	ou �j� �1�ŭ9�� #�"׊D�
���gxf	�!IN0/v�@�y2	�0*z�x�j@ r�f�o�3tO>(�P�̧`�4�R	W�r�j!{w��
M�Lb6/�.t�h�(�OW1qE�FA	�K��m�U��|��a"�ڼ�K�=KrPX�Ga��q�Y12�|R!H�s�Mb,�+��s�8X�4�O�Z�Tk�LV`�i(�FJ�Jr�(�e���`I�0��`n�p��O!^�d��k�Mh6FK�Nz�Rqڂ�(x�(�<3$`3���(X��B ��� �>Y�U�'����Gd6�b�C�?z���.|�c�zkt��7��3{���r�|?,�7f�|9t�g�^�&h��# �|fn�ه� n%�Q :D@m�m(u،��ş���V�Z&T�%c���/ <8�	*n5�Q:厛0q����`�Z�`��,3˦�TI��+��aX��s�X�z3�.B�$X��(݇f�N�D{�?
��,h���.fEnq#0�yt���  @&p�2�d7 �<��gL������i	�U����zB��A�M�(_>�S`
˼w�J��nՌ�̈���C؞��Ac�y�)Y!J%d���!-�x��O�����AQ�Րo�  (B���ؐ/�tdc�\���7C#��x� a�e�"���C�N�0�dS�� #���5�l�����vӂ�B�j�<*�<���/B�#̔�*�Y�r�����O�9N�.��X+t֎�z���=(�2��t�/%ǀ�RߴT!�wK�RP�yࢬA�a�8|�'����@e�W�K��P��N
�VV�Y�"�@+b�2d̓ ���Ʈl�pU%�% �\8�/�y1xܪ��S]�mj����<�7��~U��KK�s\��R�y2�MI��V'O��,jW^+/�R�7㛕�tI�'�K�ʟp��B-D�<��(�"�xm���T��y+��O��0b�'��ʎ�ʨ �+զx�^��$�F12��� ���ɔD�̰�#ø0/��i^�W%(]��M�.7$̪�8�V���=eR0�`�-O���ƪLj�"�q3��@ih��U�S�1�:a�B¦�kP$�<�c�pӠTx��Y7G/l1ʱ�_&zi<j����#�]#T�!N�m��4T#౛�
C/��,�+�(5����'\j1aFCW�We�uC�D�t�Pu���אc1~p枵s�N6Ծ.��Q � 8m�D{�G�k4D�Ӑ����F����l��ƣ�?*��=�b#' o�T��K%����@�Ɋ-;DYB���%��ey����s�����U�!m��ɗ&����ش]x��4��f��m�(7KD�<�5�H:
T�[�}��{R��f�6���N��R���C�;;�<�Hý$]ZEH�c�l���oh�閡�%tP��
VH��Z���f�ǘkBt���k~d�*�)�98V��PO@U�X�c˕K���!��x�@!�!_zK�yz5��+kHXjq�F(�0�G^�}sU!M	H/�٘� E��T*S�S܀��2�R�	��h*�#u��0E�ֹZYv�'����w���B�N�pxS���?��nV���ḭ3x!�思�q<X��a����VF.'������*11� ��3��	� D�no�	{�e
7�:����!D�m�v���Z��hc��� �����5���ۦ���Q * V��p���z���xF����J@<Q�o6*�0�*ќLKv��ӯВ="m%A^5��i�,uz�7���<�4+���>'I�� �����A�.M 9:��'��y��/N5"Ů\&� p�NU�o��(�c���8<X@��̤m�@�����Oh�ӓ>�w-Q�$}J� ���3�������%>DA��oQ?˦	�=�h�dт�I6FG�sv���B�� ��OZp�2�W�5̆ݪ` ?B�j)O�4V�¡��=���M[�:A�- �k�����hc	x���,W�4����6LKh`s�%��������<�0'd�:�xP�0�<D�\��g#1\q�W�1}� �JK��,}�Uz-�5�G��A�
�g�'}ʝ� a��	Sd��ccV�`}�d��`��`�$ᎻU`��s-�%xEj��f��*]��p�O׾9јP��j�(�*1�\�u�� 0`�
rj�GzB�4q|�H�>}v��~�q�E
�>	eA�-8�\g#	z�<���M�pP$�qJN���MX�I؟lG��#��4hp��d���S��5��̙�m)��	���s$!�ȓ9M�����mf��Zq�=E�D����O�`+C$V��1�fj�|Fy���o�z<y`�BȀ] DL���0?)���$la��..����EY�[C��҉Q0�N��
�KT�`�M0m�ɉ��64�E}�� e܈��\�'Y=��p%�$�=rD�V�JK�ȓiU��i�	7�B}b�U S��'%�\թM@�S�Ogv	��mY'e��+t��.r"@��'VM����0y�� �3؋G���'�:���W��0Xh�N'�*\R�'p ��Ⱦv�j� �N�s�z,�'o�呔��M����iҮz�杨�'����C
��FC���7dV>���'�N�R�N��TA���uj׌O�����'�^`��hp��� a;F�X�C�'B�A�X�[�2�P��'26���'�y5e��a(� �A�~U���'�f�!Ü�a�ibmH�k�& ��'ɶAY��ف^� ��ǒg��s�'�\�k�*�'�SQgQ*Xخ!��'�QCTL�4]��]2\�����'ό��A�'���2�J4a��!��'{���������
=]�*e3���Ih�+c�Z�#���R�D|��'�� ��A��a[f�;y4P�:�'s��bцS�1�T����C�TТ
��� 8HZrm�$�*pz�(S�I���X"Od(��d�Lip�ΐ)��+#"O�$0ca0�0aZ�DD�g�1�!"O���:e��ᛔ��c'T h�"O��#*�^=X�"���N���"O�ġ���"Qp|��jV�r�����'��� 4��>+{
�K4���wB�p�Oغiu �y�'\\Ӡ�Y���1KJ{�-J�'������7�n�`���o�$��'u��Bޒd�p��`�$�rx�DK�;+�)A�-���M*�7Mu��lΧY~(U��/�J��<h��OX-�?���)�$G�2���7$ӯ,��bD����-���>1�&��*�>�7C��j�!�P�<�`�)ʧ��(�!�AAP3rN$�`��	�HOQ?�[�A+c{�C�Ö�-�hZ��L�'ea�T�ֱ���p��L�rܫ�#��'T�"=����p 䄸MF�0#�R/B ��|2�2�Sܧ���	�!��(��ڪ8(��PG^��pN����g}�gHar�<3�L�}��m°��?6�)�1�8����A�I^��"N�3'�m��D+��Q1H̜V�L�&Z� �vQj��2 �t�b>�U�Z+n�JÊ�7UO�m(��&?	��U����IQ}�S�O�8�'I$)���f�"�y"�i�� �4��#ҧ�:�`�P�sk�%	�.�[h�t��
��l�x�	G�O�`4X���R����N�	N��`-�M�M>!@�Od��ڰ��J�� ��.jy��4��*0^����O�4��)0B�9 e]�Z�6�%��10E0�Mǧ~��� �f3�nm�A�E0��m�'�ڜ!fK{�X�O�>�I7��

�1���* �����t2<h؉{��O���3���v(����m�r��c�/�	9P�ځ��O��HrfI6.I�JW��o����V"O��eE��P�(�6AF$J�� �$"Onk�c��!!���!�7 ���"O��%!ӠN�(%��Å�:϶�X�"Om3�n�7�&�2A"�`��5Ȓ"O,��J��`2�����
��>���"O�a3�`����A5� e��"O��K�O
7t�T���ںY��Q�"O&�!f&ӎa�ꑘ�nK T�&�G"Oܰ���"���2���]��i��"O���c:Dj�񀂈�{o���"O(yi��<j.F8�w"C�'n�(��"O"����  �֜�ẀdL�"O\A�_��񢖊�~�<b5"OBT!VK��J]�U��r?li�"O,8�')O�|
@ �'�Y��`�Q"Oހ���lo �Su�Q�C�\$"Ov1�4O�F�6�[��>XqP	�"O@`!4Lϵ}`����nV�x�s�"O"Wc�+@N Q� ���t1��"O8IPp�-!#�ԋ@oةfid��"O �a�cK�>23a�]%~ �X�"Of0�׬2t}4�U��a�u2%"O�@8%N]��D�c�W��9�"O��S2�ߐ� �`A�] '���"O�=�#+�-jX� XCLJ�/�>Q��"O��g�Y9���Tʐ4+h���"Oh@A���JMZ����
	S���"O�"b(׭	�R�[�)SҴ�"O�U����)�$�)��S�6���
@"O���g�G�b�Jr�����x�
"O"a��ᆪwgI3���僇"O�e��Ko��<��`�y}�=�#"O�L9�Q�12�!6�Cr"O� �X���Ӹx��	�N<Q`��C�"O�"�#M�[�1�.��t�� �"Ov�y�J|�*�8���X�ލ@�"O���Q�*4 �d	�![(:���Y�"O^���<Cf��Q ]�v<�p"O4�k!�>��]
�}{�"O��c����;����!�v��s"O�Y�G�e
���7FτP۞8� "O�z'�=����$O�c��|7"O~�
�fQ�a=���;<���q"Ot�@�c;sr���!.T^b�0�"O�a(4CT�} �AdK�1^����"Od�Kg��WJ�����?[[� C�"O�����*�.���Q@���s@"O֕�.J�UǼ�����G�����y���d�:��5S�~���,L��yb�*p\I!�6~~tFAT��y"o�n�^��)]�%����A��y&�/hۼ����/��ڲ�]��yR�B3A[�� S!�$l���!�yj��
�2����Q�}�����y�X���v��*
�B�C��7�y��* �^%�!i]8�����/B�yb�J�Ni�,��Eu+�<8���
%�y�/H^�)�GN�9T �J�K !�ĉ'JxR���@���Aك�3'!򤙯y�"4��b�8k�`��݉~�!�$W�3
*H�W�+
��5	�͖?S�!��޺$of	A��C9�����m_�ff!��ʨ��a���8�S��D�_X!���o?��8F�ߓ8z6�HS�E��!�Z,e��$�~h�I )�a�!򄑇a����E[=R�)�(As�!�D�?+&�̓W�שO��hשd2!�Dj�b���*�lm�T��$�>4!�dSN��� �\�a��1U�%a.!򤖺A���;0��3n�L�@�@ǫ�!�䞜�~P���p�P<;%#�!��D8MlIyb��#����Ė��!�D߼P�1�V��<J�Z�P��U7�!��
zd(Y�B�
��D0!2�ϐEz!��Y$,"B։_��J�F�[�!�d��[�.p��L���L�1�ہw����'���bg�S�<�0��y�C5 �"أ�aQ2]Ύ�ʗ�A�yrb��E"����\�ԁk�f�!�y"�1Z5��� S
���DM��y� �O�����*E��@����-�yb�L:�T�A�(�&F��}(��վ�yRJ��%X6qx��=6�z�2���!�y2�%(8H�2�_}�\�G;�y��ъ�Ua!/�6�+�^�-۲B䉒��R@�#7�\�5	Jf��B�	9%����L��O2"X�T#�B�I��4SB�̑ �@#�F��lB�d�z�2�:���
�@@dB�	�@����m
*P|!���0-p>B�I�tM���P�-�Z=фf�e\B��d ��S��.�ZS��z�.B�
��S�&Ғ���M���C��R\,P��]
$�lx�2AMi�C�	�/��x�D�I�
�JH@�/��.ѮC�	8	\� ��E�D�a����Bn�C�	�h��b�b �P-`em�:dbC�)� �գ��]b�(���ڟ	�`Hh4"O,�¤.�> �җgs����"O��A��
���g�_�?j	�"Ob�����Af��❰s��k�"O�dX��Y�4�������]����"Oj퓓l�(B��r���0n�B�kD"O��;�
=|��
�jhp~��5"O<Q�֌�~GT\�P�\2h"yz�"O�< �gG�y_���%Ѱ%4
"U"O�p����6�bͱ�B�5I.�1�@"O��Z���3��ˆ`̊ (� �"O�ճ�!F$�����:7�HH�"O���l#O��(�5H	^E�U"OZ���Ap �yS�$��8�&@8�"O8a�` ���!C�?)�nQ�g"O�ő�KE(Zt��D�
#~��M��"O���\ 4x5�����Q�"O�Q��-ſ2���r�.'�@�"O"��_ ���	�:9:v"Ov��B���B(p�åZ��E�u"O(
V,�1  ��mַ}{��Ӆ"O�Ȃ��G
p����W��Z����2"Ol Q�E�=	���!�)\:*t�"O�*��޲!�Ya'��L��"O���U�e�ƨ�`L�9?2a�"O��@���5}ߔ	�K0#9�p��"O8eӁcH0i� d�E�y&���'�:�jP�N%?R��Q2
�-�|��'��1���ΡB����/��V|03�'���D��9��0Mۣ0�.T��'�<(��$. ����1+I����']LL�j�+��0�6&�y���'�N	�'(ӥ�@$1��ׂ�����'̖-��D����:�%$|ļ�@�'��a�.�7k�E���P9lvT�k
�'��ʑ�^�Y�)���E�e�*�'����
�$�Ձ�bvP)�'\����$k�8��N��t��A
�'S^�"��6q��[`/Hr�J�"
�'u�����!pLV���O�rm��"�'�b�����?9+���v�@Ï/D���$�����F�6q�O+D�ĉgCJ�	�W$s^$����;D�L)��<
j�JRiO.J�>� ��9D�`P�`�>�@cT�Й��xgA4D�,I�"�pԮ�i#�A�NY�.D���B�@&��Q�ˁ�"���*D��1��#j��]A�
��֨Д�=D��Պ�7.B�[��Q0j�y��9D������'��$��{�Xu�5&6D���$!��0I~�W��)�*q�U�(D�tS���33�L��� �8[f���J%D�� �Y1R�=�ե��G�P�F)D��!f&�S�ѳ
M-"�6�xBD<D�����8�����o� XC��	6�<D�<c�� V���1"�ͨ�(5D���p�PX�I
�h��D#���D�%D�<Y�B�|*���A4)���Gm9D�� cN�^Y�5����j1`A%4D��8P�J�Ec�8�e��u.���'3D�h�w��G:�1��͓(e�B���
2D��ү`�"H��(|��%�/D�0q0@�\1���\�o��hx&.D�t)�c�([+��as
3pG�Tz�-D�� ���`)L�e�b�)\]��"O�����؇w�YY�&NJl��"O.H�-ҝ�-9r�O-�\P"Oz ARGF�l�J)�I�!?�2��"O�2ҪQ<�ܘ����6��B"OP�H�6�P��q�Fĳ"O��B�OJظ��g��G"O�bh�-���G�V N�n���"O���/^�OҕT�[��-J%"O�����zdl;��ƛ1����"O<|ېAO�-ƅ8��m � �"OD� ƯN1^P EsQ#��56�0JC"O�h�&�j@��A��Ư@�!�B"Odq������kʩRP��R"O�������Hb��&c��D"O�����R'Fu�'��4f� Q"O�����d��q�ë��`b��ȓ^X�"�kNw2&M��g/�T��9� ل#U�As���D��b��u��m~"�YC*U�y^
�@3!�+�
i��?�l��k�z<݀�BG�0T¤�ȓXJn�;��P1X��9��/J(C��Q��)�� � &P�jH�QC%-O^<�ȓ](L�U� �� L	)7]����12LX���?'�x�Ȣ*�F�H���6�Y�2!_�W��y��A?+;ܥ��{fЃ� � a�\�U���2�M�ȓvQ
%�e�A��G�8x����.���"�
!{ȊLY$	?R��ȓw�>x����1=R��dV� 4�ȓ0ˮ��eaH:�094�A:-����ȓzD��e��4?V�!5��+!�đu�6 X1��144с5 A1a/!�&I�d�'�ʥ�ћ�HӼ?!�E�22����Ϛ�}]�EE#5!���H& �  ��   �  �  "  �  g+  �6  n?  �J  S  ^Y  �_   f  Dl  �r  �x    Q�  ��  ֑  �  X�  ��  �  !�  f�  �  v�  ��  ��  ��  ��  ��  4�   L � �  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��	ӟ��eVA�:"$^l�4ڻ,����ȓF��L���P����T��$�G}��ӹ;l1
pe��%q�uF�!M�C��B|�1``���e]��S��*W��e�'Mɧ����I�Pިq���>�P�R�H<A�!�d��z�@pW	�P�؀��Owْ	�ȓJ��d �#<]����2��݅�e<�R�(�]��!��
e&�h�ȓ"%мõ��% ���RT)b�)�矀��(J��$�*Q����y�..D�x��H;b^��W�O V,D�`�h��hO���q���9WR�pk��A22�H@�"O�@�a�(Ym:Г4Ɵ:ou���"O���A�T�O�V!1 �O-ȸ�z����HO�3� ��1��D"h������VS��0�"O6���MF�>B��vm��4B���!�'��6�'i�'���B��I�̜p�Έ �(9:�'���_��Ts��є����|R�iyf��>�}��+�&\9�ā7-@T���-�dX� �O�պvjF+/��!"Ώ��M �ў"~Γ��23�G,~`��훤z�ޙ�ȓp`���m̌@�Ȼ���40>�ϓ��?y�fUGlC��U�����V�<�WK:~Z= �-2#f�Ҩ]V�<��]��
,@�-1�n�X@
U]}b"� �hO��<�"�K�]�}���7P�]Ru�'���'��Q�5�G�O
��	�a��h�  ��hO?�r�շ	����aO�7�����`�'ݜ#=�O �Y��Ӗ,F��*�6�,�K�'�h�+NN]��@���� ���ڴ�O�"nګ�� ���q��8����:��B�	A�±yG�] ���c"�Y�U�8B�ɾ�x�Xd+�-C��Pa�l'����<}���)t*�̙�F��W-�M��Q5�yb M0E�%C�F��T��������y�-1��	a	F3`rl0TLԔ�yB��@A� I��|ɀ����y���y׬���#�|ɮL#E�N+�y�`�
Ŝq�b�R�e*c/V���/�O���e�u��QjP��;3G���'�b�ar�����UΆe2�D_�D��'�ў"}*��'3Jra��C$
0�C&Rr�'�V�"k]��R"���L����1��;�yr��9R�p�5���_� �1Q�Y�~R�)���?	��рo]�8��N 3(���oAG�<���+N��s�%�4J<��ic��G�<a� �Xcf�ǋƶ=��	��D�'7?�
�̒֌A��X���B �%}��)�ӿ:h\4JEb�%�W,08"R��D{��)�#}J�P0/;9{W"�C�!�D�6 �Y��,E�6�f���+�`�!�F�B<��A��&k����O�!��G�m�@�fE34Ef%Pq�
q��'Fa|r�
X��,
�ᄡ�
5�U/�y�!Y�A0�gϝ~w��8E����D6�Ov�$�ҳJ�Dݰr��=?�(�"O�D�Pn��N�J��N��T����"O���kݔ�RCv�R3:ۼ��Ԛ>!���	G &�1���U�:l��I8�!�ą*���F��f��2ǋơ=p��>!K��P����}J�%AR<+����*�	A�C�I�D�H9�MU2�N){��5�R��>1Qj�p�Y�rzGnݣ �d�'��O�'i*}��DZhL����� �ȓu�2!k6�+kH�ah�
f
�ȓO��0����i��\"d�g���ȓ�P�0@���
}f,���=e�RՇȓCg�)ff�d�����A]8@x��ȓ=��XԦ�-h7�Pqr�J/X��Y�'��~b+��6���a@"�fL��㜪�y�P�!��!�H!g�q0�T�y�쉕.ʝkA!�ph��Y�΋��yR-�2P�!�C�;qv�	A@���y�]�]�����Vb�8ŉ'�_��y2���U����^`����%W��yR��^~,�
�lZ�����(�-�B≬0U���Ӣ9�d(�A�9�C�I�@�(��6��sC����dM&(�C�)� <��)�r&��XG�Յ{�@���"O�̣#��!`���@��X�;��Ih@"O<��U�W�`l�×�/�&``"O6D
�O��KH�y�����' �'̈����t����E��!m|0U��''h! j�%9��"eR�-ĸx�'Q~!#�A��:��	W�����'��l�!ӋQn� R�=V�����'T�]:B��+L%��B�w���`	�'H�q�SbR>	�R�³�	DxJ ����?��)�'R�r��	�z�x����[�Z����'=��)3��1��Mq�+ւq�	�ȓ���A��_���@�/ϼ��,D~rS�0�~�Ŧ%&?����,y��w��z�<��KQ%K`�LY���c@�M�a�s}��)ҧ7�(��F�i�HLi�.ڇl ��7��#Wc,�:T�2/ə�n-%����	�L�@l�-�	dUsR�ţb�v��D������ 1�KB�L�x��v"3D�\Qto��Y��	(��y�i�+�Z�!�D�1Ky���F�f���s��6>�!�$�c���杂PF|�����O�!�D
�)(.�Ӄ��F���vA�(�!�� .�҅`�#2�)�Ӏ�]q!�d���|MSFc��cΎ�A�O��7T!��>s��j�
�r�� o7W;���Į�����YN�ɛ����'���2�)�S�I�d��#�p�J����X�U�<B��1�pd�qnDPH\|�")V�
�nC�ɑA2�H�#!ی\�0���9k�`C䉿"eX��$�G\����'�;q�RC��
Z�l���@+<&��w�Q�sHC�ɇv� 0���\;�U���
C�I$!��]b����i��&�|,�B�	=;r�`����	,��i� i�;;�B�	�s��E��ߕ��!���	0]B�!�����DM2̄9#��B�	�d�81Xd�Z�Z�1coA7݌B䉐Y�0������KK��8�j�'��B�I�9���pU  ����O-EC�	6����r��?r��0Y��Q�Bf�C䉏#��ـ�MB+L�Ե���	W�C�ɲ�6�9�k3E��@d(�=&tC�I;q�6ݹd���-��rA��u�
C�I�R0���7�y�WnL
H��B�I:5��R� J���I�����"O�y�K��>�j�X��w@j���"O&���?���I��S�p�<�"O�`p��b��}i�(���ː"O.ekD�38L�MV�G���T"OXx�!N�B�|�8'�H4}���"O$��p���\" �K���M��8("O�q�F�l��Ib�AI�z1���"O���5�M�=�"����X+'u��1"OnH�E�6͒5�.G�?I*Q�"Or�5��5����ӬΎeZP��W"O�t��L�}�=���C	%>
�Y�"OZ-��*�w��}C��̕3:���w"Ol�@��w|�Ȝ^I�e"O6l���j�J�Q�I�y;"O�� ���H�>uh`�P�r�Ir"O��b���	��PS゠Sk��Y7"O~l)$��z�ԹJ�A�
.R8,�2"O��i׮дh��:���i�Je�"O� 2 �c/E��������� ��L�6"O�=���1Y8�-ىC,��4"O��AE���& ��O׉h�&X"#"OBpX��g�d�Q4�W���Y0"O =�b'�9rx�Ճw��+> ���'p�'���'��'_��'b�'l��k�d�-[8\0to�I>(2��'R��'���'��':��'3R�'-�� ͔��Ti@���*W"�Y3�'2�'���'���'�r�':�'l���E�%FF��f/�`f^1���'b�'�"�''��'""�'�'"T��U5o\d��$L͟~���'�"�'���'��'l��'2��'�B�����X������ S��`��'4r�'��'���'�2�'y��'*�!�����88$�q�-�	Mൡ��'���'���',��'�'a�'��:U%U��F�L�f�6p��'J��'Cb�'���'���'���'D^��F�V�6��y�g'�-��q�'+��'�"�'@��'�'��'%�P���ŉ�Y��ϝwAz5
T�'C��'
B�'Rb�'�r�'K��'M ���.fPx�����X��x�d�'��'7�'!��'f��'���'q�Q�0"lzP#C�ɫA��'��'_B�'7��'z"�'K��'���E���2z��ąL~{֨��'K��''��'��'�2�l�v�$�O�B"�+W�D�2�@�<�inyb�'Y�)�3?i�iߺL�E��q�Pk��v��E��K&��D禵��{�i>���M����2-���U�Z�맥̦Y���'�h]03�R��DK:�L��g�U$��ӭV%꽒���8y��U//�c��	oy��S4@�p�r�M�N\@�9��S�`h�K�4B ��<����	s��n��s�v�y��*>���N��m�>�M��'��)�S'|�v��ii�p���eO8�q&i�8l��H��x��[�nRb�T��ËJ���t�'W�	v�I�l�:b�J�Y
貜'6��q��M{���b�8�3-Q�Z� ���?`�>����c��k�I�MC6�i��D�>a�D��F�I+��5,���AaJIy~��mR҅B"Ԇ��O*ƭ�!┒	�B�ͱ:�ެ`5 'h�"����5�@y������P*{<d�L�,x�7����͓SI�F�F�������?ͧ8϶h6� 5eʡ�����͓"���l���d�&Y�8�B��x�"��KP"�I�@@�^��M�!��dsR�qK��)Z&L�'3��1�}՘D��풧o�,1�aI*��0�N��F���3M�2 �EL�	H!��.B�Fq�C�ɩ6
����2g�щrO�v�����#,\@Je�� �"��I�����)Jp��&R;t;Xq��M�	b��YP �v�d���ZB�L��͙�h��a�d˘e�v�@�J�;ˤ�jF��B��y0G�Qn�PYrϜ�|���J�ȟ3�A+�
ϥqTx,`	�0>?D���^�?���d��Q7��O:���O��)`~b�NR� (g�۾M���0�Ν�M;���?��� �?I��?)���I?�sř)XN��æD>Iψ5��huӸ%y���O|�D�O������)
d'*hb���"����eO$�n�'�H٤�,�)§�?���ٸz6`e�@�~��{���.5��F�'���'sx<��W�@�O��O���h�?<�\`S(O�g�p��U�ɲ�k����'���@��)�"`ʡ`�Kƀv����MK��T����?��X?���p��(�n������p�2�!�G[|�&���O��WJЮA%�I͟H����@�Iڟx��@H�2���/
t����9vb0�d�O���O�D�O֓O�d�O`H�A�B<*0�1��X)e�����/�i��9:T���	Ο��I��I+A��-��]X��P��#|L��6gg�8֯b�P���O��d%���O��dU����'�iD�)A�ݣZ�,ɲ��w
���O��D�O����O��d5y��D�O`��H�2�����7�T��@Cж=F��oZƟ'���	Ɵ\�C�T�'�O���q-�Tܔ�d��m�Uڔ�it�'��	�e�f\�N|���1[`��di��,�p����rx'�ĕ'�bdR��I�?�H��X=LT�BD��0_��(�y�8ʓ-�f��'�iz��'�?y�'Q�ɊR�$�Wd�_����V�K���7��O���
�a����|2���&�h��;]���5h��~�@���x��+Tˏæ��	�p���?YjH<ͧ+�|�HC2 \�����Z/�8Ӻi�ڐ�P����؟��3�	ʟ$
D�M(]a&�#RoC�d�`�� �+�Mk��?)��UvҘ2�x�O�B�'�t!8�ۆjڀ 9�/�42�|q�(�>����?�Ԍ�F��?����?�Λ�$�ꆡ�}7z�z�MAYG���'�t�;0�&�4��$�O��茕�'.V<���+�XdH��c�iA��'��'h[�\"�ϔ)ݘ�z%f͔L3V�jT�Y[��J<��?����$�O���
i� ��e԰Rz��
>:*�H����O����OD˓�:�H1���9���.)X�s��ѡA�eQ����۟��hy��'n�#���IE-8�&��Q+P�l�	�N�\��ݟ��ǟ�'i.��#8�i�,3~U��!B
8�h��N�:�n���L�	Sy��'��f���OSr�2�V�M� )4K��F�`�Xߴ�?�����DD26�X%>-���?��$O����@�c�!��I�gi�O��op�LF��֟� ����O�=@~�ᥫ	p�Y[�i���(L�V��ش-���ߟ��ӱ���%c��:RDR�$��	ku��lǛv�'FҪ̩D��)Z�g�(C����B�c^�s�H�&' 6=L�Xl�̟��ȟ��ӡ���|je�ޛ�%�E�Lˈ�Z�ok������|���?c�T�	'p��PoX&�a"�'�".E"��ߴ�?i��?�䇅`������'��OC�e�"��3#9Px�B_0	x�듡?���w^�<���?��2� QA�VjR���OfC��0b�i!�$���7��Of�d�OR��|���O�ȲP(9p>|C4���g�Δ��i�t��R��yb\���̟�������8T�
�j⮞���x#5�.#2윪%M��M���?���?��T?]�'���<��� ��T"f�~H���H�T`�I�'��	ݟD��럤�I���ZQ���M��6JD��DN:g%�X�%[����'���'3r�'d��Rw!d>�Q�EGh# 9õe�1�`ˡD��M;���?����?I��?�Qm�s=���'��Z'R(��� �� *��	e���)�|7-�O��d�O���?�����|j���~b�	6Va0��-H�K��M(s��n��@�	�H�I�`���xݴ�?a��?��'d��Pңk�;
&Ի`n�
i�Q��i{�^����������X���ܴ[�k!�д�J���J�n�ڟ��ia"��4�?��?����J��J�����LÉ0!�`���(���k�X���	�(�A�Iڟ�����~�ӄk�(�Ś�D��u�ZO��V��/W�7�O��$�O��I柒��O@��)+(]�b荎t�|�0
�#}�D�mZ4����?�g��?�u�ۓG�
0 �*ۋ.�)"a��p���'�b�'�:���Aq� �D�O��$�O����ٺ�n	.Wt�j�L�;vhq���iQ�U�(q��m��'�?y��?����[�.x�����I����n��H^���'�,*��v�d���On���O���O��$կ#�������i�hJTX�P?�I�;G���cy��'��'��'��s���g��Q�q��
_ހa��o�� ҈7�O����O4�Dq��X�l�I�,����M?1N�mq��\z��#��h���I֟\�I��	��`��j�l8ش�8%qR�ݽUیQ�sLíN��1���i�"�'��'3rT�T��3nR(�S�q�E��\h b=��m̷O�l��ڴ�?���?����?���H���:Q�i��':DxL"�b��2 �z�0�L~�B���O���<�8�2U(O����vT� Z�h@0W�@�!�)[;'�6�O����O:�d��x�m�⟼�I�|��=4�h�-�W����
e�p�۴�?�.O"�$��}��	�O���|nڛ�Ȳܕ9x��ab	f.�6��O���[�j8�!m�ڟ0����$���?���>mq�U(s�Uh��\M*9�1©>i�@�0�������|�H?ͱt`�H����a�Rs�ȈeadӔY���������x���?=������ş�؃�ɕy�a�dD#6���"'�Mk祊��?A����4����J���<뤸�֡SG,���!S�f�>l�ğT���4 S��9�M����?���?��Ӻs�-'O#2�ڐ
G2Y(A8���Ҧ!�	fyW�yʟ�D�OX�SV�d�q`oD6~XpR@U�,9�6m�O� *1����	���Xz��f���3{詩@'G�2��̗��p�4����D�O����O��d�Oe�C[���)X#���R6�U5�|l�����	��������	�<��,+����)�Pr�!J��� ��(� ��<-O����Oܒ��,ZQ$��|tȈ *P X�J�����!�D}��'4r�|��'5�H�+��dڿ��l�nO� "�g����0����'�ȍ"�)� $����fE�:"U�pg��0�n럨$�d�I�(d�(��n�l �sn�:(r��In���7m�OF�d�<�7l̴
5�O���O�l�(�j�0a��dh�	��8���O��
:>��'�9ZvaF s�.�����
��Ym�bybM�)��7�U��'r��=?�G�Y�8�,mY4싫/��C��BѦ9���袣j�H$�b?%b@�<I݊9�Kҫd��E+y� ��i��I�I㟈�	�?M+N<��d����=-Fv�ܻG�F�a�i�����'"ɧ�j�Ć/�!@d��wU]�� �_���n����I�4zb���ē�?a��~R��j��,I��Êjg*h0Q(����'n�\R7�|��'MR�'�)�W���8H+�m�� Ĉ�eg�L��W�U�@`&���I���$��X�Ut�ْ�*ӳ�!���R&]|�D@����$�O"�D�O��p��E�#Jn���7G�(txި(��'g2�'�B�'��'�R�'	�U�,��sS܌�'͛z��$��S��ybU���	���Uy�O�.y8��WAr�B����d����
$�O����<��?!��'�i�O�H�`���*��Q�eQ^#�<p�O4���O��ġ<A�$0^��O>X�q@̘w�bL� U,2�x�+q�|����?���O����3��7}����-��㡋D����E3�M���?9(O���3CL�ڟ����#z(���/�Y�D�j��uhK<1��?��
����ɞ(	!@��f�<f���:g��mʛ6Q���&I׋�Mۤ\?A���?]��Oh�&�+����L@'��i	�i�r�'�D�r��'fɧ�O<DDjvbכ;n$ ���ǐ8���4q��8�ࠂ�@)�1�'�˰@�v8�����>�l	#	��� �(c��V68�:gH��� ��7|<D�@ߤy�����ݤ6��#�S<����K>�=ʡ��=h��a"f��i!C��f �x@�2� �S�&l	��`��� r�X5�@�Ӗ~N�9(���} k�6Oz��p�&A�-E�Tऩۧ5�p�r��OD�$�O���������O���[7��ykB��>�0�'�\�b��Nڶ#(�Aڳ��3He^��F�ص;�L�Ba�I<-/��BL���Jp�\��\ŋ
���I� �ڛvl����CZ0C1����C5ʓ[;T�$F@�F�{7FI4�)��	���x������?����'Ppɦ��#;�\D��8k�"����6��]�	�bh��BO��j�1*�)V�	&����4\�v\�,�6�G�M�ᦝ�	�c�t�6�l�`d����p]X��I����F��	��pB$հL��b����F]��D ~6*�(F�3q�j�����8�6�Ʉ��V�ܢ<�,/aݦQ�rlҏ��P�%�*�ED�ν�]��\+SJt��T�u[2�<A�%�ݟH�I�����D����'Z�N��!�S�D�d�O��$$�IV����@�EC�^kv
Պ\�#�eDx��i>QK�4f�4�����k�.�(��p!P���VX� 	�i��M����?�,��Y�#�O��s��_�s'�w��u�R��O��ē�7�`zKT=r��Ejz�!�K<@��˧z:�	"M��L�*)�V��5>�HY�O���1� {1�5�WOÒ(|	y��پ���͟�+�@�n�MxP�D�����ӗ>�Р�����_�H�? �P�G�L�K|LT�BցY�b�D��Bx���� 9�� n�b*��v!�Y�����=�&|�0foZ�U������M,5����ҷi�B�'GܻH��$#��'�2�'��wa�X��g�;%*��"kݣf����䀈+�@�r�ŞeJ���=`�O�T�C]w�*�	2dL0[�זu7�xpe�J�,���U�.Oܨ�`tE ��P�0��;70��Q�>O^m�ꔟt�N1��fJ�nh�Э����c۴�?�rÇ�?�}�'����������>U�� ɞ�<���Y?f����鋤z�r�soTzd�D�O@�nZ�M+-O��$�p���<��n�i��p{�h	�x��RFꞼM
,�9�K6�?I��?Y��e���O���O2m7 E: ����Q��1h;�E��Ħi�Tb��<Eȉ�hLm�%d^�[:̜Y�ė��r��Aoۏn0� ��@���=�CbVe9ƍ�-�qqà��M����I,�M���iWr�'8b�'���'�ӟh��}	���'��a��jV�C9���?���|����?)M>I7Ώc%x�R���O'2���=��d�O�`o���'�@R`'{�b���O��e�S�3��	�B�!&.�q.�O��Ǡ R���Ob瓖���[ ��86f���[Ʀ�s��i��������H�S�:O ez����*r�C�^��7���2�2gdpH ��%O�qp�x��?a���򤌗u�@p��M���1��r���O��d9�)§GC0b��L8�p%���I_�td��8��6
�7���84����G�9�yb]��B̙�M��?�*�F9K��O�Ł����we4qAt�rn�I���O~�d�s9���'K�F)u���ݚB��0g#Y�Ealʧm�D�d�>���إ, �8�O�)ZR�U7gj���M_��!Hf[��Fs˟Lx���T��h�"#�7N��bӚ>� EFџ��4d�f�'L�jL�S�W�u>Q҈ГW��=�E��O��O`㟌�0���]��D�S�N.4��x�	Ni���d�h�
Xm�M�ɤG'L\I2���&����Ø� ]HTy��՟��ӟ0���M�YvDl����	ן4�ӚIP&���l#'Ԫis� �HH��O�Oʖy[�D%[�Yi�h�Z�ӑ5~� �l���Ą�jeqꕦ[2p��hjׅ�7z!(�:��f ^��f��uT$�>�2A��|�$fʠ	��C-"x�S��s-m �M�����P��4�����
�KT*�N�Q�BQ�/�t�@��&4��2��8}z�*�@C(URҍ-|��ǟl�ٴ���|b�O��4^���-R>I�L�߶V��B �� � ��f�������ן��I���	�O|�ӁQ쀵�1��
G��5K�n��s|%�����T�p��(D�B�c �^9F���ɀ� �2�ɐ)��㗭��f��Ń�-�Й"��N��$i�%@�u{r�	7'��`8a���@��I
��r�Z��pb�O>�d�O����<�����'`h4:��R�zpR�4��o���

㓪�Y��BoI�(��	���6$�Dp�<�iI\���bÁ)�Ms��?��R��j)a�lX�5� �S��'�?y�\�&�9��?�O���`v��#T$��p��/xT��"��Z�r������RJ8@Pc��$9�r�DNQ�'��8@A�Zy��%�D� ̢u�vRZOb���A�	�����O�{dȡ1�#�S�'?f8�����>I`b��5)h0d���c�\$�rL�<��?!���i	�-�v�6
�
�� Xg��Ns�(E{�O�N6�W�xd|i��%��1!#lX�,^|��0�)��<��F�\)b�po�6��]���n�<��IѺ"�%I`O6q�P���h�<�6��()� b#�ϲer��C0,�a�<���; 
�`�A:z$5�t,]�<� 6}Ap�:;{�	G�\v���"Oj$���N*H�����irPI��"O`|�e�&�lI�,Y�3�"��6"O�����Orb�b�� 
��Q"O$ӂ
�))���٠��.�x�3"O�� �,Fs��8cF�A�T �"OBX�"��n��E�&�4=��"OzL2R��!n�z�JwdW0	��ݻ�"O� �3d�y��� 2�� M�0"Ox48!�N,^x3vĚVJVQx�"OTDj��>Dg���?�ؽ��"O��1�f�Ppp��
�2Uó"O6p��٩#���z�ϗ	=+���T"O��	���K�P��'��&xz5"O��3#"
:j�d� ��_X����"Oֱ�f�/M挭�¡]�Q��� "O:����H�$�61k����X�P"O����]� ��1���6��pФ"Ot}���[�v5�F�F$4��͠D"O �(���8������D- ���"O0���./~��H !Q/��"O�̣o6}A����)��
�G� �y��J�Nv ��͗G�0cc��?�y��#W�i�U$�-��j����y�a�Z�P� І`q�E�Q!�y2ř'�x�b�N[�`at�-�y���4�B h!GW"�Fy��R�y�J�z\|� R�ҹ/ϰm�Ҧ���oO�lGx���H+Mb| R&���w��H"a��yRˊ�[ ��	��B��;��׿>5qO�X��O�g�I������L^�C�ͮa�B�	xo��2��,$���Cg�C� �	��{�̄�ɕg���PfO�zY�5��F��'֒��d_�:��4��N=?	��Q�.��Q�b�H+B=i�
e�<�I] ��d�̜n�R�h��G�ɼ.	R�j��g��<�����&�F�$�dYk@��t�	*lUIE��� ���KJV�  �ERpA�H>j�`@���x�*���'
�-�N|GJ��n�2��B9j�[�O�EH<��Kڸ-���24C��nż�Xc�ۻ9��� c]�x��HW�)��f^)c�ɀ3!�4ؠ�QC�0Pz�і.MYx��SG����'E�� o�)�@���� m?:)K>��� -�:+W�O(rq�Ȓ&�mܓz$�Y��� ��ӫN�%���ף1G�N�Cj���?��0�I
L���j���7[�<�b��'�Τ���ʎv��}�1�S�z��*^�b��`���N�0�w$4���A ֌O�6� f�'�:$?b�ݜS�+3�E/9ʔ���:$��A�).�f��6�"W��r�����'�1O�yC��"#U.4�C$Dܸ�v�D�Y7 ���a�,D�����'3nA0#�Ӫi؈M���aX�h���A�.�r��t]��+U�4扥4ݤ�)Q焦��g�7�b��7O��<zA��8�J�D"� m�p5;�h�$A�@a��!����O�XBᛄga��( $Z�ҝ��oO�e��HjtN �h	A�a�'r��fA�1S��łb�W]���#O?!�T1��Kh���DX�am��J��/�ܝ�S.���C�ɐvr���i�nlisaC����A�wO���4q�P��|�dC�+�yRZ���d�0x���@�GQ�4 ����0<�bO$R�r�02�&m�̽3f(K��)@)�LD�c��o?��	������'��h���'N�v6�i~�ދJ�QQ0Ô* *��%/�~B���Y&TxU��myx��T�U��?�|Γ4��r�F/:��!�f��d�H'�g�Dao9��m0�����0<�äӸ+X��a�2����`�C.}�:�������M[bɀ<��yș�yʟ�OlT0V�˳2Y�$ �44�(�R®Q%�0>AB�����	�-c��R�o�[�N�s�EA��y2���<���t�d��T�6�u��*I�Ê}zV�2RG� ���F|�Ei�X�c�Gߪ��)B�G��u�4e ���6/��y��t2��S�����I}��c�j``�@}LX��CΜ�ugӇ��D�2j���a�#��9`'��D�)�v@�4J�CvNXz�A�+r�����d�?0F�)_�|���x�$ٹ	4va�kT��ɖ��2V��%93�6O� �Ȑ'�ߣv���a1	�uA4�����,9�<h�4v�&ʓ�M�sӂ��5��iݵx����h�xQC���E�v���K�9�}���<I�+��6���V�\�Tf����>�v��TYEm�O��'XJ�ӟ�<K�#�> �
- �	I�^]��S��S�"?�P`��2��6ώ�M����<�Q�V`�N�`d�5%�(��P��>�ܴH �QB�KU��Z�����'x��s&G�:.-��NGVʁ��':��s5`Y�.�Z9�V�|D�8�_�(O�͉��ŘAw^,I�-������@N˼x\^�p�ղD[b؈U')<OL�Ѱ	1K�A���ظ`�"�D:M0��槅N�@���a�Gݳ��(IR̓1�,�O�x0�ƪ�g��.m��A;u�E�o�T��R�h���'�"|1��F��D�1�h�17�ո��ĩNA4A���E�?6�">1�ӟZ7�:�!�h������<�m�]z�A��(��,4��z�K@񀶆K�Yv���K�|�T�%������j#�t� �y#�x��`v� �2
^�K�3j��8�f����$�=�H�2 c�{_6�+'I.+,�9�W�C��9��mC�2���
-O��)�HVz��xP��.�j@�&`�Bd$�sF��>���4(U�'�7ݟ�	�CA�d����x<H�B�n8�9�;�H�b��6l�ā��>R B@ƅof�)}�=���kܓ��9�v	�Č��j��M��-�O_�8�'��|����X;bC��E (J�❘),���X�=��H	M>��H���T��T�ވ�Ɗ����D��]}�ͣ�(�T��[a�۹��/��M��2O�q9��A;����@\�������y�a �9(��B�L�`\09TO��X�B����a��e��#uax�S�7h�႔I�5~gҠ*��C2	�:Tz��Ody��&�R�:%�0O�ဘO��Ĥs>�X�ss��/F+6 ���T�_�7m>|O������bg�,���.JVt�Q+�xxF��<j�^m�lU^5"�!΋�c��4����o���i$��^l�S�A�=���d�#5�F���T\�''���(^�^��6�uGF���'}��'f�'3]�u�AAB�B�P^�XWO�,�r����~��Ӛ:�f6�ۙ�u').扬QX$��\�
ي���KrGp7-�$�ؐ�S)K�-�։�12"�D6y:7�Hu��E(JgV%
'@ܺP�P�f��	���dE�0��b
uB�:��$OJ��6KLRT{5�R;*7>� S��n��a�H�|RM<IU�D�"h�[�3'���!�]$L8�-���'n"`��wQX5�W�ǑI䮙�g�RRR�Y^��'q���$�OHHK�oi�5��k�d<.�R�1�Tʠ#����Op�����`�"�tEЕ<O�)d&� z�Tqg��x�8��f�0Q���Y57V�H�K�0p5�E�t�()�Ɇ�Z�zD��.�O^IDϜ�l��W(h21r1�>�Tc!}��_��E�vgڊP[�d
u�@��?QtcH�+���
��^��U��ɾE�"e��CB�)R,A�G���R�Yp B���	:��'Ѧc��H4��dq���ޖ}��6k�3����T?����_c3��*F!��?4j�A�X�_t��7�!ʓ��'FZ��7N�a�h���R�^�����+��ܢYj�ȅ�~�����'��R=�8�UGm��D���!?�kTR/��˖�S�Z��C�OR����'M��	]l�U��+oj�d�Ь�@z���2�@�ӑE(���	4#� C@X*��]	P���\� �2�44O���^���\9�A=������>-���h��ߵ#����(��9�ax�`FD.J���B޻3�������%�f$C��d6�d;�Ğ*M�:�I%F��W�D\��)=D�����'��������y�)ռ{��YH5�
#�^D�0���~R�';^E�4��%]R̹s�P��"2�Za��:T���(O��p�@�D 6�J6!p�8PZ�������|���
E'c��!�!�s��!����y���FZ��'Ϫ	�,I�L�0l�4H��[;������KA��� �6T����Oџ`ʴ��
0e��1�f�.z�R$	"@��8�W��<S�F�$U�`����ă�lL�Z�I�h�XH� Ϫ7�<Yh��'�D؅�	��u�"@̔LP�S���7"f�@Be�'l�1�������G,Qq8A9�(I̚�r��ԝ��=�Ĥ�L���WM���S&R!|�tcu
jy���$� CvQ��\�V������0FT�f����ǥ�1Z�ۃ ��,�Q�Z��O�T��[#4� 0�Q>y��X򧜟�h�͝.@94�@��Ւ i�u��S�f\��O)tx\��H<]0�\��dY��y���R��f�N��큇<��@0GA�>ju��i℁+[yʗC$3�$��ɱ_^��(vk�,6߲�c���7���aɫ��a�!��|��'�^4�7N��McJ<�0t�``�˝V�p}#�b��{v(u��+,O����.�(77lQ���h��{��n=�0 X�c%V��'/�ajt��AAz#<ͧ#�V�gA�H�6-,���'"]�uHB�H�A1c.J�-�tQYV䖾|t`$>i!���F�$�0v�µ.�ݢ�%���tB��F�W�y�H e�ڥ+��'�JeK�$T<+������]�P/v8ҡM�d��İ�GH
z����j�e�)D+81OJdIČ J�m�v��״�b�h�L�� ��.�n���x����E,e�&yb7�-y-�iX]<�\�P&��bӼ��{�Oq��M+kL�E�? �iS�ψ���q�`�rr�' ���Ǐ�kL�(a��[�E�A3��*k��$���(On�I�o�@1��
+��� ��Y�6m�"e����fH(Q����e^(�Q�� 7g����nX+���mNR3-P"�)�Z�kC��Rn��< ��r�H�pn�� ���'��Gy"ˋ���  ���k�����Ԛ$���H!02ɸ����)_�N�K&�'P��'>�I^��B$5U_>�+�DY<Fぱ��AE�w8����քj�8eC�NQ�2Py"�A�jlL���?)E�Iy?y�w�.!�qo�:��mA�G/�E��L^Չ�i�d�T���aW�it�s拑}P�dY��d�}��$O�������o��d�U���B"�%�ԭ�%v�����Y��HOB�c���	q�R�2�����T������|!Z�[Bi�o7P`qR%��_ț�'T+=�(lc��*���j�'�&��O
�H�Lcw	3a��Y9�4]��H!�)l.@b"�kG&LF~��G	HsI��G�o��`�P�y�Z�.}[P��)��0sTc�	Q����֏QQ�'��}#1��:&jm0%2�biqҥ�a���j��O;y���Ҥ�'FZhPC��n�̀fgC�d�$ٚ�-�d�m�4PC�mʖ��s�d�懜�b��G~��	V��5��ϵF����C��O�� �bN�F�p��Ҡ��Y<q�<OΥ3�X�k�aw���7r�1;��LS�T�
�> �`�	 r���-߂sĔ�	� "����
Z�,:�H���=}J?����֓vr��ͪ�N+��"D��a2.{�( L��x�.9�fF�;fs�扠B@�S��%"���@�9�y򤑽zjd����g��c0���0?�Df�g���!ͶG|���B��I~ �r�BD�ly��[{≨�"�G}�ͅ2/��0׏��O��墔N��O ��T�?_f�Ps�����11�p�"�i�A�M�֬ї3M�����?���Ȱp����1a�cgl�7���	c��_��3r�'S�YE�4��(���Hף��ck������f!���xj����	")�`9�sE�5`��7O�0C mg������O����	9P���N����""O�j%��)�0��Ƃ��P��"OD|����=s	�h��&��p@F"O��b�QX���c�Si>�0�"O\�]8k� ����b����!�H/
��-�'�o�r��Ř�!�DS'.��,�>i��K@D_)C!�D!e�rB��16}�T3�D��!��o�dp3��<��Qd�� �!�T\2	d�=V��R�	N(j_!�]0r�������S=�\kЭ��I1!�D�
0~��Tכ6���υ{-!򄈋g�p�D��.VUՊi,!��5Ԓ�
UO�(�k�P�4E!�R�tzh���a�D�k�V?!�r��e1��j�H8j�ҋE	!�ą�?а�cƎ�+�����܂[�!��)<T8�b�(x�����i�!�O/@9 �ie΅8q�:�8PJ��`!�$R�Sl 9�BIP���]QWJS0)"!��_� �YA��Е��N�)A!�d��e�t\XХ��P1}���:!�$�3��vh�s���F�.!�dܿvSt����E�EԘy1�v��'�T��g�Z7{.�	ӗ/ 9&����'*�R�E)j�a1�c�!J�dK�'�0�2Ɋ0>de�w�P�H�2��'��0Iզ�C��Eq7��w��Ē
�'n� 0���Y�5ʜ{�xm�	�'��IR���.(|��0HLY�=�ȓl�xa:�!�:p�(ju�h@�@��Q� �r�),�����<�L)��!}n� ���T�� �@�_�<��k�,i��nT�S�U��7Q���ȓ)/�dk�J�Ɇ�K,�-�@�ȓ^�H�R��ޙt���5N��T��S�? ���+̒}u��r�H�Ȥ̚"On�����_�����ݐ	���H�"O�|�w R�x���A�R;F`��"OX�խJ:9"�(�j��N��)�5"O�I���(Sh���g��=}��"O��!T��0i��*L\<��"O�m�bI=n���1���*0��E��"O�d8�%L�E�d�7��i���"�"O
��CV � ua�A�|�^��"O��t�X�@�n9J�Ϝ+G'�ۅ"O�CT��0=����E���h���)D"O�E�e�I�o\D04M������Q"O��ת�hî�r�ֻC⮰�"O���m��X��Ԩ�Ē(1,="O~HrR�W�e4 ���w)zQ;g"O��Ѩ\�;%6��-IO��!��"Or��r�M@��`b�2Q����"O��Y%�ؿ1֮�3s�S$9� +�"O0� UZh��9@�.+H8h#D"O.��$c�p���fe��@��"Oh���Q�Jj`�@ċ;�@He"O�K�'I2)��%`eC�&m���r"O����Q�=�t�u�ƒⰁir"O���À�˲�#��Z(Z/���F"Oj-��J[,�&HS���'¨V"O��Gl��RB4�2�ލm*r��"O����>1��rƖ>'���"O8�gBΒSx�i�F�Z9[�"O~�pQ� Y d��,c`.! F"O�<��(s�$8⭗A>�M�"O��@�,��i�eL��N��1"O�5���*	��-� ��W�N܀6"O�5�Ũp�(d���ސ9S"O���EME�^D�LEN_8T��"O���k����е]QLl��"OD�)���5(�l�(d�����%a�"O-[F�����peB@
7�lZ%"O�h:��OH�L[b��pQ����"Ol�귫%GΦ1�B�$�١�"O�D��Ȕb=���D�\�$ʚ�ۇ"O��$[�:�Lr1G�I�IS%"O5�4� ����OV�\@"O��8�E[�U�4�y�F�t�R�"O6�h���@����Ԝv ��d"O� ��$j�,q+%bV��BU��"OJ8J�l�#��؋7��A�P�r"Ol-���(GH�h�V�;%��! "O����$ǼW8Jv/V6O�(�g"O� {�&��c�64���N):�D�"O����s*�q�ć2�Ƥ4"OlȺ�&7`�Y����,��b"OJ a�_�F2I�BV�s�B���"O�E[����H��6a�6p숱�F"O<��.I	*1�T-ג!��m�U"O�t#D�jt:U�\:d8�E{�"O� ����S���!�ŉ�����"O�h�t�F�s�ڐfj��t�ĝʕ"O6IRu��1 4�!HIn�(�b�"O��颀�46d
�Lʘh0\µ"O*�rF#[W�0���E��[$=��"OV� ��R��J����9��0 �"OJ�"�ʇ� *�	$!Դ� 5�"O A0e��)�X�#����R�����"Ojp�#�tU���ׄ��9�l��"O� ���S�T�)4d|����qk��"O���-�^���
�B<[�y{"O�@YB�E��8��.�<ɒ�1"O@,IքדU�����Z���J�"O��#Xg�L����FSν��"O4-���7Z49��F1w��)�"O�щ�AP01�DkB+�;0�~�"�"O���r%�0�����]s�m۳"O�wE��}�n��ED�\�(R"O��!*�5)��d����>v6n�ia"O:��'L��&	��
 ^�0�"O|<���,l���f�&�u;�"O��r���w����%֥��YZ "O��b�GJ�v�)�A�1JmV���]��s�I�Pw��/X�i ՗$/Hu��	u����4�)u���>^�y��kR�`�!���DȢx$̠9�M�B��!�Ď�[��Pa�L]&,x��2�!��"{��ܩ���:�����F�'k��G{���'�� js��44�&	 *�J����
�'��J�I=^������TEeY
�'UN �j\�p{�� `��~0�Ei	�'(2���fL�4njp@'dOL("���'#���5b�+Y��4@�iE,?� ��'MN*�:KH|��D�4h�H�b�'"�lSuU(}n$25"Qx�؉��'��5��C#p�(�y񃙝n����'d�����>��}� �Pt�t�N���I{�[��_�=���3��А[�JC�	�D�$��싏R��yڐ��)$C�	�p������.�daCW��?�&C�	�Cg@���A=Y�B��4MG,q�C�I�;$�����K�Q�� ����B�I�A��B������xw'Ё4��B�I#S\r�YG���=�$�˟��B�	z:�����~��YX�/<p�B�ɻw�$;�E�3`�Ѐ����K"�C䉵M6���������TC��=��C�ɠ�"�rš�>L��,Yd���`B�I(_(6|��$�R���@�Un�@B�INL�x��FN.c$�`���+�B��%D�`��e��i��Es�u��'ƨp�DQ8b���lE�< ��'P����ߟU�ᡇ��6w!��0�)D�`�MWc~�4��F�S�v  �%D�؊Ǝ�9R��y)���.]�j���?D�XY&nQ�}5���0�244�@A?D�t聇�3�t違̍,Y��z �(D�<r&c��rb�0��mE ��t(ԣސxr�^.nDKF�O�D�"�T�le���2T�tڣ �`��D��"p��ȓO�N�Y&� jmL����܇�IH�	D�`�p䉍	�<�1�&�8��C�	��t%H��_���f+ǲY�C�	�
�^萖O�q�YP2�ߵ(�dC䉣����/u	�Ya�߿*fʓ�hOQ>���'@�~��%*fA�4���dO#D����)�6'�x��
2>�%kp!/D�P�t��6*`�ɒGU>�����-D����� ey)ңA�?"6�Q�!D����%���Y��LO4��&h2D����ى:���A�O\֤���/D���З%<�4*�eL,x���YSi-D��: ��KJ(@.�5�\چ�+D�� t-:�G I
�yzG��� K�"O����TfN�2��T5Z�V��"Oɱ���gy��kC@يju�0�"O����[�q�j=Ҁȅ:2�䬚�"O�$Hv�H�b�Yn�F)��"O� �b�-+��}6`D�b���s"O�=a�
�s� Q�O�3 d��"O� ��G^�f��i��/b���s�"O���Z�=��ݳ�$'����"O�I��ȹLZ�9�?*;92 "Or)ᆋ$y�n8!�Rr��P5"Ol@ ��.��ĪV���F����"O~�##-�=$���Bi)&����1"O$$�%W6?(�a���H�C�p�5"O��!4ҫ ��)D� D�5"Ort�1K[��*l�"�v��)�v"OZ<`U(gE&��f�B�p��� �"Op�����3<�q���M1;�6�"O�(��U�d6�$r�}�"Oې�� �b�ҐB��C��(�"Oh�`��0�0�ӫJ��q�"O�`S Fh%���]+V�.	��jEJ�<��$��zd��螧~J��aT-�l�<)3����ѳ��V�(�9��@k�<�U�߅��=�g)��Ulr��Q�<��N����i2t)�8 �Ѐ1V�<	#�ޝ8����F�}���D�G}�'�F�*S���_�&�S���K�s�'T�%e�+,��9 �뎌@���Z�'�:�a��������%�h)Q�'g�M"�B*L�k��	��qk	�'$���-�=e���+bm����'�N8bnE(~z�T�W6(Ǥ���'�H�P��qb(I��	�&U�*�'Hڨ�ӳ +0��B/ݞ#bN$k�':J���Zz�-�L��$���''>0�C+V���h*��M�����'����	Ò�^���`�.8����'�^�I#��)x|B�dE�{$�s�'��A!���	tRj�q��0gJ59�'[�0�fۍ
���*]6_���b
�'���¶N�9Z$����C(\���	�'��)��Д>BL]���նC6�1J	�'�d4k�oR;_C��Y����'�p���'�X}��- ��J>o>� �.�y���x��#�`���$(Fn���yri[�BS��o�)�% ވ�y"]9
�qF_&��VK��y�ɓ�g�A�!�+0������y��A
���)���'�T�� �y�ɥv�8(���Mh�Ă��$�y2@��[��AF�E@�A����yBj]��&0�6!��:��I �̖��y"�e9K�h�$<�T�&	ف�4C�	�¨�+j�^đ��b�l���E&D�����ߴry2 @�Ø"P�b�ۢ�%D�ܹq���b����*p�8��&D�(�r.�bה
#f��	(D���#��&�����m�B�c8D��3F�14q`�1B.H<JV �kF�7D��Bϖ}�<�y��D:}c��B6D�(��L�)pB!���^#r��m���?D���iM9W��5f��>O�I��<D�T���B�#�� ��.3�	�Ī7D�� ���!d��kfA�
�CN���"O<k�dS��4��o�1i>��"OP��A
/6�����%8]05'"O����݅��i�p�l�:�k�"OЀ���U�b�00�߀@�x�{"Oq{��� n���b�
`�p]�"O���Ҹ!܈���"^�B���S"O����-�bA*�O��Dj��@"Ov����ɵ��I��2tS���f"O���vi�0��E�B��(-PX�"OH}�V��??#����W9j8��"O
�Ʉ�%�r�r�nҟ?�A��"O� ��Q7z�����F�0����"O��!k��u�.�ƃ�#C�b"O�,���=Pl�4�+:u��"O�PaF?3nh��v ^!=�N� "O\� ��0T��� �Aөp�حҶ"O�,[�K�,[!�>"����V"Ox=��ƞ�oĺ�򡝗h����"O�	I�M�,��� ��,.x�U�"O6d�P����� �86���`"O��Y���	�2`�B���!�l��q"O6����V����1��A) -q�"O�Ȑ ,����]3�o[����0"O(�Ks�O�tH|(��.��AX�"OfD��ؒ0'O�? $<��"O��ig�Y,Uo�����q��"O��������YR
4���b"O^�
W��������K��	(V"O-X�D�+U��yWKɧ_�ؤ�"OH���@Y=P8��g�XsJE�f"O�`��C�[�-������0"Od4�G����c��=UON��"O���/He���C��M��h"O��y��;�l�"����9Ժ��U"O��P���J���䞰O�f�K�"OΈ��e�}�1q�dV	Kt
��!"OD`�FZw�Ɛ2�"�/	SD�ӑ"O L� !��H���#'a�5G�Q2�"O62&͂�j-q���Z"��P "O�`Cb�Z�sL��Ac�';:�q0"O�D�F��'X(�j� �""����"On�*�O@��J]��R�tj��d"O�L�+|-�"`@˳_pZ�"O���jL8�Du �Ηhaji�g"O��ȁS�lP��ζ4Y��"OF@��W�1�E0n�iV"O贫S��/�6<x�#��bS�ّ`"O8��Ȭ=qh����	4J�!ɑ"Ot]���3o�"�s�^�*1�P9Q"O�p�R���?�����%Q�B�"O�蒈=l�}ze��9X:,�*"O&	J4h�+��p��Y�D�1) "Ony) "�+\�N����.FPQ�"O"9����U:M[�� �<��"Oн ť�:PU`�bͩ(���y�"O��R�d����]Z#Ӕ$˜�{�"O\|�I8Ԯ�����D��d��"O��8e������+�G���$I�"O�-��	�t�l�t�W�q���I6"OD�&	�<l��PD�B9�Y�'"O>ະ%ױ �L����ݳT0�hF"OU����:�ڵ�Ra�~:�m��"O
�!�	�N�8��!
��3�"O� z��Ыn�|�ׇ�h�0"O���#�"Q�"���/R�����"ORUiЌP�j) ق��p���r�"O��A��<����+�<��"O�y3�Z{ ��*�Iw���b"O��0�(�I~h�5��4~j5:�"O�X�M��N�	��� }���"O����hG,$m��I1O�i|b̑@"O��K#�]�]�z��-�*`��p��"O XsO>- �� � �|����#"O�h��fU�zd���³���Z�"O�U���Џ]���X�+I�dT)C"Oj��5�9M�`�)=@c�P;"O����̂G��,�(O�CfP""O�x�N�;�HHɂ)M�q3�m�"O5
c�Y36�L%��L�P# ���"O�H�5�3Y]�ݛ$Ȏ,^
����"O���P�1��!���?sb��$"O���o��;�H�C���<]�H�(S"O,���B&N�8�ň�:��L��"O|��W#���sE�ܧB�2Th�"Oh����Nd�[���%�ZXK�'fjqRC)�9X%���C�,]>$X��'->�C����'����韦}��p�'h���
�1��	�qc	!	N���'��0 �@iU�T���7e����'r��pc�$GofI������(�'j�4����AQ� h�����'Rp|�թ݂8y�Y!��	� �{�'[�%GM�3!�R��!��j����
�'�����ٟ��-�U*Z�*
�'Y�J��k�E�eK"ep�	
�'72��]�g���% Z���C	�')�X۴�	�*�����rςT�'n��@���V��D�� 8Z�'���e<5wVP�d�_/]�k�'x�<	��68��	�$j�-^�V�	�'ad`��Ȩs��fP�%Ɯ[�'좄@	�{PĊ��١#�� a�'�8P�d�C>�hdC� kR���'f<5)Q)�]c����L����)�'�bT(�ϗ!u Bm�d���=���'��`�,1Y���Ѻ<�0I��'c�l1�m՟K$����P��f;�'2�}�F�>���&��`<`�'Šq[.��*���b��~��<��'n�]���$th���E,p�|�k	�'����gƣn������<n�J�:	�'��A�a)�!wmZ���G�0gR�Q	�'����D�� Δ���HN�'��|q�'&�6��D�LK��[?���[1"O�m遦9�)�H��o�`m��"O�)�B�)z���+%���� "OV����U!�>�P�iY J����"O* �7~��Gn����j�"O��� �9����"W����"O\�# �L��`��)�yE"O�)2d.�%�E��(3v�R"OvL0��Y"C� ��W Y��l�V"O�д%�0�0�����F�lAP"O.1����ƄI���X3�"On�0���Jy����'O�g��b�"O،��ƌ�#�լ=�\ 2�"Oԡ+2��'ep}�C�0<���j�"O� N���1O:��k�D_�p5"O�8�6l��x0�A�$ �ZA>q9�"Oڹ��G�g��p�U�_�%�Xy"O�$B�L�?e.��#�!�  �\�$"O��)3�ss*L� �J�62�"O^4� b:���6B�"s���
"O��@�U�O�LT3r��8v� ��"OnP�mَ��PBc$�¨��"ON���֩V9�X��� ,~D٩b"OF����ίw�0�����p|�HF"O~A�b�!�ܑy�A��~��a"OؼpS�ݟy�lX{U >|v9��"OTQ�sK�m@2�zR�V�P]HAkV"O.�D��6t��N�	P�lȱ"O�yHpJ�xs�l�d�ֈ9�"O.{�jͻ(�bE#'�4vB�"O�Ea��@7cp���T&�nU�2�"O�9�����'Vd�`үԈ 7:�"O��.�)�L�[CiU�$v\)F"O�x��L"[;~����]�	FYR&"O��Cq�������Y��LY"O�0�!�Satz��	�S��""O%	'-��Nz��⣅��*��&"OF=H��I��}閤���U�"O�0�7+����ꃭ�4�`D�u"Oи��H�&�8s#g�,X�K�"Oj 
!��x��s4f�T�,9��"O�#gZ�_�hYg��m�4\;q"O<�"�\)o�X@�e��=%�|c"O�m����0T�qۥ����`(r�"O�5k��ß`����|�4���"OR����E7I�}��ɰR�Փ�"O�J1`�_z�ٛ�J
)-ef�f"O���� ����+��)��E��"O��@#�[+,��j��Nn����"O2���,�]F`�"'��6:Y�E"O���a��*:�=���Ȯ3��l�"O��#a��F�4�Se[$_��Ȃ0"ODL˥BҜ¸y@��?Qfix"O*�ithP�MM yi�"�G*0:2"O��K@M�sl�R`Ź!�n�I�"Op�{S���$^�[��J-,��S�"O�p�b膡$�l�*��
+!���"O,X�u-�=a�`zt-�.��l9C"O�x�G���pxR��0��q#�"O"`�wP0 0�[`�E�Z� "O���ƃ5VW��	�Ԏ0����T"O�����`�"���B{$^}R6"OT��Ҧ�=3���)�H� ��"OV%�'C��i���S�.q��"OΠk�`ל\P�{���
���Q"O��B�ȟ/W�Є��� ��<2�"O��2nY9���H࣎;.f����"O�pd#��/1�<��֮/(��R"O��Zu�N�J�Y���A���ʣ"Ol�:���}�h��,�b>�j�"O��J�*n{H�c�LN�Р�"O<aAT*Go���%���!��U"OxY�w�k
�\+q �-'}�#"O2�D��)\Ǫ���N�]Jٰ�"Oz���*E0up�b��F�3�<�"OJ�ye.��3~�"�����<�U"OIyG΃n��أ0�\'l;nD
�"O21��l�V�����v\(�"O� ��²���9��T �	6��@"Oz9��d �e��Di��H�U*tE0"O6-��"׸7������]�@�bř�"ON�Ӷ�E������F~T¡"O*8Z���`��5�!� {h�8 "O�۳�{��I�#KF�]q�
�"OJ b�W:h�=���;��u�g"O�U@cG#AT򼪢��&/��@�"OraDSθ�ä��� �p"OP�� W�L�D��7|�ԡ3 "O5�&��Ol�ѱeB�Z���"O~����G1� M[��R�:\��"OXj���/�D���$	x�8�
%"O��iW�D�(��v�C� K��P"O�<:����z�p�іC�P)����"Oz%��� �k$���p"6��"Ox��G��%'4xhJ�l��%
�5�E"O(Q��g��N�I"��Ş�Q��"O|ٚb�D	�p@�a_��L�#"O�M8�'ޗU� R��J�X~l\B�"O��(��7o�"��'J�ojB�"O����b n	���yg��J�"O��:$�PA�썊T��-(]��H@"Ox1�w�V<oK`]��EKL�}�V"O��aY�@3�ԉ��� -�I3�"O�Y�c�ǨP��Ţ�{�=��"O����)[�WѦ}+��̓G�U��"O�a� H�W����ǆ������"O ��`I���er&kY�\I���"Ov�k�n�d���`ιqD��W"Odm����0EbI@o�'=�q��"O4u�b[ �Q�W�<@��"O>��f\�&_�uIG7]%�D9�"OJ�u���hZ�S&�>hl9�"O�����дv|T���ބs�E:4"O�#@S�V6��U䚪\�!��"O^(�e��, $�lڇ"]�Elّc"O�)q���ˆ�㖡I/��<�#"O�ʖ��1w��E���n���C"O8����'��*U&^��L�f"O�X�e��w~�{��x~�q"O�������0iQE*͐|��X�"O��	�N�'��9�G�El�li4"O���D�R�Pq�� WRZ��4"O�<[&Q0 �X���:���a"O0y���5mz���eZ�9C8��"O�$�F��-�Zdj����o2��"O�pKP+x��Y���:K�=�"O䠀�K'9�x�3��'-<�1�"O~ 3�j�-iPؐ��גV&b�H�"Oґ��h5So�M Cm��` "O�p'I=	��hS�G 1�ڰ��"OL�S��0�N�;�DZ�K��dR"O&A
s�/n(q��C���A�"O�PRgj�6%��ش�]-Q�<}p�"O�J�c^5~�ha;� @9(�����"O��dJ�=-"���N�c��[e"O�QZ��� z�*s�Ĝd�9j""O��C�L��+�xPBlCLe� �"O�-"4�ڋ?��]���ܒSb2]��"O�jE��m8i���kM��0"O�A��Ǘd�J�e���hAK&"Od��D�B��>aQ։ƨ)À�e"O�T)�ݗVJh��*$&�d�u"O� t(���/s�}���	@F]��"Of�;�D�sl�ᚅ盔;X����"O�!u���y�\�+s�u<���"O��at��85 ���qM��!�"Opx3���GN���g%\�_�qb"OT��H7ڬP�'�M�K��"O�U#j� �"ɩ�lY2l8�!�R"ON�	 i�!k�v�yҋ�.l/��"O0v�̕9�v�j��9�PJ"O��I� �5Vs�(��J��nI8`"O��A��$d��!�**D@H�"O��
sg��!�H������[�"O�c��9��
�O\�X��"Oxx����(��1�ۂ=��"O��0#��B�8Ŭ�4^�dL��"O(L� ���8���@���07�|Ź"O|`I��۪GLX	��AI���q"O6lQ�))PM��l��AA�l��"O�и��P5{�������K!f���"O���!� �g����ۚy��y��"O`T��`ˆ��pcg��mк"O��:�!S��zM�s��ΰhKR"OL�)Ц�"�8����M���;�"O������ 4�\��� .���ä"O�d{���\N�qU��Txn�� "OT�"�JN��(x`��	�2��"O����ϞiO��a)YXP��&"O�DЃݞξ��Ei�Yf"Oles̈�z
"�Zp�MV�E"O��C����Kgɒ�<��"O�u)�\;����!M�8su"OT%�@�ߌx"�u�eO�WE�ų�"OX��@�8��l�L�1���"O�8��*�E�e@�)2��"O�I��I�C������ਈ:@"Oʰ!!��(/x��J7-��0�"O�=祔����
�#$�[�"O��eJ<t�p�*2G�0N�@!r"O�����\��CF�<[k �h�"O�����_Y��Щ�d>(j~8��"O� �o�xV1a��+z�}A�"Oԑ:e㈅Y�XE�P��zm��*d"Om����(â%�)Q����T"O��P7UǊ0�V'�G����"OXт��Hv<e!0A�?BY��q"O�u@�)�3� i[�F_(vL���"Oq�mݚG	���u�(1����"O�m���KsK��:�B�"{��X�"OlA���t���a�'����"O��B��XU(ယ���K�"O��A����(�����a�4-h�d"O�(�/�7��YH��Uq�"O`�v���!.HiR���T�R���"O����̹GX���j�#+�nx��"O��
��p6��z�ǂ�! ��ZC"O�`"��X�+���Q5���s��	�"ORE{G�=�pbB�'�p�p"O~��i�7Yβ�8mW-.�ƕi�"OFģW�1�ñˈ/OV|5"O8��r��c-4|�"�	Tn-ڤ"O��
s��}�r��	 `pl�U"O,$c�ܵ'�H ğ�EF���"O��f�Џ[f�sfB�iP�P"O\H�'��j	��JNX�Tb$"O� �Q���^��e@�h��L���e"O��p$�C�#G��y8����"O�x�#Ӈ7X����I@U1��"O(f-��<��!��l�Lr5x2"O����6�^�9W���g=|�!�"OT��ꀂ*t#�K	�8�<���"O�y��pa
�0rē�N�
MS�"O��i-?	�X���(@2�!��"O���5������u�� ����"Or�a�畜�:<�֊�6��x��"OTd*B�Z >���hO?"��r "Ot��RA�8�p������L�v"O�A3ck�*x0T�� ��`�
��"O�Q(��'
��u:��"S�-��"O�����@�H��f#Ə|:�]z�"OT�(BB�a�r9xf�� E��C"O,��F�6h]�$
�24$�9�"O2�[ӥ��?1��H  �H�0Zv"Ov-I{dqJ�EUX�tG"O���o2w�H�95���3"OH`f�D�	 3�$Y���"O)� βk?H�r�BA#���2"O�EC�ō�I��4�#dT���L�c"ObE���U&gvAR���<��|�"O��Y��?=pt94&�U�4:T"O>��E4�@��7��A��I	�"OБ92䈳B)�U�f��'��"O�Ձ�=c��3��6���a�"O܍0�$L�Nn��i7�y�(��"Oڹ��Lٸu���1NE�r�:,QW"O�0
���1�|����S�u�"O:E�3FR.G�i�T�W��!��"OlM��)ǁx��q�A�3߶1б"O�H �P�d~��ǅ[8Q:��@"O4�X�j�-\\��Rd�q�juk"O�"�_'b�$�S�#�,v��]k�"O�P�dJ�N'�xQ��	�
X��"O2��U���h�ׂׂ;8�@	Q"O���T�_�b�l|�r�p{���u"O��#&韼~)I 皛dQԬ��"Ot����<>48x�7#�xX��"O��ժ@:Ϟ9K�$��m���jC"O�`��%�X�
�#̷Sqҕ+�"O�9*sCߞ�>�+�"֘�d�
"O1zs��E��X6'�[�`��2"O|5(��%7��H�a���[�0"7"O�$`��T�U��'fɪ"'��b�"OL��@O߬pR�E�0 �v"O��+�ȅj���`p$�,<��s"O���AewC����>���A"O`\;�� "#�͙�/�;��X��"Ot��Ǩ�q�������,��"Od�����L.ƭ�&J��D���"O�T�%I̴j,�%+&��i���A"O4�R0�ɰV�cf䀦	�B��"O�	`��3��R$�&*����"O����k¢Z�@���ωH�"O���L�)8][��A ��tJf"On@�r-�=3�i�_���=�R"O"�;V��0_3.�زDK%)��� �"O��Q󉉮7[�yC^_@����t�<�Va��L3�T0s�I_ep�P��n�<p%"C������x85zWp�<)଒�L��8���XFp�Q,Oh�<� �k��9~_���޹+�&��"Oz��ĢD+:���Aޫ#�*��"O���p�r�ju
N�����"O�hj�aY�n�� ��GV��y�"O�$Z��R���2��	�/�V4�S"O,ث2JL91Pvs�F=:�ZA��"Ov�]G��ǋF1P��d�c"OQ�t�G�o�|���Dxڼ�e"O�с$M-w~�|���@C���Q"O*�[#��B�.�3�m�&2Ȱ��"Oҁ8EQ+ �6}`B����B"Ov�@%�m4��C��3IP�P"O~��e�V�	P)�eH�z�α)�"O���t� �Wg�������ְc"O�9b�KS!7���UZ?!�N�Q�"O��k� ��X��K�*��Z���B�"Or�� ����Dj�	 ��u"O���Bώ)K��4	ύ$,��"O���0�ڕg.̀�(
���,h�"O�-l��p��HК����D�d�<Y̚ ��0�쇎#D��,�c�<�"e@b�95�G�\�d�3��`�<q��	EF2\��S�Şd�<q���b^
ݲd�ŝ;T�[Udb�<au� 0=��=�֥Y<�4슑g�d�<���N��̙��Tl^6,SF�E�<�׫��V�$���Z�6�,	�Dg�B�<��DF P2@�˖Gk��Z�e�s�<��m��ki�t�C�P7.wҝB�IH�<�+�,L�cw0G�F��ƌL�<I0���@R�)4��#��H�<�4MI���<��HN!X�N�B�J�<���T e���&Op�\�/I�<AA
ʰ>Ev=P���O�u	�*�E�<	���v
Rx�,$({4)Y�)�j�<��3jZ��P�Q��䡳^�<1��I�	���!B��aU9;�\�<�(��iPC�O�:�*���Z�<�$�ؓ]�\�p�B��#[Pջ�ņ[�<�b��}u,�bc�L�D����d̓U�<4�;�(�pr�LiF^hs��
M�<IE�*�0����J
�ۗ�q�<iR ^/Tfjh�@�D�z!i�o�l�<���5XM򝱃KȉoԀ�`�j�<�C��l��1�#	e�I@��Lf�<!��"�:�R�(��MX) �Eb�<ׂ���!mJ����k�C]`�<ɤ�K�8�@[e kb���^�<IG��%���c@ f��Yk��Z�<!7m2PD���C�;��P���m�<Qц@1�R)�)U�Dpz�r��O�<Q�aU@G��s��I�q@�	%D�0xs�W8���so�TW��b#!D�xV�ҢA��!FɦcQd��/�y�k�G�XD��+��u�Ȩ�yB@�DT�k�"E� �p��G"�y��ɗQ.�C�݄G�f�a���y₄�,��h`�ٞO��Ӆ*��y�I\�L+l�x`��N"iS5�Q��y��ν���K���C�H�a��X
�y�m��7�|azԢБn4)��`
��y�c�>�Lu)%�N)5�4Dbq��y�MN�@UB��/�6+�@�"���yR�@  ���4`^�*�RԨ��Þ�y
� ^����J#�Ñ�A<Y�6E��"O��s �Ο+��؈���B����U"O�٣�"ͤ ɠ`�6Dؐhju"O2���ʖ ���OLŬ	�*O
Qi �W7�<����`8�m1�'X�C�AF��S�ذ.�~��'"O��@V�q�L�*��]E�<�F"O*Q���T26�ԸF�áf>"X�"O@��3FY�l\�u���>3]+0"O@%pU��b�^<	�1(��&"O�0�� ��8_�t9A�	
%>0y`"O����4�@����~	�(�"O.� ��K
#�����P�^��"O�\8���c����Dj	b��SU"O�1�,P*U(%�'�?o�,�T"O`8o��:���k��j�"O�d�� ���R���ϔ_���B�"O*��MV/\��e�EDR��>�jF"O�y���/*�P�B&G:Lg ��"O��p�G�~��ő	E���`"Oj [����Bf��"�%W�@5�)H�"O�z�.�=u�"�8kI�:v��"O��;�k��A	��Hd@�"O$���ͪCJ�m8FlW� p�y�"O�s�m�<z�ȣ�L�Z��#"O��zlC��@���G�{�iC�"O�06��U�.H;Qh^&��t�"O��&�	X�w`�MQ�v"O�\7L� ����i��CW
$�"OְX7f]�NBJXq�J˥l$�9�"Oh�qTÇ����ƈ�V储` "OV��A� �,�e" �u�2H�S"O�s �kG�i� (	.!��!�"OPP+�O�'f����g(G�ƠC�"O�!$���U3��c��ϯ���"OZU��gƳT�R�2��L�vnr��"O��eȜP4��A��6^�P� "O�YI��g+�jc�9�l��P"OE�3�Wx�z)��d��mF��q"O&+f@Θ:�B@k�B�f�v��"O��8��,C���fH�^���pe"Od�B8� 4���6�u:@"O�i`&����N��]�h��"O�dr�--wf|���C	.��$"O��ztO�a*"h�eKĸ/��(�"OTpag�;+����`L"�Dm�6"O�Ir�o��,��lJ�X���#$"O�,���Cj2-�� i�UAW"O�4��P#~��L��ST��){4"O��1E�6� ���B�|����U"ORв�Ӡdo�T�'䖪.���aw"O�`q6�Qɖ�c#�J�-I�"O�Qq��Y,h�(1�p�]�c󼬈"O��q��s�t��DZ@=	�"O�Xr^�XIJ��BRl��,��"O����jU��r���f���hAq"O*��)�BG�<z�FA�uԖ<�'"O��)殁��.��օF�g����"O��ɲ��.B�Ge�&T�
��U"O"���L# `>Zdb�B� �9$"O��v���cQ���/�lb���"O��`e	R1:�h�-���@�W"O����WKY��bt�M~��"O$ar��ѱIO�qi�.#@��J�"O� x���'�lD�P�B%���"ON]X�A��k_�u���8t���"O�buAY�P_�90�V�4���B"O��9��'-0H�����`���"O�1�󉐆B�̀�pO�ZwZ�! "OЗ�Dd `��.Y���L�ó�y�)��\pB�IGm�#�(���R�yb(�4&��-��7)ZH"v�)�y��Z0;�8
�i�!ò雴B��yb"M��DhrQ�G3H9 ����Ǩ�y��^ ����W�8�@���y2dGF�vMJ�[ZFY��P��y�#C�U�<�9f�7P�BURs��.�y"�ĔE/,}��3An@[!����y�c �����;�>��CV�y�����>��O8ز���&�yR�B�]j*X�eI�4(-���yB��bɸ��BG"2R�E:R$�$�y�%��D�¬0è�0W
	�q�1�yb B2C�1$y��Ј9� ��ȓi� ��B�6u�t�@ԩ^\&���ȓo��C�&�Ak69FӠ�p��{�N�+����|M��]V���Y�F�*q��> XК�Π
����ȓ1������m�p���o����ȓ@<��rIM0��gψ�l���Y����.K/l4Pc�
�.uNT�ȓ)G�A2@��0RtzL�RC^Pm�ȓ9�x聐"���,;�͒�Y�@�ȓ�B����o�aȐ*ʊ8��$�TeaS�]1�Jh�5�S��ȓm����E^�2��D34�ʕ�U�ȓR��*�l��T���vn�
Q�ȓ%�����X���y����Oa�هȓ.z܋t
�V�0�72�������ثK�����6?\=�ȓ!��" [�-h|��G�S2�|���&2��p1d&0Y8�qGgI2#������L�A2N%1 r���)_T��k� (������$ �AC��ȓ3

����U4��l�ºӂa�ȓl����
J�y����-.e�̈́�)�ȁ����zcd��i��Gct��ȓ%�v���A��A��qX�}�ȓf� e{��ڣ7u>���n5l�ry��hPs�%M�k�Nl�Q��6V\����vrv����8 �h|h���g�ąȓ{U.�B� ��L0H�����3I���X�� �F��0ܢs� �E ���>x���F؁0huJ��͊(��m��c�����u��Ub�DM!
�м��xoL4�@����-2v��}��a�ȓ4� �r�[z�fZEO�o�� ߮�kpND�|}{ᧇ-^�Hp��SV5�Qg�qfN�x��t�y�<a`�̺0�H��	�%K����z�<ᗋL�I���E�E.1d�D��B�<��4W�b�(�Dk�8�s-HF�<Q2b<����f�*q�m�<�$E�B�@��C�ջX�Q�2B�<�iV�t"8����=d���r�Xv�<���)"(1�Ю�;32�A�r�<��i��Q���ʴ9�JV�Lo�<y��	}�p�;�.[��m��i�k�<� �ȲEO3,a��l� �*2"OجH$�P8xa"���Q$d�j�i�"O��kWd]�dZ�9����3E�Zt"O\1xE�]��;��6d��<�"O $���/7�U3'�ř)E�y*r"O)Rv(F�(��%���	 PC�؁�"O���Т	8M�F\ ����1�<P��"O�	�)E���zg��� ���"O��	Gj�Y���i�/DV���"Oje��)U+Z*� 9��Dܒ��"O�PV ,!�|���F�-9 ʀZ�"O$�C���K0�jҦ��$��"O<y+���uK��/�#��Ac""OL��R/ɼs�M"s/9#���3A"O��cJL�:_�����[B�[ "O�캓��x��k��Ɵ7�yp"Od,FN�c��1A��{��e"O�3���#�F�3�ǘW��1 g"Oڭ`̗�\x�M�����`�,��"OF��3˵4?������|�&���"On��T�Q-M�$c'!U?Az��� "OZ����,aVQ��!�uq��"O޴QP��!M.�p�N¾+��r�"O�58��8=��|P`NT}�e�"O��bpl��<6�\sG�07Xޜ{�"O��Sց�!X��u��M�r'��"O���f�˾1((%+P,���I�"Or�;5�N�m.�I�J �;��"O��:C��v~��`VD\6 �5�D"OҼz�'I=%�h3�V+Q��t""O��-Q6\t���!E�C��P"O>�֯3ԅz`*�b�z�hF"O<���'���iEIW08վL["O�����T~�̂���L谭�"O�ؙ �V�<O04��ȟ��@5Z"O0�c�¨��X��)%�bT��"O�f�:m�0C�P b
��"O���M��� �sLL�5��<#�"O������ed�qXA&E-(����"O�]CH�$W��:�䁌HD���"O�p�D�������Cχ~ 
-��"O�e����hHe�.���0�"O�%��V'xx��Ɨ�l�7"O��It��4�P�V�HL��"O�5xFn޳G�UP�$��.
�.�!�d��3�D�H�Z=3,D���+,�!�+4�r$r3g�
B� {'뚙Z!��t����O�gv����q.!򄂣Xa
�k��s��ɴ��.%!�䍠-�D��V�z��h�%(�&!!�����X��{3V���ޝq�!��VQRVѫ�ݵ.+^xI���N�!���F2�ek����NwF�б��A�!��; ����,O",v��#WI�!���]�vH�c��
B��:u!���a��) ��Q9A���"G�R�!�$�G�`Ej�jɝ9��X�'Z�v!��הe��
�ΐ�=�B��FömL!�DJ;��a��M�8��b�[%5K!��
/]��{b�	yr�w�U�c�!��O�D�0�\4�B� ����!�$]s�0=`�DFV�bw�,M�!�ā0)�4{4G&@�$���u�!���"�Xdkċ?0�5��/�9t�!�� ���`� �fԒQ�TP I�"O4� E*M� �D�0��^T�E��"O>�a��[�*��ț5M�%vP�5Xw"Ob��膢G�\��q��Z �Tp"OZ����^	"f,��a�_� ���"O<�c2�G�J ��@ƙ�x
,0��"O�%s�J�X� <�U۳{"�"O8�0Un�`_�$MүB|��"OR��"/��o�`P��
��pr""O�A󀭎:S��Mn�/��e�"Ol<��N��B8#vǎ)�~=Q0"O�Y� ���,��Dl�-3^�R4"O2Dp2ѰS�xE��>:+��@"O�<�VIE;P8��j��S7)p]�"O�Ԫ0Ĕ�|8n�ҴO��ou�@"O�u���̜:��<��I�:��C"OБEE�G������ELr�z�"O>��MpW�$���Տv�Ʊ�"O]Ƅ٨9��b!^�_lE�"O��s�����C��.]Pl�6"O<p��K�0+q��[sab���"O� �a��7p�<��U\ *0"O�	�Х8^3�X�@�߲l�^��"O 0���� @�2R&˝+ E�F"OP)�M̡!��yF�TX*�I"O��3q�B��p�p#d'C�`S"OZ� 1��]C ]y���z���s"O�iH��V,/8j`+�@�n�0���"Ol���bЀЧD���&eڥ"O� I(��_�����S�=2��"O~y�P�Ȅ&xj���bʡ~�d#C"O�`ea��X�H����|mL��"OP99��&�]�!O?X�g"O�Í��N���
��jF��2"O��\iz"�Z��)(i΀+r"O�a����\�i 'N*uQ���"O�<;W#�
���sgfӓ�!ч"Oz��g�}�V�SW���Z�"OX��g̀�Po�;a$_:�>�Z�"O�Qس.R��z�)�9L�ʜA�"O�B�K��H"@�x�	��ꘪ�"O�`����iܤJ��^�a^���d"O�t(.�,u,�AF�At@ {f"Op���yI��@�� +o~�؆"O iӰau�~$[&��	XwD�
"O�H���E���[ k٠A	��̥w�!�L79Y�h�%#ƨB�zxУGʧT6!�$�uL�MJg.�$?��ᒰ�C&/!�$�u�0\X�J�?z�i�M�
=�!�$�,��(�n���*��ސp~!�D�:!�ڥRD�� $�  X �A$u�!�$�& ���+�^U0��&c�A�!�93��]a��TI��e��gQ!�R=UۜͰ�#OR,��Z�(E!�I_�9�󋘘Q%�p`���,!�d�,4{��x�'�8i	���.�!�dѡ2�@I���ǔd���á��!��A�z��b��L�q��
nB!�Ӯe����I	�"�Ɗ�H>!��4nQ��s�!S?��-h���h�!�I�l�eH�@E*�1O�8�!���.)���Sƃ*E�h)Tn�+"�!�dA'7"��X/?(Le{խ)d�!���)��la�"{�|!rgH��!�� �h�初�^�&<���]lL�W"O���Ƭ��P�<�1G��/bFq�p"O��k a�/�n�!�f�Ld�Pr"O��+�c�Vi`50�e΍l��y��"O��R��[�V�H�5�ȫ(��1�"Oh�0��@c��#`BYY���	F"OVHf��@����j\����"O�3'�Q��V�{�c%��t�5"O@(Ҧ(�gD`����(L����"O�Bw��;06�h���� �t�C�"O��!Ѭ�&:��ʔkV�'g�@7"O����"�-� 놝nG4��"O�m II0T5pԻ��QC*�`"O��`�Y&���sp+�6x.z�!�$_:,4��5펄@��$�`�p�!�dø5��S%*���P�OF�Z�!�$�]�
��!�D5)��5���
�!�D�_�
$qg�����,	5�!�DҪf,գ�	�L��=R�+�)F!��wL��X!��z�$5bӨ[)3!򄄥Μ�@"� O�ZqԇP��!�D�(LPa�j��2D�ci�.(�!򄕤g��(��C^f�A���S !���l8�������$t�!��>bDzГ�L�f�uJV
�/b�!�Dŗft�Q6i�<8L�h/s�!�D����ٰR�R�G��N�!�$̓#�H3CA+o �m��B�!�d OvI�%���$�RdD�u�!�$ɵ&�|�K�87�j	��R��!��KW�V5["��p�H��"�O�!�λ}��i�%7v��ϡ�!�d�5��<y6�H/c
Hдm��-�!�d 9P����]���Ʀ�k�!� �yK�DëG����[�!�$	-4|�|���	�Ȕ|����<,�!�G�-O��s�_�K��h�3@̗y�!�$�*]�4�郋��eɂ�E2B�!��Z�D�9�tK=7�)�0kL�x�!�dA�.u��B�^�HJ��p!���hآd
@$�7>Š)��e�I�!�DP�o~�Y$�G����	�+U�!�d�9G�� � 	8���1U�D�@!��\�VX��G��(,I�b	~�!�D?��`����|����ٕ!�T��p�TD�?d�]�.X<a)!�$� |sE�M�8����g��!��t��v�� ��	�H�3 �!��̑bA���P`����xM�!!���'^0��D��
��E�"?�!�E�{
pdr�ԇ�����L�!�dK�b���S�(	���C�a�!�Ć$294yP�κ�"�
��B�!򄄪>�Z��(N;B��!P3&N���'@nKvA���ؓ��U�/Tbԇ���%0��F�b1�pb�@XX���9�����J�'��Պ9[�����:����&���F�C?\5.ф�50.=o�
^��{�Nθv�P��'ٞYQpmKU�xp�]6g�@q{�'x�!؇gF2Z>��P#�\�<��'\ �R�NA)�I�0` �v�'��$S荥oj�@p�!~� `"�'�芷�2H�����R~�ry���� � B�ĲP݂�H�Ԩy��`��"O,�sCl)�d!s�h�\��٦"O�mq�ל>JX�u��4-F��:v"Otx���R�z��,S�&�3b�qI�"OjwI�-o�X�c�J�����"O4�SvC�@TQ�%�t'�!��"OK�RR��!�::~j�� ��y�9&f,�
�H�>b�h�ZP/��yg�&,$�D�T����`G��y2=}�} �΋9`�����K��yC�A.|����Y�p�կ�y��'E�V�8�ƀ�;�҈��m��y��Y%,�V��bF'�h�J�y�l0^����VD(\֬��N��y�Q�U��zN|�Y����yBE�/^x��Q�\��Ґ��'Ĩ�yRK�8g����pk�hѲ�y�ę��y�5m�z,H#ǩ1����%�'�y��%��1���I� (CR2�y҉�3i��u��$ [6��V-ސ�y2�\A+�gޤz��4J��Y
�y��ªg�h��쌌nSIz�A�"�y�f��t�$|#G�X&�q�U,.�y��J9ni��*4Dau�ě�+L��y"AI+gj�%� �\̦��1���yR#9��I'�V�L1�aj?�yb�8> qc2�I�^~P���l��ybhQ0'�����[�W�S����y2M�]�^�����('D� c��=�y��%F�#өT�F��5gP3K9!�$x����a�D�}Ĩ�n!�D�xv��a��H�^	J\21H��S!��vM�`%J�m0����F;p�!�
4AD�˖"2�P���FVX!�\9:mH�����f|SR�82l!��0�.��w �8���3ņ,$]!�$�,{g�N��\��c�{P!�D>Yߌ��#/1��q��#F!�دW`"�GS/b/j�ꣃӐ0!��	�N&�3gV-�m��P��!��#0�0��X�_�����i�
�!�$��.\ђB��L���$��G�!�$7mh����a�4\݉2��I�!�$�rOHa��#n�I!K�\�!�DU�'�"L��Ç�d2@y!�d]�'�yu��=(�Tq�!�X+!���#5��!�"T#~�R�+g��+�!�	�v&Jd�p/ڙ)�p��f��!�D�4X�aб��s�(d'؉\!�d//T�0&��6?6\)U��/b�!�d��x��5�j��E��`Z�FN*P!����[�+ܝfn����Ee0!�dĴ9��t{��	`��s��U!�߄?Ò��� ?z١�LT ~�!�䋢NS�q��/t&DEZ�,S:�!��'1�xlq�W.���,
`�!�I�.Dh�2��Y��Q"v-�
%�!����-�&�67���pMe!�$ҵE��H�#��&�\sS4=�!�'~�e(�W�x�[���Q�!�D��7<��V� uq�=��(W3r!��d���H�$Pjb����E� `!�;	�� ��X�d\�iX�#,(iџ,G�D��7s<��q���,�P����y
� 
���.�"Bab��S�Q�S"O�؁��Z;�NT�#4�Y5"O��
���q����
ݠbf"O&�;��- 8��E9ª�0�"O�aꓭ��V�BA�r#?D̙�F"O�� ��T�tLc�B�d*��"O���S/�=T��e)�+��A	�@z`"O��s��9�	J#+�M�=i��D8|O�q1l�(B�ܵ��)�L���"On	�Ɖ��[�D���-�+��E�E"O|�#ef�x���d�Z8��U@�"�c������D f4$��Q#}�$�Z �O0#+!��J�� �G�
�J( �m̮!��M��M��NP|�����	ؼ>����D"�D$ �R �ѯ�`܉��Y�V�!�Q�,���-�|�Ö;G�'��L�S�'�*����.Hm���!B)d=�ȓ� ��=8�|��Νd�=��It�42�D��Ō�h�B� a�'W�C�>�0�b�͉�i������m���<���T>�k�.��X*��FməA�J]��:D�@�Ë���@
�)	�wj%s5+D��� h�����V��"�-D�@�)��m���)ڭp����$d�O�B�	
9X�-ȴP�l~4�bu�Q?[�B䉷��)�D�|���*�B.jB��h����ܐ(��:B�I5)����U��"�=�W�ZB�I�;��P�D����z�O,3Y ꓡp?��K4"^,�I3%�2F[v�10�E�<�@��U�"�h�-B	f�
2�Z�<ѕ'�5<����U*H�L���Y�<����@�΁��&@05��;Q��[؟�2�'JN� 1ϭO�����̌�p(J�"+Oң=q��D
PCN���k�$��@af���Q�QN>�M?1:'�I�v��j�n�>̖(9�9D�8�W$�x��;$ �X���;��#D��q`�Ц+[F C��D2�M��$D��b� �?Y;�)��A�*u���0$"D�T� �I�yD����N:��c�#D���kD�[� �ˣ��d��!�4H#D�,�Q�� a�Ւ�����y��&#D����L6ͦ��'eU�m���;��6D��`�
Tk�8�D�n�Y��8D�hӕ��O>�A
!c&Zf���6D��
V瓄,��I��(��B�$4D�(p��)�"U~��g�0D�L�C$24��+�4���V/D����܇�����ODF��!vA!D��1d`�8rW�<Xg&�,z��0�A?D����M�/r��@g�<^���s��;D��Nѕ\58��	�v�N��CH8D�Ԩ�!Ǜe=R�!$���8�Z�4�3D��*��m�jE�Dd�.����n�<y,�/=����T.U���k�F[��ў"~�	�W�~�k��P�RxJ�q�lXj/B���0ړA�H��K7+����c�������hIb�	�\��ZSs/ X�<�ȓL���g�&Zǰ��3���*��ȓ@H�%H�� C�l�A��)�����H��ͪ��2cfi���;���ȓn��y�R�6R��4��8����w���P�A�8�ر5q��E~��S`h�YQ��O�~x�0O^��C�)� ���2���@��m �aŢ��"O�Es2�	(=���M��S�6'"O�(�b�X���쇖3��YS�x�',9 w�Ԓ���P�E��\k*u"�'��Hi1B�M�|�а�-O>&`�ٴ-��<E��4]��b�@?@�̥��gK#1xZ��	t��^��)��V5�5E��l��?v���D=hQbsU�[��Yr���Nx�$�'�
��O��B���� cքq��1�	�'#�Q�*��>f��d��{������6,O69q��I���(� S�J��%��'��~,F@B�@�F��\��B/���'dҰGy��遨-�a�H�$��=f+��<��x��ɺv��	�֡�35Le{$�,\�H�O����?(�t���GS�6�����`ٛd""B�ɝ�#˞�1\�	���"<�
�Z`��i��׶zX��9f�� d��'��}�®'�j�`��-Wfi)a��y�m��`nt9f@-`0�Y����yl�8d)�K��F1 v (�b��y�/E�V[�x��A�;��0A+���yB'P�6n�#D�
��ɪp��6�y��)z�6 C�l�tĘ�J�/��D2�O�к��Da4M��M­A��W"O��Gc��,)	���=9�2A""O��鳆A��6(��� v�L�ʁ"O��@��l5�1h�aˍ=�JU�D"O"��ąA�q�Y�AA��/5ޙ*"O�8H�H��A��%O�b4���"OX�ĥ�|SЉ GY*���Ȕ"ORX��	�U���̕�B�*p�"O�\
� �b�H�1g
�hל=H"OF=Q�k�<!�̰
��8�B}1QcTF?��Mc �{�<E~2$`�p�����<� ���G�Px�A�',�� �at��aD�4�j-x�O> �E�P�V��9��K�+<3(!�b�|"�D�O�b?qRd�S�0dlL ��љ�N�{ֈ)D��9�N%w!P�;�L�!�6D��&D��q�����B�6͈&7�T�E$D����+�Ls������
�M !D�h�2���VF��HFO�@�C#9D��c!�R8:���qs.��c�7D����Ņ66�L(P��]���k7�II����;��]Iw��x�h��W�BC��1O��!�7�]=U*���$�x�&C��=�D0ZR�
�l�n���ټ/��B�ɠ:����(��W,D����$u�C�$ȁӀ�m��:��(C��C�	.<��Uk�
٨���i0g�2B��&�&u�����R���`B�I�(k.I*�ϕ'WI�;���8��C䉐"�l�֤ՠ�	&W=*�C�']#,���C�p��ÚL�zC�5���CX�<�sa	�<C�	�+�~5`�LKY��ɔ�pB���%�G�֍��Ig4�B�"O�M�e��E�[T�3j� �B�"ON5��R'����N�2�"O�|�W. M\h͡T�ϭ6D����"O�U�D�Gyt���ϓx��J�"O �K0(-I&ƴ�T~���Ȱ"O9�n�,M��`� �� 7_ܳ�"ON�h�F�0y_:��fX9{���7"O@���ݥXdb��&r����6"O� ^5����U�)���ӔB��;�"O���4/�bHUc�YҨ-��"O�;�L���ED�4Ĥyr"Oέ!�&�zP$X�s`H�H�r�0v"Oݰ�e�9�d�u.�.A��	3"ON5��ā�NL�R�H/�PI�"O��qJ�]�6I� P/M�L͂V"O =�D��2l��-kR�&�T��"O�ͪPg���䉉W�˴:�,��"O�)���I'@4�fi���<���"O��GVM����sM�4Ќȑ"O��*�ĉ�4�`��˂�,�8[`"Ov�Je,�aޤX� X�$��1"O֕"�h��)�6q�F���Y��"OP��nME'<@�]7mv ,{�"O�]P�k�*"��� �
O 7�T<c"O"�hRf�%w����J��p����"O���a���[�bL1!�(=��!s"O"�P��	�3��A�I)Yr4"O"=C'��=I�xjeʣ�P��"O� �PdS�m:F�rV � �DX�f"Ol� QD�+:Q��h��+�D�S"On|�-@�Z�^<!�f�%V���H"OZi:��ůd�*sU3)$X�Z��䔰.+F�"AT%D�26N��1Oٹ#4&HtS�	Wtpu�b"O(=�0���UM>�8��b��D
P"Obʁ˄�e똀�0I�6�$�"On�zk�0�x34GH�>A�"O�պc�֞L>���%�?��E;�"OԵ�1nE�yD���c�;�F��S"O���ӂ�5���0��(L��l!Q"O���OC�L��%�6`�y�0t��"OȨ;��A |����R�U���q"O�D�Q	�̹���*��L�"O��N��_�z�ٕ�F��X�g"O��3�N��#�,$&	ԫ�0m�t"O^0`Cl֗1��<S3�Lr؄��"O�a��4��0����KRP���"O4�ٓ�9���rm>(\�0A�"O�t;P�P4|L���f+^G�*p"O�d�˚�:G�`����9��KB"O豺���9 A�˅W�N �B"On��'M8X��a�)2'�B�A"O�K��ĕ3��q��b�N��"Ot�P剋RȢ��'	8��(R'"O0�6e�B�p�J��j����"O�6(5y����[/1�^S"O�xKq�:"�v%+t��W��u�"Of�i��6:�6�1!cۗL��aٖ"O��j��=��a($j�"O���L	5<PҠg��B�Q"O<4bECQ��İ�O=����"O��篁�V�@0����:���q"O�{���z>H����5��8"O���Pn_�8����1[�^躥"O�`�A��70���{��L�e�n��b"O>��&�K9B(h�HE���h�����"OH�sf��>s�X*��.q\�%{�"O���f'�Q��K5?Ox\�'"O�ҶfƊes�t�F�J�<#BUi3"O(M�`�Ń@?��Y`*''X=��"O���WDA4�b��'i�,+XH" "O��+�%#+��N��9/���'r\�K7��Qsn",)~@��@X����S�? �Ms��L�o��x��L�Ea����"O�sdk�9��Y)��J-��:Q"ONE��ɏ�J@
Yʐ���t���S"OV�c�˄u0�eZ�"Whm�`'"O^��E5ܔ��a Ğ{0`�B"On��B摮�"��"��M����"ON�����t4����� ���sU"O@5��%T>n�f����`���3�S�O���a���X0�d�"Sv&B�I8I^�i�Ɋ"�rPД��7��<q�j}�x��f�\����҉��*���ȓA2H�$�Ҕ������ٵ#�`OB 2%J�!dQ�=`�jũ=�B8� �'�b�;CD��:�b�fI�nXBQ�%&D�4 uböds���!��#(B����g3�#�HO1��e����S	�U�v���)P��"O�݋0Ƒ�|�b�2"��3+���AW����K�<��>���I�Kc��xVᎃIc�u�`��!
��B�I�r�����;�q�e��"�H}y�OF-��+����<�w�.P���"e_�~"P����h����O����֯t�d�A��-�ZQ%J5b}ȕR�'ڥ4 �
�J,C�m]w���y�=?iW˃5J�?U@bD �;Z��y�ˤuH���Ю1D��Q�F?t���?]�!� �>	�#�}[��DI|~J|�'��Q�rM̮��� �拈gl��
�'�\h�2M�%:����׻~�B�K��%?) #�.t�T��)Nւ����5\��aN�-fQaz�+}2��OԲ�Q( �XHP!a��ܠ��'"O��aP(J�=I�ؓ!�[�_�" �����Y���O�QG��4�����"�:��'�t\� �6;�m	���vo��8����pX�0�` U=(��j0#�"7}b�h�l3D��[�@��7 ���
%�cԉ>��C�	�i��a���J�����1x���2��$y`�\�D�2�j�P�o�&w|!��	.�����D5�D��!c�qO��=%?=��&�3^�2�ա��&�"aK2D�0B�/\�v�*�ψ�I:|P$7D���ӵ4��SU�	�Y�����><O
�Cu��� [��'|���@�4����%	�o�P���'�>�3�N�=!~�����!o
`E�N<�5���A�ЪTMRg�O�]�R�?m���#jS�eD�	�'���	�)ަnװ�kPG�.�X��0���*�>��K�?U�>�>�OTe��.T�v���٦��o��9'OPi��N�>
n�'�,n��DC�OI]��� ցy5B����'���AW�U�6 �&�o��I��$��Q<Z���YK�a�g-��?qiD%T�9�F�pM̹��H=D��y�&3z�J\�FNC6x�Q���<!A��8	[�����ޠrgе���>ҧ$쪑��! ���G	�6Q�
M��>�4MہN iY���j�0 @�̈C�6�����m�,[��O�3�	D��ٺ��,ڌ����ց_ ��DG����bo�3*v��2�e�-O����R��(��۲��.6Q���T�'e�����Bk;�����+�J���FN��@�D�A2��!d���}mnj�Hܭ%��yR1̘)�4�@&�`}���`�`D	�ř3�q����l�>�O��X9��sG�6�*��_\y"OݝMB,��J�x~&�ە�Vv�1�8ዥI�v*Y0��&F�z�����PPw��<qR���E��|�1����O�$R�/�W�ֱ�#h�4 �J���务B��59����9�"X;���}Q��O��U�ک�c�B�"�\��W��#F�0ՊQ	C�}3�a�GB�I�qT�Ӭ�:���'D:݊A�d8��I�)l�\�e�bhHTF �]�&����%Z"f�2��D�c,-�u	��X�e�k��J�_g8�X��	���1e�E��0<)��F<F|�PdnX�]#ʹUȁ�
���JA��;h�<A a#Ϋ$%�4� H^� Ԩ�6�R�8�B�"K 	���Ba�M;i�:Q#�) ,��`�i�Y�,�*"�p�І�	X�(�N�T��a�*��%(���3`��a5D��/ܠAK ��	�_D��a7�XI�5J�lW����!d�ːtՀ���`�!1�`y�P힙A�Ez�	�\��CR��7
,@��)�1w�z-�u�]�!LJ,1� ��I�R�ɖ _ ��#�$��2"P���㕈6� LY�C٣*�����E�HcUf�C5���(�@8��H�a�  Ӆ�	Z�D3�C&�(qNC�_��h�E�c:\9�C��$�;'h��M_Zl� ��4�F�5�Щ
(���I�j2�y"�(	<0��#l?�, #J�_�l� �W���풂yt�����
�h%�;�&1�W��.X�HCp ^^���GSf�nZ2���R�	�;}����.���O�����χ�k���R����S�ȉ<��px ���M3�cF�n�P"I�4㼌	��K*=��	���(�0�.
V%��JA�ڜBΑ��8�@F�
F|q����Y��+p��
7~HӐ$֤~�	�E`H>�~�P#�4�~���,��k =.�g����%js�A'*֘)iI��u���kbX��'�Mo�r��%+Ӥy%�	�1mГ����NW�[�6E�g��	Γ���R1�V'J�X�c�[""�,�a��
n��(���[�DԘECS!�\ܓjͦ���c.}��$G܌i�AƟ13��T`L	0�����U�wxL�B�Ƈ٦�a�'s
�걮O�X���@��k-I���(�U�̌5��IQ�}��\�W�Ƙ=@Q����ʷ	�<	u���-3tT��%6������V^ݙB�ǤB�詫pmLF<�8�b,@��THGn8��4CM .�����p�J�Ӏ�-ғlnT���0	#��r �0^y��%��!Z(>5��BX/ �F=�E�[<WL9��2(��ΓYv��o)F�H���ᘉl�^@��� �✨����ж�ɶD,4��stFX{>O���B��]�v��$�P����{rX�a���i`@�4k]2��'�P`ʖ��"�l�BA��F��F�|aA�%�a����.}��K�(��i�+=ڀ�OU�
���?v>�yu�&N����_�%��u,�$38 X�O�= ���d�*�qa���l̘5��p�Z.Obe	Wk�=�j��b�X'+
,��a�t��}�Ë�O�}��A��^du9'kߔ8�pċ�#�.0����w�����[�&(<�4A�|�q�a [���Ұb�J*�����D�=pf�1\h�)���d�0��Ύ���T�&\�o@�E8f��m���@(��_n�9�Ƥ�f�(0�f��@}�N�S��b�ég�ơ�8S�� 5K@i�'����X }�]��.?y+�3XyQPAA& �ȲfU�w���cT�92��
-h^EbǬ_>BI	��&��Ɣ&�y������)܌����T'���8 ��%�êH��ɰA1�ӧ}\�l�0�E����a$i�?��� LD#l!R��@�D��M�k���^��"����ԉ�8����\��C�g�Uy�X�pA��,;p!CY�"t2h�g
�� ��c 9��)�V~�t���̓*1l9aټ#p8�У��[=< �.+��Ѳ$�:�he�U������i.Od�D{�Î,Yz�\�VG�X�J��#kS� ��ݚ%gO�my)��Ȕ�b�R�p��CG
5;�
��
�]�$`��:|�p���ȇbT�zv@ʼVJ$(�s��([�tD|"��Q�l�w
�w�du�'?�L�0*�Mi�f��{u��{&C�'��ĳd���n���G�X�b9�T�P�>Om �VL@�x}���w�~4�q�5D�X�v闏u��M�� -.��Yk���5>m� �^.����o[�~��aj�F/K�,�%BZ�(�@��Q`�جL�:<�E�Z�*�����(�%��W�p�N�G�1Y"��2.��Je�@�Z�д��!L��XAm����2�f"ҊQR$X�\�r�`J�J���� iU��W�H�P$!�a��zڈ �v%
yg����ɑF/z��W��K �ɐchњ�u��"G�~ ���D�<������:+`����H�N�7�#7<�'&�@�a�).N�BS���]�R8��I(,H�Zc��\��	��\]fC�k�,���-��r�Ni+l�e?|tҶ��ل�B�mT��ZMF�O�"��MI*w�@�x��I*v���j.��z��)7Q42���ԛ)��L��R�¨5S�NĦ|�����jF Q	5)`�G�]���ݡ-�v0ՠ>h�"a��J���R
�A�'�r�6]lX]8����ER�{��
�,%n�#�L�ufP}��+Y�2�� Lav�A�TR(s�nIz7�@����Y�G��N�$���G><&mzlR3}�.��r9:[d��#�il�e2OUr[@�gJ�B0��%e�RQh�'ps��<Y���G*@�S��L�4!2�`B�%r|�	�hB8ۜ"tLQ�,�P:��X��,��!C�A�"M��S��ĺ˶� `���bq0�QG�լb`�0��B��k��뉘&K��8��'���D��5�&M�SL�64&��Wd5Y�|�H�>Oдy�xA~\�e�'=VT�a�H�z�r�HjP�x�}"b��U8�O��jG�)��@ӠÜ/���REfNR��V�58B�I8]X�q��9�Z�Ʌ.Z=}�^C�ɇ2b�q�Ǽ[�2��͚�E��C䉶/,Fz�O���P�MU� ��C�i�Lq�:��ؒ�	
?���)�'���*�Lӆy|�����)��
�'��	&� �4��\�"]�a��'ژ%���[/c�X��Ed��M��Q
�'�� ��"�� k�#K=�F�`
�'4����iA��@ �Ǉ{�Z�']0ya� �k��\)G�N������'m
a��0j��(��PzÔY�'�6�K5�ˮg���2 N+��\��'�$H'C� I����mJ(	�i
�'�<�1Cj̠D���$N��L�R�'ꬕ��-V�pZ|���	�rŠ�'}ԩ��a(\��J4*Ê?J�Q�
��� ${DA�~`��e�R�d�<°"O�L�oΝV\0�A�'/����`"O��:6GE�.�P�qd�;k�&�ʃ"O�,r�G�E;L�`잸+��Ŋ"O��8"���D����v�N�;�и"Or)cd���^�FA�@&��v�$�P&"O��b�?�P�b�O� Tl�f"Ob�2s���Fr¯�|NZ���"O���!͔��֡���9<^���"O�x�IB1�dX��'3"��"O�����up2�@�LW�o�(Q�"O6�[u����⃊ͅn�t �"OF������)��j_N7
ɈP"O"��BH�*l��p�'�?��"O���b�A�6�Q��<i:ʨ@�"O� zb�S�ޜI�5�ɏ��� "O�X����;s�zh8�bܸ�:���"O�	��׀{���c��G�ܐ��"O��ҷ�2�JغaN
�B}�p"O�ec'�S�3t(aYFtp�-�d"Or�k��
0�`�d=s�m#�"O��y�EC�+ӢEBh��o��)�"O��vF�j ����VgD��PP"O����D[�=Pb�Xn�t�"O��se��L�AƘ�ؑ��"Oޤ�FŖTm��I�nP;�JA��"O�K�bW�s��x��j�
����"O��ӳO4K+ٱؔO�2���"O�T��k�A�b��!���`q"O@`��PIPe�rl;����"O��p�"�/>*�:��[J���"O
0#�H��)��Myi��3�8ѓ"O�)�6J��5;L1����/1��A"O�m��߹FKr�A�UF��I�"O�)r�F�h����R��I �hF"O�"��Q�!��0����0mL��w"O"��͘�(�U5}�T��5"O�������ÇG��Vu��"O|u��`ˆ"����K4P0�"OF؆����B��ˠgX��"O֔���x����A���6P�5)�"O.yC�F>3J�� ƽ3�r�q�"Or�0���:Gg|�J�����\q"O.9��[
tv�Eͅ�#"���"O�Ii��[8k�~��q&Q)W�"OhˢiOV���kĥ�~���F"OZ��t#�:�y��DA�5�}"Ob�Y���5N�q3��a� 8�u"O�᧧
�眘ʧ��ߜ��"O�cc熢.���+��É Xe٣"O|�q����"�>���O�
4�q��"O, ѓe�6<�8]�3B��!"*��"O�)�/ÑZB�aZdc�^��
�"O�T�pa�,wV1�b�
�6@d)""O( ��)Q;w��*��zCZ��q"O����V�$e���AL1Q�|��q"O����mH�E[� �.{����p"O�`(�k��	h��_l�!"O��3��&�ޘ8�n^>:��"O"4�T�O�A2��HG,] k�J��"O�%�'L^�1�h�k�j�a�"O�RqΖ9�Ji ��-k�@�#�"O���t.D���d��'Pe+2"O���㘮0Q��t�
�BL�0
�"O� �X#pB��.Q��W�j0���"O}*k��j�N�ɢN�
#���t"O�%3�cS(^�м���Z��6"O����Y�7v*a�W-ϼ>�)�"O��` E9y(JG��*�"O������Ts���$Bp\���(�yR�E�N߰�iFm o,�;�
���yR�L��Cvg�&"����F)�y2�`+<�5+�'�P�`lU�y�e�>�0dC: �l,Ƞ��4�y�&��T�Ґ��o�����:0⟙�y��jL�J�+�(����͓��y��O<>�A)�xъf��T�<y�7[ ����T2 ����̓u�<i�ȀM/p�	@�ȭ(E
��g�v�<�t��^$���[�:�0T��z�<��I����ZSn[&����\�<��b�+z� kPQ�"0�� �Ȇp�<�N�MS {�AG�C�QP��z�<�����.\�� h��ᦃ�<��ȑ7o}����)Ze��( iPz�<Y4���N��Z��O`T Tu�<�qQ�m]$�р��#b��Y��\d�<�S�Ԟ��y)#!�R�S�Ȁy�<Q�C�5d�B�A5
Ԛ�Xu3�(�{�<�����i����s�J����R&�S�<��-ӿ#Xɪ����ET($hu��M�<���W�$�(��[vO� Y�n�N�<�S)7n]	�����z����EW�<p�ʾT�P��1B��<Nx��V�<	��R[����CT}(���AUW�<$L�:�z=¶"j�n��DDX�<�@ʫ19*R��n� �C�#q�<IJ����"�H��"TԨ���{�<�#°_��K����7�콓5�Oo�<�1�FI�����4�Xā��d�<��ߏ]���(�AF��Gl�e�<��b�Ny>M���*q���Ir�e�<	�����i����$:0�(jCg�<Ɂ+��u�rX)#,U��	&P\�<�	��~
~}3��	�B��!1F�Z�<�x(�e�Ժ.����uŕQ�<)D�A>7֐yif���'1`��#�Lx�|aF� �&3d�(O���GBS�H�����6��U3r"O�5)�ݸ��������_.���f�x�g�11�T0!A�P��ȟ��P/rp\��V�͒Q�"Oj��!	�S��.Ja h��@�5�H��Or]*S������}��ɰq�=E���� ��Ȕt��|����Bމ}��x�&K��'����GnB.m&��gKH�k�����Y���5��
HY�k\�R/N�?CLV�"JA�DĬuF� �O��]sWb��i��=��Ξ=���{�'ޜ����0t���{�X)	8=�,O�U˃�.f�2<�D蒵d�.p���	�x���Bs�����BB��,�!�P8 �[R��
d�z�ԠC�O����O;&��H*�C,�����{2�ɂrr�j��6S:��������?yv!	���A��?5���{]pD���[���9fM�0���C%�t��a�iʃSa
��CIT8~����%#4��(B�a�ΦV����S@p�b�����BdĔ>j�9C��%��ɐ"!��Aӭ�<�t,�}��L����nϮ��v��<���j��Q&�IY��i���(b�X��U��h4��|���۲q�mI����B��T�ּ?���c`�Ui���	5h��Ӊ�u��>9C�	�@�zi{�fR�������;4[��`t��4dn�y1ʙ>�|���
A�pqK��Q���P��91R�����U;uo|�^`�X�/Z�iz��ʠjݻ5=���$ح��]:S��M!�`�%NغK^LS���'7>p̹ĂH�^k�d�5V=�qR��H)�H��J^HC���0����
����C)D�"���'�ND���O�J�	�.]RPc
� �pK��ݕ }�����D,H�4�H�.�M)��عY�N�BĢT�Nφx[��]���ӕ�կ@%Z�۴�������C�Ua�}`�)��3� ���#}��S
`�%S�q�.X ���<�07��lP��wo�����x�����W�7�L�y��;J:ո��ьk�h�"��rd򤻴�9_.2 IT��	+���A�ηv������C���2	P��xkwJ
8\(< ���-���(�4q��N�
||�Y�L&rIx}1s.ʑ ��a�g�S�K��&��|R*�ZMv]*1$)]a6���Q��e�5��Fx��u�Ӭ����^�\OvY:��p��T���E{H���E{(t���M����u䍸hR����1L����ń�;o]����X��(+�`��T:�剓���t5^̓��1���E+����W�I����Ҧ�Y��F��q��z
���!
_.�MK�_�I�j���J�h���[P�I�K�d��s����%\�~���_<�Ժ�DX릵�ǁ/Gp�x�E(<�V����H:;z�Z� QTڼ���D+o����ӧ���HO�T��M�`<�A�O�>
*�lk7�_#��p6��r����0�
5rȤ`�5�L?�7G�O��SEî6^��5#�-JG��0䬗s`d�Y���X9RĊD$.�O���0	ۅߦU���ϩg= ���@[���E8�-�
���b��r�扴	%��I��1������JV q%���-J��e��hדe�bE��c�} dqp$�8&��d[�cUqF��&�_�q!�7T��?9bN�5[�
�;�9vAZ�f�)%�t�լ�<@�X�s��Z�ͪg0r�Ƶ��Z>x�\��=�V���g������%ߞ�#��T�j���;��.s�x�@���q�r��F��5�ᰆ�A���mc�Fj+ЕC�#_o��8`.=�%tJ��-y�X3���f�!x"G��g�W:j����NG�5�٣�A/wSvŰ�'�p�H�4#yR!P����[�	K7_�:;d�ȶq�,]�Q!�O����1R�|�qaP1T�F	�Fk��d=sŨF��oZ(`�l�V�b��,�R�X5���w�6|H;N����*y��p҅�'�V�#�DS/ ��bDdрo�48r��[Ԡͣ$I�@�O�Ȃ�_'NQ:DXB��{ �7I�l��e�,O�!X��$ �6D����=��L"T剤B�1h��ڦ%�,p�JU���pZ�@�RW����#�;-
&��!� Pl��j~6���r���0\i��ר}���?�Pc�l��p�
R�XZ��5F��<نNށT�4��u�@�Yl��蠃�k��9u*S9[S��'�6����2O��u�ݧ�����8	�������pK��{�a�;v���#�f�-ddJEpG�80h��/?dn��b��vF��ƹt��VFL�bkT�]�fM��˒-4�J���M|���$��J'�ڲgY;��e��Ӥ1������כ,~��Cn]�i�0Y"�蘊Ab��b�����Y��i'6����)O�c�_�l₁�G�%h0P���	|��S��_�Q��m���OD�ޤ�H��~Q���tn��x��8�p�V�Iz� w&]|hM���D�nSL�[�΀�?M����-��	�C���
F��&��c��ȈK�D�x�x	 kù*1�Q)#/�<Q@�!�p��;l��\2q+��1�	�'���K��i!TAp7H
�1�v�c�N���m���p���z3�F9S����q�k%RIxȊ*2�d��w�.A 3BJ����,S���'�(Q+v��7K�e2C�i�j�3�-�E��|CD��T>z�����t�K�2@�Ij�#�o�tO�5�G쓻(2�9KȤn*~A����1M��0D��%�����)y�-˦��yFAkg�/G���
j�Bҗ��w4X�b�>��<AF۫IB�sρ�@���Q�O}2�~0):�o!�r�KM'	.���ߴD
��)�탵Ș-g��q�'��K����"O,Q` �����z爽UF����� ����٪`z��kU$��Kh.�O��4�G��3���]C�4|���oIظZ�i���$ ?��A �oS�u��E�`a�Z�-�(�Rћ��}Q��!�/Q�EP@ˬW� �F|2��{����J;U��XQ��V���O��FB�;�j�*<��%LM�����w �%>��&h�8~
X!�IOU�	�Δ��@�I��$�)��
��)�'N���!�;=̦X�u,�dMnA���
I���K|j��D�;�0�;���*�.\IĀ_�<iP�Ex��h�K��6qx�"�ږ�M��ϑK~���f�/\A�D�J|·O��]���B1f��A^�Ct R�/+m$��ɒC5`���2Z)�e�ׂ��6r�#�	�%ϓ.>H�!���2��Ʉ�	�jL�L�%��>���
^����Ǘ-�9q�M�(E >��׫��G��e`Ql��?�6��n�ca��C�*̉CA@	��T�ȓ ������V�Xbl���9/���ȓiR=`Ŗ0��9� I�	��q� (�ᛯb����k��% ���2�`�`�I�mq����=m�B5�ȓx9�5[�L�40��	�&�[�:U6-�ȓc��=��¡+d�b���~e�ɄȓJ�T�AG��z<z�i6$�0G��	��U`\�2Q`@�H��e�5"�*e���ȓK
<�EN֊�����E��Te�a��P�0�����r/
@���nP	pd�8s��T�7]v]��S�? Z�JP���i��bO׮Ȕ��"OH�S	̜��]��.�9A����D"O,��*�f���C5���i�"ON5ڄ��*��p����^e�(ӳ"O*�kRI��$���N? f`$�"OX]�cЎ"�����[�"ք�b"O�Qs�I�+ER�KF�m&�y�B"O���� X086P�+��F|ڸ�$"OԹ�#ąw�d��l�Of���"O쐒�kD�+ZL����yF �C�"O~y��)
�V��1Bj�hK��b�"O��z��F ^�Q=NȀ�P"O�{�k��EPp	�3��*Q*>��"O����NZ#�$���b,>��"O,��C�	 \B�9W���\	ڸ�#"O�����ؓ)�R�@�m
ڬ���"O�F ��~`�����U�r�U"O�1fyk����e��ѩ��^�!��Mh�̈�GA�JT�I	ui�!��!��d�7�Ԇ{_�9�dgK!kR!��3�N��ㆫع�g�5$!�H� @m�3D�>%�Z@����	�!�ș5��U �.�m����K m�!������3I�^���q4
S3�!򄑉= Pi����a*�(�\�!��IL}���<ml^�+@�R�:!�$�6.��K���
I���ńB�Y�!�MSf�Y'ΏR��`F�%K�!�Dɤ
K�8��d��!㄀��k�-Qv!��6r�A� 
5��ғ`
�f~!���/\V�K��S4�2���Н|�!�dЁ�29������9��K	��c��&��
�5B�A��@���3õ>Y���O��jWAӱ����fD��P:���Ԏ������<�����. �d�ы>}0x ����۲�'������?�WM���Y���ԟ@�X���or�T�#G�;.r��3.�����'8 �y��W��Ov�'d88�Ze�r.x�0	�"��I�S��{у�!XI�o.�矌ap�	�j���נdiȄ�ql���0�V>�z	B��>��M�|�w�E�Hr2Ŋ!���@��uA�h�x�X��4�c��O�?�3Q�ފC��!#�	\ޜ�s�ź�0��9��%���p$l��|�Pà�'\���a���	�O���#�p {��ĢXE�j[4+���Ě>��g�6hW�9�xJ|j�'���1ҏ[,	�J�2�K�y_�E��O`MxD
թ^k���|n:�ӈ<�b�I���y�a���]@7�,=�01�>	�'i�*}(e��!�&�0��|�a���RwŤO6ʬ��O����\#����bР���H�8�<���y�hU78�>��=%>�R�՝M��t��S<��pw/0�$I&x38)�{*���(쀥&�Zc�UB�V�6��'�����RJ�S�Ow�D9A�K����Ӯ��[u}��4(&jq�3�1�)�'T>���f��E�<�3��'!IPK�c:Z`�'C���'05�9x��ٚx��b�/�N�8,	K<�զ��uPJ~�)�	U�w�ȩ�n�~��x9q���S��d�w�j�Sv�	���S�O���2���}�b�R-Q\����4S'ބ��o�Pˢ!��Oeh6�y��Z�+O��;G�./X2tٖHT.U��@Rp��0s�N���m�F��i�&
㞄�b���z�6̣����4h� �'�ܣ�K���O� �B�L�0"�����7u#���'ʆ+2���~�ͅ��$����Y� z����Pu@C�,{Htk��_`�<i�M�B����B�
�Ā��nD]�<i��F��\���b�x�}Ĉ�c�<��l�0\�rB�W���q2�	[�<Y����Z��U���-��5q`�S�<I���0p2�+Gf] �"��	�L�<�G��L����ղ["x"4��}�<�劌�|��1!͈50��X�FPw�<)fP4� ʰL��B�6 �$Yt�<� ���`'�)6ݱ"7���C�"O����h9zغ�9�!J30�`T�u"O�!����dn2EӃb6(�&��0"O�أG��i�l32�Jg�y��"O�(B���%X�=YƠݹx}*��"O\hkG�L�����Yl�A�"O,����2f�W*m3��Z3"O���0!ܛA��;���=5\x!S"O$�sRϐ�/��)F�̉):���"O��H�mJTqd0Bj�J�*Oi���A-����Ҥ�6�0��'�z8�@A>�:Yx%�[Z��
�'����p�6_�z����8f5
��	�'j��i#C^�"�$`	�'I�[����' �8��8}�� ʀ� d�a�'��˓/.er�����%�FS�<�R M�4��0���.��a��N�<)e��#C�<��Uj
<j���`�GJ�<�R)I�i�m����P��b��I�<�叙��q�"�5u�u��@~�<�Ӄ�I}n����%z`��Op�<1�ն�B�(����l�lȡBMp�<� $ p�8s�.B�r�NdᒅZU�<���]T�N����^�=��IMQ�<����u��A3���s��� IQ�<I�C�3m\ɂ!i�9*lpR�P�<�HW]�C�a�"���NJ�<���<}9kC��g�j��U~�<� /�9BIQ �?{7�5��ƕD�<��Ѝ>'8�p���T�9� �J�<YPP�ߺ�����7H�M�ȓ(P��UNW��z{P��F�^Q��9T�'L�'��z�C�	?�I�ȓ]�2��!B�MS	�����QMtl�RE�0j=�e�To�E��X�ȓV=��p���s�"�R�2���ȓqI�XZS��  &*aj׃ٓIj ��ȓ?p�1�Ń�%�2e��AD�]��{�� ��H֫`�4���FbBL��tuę�퉮Vg���D��

�d͇ȓ:whER�hY.~n6�`�M�b����5�r}q��6XS����F&r��ȓKa|���BF?@��*#�?�8؄��ne����-WԠz���?k�8D�ȓ6�a��D�L��!��.1Z ����ͪԙ!�	7zo,�I��߬Ax�%�ȓst ��D�t*^�����mTH��"��Z�MB�r��RQ(����ȇ�6h�i��#=�}뛎k�\��~�tb��D	-�5�@撥��ȓҰh37͓�x�
�CaU�����ȓhđ($�_3�QB��GE����JD��Y�&س������%�hd���l����]�j�b�k%ѕ/�N�ȓ����t$B�84��1"C͏.����; b�zA�S΄!�I}P܄��B�-�B@�*1���G��Gb�}�ȓl�	;�Nf�yL^��Gm�<9�]�^sR��&��%N�Ȩ�	�l�<)�H4N݆�8�` b���d�r�<yu�_������W2`��-�U�<YǊd����	ljX�� T�/SrB�	"2��RC�	:b7����ꑫ[�B��bu�s��G�N|jU	s��y��C�)� \|�C��&U|��SD�8ξ�"OXQ����C��0	��ǟ�t�#"Oh�uB�/��8��$5�
�÷"O�	�AN;G�r��hΫ?X���"O�Ĉ`@܁E����e�16"RA��"O� ��Y�ؽ�0N˪l�fy��"O8�S�
<��"� �L�hy��"OB*�'��dFJL��ʛ�O�b��"ONe�7��<0>>�g������b"O��ȒKU-�͑�e�:��"Oe���R�2����/�ei�"O�u��F��f���s���Z��+"O��*čƄ4�#`G�B���D"O���ɞ.>]���!�<A� ���"OP��q��bd�yz�@B:O����C"O( ��Ǔ�0�<S1������3"O�@�&���c���_��u �"OV��H��4'@A�`d
�ܾTA�"O���r�[�N�2T��
����25"O��I�R��A���"Or�z�쁄o\�- ��*��� �"O�Y���f�M�c���9pА"Oب��IPWH]�ԃ�� 	�""O�X�Fa��S�d8y$#׷u�d%��"OZ� D��)v�֕H�bP8pꤔ�R"O0ݹ��τX�h������K�"O���@�:��12�m� x��*"ODsŎG&?����w� ��Y
6"OJ��U�ȫV�X�t��24�6���"O��k���~V�1i�@!I��*�"OF8W�B�tMԙp"��
�j�[�"On��%��/J�YpnJ�����"O��9��)HRE�a������"O�d fl�/s���;#D#�J "O>�A���D�I�g��3�RUk"O��'J��ƀ�4������	�"O��;�)�"a�>�ym�[�����"O��[%D�.hV��k�>��q�"O �ф��.2��H�6�P�!�Pã"OJ����:������ZQڜ��"O��5eͯ1�j�1�m�$}A H�D"O���`�[#^�v�q���6;Q��R"Oέ���"F��R�F(D�rT"O�U[P�(�M��W1t��"O,T8��^?W��⑯�&!.��"O��;1j�P ��S�>1�L+"O�]��F�A��9���.��\��"O�ya��DN$q0j�Q �P"O���W�譛���2>�$��"O�8�#*�#l:�8&��֔J6"OĘ��!g<�Q��8�Q��"O�y�'�Y&��H��k߹h����c"O"��uj�aʙ�Ԥʡ$��|��"Ot����<L��0�D�I�f�j&"O"�kեߟ<�Z4 B��$�F���"O�*�e�v�%������I�"O"�y@��#R�@� `Ã �jј "OD��A ˵Tz�	�5%�c���be"O�T���@(9Kd���[�*!�ն���BbO#u���ʥ,C�s�!��[>1��0�ubU-�*)B!�R�&�!����B ��b�����*�2�� "O0�2�eC�'���УJ�&({���r"ON�����kK�'뜮ix,P�!"O� |X�G��~�-�sǏ�P`��p"O�qa`F�ec�T���ܗ�d�"OB`�a
Nk����L��l��C"OXyx�+�S!�ȃE�$�\�BU"O�|$ ۶ U�i�qgāpN��q"O��vbȼq�n���OJ#�ج"O�QH�L�+t$�D�'�vdC�"O��R�P�f%
"T�$W�(8�"O`��ƤR�Z�6�s8�)#�"O���@�p��&&{j-6"�kD!�.*�6��� 
-P���f*W�~8!��O^�8���n�ͻ`j�jP!�d��N�LbGl<|�8����hc!��&�T�r@OȳH�Z��R�ʥg�!���m��Ā���AR2�����"<{!���(W�U�4	�Y<�\��7?r!�ԻF���u��>e/�Mi%��BR!�D�w6���R{@8�y6$͡h�!�D/2*��gI�!"|{�K�N�!�D�q��TPҨ���jӂ(T	!���L�&�8��ӓf<���ԏc�!�"9�<�u�C�oh,�%��1�!��6��}��4u�Lh�7M&�!�$B/�(#�)�%��bTi.}!�d�e���㑏S���'h!�9(*}��ℎ+�6��0�=/S!�ċ�Lb1ZC��	
��	 �L�iO!���z�:���F�]�ؑ�7,�5HC!�F�X��81��B<	|^4����-!��,s�8q����zi�4;ቝ��!��u�H���d��{����h7�!�$0K�\֍Ky��A���#!�dT�A�%��t��K��n�!��<�쌓��C'P�Z<z�A�;�!򄝝f�����)�j�b���~�!�)� ���ӰA�$�ȆK*S�!�ٳu����@R�Qs��K�J�F?!��ӑsH�q�C _XI)�N=-:!���9xU6ݣ��y~V�ZBmX&u0!�d	�X��H��R=R|�T;��
�D!�$�|`L�*h��H=0�r�lM2:!���m 0���]�4�Ċ	�p�!�$͜|
2�2a��sb�,kh�6�!�K��A����OH�ܺ歇�w�!��z�l<�CSGa~��*�)P�!�$�5.�j����@n�P��2T!�DN����f�P��(3�&�!�U!aRx{,��k��HP�*0 !�->�L��&B�t�K�)�r!�F�s���q�����X!�DE!?.�{�ҵ	MZ(U�ɟr�!�� b�ucE��#LE�1Y0a��u!���AH�`i#gR�V�7�	:	t!�Dʈ{���eL�m��a��#N�jr!�䙿"�$�������Ë)`!���q�3� E�ے]���^5[!�Dָ!�4��ᙈ`zRH�����D!�� @��	�DcE�)Rrh���3fS!�DM�5爥��A��:PUc�㎲,O!�Z��F%�7!Z����@�-�!���:� ����:=�|����^�!�D�b �  �`     s  +#  A.  v9  �D  8P  d[  af  mn  �t  �z  P�  ��  Ս  -�  o�  ��  ��  R�  ֳ  >�  ��   `� u�	����Zv)C�'ll\�0"Kz+�D������b���Q=�y����yb�҅w+BlyDn�?b�ҐY7�I�P 9i��!o�`bU��B��!��4!�Q&T*��	]�n����	o��D��΂�iOdM������sge��Y�гSgX���[����xf@�J�mڀOf�L �gW�T���!���i���A�)��CЍ�fiaK�t3��i�|���'���'���'X`��B��[���	OhِT����?YW�m盶�ק�R�'?�$b������'��A�>ٞ��2*�$(�`hq3M��q���'�&6��O���?a��뺃r�)+�z�P�gW;N��}@�BI�<�死v�؏%�x���O��$�h�Ì�dK<H��yx�'M�J�P���־gT�уµ>y�'��'h�D�Z��<&@O����	�H����kS�|3�K��?��?����?)��i���'��߼sf$C9r\�P�,�G�jR�I˟��޴��ja�ƜmZ՟�Z�4:����B�i��I҇�&$Á�Yq��b&��<���۷F�<�޴&����'j ˑ��q��j�dz���o��?!�Ȕ��Z(#u��o�x�#a ��(��²d�d$���צ-S�4����O��	��i�,2�%؅M����华5=d5J �-dZ����>P�@�1�G�FA��b���HQ��	�x6-���ڴר����ܟ^���%�=!����u��H���Qw��=����}ӶTo�|��3�ΞA���`��k�v �D�R�64����=p��PA&'�O�(�h�AC`&,|	�4fɛ�s�r�)��D0��SԆ����2KQ�9��AгhKZ�Z@O*7!�Q��&y�	"Um]+m h�&E�Հ +���O�H�D�җHzMჄI�H�L8���ʟ|�?y���?��O��F�'2,<x���a�ޓgu&$z�a�a���'R� X��'2�'z8��CɛVX��S"��q�Hh*�@)Q���A� L2]k��i b��(��(v
��(O��yF�)��4G�؊�H([�`1��eǞp���FgU3	��c��(K(�Px��Ċ�G��I���K�"��i���ҸG|$E�N�C��'���|b�'�rV��	.b,h�b�)C�\�2�	�U�̉�IΟ�ɓ$JObN�$�T�s��S��?�G�UZ�M��D��ZFD��Yޟԕ'��(��r���d/�Sݼ��#�R23�кL��HQ��ן��	$��1�,����h��	���Ю�'x�b�':q\;S��mR�e�V�]��s�W~`՝^uMX��O0>�ت`��V7X�q�#�F�)E=~��Q:�i��m�.#n����
Ҙ�����Y���v>H�l�9^��dg�;s`ne��?��Ox���O@"~���U�����&X�
3�G}�'��	v�Lan�L�	�6��H��CL���x�OB�e��c�4�?	-O,��P���v��O���<�! ��U�8�b�DO�PQW�Q�|QJp��zK��ʖ|���.�L�)Q:���O���b[�C{�tz��[!S$t
��T�`F|Y�'aż7?�	J�aK�T/1��C�F���~N!����-޸nHF��W�M�V�&	�<i�E����V�L>Ң�08�=�s@E�;����@���?���;¥�7n�\i��gɜF�i�lZ��M+�iyɧ�D�O��4A=����L�o�J�Q��q�T9�!��;�����ʟt��矸�Xw`��'��(�T����ӏ!� �JĊV|��qq%�L��}��N]�O%p��V��#p����$O�A����cH>�
3�J�Li֭�_e�*H��I�6��
�ށu��K�h/ʓw����C�ރ��i2'� 0`����������48����ExRJֿw�^DHċ	�8xpȥɱ���2�OE)��X}<x� [�.���  �|B�y�`ioZDyR�TB�7M�OF�d�6t�����
��]��AT(W>r���O�5�#��O^��O�ոR�T��jݠt{�<,pc  ���4K�R@x4�Vf��=�z����~�X�<����;f6��ؤ��#
�:[� �x�E�AŅ��}�1Cק^`��@A��=�X!�Q���<���I�Mc�i8�/N#%�$�e	����*��ꦝ�����?��}�	������jþ%z:�
��C����?�/��hӪ�A�TM�2#� 2����S.�Q��:�M�R�'b�R��6D����៴�oZ�?�Dm�j��U`p"R�?Lx��f	ϟ��	,H�!j��Z#H`��k��X���I�,/��z�͝-%�\!���� �Z�|(|ce�}R
)Sc�mi�i���]�S3���gGP����)Hl�]*R�ߤI�P3�~B�޿�?1�i~z� c>q��ǥN�<=�E�V&#\D�`�/���O8�Ov�D�Orʓ^́b�/�"����O�(�*��@�ɉ�?Q�4�?1ǾiA��Rڡ�H�L�JP16��97��O���O�����ǃ�&�D�O^���O6��M�ȡ,ܓ�d�A�o���؄����l���ю�M�CDWC��O�L�����
�~2��� b�rcN�Wb�y!�׸1S�8Q�J����q����M�နE/�ʧg
t� �ļK���>7cX�R�g[�,�Td�6��MC�\�hɧ��O8c>���O������ ���R��+B�F�?�f�O���$Y�}�$h�# eZr����7L��'6L6-�U$�0���?}�'��DK7�²o�r��%b@!n(5*���6]϶���'+��'�2�O���'�� -gJ̈�w�Zw�(��˳	|ęp��jhfE0���=~<�C��3��=�2T P�ڀ[�h��A��gb�e�2I@e
�+݂p8�ʍ�C&����g��<j�j���d����aL�$&8XBi�"��u��H�����M�'4�,���CF���+�gn�c�.D�<���@�+V^��Ī�=@Ph���0�D¦���gy��&r�6��ON��ČR�%2���SON�;���7�$���OR	!d�O�d�Om{d��)e�+f͏��8P)�=� �+*� JO����.F[ܱ�D&�8BՐ�ӏ�� K+V��t{<HG���p����,� g�,��Ɛ�oG��@2D���L�hO�E�'��7�U�4,�4�������e9qS��u�IBy��?������$u
�9r�~(P�&%�IN�����i�T�#�c<6���Y�,�.*:Rh��.d�H�>c��@ٴ�?Q�����G2:{��ć��.E8Ӄ�:
/rM�LĐ6A����OH���ڟᘔhR!W�5�N�����a�4�?a�FK�z<^\y�mX�X�&�,?!���^R!�ϔ��(!u����OM�#`�[���I�� ��5H���OLq�$�'�R�ڟ�2@Z_�P$�R�"f-"�)Z�<�w4RN�����F�>ZԨ�G�_R�'/��}Z��4װ=׮S��L����Mk����1E8���O��$�Ob˓ ͸����%NXxz�.��}'�Ȱ��߸X;Pњ�g֠�C�$���i�\�B��	�$͒>	%�.J�r���6G� �p�Ή@��u�E�(_�K�C	0b�ʧ�ذ��U��C"�)&p�"'BP�Ye"hh�@ˉ�M��]��2��O���7&���%�T|X|���:Jr��qEm��d��ey��'����
T
(�sO.f���!Kw(�	ßĺ�4R�v�'�l6m�|*����ɏ!�@����JZa��9�ȋV� �f�'*"�'���n�47��p��4L �H&��k�A�Ĭ�>e�B�XӂN�t<D�5,�u��TZ����(O�g�n�L=c�kc��H����qp����!M��hf��zո��C1~À�s�L��|����T�Ca�<��1L� >�0Շ]џ�
�4Z%���Fx�"�Z��Q��
�:��$٢�(�?�ϓ��'��C!�'H��U.�:L���
N>��i!�7��<!�ɕ�)��'��.��V�đ�ISJ�X� M�o�R�',��+��'�9��x0P�V�5L��T�@�����6��GmD�.���S6BV�U�ԑ��(O��q׋ɚ>�pcd�[�E�9`q ��
�@�0a�#n���zc�.7f:��/I&�(O�hb#�'��7͗_y"i��?�$T�u.�		�H� �!O��䓀0>���Օ0��9H�S>f��l:�_��Z��$��%�����r�va+e_&c0����fyb��O��7��O ��|�!�ʰ�?!v���8�{��Y�t@:h��?���/�ޑ��Lôs���� 
V� �!��c���3̟`����fH���ny�lP"���+���	�,��S"N6gXhyF�)"A�9Y +H��(f�x�0���+K-�5,���2	�E�	'��S�O�L�ȥț>Zk�����9R���'��ht�F?U5���_7z�`���Dz�O��q/��b�:�3&8wL>�ґ�ib�'(�NB|`0�'�2�'�b2�R��B�h���ؗ�B=*b����b�*��
0*��@r�ؾ"��?-)L>q$c�*X��� �]�����ϕWsx�&M��=t�e��)>!�U�|�������^�7޾�hȷ{)� )+V���7�Xy�eH1�?i�'���|�퍬d�Hr�P�H�|�{#��O��hO�xA�B΄I4=:�+� h%L��_��I�4����':�6�|�����I��?��S�:*�8�΁y5�޶
�*Q�'�r�'��c�d>�4�)��ԟ�4�&�5g�lY����!b�R��2�C�l:Xs�h?E8��+�؂�(O��S|>!��	���J}a��(I�(���'p����ҍX�tF>����_�(O�I�&%�,r=���V+-g>uq���Drjq�YDz��$�7޲%����#;ø2�N�^���O��D*���'�f�q��B��.)K�Aº7Z܄QM>�1�i�<6��<��O  ���'���_��V��� =r���֮���'d,Tj�'�8����@O�_�MPpHZ�5�0Aj�k�m���F�/5��e��^���H��(Ob��@��4%�H��k�d \ҵ��h��T�t���Y����^[V��ō���(Of�g�'r����x&.Ϧ ��!`vh���Q�M-���O���d��G%p��χ�t�xK�A@~���O�p#�4�NU�/Z6����$�'��	9;2�
ߴ�?���	�=r�&�D� QB��Ҋ��J�Ԃ% �E�2�$�OI�w��6o��hX%��6q�����?�@���G����^7V6L��I#?��B&YH�Щ�mۛ&D���N]�$6����R ����qb�wt�����8��O:��3�'�y�X5-��ʷAݹ9h �m�&�!��1p=V|�W&��h<� �`��.�џ�����s���.�(\P
��G.�b��6��O"���O\��nQJ�N��O`���O��]&@�.yەM���pDڗl�#v���O��k�"�IB�)~�p�kG�|���$�b�H�z?�4U#gGV�@'þ<��w��a��s����l��J@�Mc����X������3�%��L�!ܯe6ă7������.Ot!�p�'���?�ORE�nG<	�}s� �y(��E��Oz�$�Oh�D�O$�?�'�0�!��$U%Ni�C�I� V�+)OD�lZ%�Mk�'���S>���e�D'8 �~���*ؽE`��	��E�0�p�����'���'����'y�9�"��#_���$�W\��I*D�^	�>����E&e�5�6��$q-�?�T��� `��.�^]�%m��	yHE��
�C~:�:�j�l��L��/H��X���
ۜ�O�T�@*xY�	�UaI�Q��"J-���'$ў�Dx�	G�,|�p��8"a<�Q#�!�y�O,!>|��,.�J٣c�;��Q:�V�'��7���ҩ�z�$�\"�8Ă�45��!��%��$�Od�h�h�O��$v>�ASc��ʭ�4��޴F[�|��-\�m�n�	D	L�qV%��I�Z����ua�9Z-�4b�
D>�M����d��q#gU�h��f�C�8�D��O��d!?�E�4ޘ�G,Yi���@XA��U�|CC��-&���s��^-�u�?�O���"(S��[3�M�Z�<��s��0'c���<�VJ�B����'F�S>�aD��ҟ��5� ;#��к��>�t	B��՟0�	�c�L;WO\Ĉf.N:�4�W��
���O�( Ҫ^��<�W̃<
H���O�hؓIi{\��E�>!�QJ�dΆ�X��L?):���%/�|E�W�6)�a��� ?�r�Ɵp�I_�O�ߥ\44Q#m
А���J?GQ!�$)4�Q �H�{�8��"� �џ,[��iF�;?bтlZ,>Ac� �5G���'���'K��{��9.��'^��'���DS�!8�&B�eH�P ŏ&%�Tp����bBڋU��SC��T?;"ʓϘ��s.?Bx�����~.(򎐡	��H����>��@�$0�|A�(�|��cl�.ۆ)�;�˛](6��ӫ�!5f���p`S��O��D%ړ�����B�7\�XʰU�B;�(�	�'�,s�N�&{���! �9��@k)OfFz�O6�V��YQ�� Y�c��B{v2B؄d����֟��������u��'""=�%C�H��Fr��sc�cx���Ib}���V�)���\�N|!�@��(OZ�	�a��h�>��d�<D�X���+�1�����+�h��hZG�9��o��(OX@��+���x s��Ȭ�KF_��A,�O��1+B�8U��P�i�K����"O�lq
��te�!�-v�z�˖�|��k�8�O�D�A�צY�	���`Mߗ2�z�'�B��@T�<�I�EH���㟴�'��4YT�������26��P1��=}��a�u��RK�Xc	�"-z�T�6�j����
Zk&�*5O2^�����A%Tu�����Ip�{�� �,MX��X���'���s��'��ec )ِ���ꂀ�L��	�'9�!a�G�&U�!I��3DL����s�r)�(��EkW�_�l\�(�C��6��~�J����?�����J�a�&�D��'W,�����͡��/�����O���']Y4i�FW>�p�t�T�?�Xt���o* �7�Y�%�I�w/�	$JwN9�'Q�^��DQw��-�H���"�'��uN�Kf���<�E+A��2�,�O��0�'�yb�˅3��Ŋ�A�!�X�
��9�y�)J������)��Q8v�{�\��O��D�t'� g
E(��T1J� L��&��@v�F�'u��'��cC��'���'��
��y�3*��Y��i���6��� ���
��;��6m���B��P-m�8xy�'��p4�)��m#��(6��qiIU�~j����O��+_�1�	���O_1C���y7�ĄK��०�
E^ x��"�'BV H��ҘϘ'�<��֎�?s?J4i�nշ3L��[�'5�}�d0a�&b�%��-���.Oz0Dz�OM�'�����A5Z�
uqL�	H�kR�]u�ȂU�'�"�'��O���'R�i��g8B��2g�U=���tʑ�_Q��z��Y�>��9��M�����'	�QR��� ��H��C�jH
E�a /�#Y�|�@�'��t���,mĳ�`�4�Z))���̟��Iq�'��hA�L�2������&��v�,B��:
�L�Pc���0,)��[�`_��O��n����'V�L�Ԯ�~�;f9�w�V�!��8�擗7c
�Y��?���?����D��03(p(��w�1���?�8����M|E�M2z.��j��ǈXe��#:ʓAD��vK�)I uC0g��k�(���6�80qA��|��
�ۀi�Z!)�I.���4�	��d�'08Q�8($��f&�9Y���J>)���0=�U#N�m�U��ś�#�����R{��HX�*����5P��Z7MμFU��	gy�&�&�y��'�r^>�qՃ��4k��Ġ��PEШq�����'@����	!x��+�H 6>3�\b�O
�<�O����Ĝ[Aj-sXb-�d�6</��s�r\k'+��}4�`�èYD�O�ĹJ�`Z0q2��ǈ�ra�]Z�Oj�3 �)�'n��1գ�%��I4�*Y�ȓȆ��H(0ʾ�ֲ (l<G�G8ڧ{�"=r�Ί�\4�����E����ߴ�?���?aU��.U"��?i��?ٝwDxt���"�!5(ېf�l`w	�r�x�K�g_i��9�&�F�O�l�H�-�Y?�m��K��sSID"dڕ3tG҂������C����S� \�ww4��|z$&P C��)� ډ��V>T|ٱ�P7l��|���?�dP6l����N|�u	Ҍ�kx��kq�
�#|!�䐋+�����ئs(L��k Dx��'p"=�'��{�	jvLM�֦}Ҡ �Dh���*�JD����?I��?v��@�d�OR�*
�t�0�k�B��	��QA9&-	 �ˊ=�X�((���!�d��7�V����<��F�B/MNn5Ҕ�K�be(�-�+b��lӥ@Z=w����-�u�:[E�I0T��� $k�2D��ʈc� y�)�Ofdo��HO�#<ѐ�ЊJ��� �,V9[��1r-�g�<�S%ɻq��������G5c�OZ�o��`�'cn�i "�~���g�DH�7��w�,�r�-ԥ1`:���?@,���?�����d I�=�VX��+�4ҁ[���*x�q�^�*��`j #'���c�]�>FyRm���>�C%�,�y	�`�{v Ӌ+���7�M$Q��c��]n�Ey��^��?��i��ʓY�t)�T����4"5��p(�%���$e\��H��N�~0�)B�����dR۟l��S��J+�v;���O��46��ia��'��ӆP:���-\����"C(`0/9 �uk&g�O��$֝5Yh�� �Ѯv6LpA!��%.`b]IW�n��o�n�a5����R,�UdQ����'R����*)\=r
�����S'��_�T���^�hW��&d�TXB��220u�������Ot-n2�H���S�H@�xH�DVE V�{q�Ѹ؞C�I58 L5��m��S5�5�h�?�"�S<H*�L[�5K&�	�,5sp*�n�՟��	���9�n�_�\�I韀��؟h�;9� �1$�r�����Q?fZ0���F9$7Xi�F�/z�έ�Ww̧M��*-O�����ez�	��!��8waӒ=8�y����,lz3���cx1���{�)V}HĮC��1��hA�h(I���?���`�<ysI� ��b�L>9���L?&Pp�f���ۓ"U��yb��)�\��W���e�q�i����d�Z�����'6�	�!�N-�ǉH�E\��� �U��|���ӀD������ß�]w@��'S�ϨC���z%D�"}~�hhv*�t��Uq��ɬp-ة��T��ဴjӎ7Np{��D,sUV`SD�Ȉ��P�I�3��0$gE1b�F� L�F!��k]�s��R��H*U���Pa�����$��54�n�yw�'�`7�Y�'8���4����F���RA*�;�y��8x�jBy�Đ�����r�6�'��I^��������G�j�)U��0t�a�Fh�>=<���OR0:%��OV��o>�H�.J�j"d��̙X�ї���!�@\#���&��%[�T�y���kы��5�Q��;���<$�L�ZV#X�C�.`�B�
�TͨD����$��6mE%xb�;^�p�z���Ǭ7;r�j�Fy�'�6%�h��Gp���Ξx9M>�
�f&���B�=i�(Q�a��5�2����?�F���K���Q$��%��4�`���̗'C2=r#�j�V���O�ʧ0X2���[)���  ��+�:�½9���?�p�ͻg����`)�
QQ|�u EwܜF�����{nܝ��n�?�^a�hʈb��;8�S!�\���1�á)�9�����ݔOE\��$��}ך�#D/¹:���O�9�'�6M�U�OV�)H�2��tJ��7.�D�@�&#G!��a�RQڗ ��q�~\�G⃣+dџԱ���,;���x'(�;T��Z�Bp2��i���'�2!�KE����'���'�:�*��7*T ���/#-�I��o�]�X�����
�zQ��ݸO�O�m�DW0!)�I�7L#�Ej�DОg(��
����Bz�<
`-vQ��J�Sfr�t2�Ԩ� �p.0BT�Y�t����k�	�'��D���*ȟ�'a+��fSz���31c��)�"OF���T֔��B��a�����P�����4���D�<A�׊zՆ��4��~~���㑝����ј�?����?��}����O���o>qq�FP�b�����r�d���V$^K4�#iY�12�H�B��[+Q���&$�k�2�	���<E@�1��	N'=YfϞ�M@,�WBV9`���c"�	R�Q��8�I�<��D��Ox"�3cDϲa���$���Ӌ��>�f�.�U�ǉ=V%
C�ƾ~��q�ȓ1�4Q�Pl�~�d�EcĢ�p�&�z�4�?	/O>YR��C���'���PUAΎ`����ƙ��xD���'2F�L~R�'����T�����6���рђi��#�	�8�Pz�ƄT~h�0�)��b�A����;�Ș{�gʌv� ��:^�>)5���������T�d��J�`7�Ek��d��&���aӦd�'�H�j���k^6�)�SR�J��O>I�O��9+W ��3�ܔ�ש� d^����Ɇ�?9Pa�E�HS��9�V4a�����'��h�#�q����ONʧP��e���#�2�Y�"�� ���B��3T�����?���5(����#c=L��%�F�ђ�x��B*������8��+wG��4xHR@� C��9M"�a�F9L�[�F	%D��ԀC�Ӝ8'�&=�sc�M�-���� A�U�ʄ�'\��,����+ҧ��� 8����a8��%ɸqY�"O敃6ŝ?��lc�&� Y�%��	��h���p���R��� ê8�f\��Hg�z���OR�I�|6�Ԉ���O.�$�O���p�e� �Уw�@\u-�&b��hٶ��?$��ۄH��j��26j�c�c>}C%�ǌT��U	|'R�j�I�SV���D�?[	��%$
6$��L�f�
CĈ�g�I�+74��'(����H�mv��H��H�MBx���i���&G���	�?9���!�TT�.ܣQp8(8�l�^�t-+
�'�L��Q͜21����@�1&���(O:]Ez�O<�Q��0�C�=��ـ�FQ��>|�V��>o��T���ɟ��ן��I>�uw�'��3�6�JH1�6��ծ��� ��程(���a!���~��Y,#D�pp��o��(O��Y���6�h�"�f-X��0x'U �\��H
!`� �f� p���舵�(O�Tk�
�)BǰUX�gU�#:H��&6I��dy���FzB�ɯ3R2�r'�T�r�gI�3{��C�I�����Ade#T�H��z�O��l�џ��'��Q�#�dӘ�$�O�:���6]kl�����1xΒАD&�O��DQ$���d�O��S�j�7��P�8��rN�w��ܒL��P�>�[��� br-��摦N�D�@/.ʓG�:PZ��������\�Nά= Ě v`�K� ɰD�lt�����6�@|@��;ʓ7����:��I�n��Q��:��	�n�������-l��(��_%!�qs�憣D!F��?A��4����Ʌ-�iB"C����چ�����O�UA.ߦ-����H�O���	��'�x��
ժ&��ԙ��[�	_�� �'�BF=�l��cBP�U2�+�7�6H��̖�>^��tx��A�L�4�6�Zå_�
���KJ��{����s5b@ө� �bI��Ҽg`d�OI�!���
Df��)3��|nv���O�\��'q�6͎V�O�󉌟z��!&�'eU�HK3��7o�!���0�6�q�B�y��T���E,wqџ� ���E-ery�Q���w
�؂��a�^6M�O���O8�K�l�}�&�D�O.���O��"OpL9�h�55E�8[2����5亜Y��<qs�%JQ�>�%F@�3��O8��qIV�+lp���M
�2H�	c2K��<���!������S���0������|�p)��p�;>Ry#F��,c����׆�~�%�H>ٗ�ɟ�|�<�b�t�0���d��dRp�<�a�-rЉ��E��-G�ǟ��I��HO�	=��4d�橹� �(����d��8@�Ͽ<�'�ѐ\D�o2}D2�#�'��0b"�O<G��j@,K��� nA����d�
��vj�'+"�ƑP�^ kF`�J4^(�S��.j"�%��<E���{J	�ͱU@�)2�=I�ɟ>P�^=c�Í2v��;���v���;M�&N	KBx�襉�j�PЮ�rp�Z,��SӮq������|����u�h���8s �tib��{y��'XrY{�"���P����q!\"����K= V�&Ȭ� �/P%fZHʓ`b��3��?)����I��� ���O.���T��yjf`�������O�l9��R�Q&��� �T[قD��c�"�;јOT��K0�H�}F~����4O���z�'CP��"ZkW�m�g�İ3�\
s&�J!~A�$GP�v��S�A�ó��bi.�8A*��	�=�.�d�Ov�S�b~Bj@�B�F���gڙUD�C���yr�CZ�5@J[+I��� V��'�hON!E�T�H�3s�`�.�>U��y�$��}a"�'�rG J��=��'{����ٴ.���O֤jg�
:a-d}�R��8�<)Yc��0L`f�e/�@Q�p-�%T��'0B9�K>1Vo25�J�wC��%-�P�$V���"�-�$f6��2$Ö^w�1-�Fa���>{�	 �3�,܁��պ�����FҚ!	F%�F������O���#��y�ǉQ�˖��i��f���y�[����([6�ʖK��?1��i>y��^y�AΨE	)�4�ΆU��|I�"CKɈ�"#�J���'m��'ޜם��(�I�|���ĭPd`q҆�A';]�#ڛZ9���(R2^����J>iSHe�v�Cu���<��h�if�j&_4�l�b'j�
 �y	�J]5�=#˂�D�Lt)æ�
�uX������	�[.��R F�|��\����E��EF�C���?�Y�P=�3L���E	�g�?X(�ȓI#��@+S�mI֡��b@�VL�D�'�H6-�Ov˓y��FV?��I�|T��&T��h���!1���.ȟ�9'-�ҟP�������,�D�򔀂BJ8m� :T���r˨(q%F(]F��"��8SB�� .&8��<�pe�j(�|�!�%9?�󃈟�V|T��MƯl�Vʤ�@�f�z�n�{����$(�<��x��x��*�M�A���"d|d0��܋,^̉(T�[+��8�O��zG�ĀQ=�����5�i�6�'�6ʓB��J#g��|-r����Ш�'gj�k��'!��'��әp5p��	�������O4f	Ȧ�̡�6Y��n	���{���[����lڜm�D�e�ţ!��Rc>�C����=��$:d	ηg&̪5�~�|��M��t�>�z�Ŏ�
�)r�Єڣ�8t�q�7,�ii�z�fz-���>O�,���'X򑟒�\�S�? ~��FO��T~r,z�__E*	�"O�Be�;J�Z#�"�J�P��I��ȟ��&j��a�~����_rr=�F��O����O�0Qv� S9\�d�O���OR���O֨Ѱ(�K���b͊���i�c��;��o8"2�-a�[+R���O*d��Q&�m��L5JG8a&iY�K �<(b鎼 ��b���S&���E���/ڤl\�a��'�(��1���L2,�I4�O�z��3�OjT���'�r�	�<Yb��}�"<��kǎl�U� Ct�<���[F���G]�yO��H3E�J��4���$�<1���74Vf��:f���8�k�)�T��!	#�?a��?����
��?��O��$���K���q�C���bv ����F�Z3@q�s%�p�.�M�p��`Z��Gy� ���ѪC��eM��1AĮ1���-�8��\y�w�� O�k�p�����WP�iC�k9"���ڸI�x	���2YW���B�'sr��a@�p�L�I��G�JL|��	�'��y ���>�\%�5-��m.*��)OUm���'��8�¨z�z�d�O�擱
Z7��^�z�A�
�!�`�\�H�����OP�D =j%���NĘ!��<?֒��c��G��	��c�H�$��R��>1 ���IG�	@����X��9�a��#�ty�h�Z�l�����y��$�F#�����	�o�`���f�'W2bs�)0��G��8Y(�by�<�C蔯E�R�K�m���[qx��s+O �s%��,����!_,Q�H�Z�t�Iş���ryr[>A�Ot��+5��T����C�l(MѬO�������'���Sܧ2����K�:6��k��#&t(�?Iܴ�ēK�����rk��yC�x�1(ؽ}���I��ߦ��	5�9���ߟ��S��=ThE���^�{��)����{���5��M���3xX9Q�t�B�=�����3VI}�4�;`�T��/�;�zP�7���I��1F�Ox�d~�<�к+���?��'�?	�'Z�i��G0J V�B2X�t�r6���?)��2����yܰ������5�y��y��-M̩�-�<~l��;ѯ�������O��D[8���O�R�'����'��-�dL!M�d8"F������F�O�4��'�B�؟f2��On:�ԟ�F�5@� ��L����J�
�6�F�Ӛ��ɡy�
���O���؟0�;�?q���JFٍslB�b��
�41���[�X@��]���IʟpZw�d�OrYb�ן�V�����%��V5*h�Xa�W4G����qKz�牭(h-nگ�M�e�Hi?�]w����O����t�^;h�i�8I�K�+y���7�~��Q2gI馡#�4����&{���\���Ef��ٶ�n��ɵi���vj�33����O47m�?mZ6�Z����Iј,���d�iΘ})c�!-�D���Sݒ9��O�&��u��K��#Nb�n��T�'��"�~����?Q���?��L�+�l)�d�ݾ%��|1u�/���tyb�'R�	�L����������%\5,9��Q�<��mZ��l�	��P�	ϟ@��v�T�'zb�@$P/�%
�A�a�����,_m2�6�O��D�<�)O:�<vbX�"L��Ͷ{�� Qt�W}B�|��<�f���ɃaEUl4}Ƞ��DN�vQ�$�IԟLr�� ʓ��j� ��(#rT&p"e�7=��6ͩ<����?�����xQ��S�!C�k�F�F!��P�"O4y"3���Sm��$��<�Dh�"O��&b&v6`�C�)5���"O�XZJX+c�~��PBց�ℱ!"O��'�ߵ}�d[ B�\�&�g"O���L�AW�e:��V@����%���e�r�����Q�H$Bw�#)�@AzT��(m��IQ�]�� 틚H�\U�u�3����o�d�$���L�X[���%)b��e	��G�Vmct�V0_|M+ �׎f:�ջb,G5���3M3���D��\�TM�2Z1����5���j̲A�<x��!�NH8 ��ldR���i+���/ ������СF�>2��liҪI9	^���h��^H\�3��.J��Љ�#'$�=[�l	0�Cu��)!��m���v�DŪ�N�n��x۱�ѹNl�2"
��	u�6m�!w�
 IG�!����b���E��O��$?��D2�Z�NoB��0�pN��i
5!=v�'D����M�l���D
FT3�}&����n������m΂c��sP�A��e1a\>�A =T�T�&I��|������5�R.k�"�'��>ulZ�#��l�!�ݬ�D�i2���~�BቨW�x$:P쇦s��.N���j��'�t�<)����>j���4{�j�s�#["�7m�O��$�O`�kT@U�^y���O���OW��/��t��@k�d�n-u�Pd��M@,gl��`�!N���Z��(�Sy�$m#T�'���:�ƃ`�,��2pU ��A%O���)2�1b� %�P��n\l�W,�/h��qaR��wJצ�J�vL�%�2�"S�Z�5�(Of�����d�?O.M��D4?H���4$/4�9�"O��@�Lנj�)ч��7q�����O
��VA�����',��)P��ܰ� 
_��L4P���*�	>�p��?���?1���~���O��S�p��p�Aۘ���1��;,�aK��6!S�\v�4�G�S�z��D`V��(O�	� \,	4���EÇǂ_p��h��C���@���yD0dѦ�U�p�Ҩ1�:��L>I�g�>j��C�+W�oA�M�@�Ӳo6m�	-�M���IS�}e��j�N�;�2�PE?7�\�I BA|a3J� �J��+J��R㞴1�4�?�.O<�1��A�Ļi;�l	C�\+��ԩ�3I�q۳C�O��dׁ|�h�d�O$�S�3ᤡ��K��#,�r��N �
�b7Kg�����2�
��#��6��O������X��y��z�j�҉�	{���r���>e���F���&%E~̔��?����Ė6���赨��7�Ĭ�sb�a�qO����� ˦�r'��'�<l��*ȢF ��ҿe��tIB)C�V�,8����*A�fҕ��O�ʓ.>��L�?��IU�t X�Nd�f�Z	j͙�ǋ;��6�	���I������Y��xks���'o��� �� �)�~�7$8��1����c3� ����h�I�h��|0�8A�h�K壋�	�⨂��t��6t�h�Q��!���(� ����@�U�I�G���i��PC�'�a#޴	��R�615��'g4� �زH͚�Pw���*߸���4Q��kdC��$�ipk�1&.t<��ȦN��F�'e��'@N�3��ޟj$��',����3d^5$���`���/i�6tat��!*-*�s��G6h Q;5��L��� �i�|�F���E�ubwC[�zU�i���^�r�R��\/UBl5�v��k�t�@��,�O_�$�d�{ށ؄	B�J��t;v	MSNI���a���,�<�BJ��a�L<9��Ɠ#5rd�5���On���l�W�<�6c�]p	��`o6���Q�DG�����'���#9pAa�+D5$a��2"({�v̈U$���D���?����?᥿����Od�Sw�T�p���<[�5��G�86<&�%�ȴ	Y�1��Q8-]�2���0fcb��s剺	�h|q kāk��R�e��~e�!�q/E������6s}b}��Q.��� #�ɍ1.�I��T0r8Ni��cIX|����"�O�o;�HO�c�9&��5��eJ�K��|I"�c.D�X���:�@zso/.��x-�➌b۴�?A.O��[�=O�u�Z0Z��30�Eb�j˘Fa�(����x�I�V˾���Ɵ8�'5_1V��uAt��ǩ'z}�v���rkΖuy()y�Y:\y,�(Ӈ ʓ�pa�m
�FY��7ݮnVDJ냅�}"�I�Sj�����9f���1sG2ʓ0t$��	��M�t�O�	qq�H�~x��q!�Wh/ *��'lOZ8p'MC�@�� ���p:��
O�E�֬I�esf�@aăo-��2�aJ;v͘�$�<�.�*�������O�X-JֵilKuE�3r `��̏���&@�O��"\�.D�#F�yD��*vA���ʕJ�:l����<�e@�.Y� E��ֈ,��%�@�Ʒ&y p:�&��1��<�v�_�_�PdcrS>�p�h��~5py	t�,�BdXb�)�ڦY=2�jӬ1F�Թ�2�(�a�,2���ccZ#O��k�"Oq��⎠ղ4aUa��C�V���'}��<A"o�A�j�3�,�3ʘ�X��20�T6��O^���OP��Ċ�� ���OT��O�i�4K�n�s!e4���!�G#��ݲ	�&rД0�5�v,O�|���E��|z"����{a)^�)S��C@s��L�E�/�ݱCυ
 ��d�ϱgWxz!��4�8�v�`�w��10�K�_����5����%L�æy{޴�?	&B�8�?�}�'כ���*
 �F�
2>�x������?ٌ��S�A�qv`��Z���J�F�r,��	�(�ݴ|L��|�
V���V�(R�Ė	<�RtLQ�Z�¤�"T�p`� _,�?I���?��N�n�O2�d{>ɺ2�U�NxZ�{Q�
0�� ��'qb=�dCȢ��aPND	ڲ�ct���yXQ���d��*��QxVg��ڈ���y�°��˔�@ZP]�B��\��<�$�B1?�L�y7�\�>~��ㆬ��<�i��MR4	�=;��O��mZ-�HOLc��;!�4p�#�Ì�3!����*�O�OލR�M�o����e� �m��d	�i�I|y"��E���M+@O�^����[�a�� �" ����'2�8&�'<;�S��s�T�����~�)�У-����'(60�� n\H8������(Oڕ�S��8Y�H�R�QXj-reN�c�^!&ɇ.���B F�m���8e�X
�(O��P�'v�7��L?aH�
z�V�;g䒎0�xq��Kܓ̰= (��#*����Z��y��LK�'�ў��3F<+B�
E'��6"�;QcR�x5����'�|M����\����IO�
�7��N ��pD�k	�@󔎞�Zn*,��ן�)�F�/y�����$�uN�<gB]	��gH�G��E�25%. %�F5s � ��ȶ��C��xR���^yt�E��5ҌU�e.L�'��yucVjR]�� [.'.A�;=��MQ֓x�dȗ�?����h�6��%U�4x���4v1��LʤO�@��:����Ī��ow�D�"����#�i>Mш�dU�.Y�}b��8��rWjO1[H���4�?!��?��@ªp#~�����?���?�:���9&+�5_b-R�O�_o�aѐiT�>�Ccؿu��#������O��6@ޟ#p��e�X���Uj*5p��ٹ5�L��bjlL�aM��*�8���,�a蒔�.�r��,��� �Y�r�	
�xH���ɣ[�l1�c�ן��'���j��|�����'2�aRq� ?]��4�mdJ,�'̼(X�d�'ε�3dB�S�\K�'��A*��|�����(B��p��ʼ%y8�#PgĖ?��|�񂎐x���	�X��ßx�[w��'v�)�.L��A�$�Q-&�eӸH���qr�3'n��'���K�E*7��#r1@��Dݛ>.P�B�[!$|��4C�:bcOcFRB@�a؂�b""`Ӣ����v㜔%���3�W5v��`d�T`�ԍ�:�x���O���&���'K�5��	_T���3��W�"؇�	G�I-�8i"s&�(h��X�IM+����2۴�?	*Ob�+��Y���i�1�Fτ=0R����xC �Ol���6M\���O瓩%u�������u���Y����V�F�vh9Z�� J�IPn�_U����	�l��+��R�,�3��or����9(xT!� �5�t|rd ���5�a�"��O��~<�o����dH�L�XP�=�
ۓ
�`\ʣʛ����z ��-�||��$�.����:7W4M���Pk�I"��M��?�)O�}H�kX>��D�'��CZ|nZ�]M\$��ӜH]�ó��<G`�����?	� ¥G��B�l:��j!B�p1�b �)��i�?f��`�s��Q7��44�FO����b�y��i��?�:�˷FK�t6�M�-����G�k��ЄM3��(�b�xB�	�?���h�P7mO�s �pҠ�
T������@�#[���=�Vш�MN�Q����u�˨�8L��	��(OX]Q�&�. ��yGf�/L��A`b�]��M���?��wA����A��?1���?���ߩ9�a��"!��0�J
�B����A��4y6���D�:�pԙg陯r�0��4/Է*L���+	\*`S��Z���\�$	�e��8꣣��O�v�z�N��w�2����p�'aw8��1�B06aE_�4P�L�u_�4 � ��M��[�����O��#&�X����<L���b�J�8G�<2�%D� ؑaݒ
�:����)<X,�c���L�I��HO�)�OJ�R���E��aX�0B�r�I(u#@,nƄ�1��'r�''��b�e�	����'"��qiWޔL�L����@M�p8�`	B������o��B�'��|ن��>g��X�Z�J��`�(��Q�zl%�A�bU�'&$,Ol��$�Y�]�*T�6!�n��4���U�L�r�`�,�Gz����\p^@2pk� ��9�[MR �ȓC�� �qϖ�?4 }b3����=��ib^�Pp�dC��	~ӈ��p�8`6��2�@ۓNY8�������	�k�y�����ΧBZ*����=n�ɩ�L56O"��#Ɯ� HDP�PP�J��F(��@qB-ʓ6K�Js�c��]Q�7d`93���2J9r�I45�� (��q�8H �e9ʓ#^���I��Md�O:Asfi�=ir���@�2�$�ke�d/lO�lJ1"����dJ7JT
��ub���f���D��Y^�� B/}��m�A� 4����'R剎R����4�?�������$� 6�K�d�^�sT�� 8PH��:r��P�	⟘0Є��^^� ���O6T��$Z�X�V���fIz�M��K�`��4"� I X�A���ē(OV���� A��Z0����0��b�(4!��$�q@�=_8:�HF'��٢�xBj�?� �ix�����0ڡl��F�Uڂ��+��|� ���O��OFc�<@6�ηYp�Qs�AK�uQ����hO�i�㦍۴��=X��4b�/�<YB/]�W�����``�D��Ol����^z�T!�I�O���O��D`��x0d��q���'�3d����K̅0%qS��*L0|�@ě�Y��dq��֢c� ���4w��p;���-u��K�/^;������"G�lT�Ǻ���q�Mo�'^�!q0��0��Y>r/��j�"�]���s���M�s_�����O�>&�8I�b��<������X��(D�,
4)*H�5�kCmQz�HsE��X�	��HO�i�O~�,�x�[�O�?Cl��Mё.b�h�2M-LM�i��'�B�'�Ovݙ�	���̧6�phȗ�W�h<�-��� *�����HD�	��!�*#��a�#�6Xը�ɷ�3�_D�]yd��.d�V�a���L��t˕��s��Ts��܅e#�k�,-kn�xD� �D�& R�%K�b�v\��������)�o��y������ΟKk �8�ʁgh����;D�ȑ$��?O1��`�!>�R��A�;�ɱ�M�I>)�+H�kO�S�=� �M��L@��cJ4M�2���D�3�?9��G|hT[��?�OŒ�17AK�r�r�2�@�L�ѮA�%�p��V) ��f猦$��"?�3�ʉRX{+^/ر`'@JMV<�c�$F�:��7�F�RL��2�	�+l�$�O��4�tE��H�B,b����?���=�
�T��k�l��S���U�K�UӘ��?�����[�Z�r��S`�*@D�r��C�?!/O� saϏ�����'2哶gx��l��hq3�G�!|�Tb���62ܐ��?A��E�P�Hڧ G�+Ԃ�a��0^�e���͕`*�!n����·n���yx�EHfi+<��)�Ak�v[,	i��)�� `q��
t�jԬ�4E�'��+��?���~�� �YK�Mk-�sƏĴD`�j�"O60b�ɗ5>4��mۙ%� ���'�(�<�2NϙP\�5&D�.EюHB�ɟn�6��OT�$�O��q�� �����Ob���O��Z�:�b 蜤���G2�	�tNN21�n�+3j�4x�@@�<��o�d�th~R��=���wS��5p�d�N�Nݨp)P�bD�<P��)5}��Gh�F��Ì��g�"e{b�әnZ��d=?�����͟��>�C!�d4Xy@�/Z4fB̀"��Y�<�գ���>�3L�.wG��' R��GK���d�'�	�8HjKr偌Byh5j͉3�f�Sq*�7L(��@���?A��?!f�����O��=M�%���@+G�>��ץ�LT(��T�9j�,s5
N�K}����#M^�'6  ;b����x��=��WA�.�r��Ï�0J�Q1(�Ayџ����O4wvHp�v�#-�����!=\����O��$>��S�L�p9Z�F�)	�>И1%�:�ܸ��5Ǌ�h��(i?����
��pD�=��i��]��Z0&ݗ�M���MSE`��(p"�@A�\�\�.U,��'���{p�'��4���C@͏�96ܙ3�T�dL�X�Æn�\���Ե~�	��뙊U����� �(O ��F�T�����d�t�"҅-f�;�dN~z0 ��
nI���F[��(O�J��'�\�'<ܴ�g����8�����)}�@`�'��u*��8vB5
���(u�h}��'	Ĕ�$e�:c�L�5��;uzf� F MS�'f �"�FfӲ�D�Oh�'n��y��4<�½@7L
)~YL����� m��0���'��$�|L������Y4�3~ ����	;Z��ӱX&��qA�2a� ���I `4:O���:���P-$.`|B�J�����s+��Ps���/����bO��f�8�j%�x�E�*�?��|��䡙X�ԡ�4bDx0(U�â �y��!B� ��Eʱ`�0�A�/ͳ�p<�u�>E�<K�$W�
K ����.	5�82Q�iC��'��-�}�b|X&�'��'���4�9��0��T!�͈�DdI�Mu�v��#�E?�����o	��1�T0��HĊ�?qu)�4[�R�M"o8��u�G�.ͻ�#��T�8��v�F8l�������I� 杸5�9X�Ґ��6(�p��0N�-��+�p��)�3�5+�vI�v�=gŘq���/J�!�$6u62k��P=��q!�ސ�����S[�I!{�ҵ����W�B�
�"�-IY
�B&XAr���?���?�ǲ�J�d�O��S�?]�q.	�V%J�#��d<��U�����D�Y*RX<ReA^f9�ቓ��(O��%�_;j�=	U��y?��n+lr,��T��vDRh��#A� �	�f��'�(O�m␧A�$����Dv2P��.�'0�O�
�h�n�X.D�@oDp*"O�����J��8���ܦtm<�����Ŧ�%��k�!��M���M�'$��9-Y��Ե��'�yj��'lz�;��'v�0��hX�����5�q���H
zQ��FV�W�6P�j�5q!��y�,�]{�N��(OjP�l)aNr=��R�J��o�~���F/~�p-���D����&�J%�(O�Dr��'V�'���y��#��J�̖���[	�'���ト��*�����Q�b�H��'�+�L�>�y�K&U܈���U��X$�(*���M���?�)� ycG�c�f9y�	l�3Gw�u�!hџ�	�`|!q�K�,-���@@c΀>al%J�A�C��q�O��(�'��%.rH\�i��Y���9K<��ߙ3����p��V��qGCN\0"�q�͵|�$�d]()�Bm��y"B��R�I&����U�)�#	g���&a�jx3����B�6��p�a�&�6�	�$@�Tͤ��Ox�'l�hKv�@�7dL9 pJ�6|v������9�	���ɈB<��y�jV��������La���%`����n�;h�4��R�؏qx�����`)�5>�e�O`���?tJD1��X�|�Pa��(5�xĳR�T�d�֮�%�f�Z OK�Ǌ�a�dlӚ)s2�l�4��
l��:6]|�Ru�EY��k�$\B�J����i�7M�O:4�O�7�'x��#Ó[*J��3����c��B��!�|B�)���u���h֨]�
�h��]':��D�Om�'�M�L>����Z�O��`�F o��@p�j�-az�ZuM�An�ZU
Mğ�I�P�I��u��'��<���YU^n�4��F�6zh����%@�c�b-���F#C���@��7��:��(O>-��[ 9D�JA�����qo�\�j!���ԥF�ƈꀏ+�F��E��)h��l�œ+Ts~����vs�P���_0����X��m�����GG�(�m'D����G��3��}�#� T��dx��&�ɕ�MsJ>� �X�'
�F�'F��Ύ�0�����B�!������$�OX3�)�OZ��g>��4Y0$�>X���:���Yp�H�
%�ৢ�5 ����˕��`��C$ϔIDQ�P��"�5; h��o��0�����]>3lȹ	��|��p"+[��2qB� �gQ� PF��O��O�0�4o� B��ViҪ�e"O� ��D�t��M�Sm@i�p
O��RbL0i���'/H�MF�h�b�0%ĒOd�h��O���ڟ �O�h�	��i�d�*wj÷-�:I�*"�n����O���Qy�Ya���+w(����ݙ��S��l�'4����CͶH�0���]�b�}$�|4�:����S��&��d�F]�@�xұZ>��MZ#�N���*I	Ve4ѩ6�>�dU���"��)C�cc���e.�\�w���[�!���k"��<�j��Pvfp�/��|�Q�)`�"MbA��;\�U�����`R��V�i���'���WS| ѻt�'}�'��;AJ�Qv���xEp\O�q���
1V��&9^tđ��|� �|��(>Hud�d�88�-A#.S*�yBsk�HP���S���h���l8��,��lW�@��w�r!S�"]�P*�0>\�y��/�v��?^����xBn�f�&��b�&i�\�0φ��ybi�5.�ӥ��,d����� ��.�HO��:�$
4d�0���A�:�Rl ��ɫFp�l�T$x,��	ʟ��ҟ��Ywq"�'����7'���i�}(>	�k���,�p�,�z���e��,�,Q �)L9C�t��Ć, 9��ul��|����$U�G�x!k�B8|�j)�u.��^����+�)6]=����":j��� �!J~���9r{X���'�������BͳBl��2l��o	�z�!��(8�� ���Ψ\�"x0m�qOB�oZU�	�-Vz��۴�?�ܴ"r|p�ץ�6@��"���v��(��'MK�')��'8�I-v���sG�9P�Jh1�C	�G��@9� U�o���sa�0p�\�x�΂�3x�I����P�n��!r秓�V��-a�N��g4���A�/�A�"-W.4��xV���
k����њ�E5}"��Qi�q��c�=����􊅼�yr��#A��j�G�-}tDa(s֘�Px".� F�N�:�ϝ�#;�����0i��bĘ|´i`�6�1�)��i�.1�6���N4r̒�I2m��?����Z�<u���4�7Ƅ��Ē�R�!�<��(A�GN6I7�Z�!�$�.n0$��2�3K�����y!�A-S��(zi# �09e��so!�$.xQ�}*�g\!�ؘ�F&��!��	"h���J���M+�+Y�+!�d��2E�� ��p�n�&�/!򤊔i ���#�I��}0�,�;H!�d�==���AC�<h�x��U�C:!�䈠_�&D�Q��?I�J3�֠H1!��K�T	,ъ2�J�
Ԡjk��p�!��2	���ů�#<88���!�D��=����7Q��	����+B�!�rd�ؑ !(U���kV��`�!��,Vj�4G�IllY�M��0x!�d��H:��CMB�/^j�c��ei!�DS0.OH���P��D�6�(yh!��rAʵ����O��ٚ1/�,�!�ą�a �1���ujX�d��8�!��(�H�0� �"U���F�	;�!��X�e��8�n�#hM "�EE�>�!��@#���'�0�Μ��c\�|�!�F[��1��O�e�1�6�E�_P!�D�3��QG��99�h��G�yL!��Z�� Z�eL��J�ƭ\3!���	SCH%p�X00p���s&!�䗜"�6���DæD�����l͞2w!��<y�*���@�'P��óK� "�!�$Z�;�@�+��o;桫��ߋ%�!�䚚N�,h6C@�ӓ���!�D�&�|q��#p5�蠀��p�!�Ȍ�D����U
����K ~Z!�$9f�e#���	-�ܙx2�R
E>!�DE�eJ|�mw�t*��! !�$W�_:��H����mh��l��,!��G<Bp����_6�-���o3BC䉂9�,��&���#��S�s*C�I�c��+� _��YX���XW�B�)� � ��tPx�6�R�&���S�"O�ݨ� �:$׶����djV"O��s��Z�;���+�Z}r@"O�́�Al~ޔ#B��6aԌܘ "O��	��ڻ�z�
S�I1P�f�#"O<-qw��?/�@��.�2�l�Ӳ"O�X
Ыѷ��yr�$j�Ȕ"O��ʇ�كG���#q���""O�|��B�p�H̪4��$�K�"O�p	saR��谡 ��7�0*#"OD��&`�E���a*#CQ��ɵ"O�xz��Y9�m�葟!��uY@"O���B+;{.�I��2��"Oܵ���Eu��	��h�"O�,!��ي"�n�S�(*�|��"O�0Ф'*#b�\3u��[C"O��Ie�U}ꕲ!@0=@�Q"O4��M�	o����(��C�"O�`k��ہ5��[�g�!x�PBw"O��r1��')�Ŋ�/D#��2 "O4�AƄԾr�� ��'P�CD"O�m�Wf�3^����m��EÑ"O� ���V/@4�L#1Hئ�F�00"O���/"_|j]�r&)����"O��c`�61�${$��b�d�0"O8�*SlGT^�bADוh���H�"O<�˔���r���84�T
�"O�Tq�����a��!�9~6�6D���]v���� ���)�`"D���s�7b�b��噋
��9��;D�Di o��2`8��]�1��� �+6D���R��^>h9��E[Q��ҶC(D��9��(u�-0VO8Tnj�HP(&D���/�teh<a6�+.�NQ�b"D�КW�
4jH�q�k�"h<�Y�` D�\���V�)b�9r3g�M�j�I4?D�`�����H�0B�B7.g|�0?D��C%Öo���H�B�v�{�"D����-�
|�r��G P�Y5�L��d>D�$Ӆ���r�x�C�pNr�)G=D�@�G�,3����K�}�J�a��<D�xjDL["i
��@ɭ��ѩ9D��q1dø>Fy7�Y�hT���8D� �&מ2�[UED�GP���3D�ȪC��h��}�0��3a� W/1D��z�J>Y�X"f��4�ҍB�<D���S�1=q*��D&]�}�8D�D�c*�`s���vfG�`TA��6D��Y�QtC;3o��O���q��.D�P��MZ$:t,�%iW7�ژQE�)D��8�K�0�mk��+4�d''D���g!��/	��`lP�N
�a��.$D�H#'@��?����>,m��M!D����4pO����...ؘ0�?D��pE���0Bŷ^�X]��%?D��0��0-�`�s�ē�&� G�(D�8��|� `����*��<���*D���, �J+�A��La�0A��y"��t[b๵��%6j"���@�4�y���8Dx��!�F<W�Jՠ7�&�yRB����]k�K�Y�V!xW�K��y�m�C����T��T�6gA��y�%<q1��B��G0���ui&�y�0>�� �P�UB��b����y
� ��	���W��s�Ɯ�hP8��"OB\��J�  2�ؒ��44���"O�Y�gŸ=�r�Q�"�3*bu�"O���&$ԃBD6l�g��_d�j1"O
��J�''�6��t�H�7�zqS�"O�4����+t�a؅	����څ"O
 ��O׊+��qg��I�8�"O���G�G�n����%�1�`"O��aD�;.���b�L��y��"O�yD S�*�5�#��@5��"O���C�����ƭ�/�>�9�"On��I�V;`�-�&�����"OH�K�e��m5��s��ʊ �u"O���,�����=ucJ�au"OzIr&�C�H=b��A�rR.�!�"Oʤ�a��<��ɻ3�ۺI@b�{"O��1�_�:^�|	L0;:��"O�Qţ�>i��-�v�)�� �"O\=(�� �`�	�Ȁ? �5R"O,��&Gu�F刵��d�L1�"O\��Ĭ��p�ځ�e[;3�R��a"O𨻷�ְq"i3�%�4B�e°"Op-SuH��Hl�5�WDP#H���.�y�FQ6Y֒8�O�$�ޕ��y��.ޥ��C�t�L[��1�ybA��*i^��â��0����Q��y����K�n�z �	*T��j�
�y�n�	X� ��@�&L���6+�yb̖81�ر3b �R�����=�ybB���Nu!G�W7�� ���V$�y2nW�l�jH����& �4!{���y�F_�D Ya��$}8)�^��yR���=�e�J�z|`��
B#�y��:^Nl� ��)\��b�(��yb�H�FtdH���+�h��C���y�VE$�(�o��j����Bȡ�yrJ'��	J����Լ�]�y��ƽU!VX릣]:2����G��y��Qƚ�*�K�:;j:��1�	�yB�@�CuƩk��%�6�*�-��y2aJoJ�ء"���qH}�p
�&�y�D�+'+yB"��dWz����(�y�(�|�x�܁`����.O��yү�%C�5Zr�
�`�� U���yb�!L��0B˘��lMq����y�C�X�.@��dFp!j��ye�-l�� ��*�d�6�L&�yB	]�:z�ـ�,�.�t<�%h�9�y�B�na0r�D�|3��"p�$�yB�D
M\�x�c��C�ɋ�+���y�JI���p�b	>=�)�Uօ�yҧMiR��wo�7�F���/�yB��W��%�Q%�$J������y��F!QH����׋!B��P�*�y2�/�IȠOB�����u'ٕ�y)��\�y�՜�M�����y�bO�!S��2L�B�褩�)�y§I5V���EA�0m��*����y�O��p��F�^�
X�¾�ybau�9a� �AY#F&���yb�C,Q��*w-�0n2�ieA���yR`P l\�����e�v¤O�y@�=��Q�.K�[�1(�8�y����3 ڥS�>>0��1�7�y
� �]Xs+̅'H�*gDK�3��B"O�Yc�䓓uC�M���>
$��"O���GBI,R�r���aV\��"O�f� Ƒ@Ԏ�<���a�"O*�`ŏ�ޞ�8'�JQ�1"O:�bR��A��,�V;`jP� �"OjqkW�R�����I��SPU��"ON� �N�[�n�)@I]:��1�"O^�j"�G"58b j�n7f��Z�"ONa�s��iqFq���H���B"O��bE)KD	h�S ��
!��05"O�uAw�D g�.x(���J��D��"On���>=�T��	��T`�0"Or�1��R-h� ��a]�z�����"O�5����>S��=��I1 M�TZ"O�)�C��ێ��g&�|��Ek�"O*��j6O���� 1P�F"OM�v��^Mb4�͏�6�t�R"O0	+U ���n�"Ўm,A�"OHS��X�֎��~��@b�"O(h)�V�S>I��-�	E��s"O�,T���Z6��Kqb����"Odu�V��9��-[KP�D|`�j "O��I�ɝe*������)p�t"O$�#F"ºqÎ�Ξ� ]
A� "O�u���� ��v��8[���p7"O�ݩclG�Xv����	:^} ;�"Oec�\UO� �@4pޝ��"O��㢁�	� L�������U��"OnH���H�Y���Z��l�p-Ip"O�,P��$-@�;f`�_��q�����?w���`b�:'��i.�!#S�'���Ӂ\�$�4��2%���1#�'��h�5��&�ەL����I�'m�}9&���XKp���kF�
1,L2�'�6�i�˓W��̸��"���c�'
���M�Yy2c���;��QY�'�PӇ�#ZP��4@I47C��K�'���'B�����K�h��E.�X	�'��|q`aF+�:YǄM���`�'�Pp��Y4^�Г@;GRE��'
�	WnI�h����d[�*С
�'fh����+�X 8q&��M3@�C�'#�{��u�NQ�@��x�1
�'�����N��x�Ӆ�A3
�'q��!�C�R�;�	���0���'�TaH�1�X����?�X���'�XJ�CQ3`�Y��ƈ�6�4���'��yQ����e�\�U�86X�Ha�'��X(u.�_� p墂E02A�'�Rf��R�Q�D!T)�H��'T�uɜ:k� ��S��C���	�'T����㖚DG�rs���&����'0j�����"`
��N0�|��'�hݹC�G;��d�nY=>�h�h�'ʠ�U�sr�0�M�66�P���'rh�s����*�]�d�ޕ?g��
�'i���g��(r�2q�#<v���'�Xl�Da�|�8�:�,݇���'i ��(�?�!rq�M35 &h�'n	�0Bƅu(ҭ{�B�/n���
�'���#�(O1>^Dr���,�L!�'\�8����k�� 4)�#
�'�#�� ~���E��n�ڝ@�'��]�%�z��c�%�d��(`��� �q3�C+f�D�ҁ�.~�$��S"O�m�C�;�t����>��@A"O���BR�p�NM
lb�`C"O �"�"�,W�(\���)c�r06"O8%�5{,E���Z�"Ot������B�3�� Uzn���"ON�	�I��q�P��LV��1"O��r�&	� 7p�@����lM�(�&"OZ�h�O���]B���64J�kS"Olm#��G�R~�ĠMٓ<���"Oh��vlP�A���+����I!"O��x�M	b��2�S�Nx��"O5���B�*�(�����G�P}Yw"O8��4C�)XTx2�J����"O`J'k��>��hS	K�i%���D"OZ]��
@�6������$ ��"O�m�u�5T��;&�y>��"O^��Gi��pPy;�ր!J�b"O!�GȆ�$����9P��#"Ou�0���x�ͫ��B,Ojȧ"OPy gΓf˶%�1b��"O�M��II!�΄�����Е�"O썓f��6A�ꔠ?3����"O��I=|�ȥcPB�$����"O��۲�̤,熄H��D�2�pի1"O���a.[KL�����V�>�P�"O�a�Ғ.hހ�W�ɵ@���a"O&d;ӧ�7_q�i�f��q���y�"O�iE�G�~�NDH�������J "OJ��'�O�T�&A����"O=��@��/>��w��i���3�"Op��XW���C@"^��
<J"O^�"4�*r~.@��`W�zeR��r"O�-�F��x��\	!g�K�����"OF!��F��jv� �d��|eAT"OV�9�fBI'��q���?��sq"ON|�*�%aî��-�?B��q��"Ot���!ֽ[�bm*Q횔?�bj�"Ox��0&Ȧ��b�n�4'��I��"Ot�3K?K64�#�9)��Z"OT$)!"wD;��[�1���h"O�0�����(ޠ�c�I��:J2yy"O8�H�)�E��K 
F3L�	q"O� ��D���@�Q�Qv�06*O�X ፯?Wz�7�Q8�Za��'��#�'�fQh�E�/;���	�'m�D��ڀ\sZ������.�	�'p��ڣ��HN�!˕ &(�HC
�'���:O=]�t�(��A�\q��
�'b  �f()-~���Jұd9���'�����!�f`���$RN b���'XUi����p�%O@�J5�(x�'��t3Ǧ���HB���A�Z�!�'`��Q��ՎS�(��*ڻmR��{�''�9`��M���
e�i�B�@�'Tĩł� %�)1�(G)u҆���'�xC�o� +bl�s6(e-ʉ�	�'b@����:���Hf��oF "�'�Ve����
����I��D��'�ш�?����@O�@]��c�'U���� ��uS@eZ�
"�Ļ�'=�<�`��(I iO�Pc�TI�'�Z(X.P:Qp���b��=B����	�'$̽ʤdل;�2�"
�{K�p���� 8(�a�UB��%:���Q��9�"Oj�	�J��1)Zŭ���C"On����]$7����'��0C����"O�E{`��o�2�[F��~��b"O��7a��P����.�\�:�"O��9�-�0%��Ph��L+=�>��6"O��	��QoO]ZA@�*l�x�t"O�,`#�Z,s�P�刷Z� `�w"O�!�wG!a�`�k�+@8�"O������=����@�?�����"O���'�,�����A"t�$�)�"OrQ�ӭ��h=D�p���b�(���"O�E�M�y�:K�A8��|��"O.X"̍FZ�tz7a˖;<R(�b"O:��KCm�!�v�p+|5	�"Oj�;�c��ҕR����ly�Q0"O�t�J�:�ѫQr�@�s"O�h ��L{������0"kޤڳ"O\�R�*�*J���}`��aD"O�S�؇kA�����5(#戸�"O����?(0�b��WV� �"O����$�{�p1��J7"�1`C"OJI�Cb:G:͂��ֳ\�B�(A"O������;QF����)D�=��"OH%	⤍�.:��#��e�zl�g"O���`A�2��F��r�|Q�*O.�)ĉ����">Ej���'�"Lx��ȥ����B�(���'!�d�F��i�
�Ř |DB�2�'��}���7�!y�]�=�B�R�'�ڔ�,�
J�0@j�l��H�	�'1^`��O$�x郤)�q`���'�FE�-n�.�CJ��h����'�p��!˱3��	!��_�f��4��'��YYv��27��0j`OV8m"	�'������1��5*�E�,}q����'���H�%P�:�:I�F����T�
�'�N9!��^�:�Lb�_� ���'�0��3�)us��Bt�d��=r
�'����R�Gu�\�wE�(�u(
�'�>����3����	�Ip� b�'f|�X��V*��YGǋ�{b����'P� u,K�(��vJ�x����',$�)��^��P���%]2���'����L�:a�P�Qb+$����'�:�	�IIt��Q3G
^!,��'���U�K�JN�Y� A8O��e��'J�����n����/�M�*L
�'A.�+pg��3n��/Mk~a��'���W߾6�:�R%D�.]��'��LCE)Y=x�@���w��b�'�b<�Ȑi^�)���Ot��
�'�l���Ö>����N�W����'f���dB���H��#B�֐z�'�L��t"�&m/ּy�s�\�a�'|Tqʢɇ�B�����K�Z�J���'�0d������,��fSM�D��'�������c�|�v��1Y�d�j�'l�u��\}��P�hG�Q`���
�')��C.ژY�����X�Mujd2�'	"� v'T.a�ԹځbA&\a�R
�'���k4iI�yĮ��j�UQ����'K6"p�:b�pX�ኂN���Q
�'��9 �Ɖw�(��^�Iۂ��
��� �4��d�:�p��ԙ>ؾ�;�"Od`9�a��RL�����>KhvAs"OtHS�^0Sr�ɵE\?c҉�"O�\Qj�p8)�#T�Q���"O����a��zt�Ւׂ�{�����"Ot=�f�L=����{;6,1�"O�$j!���p�zՠ�JFj��7"OƩq��ہ}�lR4I��?b$��R"O��R"b�jƸ�Qd��CG"�Ȳ"O�}A�&H�Pq�"c�.y�����"O��[�k�,M�:�b�'?4N��"OF��C�Ӈ;���Bf�.D��!�"O�d¶�̙jXX��Xn���"O�l�v���}���""� 7�N�р"O����͜1a�NT7�?&:P�u"O a�bh�CQAQ�Q���"O���P�?-��Y!�� (PQ��"O:!��,�eW�7��5���G"O��`ҫK�u�|ՁF��>}0�3b"O��cc��V�B�ڠFܽ��'����ܙ8b���G�.r��
�'�z���K�=)�qsu��$��"�'m��;3��ym�|j�hX�\��I
�'�.H�W��lr�-R��RNA� �
�'�T�T�;G��@�EV�a�'��:lΙ9s���s(�{�洪
�'Q����/���u!ӊ�6,�R	�'$:�ir�ҵ-5�Hi�$�# 6�A	�'}Z!�',P6%q0L_'e
dq��'ς�ad��<Laf�c�O��
���(�'#�0uHt�*0�@ �9�,}�'p,�;2�Z�R>*e�G4��'�X"�L��4C�Iа O��ia�'%YW��jܮ��#]�w���
�'�ȴi��{#����n�x���ف��\�dT���D�f�>]��6W��'L"��ǜA`���*6a4<���'j@��`Z�#0� tɖf@f���'M��2!�܅9��h���%p`ʵ1�'��M�2�6o�D1�BU$����'t����Ŷl��rb&A�E�\5Q�'4�x	$��
�~d���Ғ30.���'�~�r�a fحXѠW1H���
�'��AC'��!_��*!$�!����'0�jJ���C ��=��R�'�ĉ��!I6�iA������	�'+�!pB�hiF���������
�'��[s)@�	�@���$4���	�'�6<�&n@/R��:0ȩ:+�e��'Y�ݓD!�Oc����?	�&La�'�d�B㤞5S�iPǫ:�|P�
�'���RF�AXDq9�K^2]���	�';�%�e��10��|ؖʛ�{a���	�'���YDb^0[h2`��E^�A�uq	�'�j�釂�!R�
�$-�u+5 �E�<�T �[D�%��JP�+o��jW�Bk�<� �V\�H�C�B�V�d�<���+a�ޤ�l&'e~`
a�W�<��^�R�n��	�=�+��N�<I��)7�J9��@�	�<�(eg�O�<����񔬓Ҡ[cnB⠜�ȓs����.�������a�ȓ�D@p#��=(����b���%+`}��d
8����&_��­Ǽ@�d��7g���&�4+ö9�rm�R��q��S�? h��C`Wo2.Qp�M"
���rC"O6m``ʈ�'ypXyBom�R��"O@-�3�ۍz��Q�blE�M{���%"O ��'��C��q:�E=s��P"O�@�@�_��9V��ya��iU"O�)Bs��/B@+E�)
GB]��"ON�27�E���(=���v"Of�R�Ֆm�,�47(�(�"O�@�a�H��ٺ�#��W&����"O�\��H������_�C~�@�"O��"����#m^�f��
~�:�Q�"OL��dϰ�8�2S�՛K��`�p"O��9S�X��uR�f��X����"Ozd8�-ՋC��I��Ǆ<�|9$"O8ؒ�@ߤVˊ�������q�"O��e̎ x���5eO==���;�"O~�uf];F�"H�-��dp:�j"Op�0Ў��\�$!�#��
YrHے"OڅWS3d#�l;qo�_�<AP"O��{v&�	�����:@�%qd"OT�k  �nz4s,�2"OR١0
Mn�t��ӑ+�̡+�"O�9�1��Z���_��@I��"O�� �E���gI�\�t];�"O�	i�-K�&��[a�ԻG���b"OV)c�-���F�c�&�p"���yB痒z~�;�ohY�8��b��yHő4-�)���N�[�� �T��y�E�!�x��
$Ԗ�A���yLT9����"�
��-r�g@��y� ���xpa'��l�4�����y���Kl0㥉�gE���Dʂ�yr��H�M�%���[�f��cH��yʁ2/�y���ZSA�r���y2AK>��QH7�݆	��Cw�U8�yr
��P��Pl�lU�Y�v���y���<�b(z�a/49���F	Y1�yBʅ�S���:RhȺ���r7�.�y��	�A���HŎaY&(��y2� �K��� ���)Zv�5$*�y�L�V&���Q�Ko`�Be(�&�y�'%/��0�I�F�J��m��y�"M�l�4�(�n
m�ܼ��OK2�yK ��09x3%
�bft,9J_�y���'59Z��U8X@�8���O��y�Q9R:ܲF*��Q����'�yBN�Ic|� ��R�6� "�^�y�ĞB�4�F����x�q�K�y�JЄW�T<���Tq�f���yr"�$T.�`"��R¤u��yX�R��V)K0 w"D1T���y�ƛ�%���
߲��|��F��y�c�qh�b��Q0�!#� ұ�y�FբǬ��r�
�)�e���ҧ�y�أ:�֠�q���)IƬ`�O!�yŻ�0���)}�"��y�IS�X:�9�vE �&�H1�
?�yR��%n`��^(`�@m��w>�u��'IKY�h�:hǿQ{| G��E�<�g� @�`�PO0DG8�ypoC�<q��	�e�w�Z!Y�\���s�<	`n�\293��Z|��m�k�<Ѵ	�6?�D�8�C\�h%�2E�g�<9�־-H{6��42�"���Ti�<� <��� j�h�B��K�B�0��"O>���I<�ZX�ɉ5f�����"Oҕ��i@�3/�<1�:�a�"O|�SթEl�r=��όp�����"OLP�@L�P"�����D9$���"O8�� �jq�\"%�I �p�"O.]{�@l,J\�� �o�����"O<�؆J��c�l:��7���"O�?�p�qk�^��-K�"O"�ۖ(�8폺P�Z�
c"Ox(C��l��x�� ,���C"O���e�X�0����>��m"Of��N ��աAH�-B0}Q"O�`k��?s��Ä��7�+W"O�a���)SHV�;G� �r"O -ZC#�EԴp:E��"gZ5�Q"O<��GF.��őe���N	�"O��@ �
�e�C�M�3"O�U#f)D
�pmx$l�b���"�"O\�4�ƕ�Ȑ��d��Z9	�"O�,r�BۄAg�=�q���X�(�a�"OJ�yT@�F(�G�R4�f��"Or�R¡�"|?��0"Ó)|xb�3"O� Y�L�7R�N)���W1B����e"O���Cفm�})1�ŚF��Y�1"O�:��Q�B80Ö!Y�!���g"O
!�%&D�k��Ӏ��E:�B�"Ob�C$��>�Aid*�D 89�c"O^�)��B�Tw<ڗ�]9\��:v"O�I�u�U��]���H�#Y��s�"OL����,�8`J�o>8 V"ONh��i]S�и)���&�0Ep��'ў���H�Xz���"�25 !�p�%D��5��VrhyAC�� ��4�&�!?����S:���ѡ{���yCO�<C䉧e��dP�Pr�;4@őY�:C䉛P-p��CKpǆ��B���8C䉸5���@*�,�X%Ö,7J�B�I8>���ӱ)ll��ژ \FB��*>��щ2ʙ�;d� �A4}>�B��vg@@��]
j/4��T()�|B�I��j� ξ=5� 0���c�FB��)�9z&����pi��4�&B�	�bS��P�'��=s0	��2N"B�2-"��GmK+S\ �[�\�a��C�	?3z�"�A�F��Piڽ.uC䉰�Lik &L[H񀖖V��C�I��|k��e�1��Rj1�C�I����$��SPQ0�<1�lC�@��%�Vm͡|zZeqT�N$9�HC�I�}<� 蒈ù<��u�S�H;ZC�I����b�Hٴ�����E,�PC�	9q�^��WbD Nʶ�!m��P_@C�	�<=Z03�1h��!��oH�3C�ɦS�� 1�銘2��U�"��4%C䉅�����ɠ;4d��0.A�@�C䉓�"!�u��2�f}�j_�h��B�Y.Sk[�n��E:Rn�![�B�I�nBP���U*�~5 �$ė;��B��(u���5KB�z��� �k�8B�IH�HHX�J�SFms#�5Ih"B�	�;h���ҭ!���p�BT�XC�I.SItU�E#g�LHW�˒a��B�	�O�H(bkI
Y����ǉF2p�C�)� Έh�əV�P������!"O�1��G_5U2�xsҮ��D�ձ�"O�T���;o�2�s�K#(R�C�"O�|��"Q�,�0�B���0I'ZAk�"O|�Sc��<����&(�KHċ�"O�(z�#�>�H��G��5���Z�"O��Qr/����,�LG��R�"O��r�U�Fв�8��}�G"O4����S���Q�s��)(��л�"OD�'`��@�|Y��˨y���@"O�	��ǎyP.MI��ƥe԰"�"O>$C�o�/R����,�O�(�`"O4��&A�lI�0��k�+u(�S�"O&Ź����8k�C��t�6"On0��Ĝ3xy�@-W���the"O� *�	O+M��F쇱/� ��"O�)�a$k(��7KJj����"O.$���C���G�؄1MB�93"O�yڵF� ��-03BY��u@�"Oz��`��;|
I�0߀�.�K�"Od���W	�D�e��N���Z�"O�D
Să'6�蝻�_0���"Oz��d�@S��{��4r9:�"OnкU.X��Z���NQ�i�Ay"On���,�$�t�93n9/�.���"O��GO��*P��Y)=B)���O�<�ܖ�B�����<|A8,�o�J�<�7@C��}4@�8,��t�B�L�<�8�ޔ�!���B-��I�<	SI�= �Xa�e���p�s)D�<A�I��Ѹŧ�h���y��E�<��D[�V�v8��̀1qy�x bN�<���R.O�LP3.F=KW�V�<� H�.�J}��I7]� �����Q�<���
�r�I��@�1��K�<���"t�Y�VM/3�v9�fp�<��I3?'�ԛ$&�)sw���ŉ�`�<->�@4��|�͂E��	G\�B�I$(���������:U!,|B�Ir��y���4���Ȁ��"Tz�C�I{t ��-&W�@hG+�w��C�	�`��MĪQ�;�j��'�$�^B�I.v�>d*WC%*$P�ҳ��["PB�	�&z� C��Z*&����]	��$�4.���1�D�%P��{���l�!�
�M���y�&о:� a-��!򤕩A�����\�|{�%ҕ�7�!�yq&��v�����p��c�!�d�>�hQFA�7� 13L-�!�dىflq!Ĭ�t��]A�Jç�!�ț~Y* ����*hml5�b*]0�!��Ѹ0�윀T$�Ta�� ��c�!���%-�jCCň�/,vQhҠ�?OV!�D��a �@C��LH��P/:<!�DR2�D}!&�����9�a��!�V�[jD��Eě�fL���w�!�p�G��e����4%�,64{�"O�#J~� � �@�  �(w�<�3��V+�h�!��e;JI�@/�]�<!p��%󘜠 �r^�0�T�Y�<Q�i���;'!L�Qm
��A��S�<�2�ǁ%ˠ�E��.�	��NOY�<ѡ�I��A�B�.x<�0ƅ|�<�ĨM�k=Ҡ��<#8�۵�n�<� ����朜H���wN@�st4�[4"O8�a�Ȏ~J�]��5?���"O�y�l�x�{3��*U��*�"O�+#	:�b����ӑ(R:��G"Orq+����8��H�qFNܱ�"O6��0�.e�f�F@��PW"O���@����i��I���	�"O P`�(SJ!�f*� �Q"OL\�4��;k"�jjV;�5�T"O��q��ɈO��G��0=���@"OZ�d��g|N�y3@��0�2g"O�}����L�p5��o�d.��Q"O�����L�r �0A�.�&aN���"O������Ho�	��랯z0���"O��Ђ�ŜLAѫ�:3&�4;v"Op� #̬ Ά0 ���_
X�R"O�x��-����(�'N^, ϒ�Y"O�ī@��	o0��.�2O�H#d"O��XG�?H�r4��)F��@�"OL�۶k�0b�U�rڪ}�l0B"OL�[��>I�H"
��0�5"Ov�Qtl\2M��i¹lz6pQW"O�	�f��N�R��Q��hx�a��"Ozi �g�+]>0�J�D�T�x"O�A��о5@T�#��(Iu&x7"O�\�r@= ��!�!\o���"O*�pѠM�h����ϊ)r\�88A"Op�Bf�H��Q2�ϐ>^V�u�"O�|�qkE-�5ôo �DLH �"O��MR�=&� �T�
2�9 "O"��C¤H,�Sw�θQМ"�*O ��",��<QE(6$���'�x���Y�J	��E,�}f!�'c�P҅��1�U�s�	/y�����'�!q%:ͦ8s�� G�	��'���A��oS�!�I����S	�'�n@S�̼8��=XS)�������'�bT��U=*���qf�I�����'����-c"�Q�P;켘�'�<�rdO�K����K3�څ�'G��-��\�R�΄#w�Ժ
�'Ɛ��%LI.(�\I#HO$08���'�d��8p����!�#���S	�'6�@��D�1uT��B����Y�	�'�(����tĐ��F��CR<S�'��a��/Q�7��1ՂC�5h�A�' D�c��YI\�Y;��^�&�l}��'�xxz��<D=��ӭQ���	�'��p"q�D�@� <@�'R��D�1
�'I�P��@DL�����-Rר�*�'�@ذe�n�~<��lΥE~��`�'8��ӮL�W�B[�&��>ǔ���'��L赆��E[�����5j��+O��=E�D��#YB �HAQ�]'n��\'�yҦ��y�<  �ޓ&y YK����'�����n�D�A�̸h �V�zߡ��~��!�0)ڛ\F6�I��#M��"OF=�W�Y(;���ֆ�&?�����I1���������H#&�2eŌ�"O���%���P�T����\�O���1W�PG{���G�H]�B�K�g6A8�K@"I!�D�0}]D|x�� �hW
LbJO�P�!�䗷0b�a�΂hVDr�JZ�N!��0]<vu2�l�R&2p��/�,e�!�� ����,��/H@�Ҁ\?���"OP��&��/3�!��Y�(Ѡ5A�"OR�[V��3�\�����Л�"O8S4�G#�4�̊��ؘ "O�5���i8�S#ˬ~�<( "O���Ç�U���r���f��b"O"�Jƨ��_e�tqQ�ڟ{\U�@"O:����J������R$�����"O��Cň�M���r7c�05�
��p"O�@C��ȡR7Xl����V����V"O�,�#��cf�쀗��3Fg�pj�"O@�S eƈ�!�'�1�
��"O���L�5����F@Kb6y��"O�|#FB�sP��*���-|h6"O(C1ʐ
���rA��}$�h�"Oޝ+�Ȋ�8T����J$b��噳"O��`[_.��:�ʛ�z�ʌ�@"O$󗎞�_�>�R)_�U=�y��"O� AӇF?[� �h��ٴ`'��"O�]���9$X��ТJ��m v�*��'��	 :�y���:8m�lY�C�g (C�	pd8É�<�ං�rt�B�{�.������H)��B��_%H�B�� @?��X�o�]�C�2nƈ�1�@+�4a����s�,C��yk�!K`��7.�)
���6�b�ϓ��<��-�l\�}��L�)Q� ��S�����Ob ���0ih�!�ǩ��nD5��"O��+1�ױ`��|Id�ؘZ�4�r��	%EYtF��g��@-�ֆ6��u+c�Z �y��G؁���H=_Ì�8����yR�Җ�O?��󥁍O��bP%ɍ�d̛U�>D�ؑ�D��K�Q�!�g�J���/ ʓ��<�� Ř"��rB�S�Y@ȁ���~��T�'h�,hh�G	O�V�)u�C��B����y	ІN�v�LA	�d"��#?����Q>b�X�����K�P�VS�C�3Sߜ\3�䅧yΑ�w�����	�7�6�)�'M$�}�
�F�RP{��>a����ȓ^(\e��E	0�@�R7g2kt��&�X�$�'{F��g-��kH��Ӧ��&6����,�j�D�"���P�!SZsҽMB�E@!�Ę8J��(����:ZjM`d��k�ax�퉷4@NX��L�%t^�d���Ȅk��C䉏@+�h��LR'<j��w��1��C�	,$�T��K��W
uY�/ƊS6�C�I�|���ヤ��(�U��b �C�ɽ+e���A�.)#��Ǫ˘r�C䉧E�p�آ���;+�Xp��I� `C�	�fyy� ��ᴐ�`H�i�^C�-{��H�B*V/-����s#��}�vB�ɗkڰ�k6�VF
|�k��%T�PB�I#`�4p`4��6|D���_�CfC��;N��1K��t�:se��P�B�	�7��dIP�s�`0ʂ�E6~B�����$�12���+��;�TB�,(w�0��Ejn��	�ڌZTB�I$q��ƭG2x�2�U��3x@B�Ic�­XcaM�(|j��fg[�-�|B�	y8f@ ��A01�N츣�Ĳu�^B�I���9P�F�e���fA�W�vB�	 Gp�Y0�!hf�А�61.�C�ɒ'��41��Oݮ�u�N�J&�C�ɻ0�f��ԈN����1G�?[��C�)� ��#"Q�p�JW�4K���U"O��� ��5Ca6MJ��a�F��"O&�@���vH���
דt��Y�4"O��;���-]��񡃏3x|�miu"OJ�z��C���1��$��I��S"Oh�ҏ��>rX�k�߰(a���r"O��FBB�}�0���CAw=���"O����(�[�fhI��!��U�"OB�b���2��9f&�,G�H��"Oh�:��7��D�RA�,p�"O\���F�Gv��O�>�^�Y"Oȍ���C�H]�y@p��$5Xd��"O���7'��7CHB �rD �B�"O�d@6�1o!>�� �[5N:�t[�"O�3i�g1�菽f!rP��"O�Mw�T-�J����z&%SP"Od{Q׵d��̠m��H�h3"O-�p��
��t�Sf˖!���J�"O���ᮑ�X0��ղ:���8�"O���@�P;MQ@�h��8{�DH�"O�E١O�TBH{5�u&dr�"OVd o�t����5���2"O����i��=gL��%�)3�l�4�y���'����^�]B8	���ď�y"c����1�ri�?,����� �yB
6��!�4e,���q�L���yR3|� ���^����/N��y2�E�<˘h���492�\��yB	�9]vp�`hH5�$%[�œ�y�o@!k�x��g	�%#����S%؝�y℄�l��q��!��H�nܵ�yMK9@r�s��-� -a��P��yr�[&
M�9��lK�}�:�	��?�y�
xn����̂)�B�q��:�y")�))4��%`����c��y�"0�(�6�H�X��vo�yb�V%�zWo%�����P��y2�RM6ى�a����$�t�C�y���-k
$b �w��4w��5�y�d�E�(B"�W�v�����N�y��S�j����! 6� �u	��y�C�{�x�hkē�
����=�y�h� (��}��σutQ�kҸ�Oz��U�P���޴�?�����I
/6�̅�p�E.P0Q-�z&���bm]˟��I۟,�������cDK4`� R�ʈMH�0���X�B% *����,}�O+@R�<�6Y#pޙ+��ץ<o�����C#vv�]��q�&`��ǘ4;nH��(�+L�Ł
�}j�&�\�)�O��n[��'�M;��Y#2���'����$W�C^r���O�0�RJ��c�Eq� ;`���>���Iԟ<�ڴ}�v�iZ�7-B<Y���ѯ��t�#�'E��wkuӊ��O ʧF�������?i�49�}����h<�3*̐�ډ���ZI*(���8�؈Bl�0wũ�$C�_=�S�?y��<_�=�0�;32�i�3�أu�>�nZ�}¤pfË(W��J�,޽oYV�Bq'�C��&?��[�b����ƭ*fD�	BڊQV7��,w��n�$Q�����i���j'	�+�يcQ����'k��g~��O��v�(v�X0b��kV�pu�ɏ�M��i��e���$៊�]�k4��q烪Wň��A2pR%���?��n;]���?���?1s���l����D�9��&��3��<a1k�/-ܭpb�ͱd����P
�
��������%�%�$cvppS��;U5Ƭ��B<~��,���-����5�E���_?�P��Y�)C:x��O(�s�4&ptɀtc̡[Lzd����\sGW埤��4 ���gyB�'-�	)�n���'y:��Af��H�ؐ҈���OHQ�ul)^b����-$LB����Ԛ�Mźi}�'�l�R�O��I�0�d)�u��4S�0*d	@K�V��EN9��I����� �ç��t�	ԟ�ڷ�ۛ*+�2�,�.n�k��"l��1��U��l �!��q^؉��	��gĆ�<i��V "�,ة���%(�<��ՎJ�o�.��pLG�s�r����e�f�jݴLsPQEy'�?�q�e���ۂ$تh�꽀�hQy�vPڗ�iZ�]�8��q�S�� ���P�(_Ad�h�]��r�Of���_�^8�g�%!�"9�g�\0H��$��#,8mFy�G@$"L֝ǟ��Ia�Tœ	&S\��A;PE�� �䁳NUT�����O0�D�O<$�B�;~ܠ���O;fe�aq�#ͪy4�8�c��o�>u����	E�|MZ'�êG�Q���K����Bցu���[w�2t� ��^�oXf���.9�@��d�P4Q��E�O�xo�ħ�M;`�L<�@#"//V��幨���������\�>�����"O���zwJ_$��w���	s�DMnZ��9�@
D	,ΩV�=D���¨����o[�����Ojʧ?�������?��4N)$`⧗14\�RFEo)+f�'R���R+��;��P�������R�*���)g��r#&��(� i 1DP3��y���n�b�+0��:Fƀcǟ#8[ze�� �9����\c�@(K����Lhy�c��r�����4d�	����?Q�4�?����i�(����F0
E�B�j�|��'v��'2f����7O1�T��9KP��(�{2�'�6m�M'?���̺�S[�5<��+�E'c�j2�oO&?N�'�a{�A�<v   �j�b��X5*���(�����矜��'���Q�xǆqZ#��y�(p��lH%!�8s
vx@���,{iB}�K^�k�O~���c���� ���^�df��ёG�����'!"䟠Q������'�b�'Rb�d���	�.0��x2Y�dߎ��f	i��Ŗ�?�kV�X��}��dx����T�v������P�^�:�[����"�L�O��rCE�C^r%9��?#<�j�(ީ�� ]�>\jM��B�w~"A��?	��hO�牢r:���Ét����5D�?e�C�ɾxȊ����ذQö VBH���DGe���d�'C�!�nUk֨��r��L�@����Z������?����?AǼ���D�O��S��
Wi�:a]�`I�\YIR���h���4W�F�r6I�U��:}�~]���	�T�sT�

]��I��K3 "H�7eY-[cR4�Q���2cb��F2~q����6mP��B�nUA6J�	�f-h�կok��O��F�Tț5t�<m��U�<(IiQO�!-%!��,U�
���$.�n��'�ٵo��	,�Ms����Ĕ+�r�O��9�֕C�G�>��֌�=%��0��'�:P���'��'�v)�O��(��A��Ʀ�(0���⺣��՝M6����Y�{�]���Qe�'d*e�@�?`�@�e錢���㷅r�����e�(��f	 �xXš1�����ɟ��|�5;!�l=�e"�U�b�Б'�sy��'�ʴ�DӕV�T�c3�f���=剞h��!6&�0Ű�c䗹d�<�2w��f�i���'u����������ʋ�6��8q�	�$��ҩ՟�ړ�$���cN�2����
ŵXq�JYQ̧k}���SDI�^z��0���X_N͓*|��FA`].��6��
X}Z8��bE>jH��6�F�����68_��@�  �<�1H$N�86��DIt-��'��)�)<?� UB靵J~�r�� >l�M;�"O��Z��.�� ׂƞ���Y��$�O��Dz�Oqz��4�`
�	���r`C��'K"�'%>-1掗"���'jR�'�p�꟬�'��0��ڢwzŘ�Β�89��_�z֑�w��n���ȣ�?"�i��/��e��:�	��v�0�y�ٺ�0UX�J�5 �������1�-�����&6�xaG��-hp�N	Z�bp�Z���ĤX�3��ɿC�f���O�=Q�'���AoУ)�>��P'18h���'9��	��F5W,�A���B;g=҄���'3�#=ͧ�?�*OtP8���s ����9y���X6�-o�}� �OT��O�����"�D�OP��Xi��Ht�_׎e#�g
]�贲&�CͰ�I.�=�l�0kS6d���IY�q�򫙘S�M�� ����̔*�(�I7LP%G���P��XB"�Ё��C���'��ȁ��O���0"=^Z�����F�ByJ�h�O�=����=iV���!ӫu�v�!�t��y��	=8�2�T�Bݩ&ǁ�nB5�]�,ڴ�?�+O>��@Ц��I՟4�'e�T��3ϓ�_��D��L�)EYZ���w�4��	ן��.N���p6��v�F��L�w3�8{kٍ^ǀp��>��A%O6 U�����%�A͎�q �x
��B%ˢ2?x!�e�ɜPl<p`�n�.e�"�(өS����B6 .�f�$�'8�QvM�eV`��t���7�d�2�B�O���"���O��d�<���?�� ՐlH��"m@?0�����jם�?�pKN&n*�	0K>Y��<�'@P��:b��ic�/
�tdr4Y�����0'��	֟��'R�Sٟ�_�|Kf�އd���!�a��'���O��n��)�"��`+1h֙Y�R4
4��[���$o�W�	0x+�O��ȔD�N��tX�؍�v��#m�����K��,Ww����O����O��	�6���30�d��e�05��@�dK�̦%�	�l��U�	��?�G�ynzݥi�4Of�3EQ��0�N	"[Z=��%@�l�"(S��'�B��r]��c�������֟@�7�1x���36⒝�hQ� V�q��a���x���A�$����<i��Lnz�A��5Oܱ:���>xb�M�l@F����O��a�'�bd�<J�꧔?!�����4nP� mK�t�+���L��4y��'Ԧ����?�U�.�?P�'q����Ms�.D��|�̓=b�ha���l�(pB��i!�����B�'.�����Ox�ߟ����?��FFˬV�j��[#s���rV��ioh�Γ9�������D�^w�B8Oʙg۟��z�����ʇ�T�a�ֳnْ���lӚ�	*2�n��M�7&�G?Y]w��T�O�� ;�JR�Sp� � ��03����@ir�RA�AEn� hVF����4���	����?I%i�r�¨�ЅźAۢi�'*ԍ%�����X�h8���M�p�O�������a
�I���&땲o����R/�a�<���$�8�#�/Y�asT��hަ!��dyr�'���?���?�����1��l�8)Z��*?'h��P�T�'n�T�8�I����IZ?��l�D|�ǢT�H�\�	�%�����	Ɵ��	�������d�O���'�{��A =���:�����hӾ��+���<�|�'8����i�M��U��.N�-�O֒O4�T�O�Y�I� U��8��B�`��i��՟x�����g�%b4���@�#@�z����]� J��D~���l�� W�T�)���`AFB�a�~LX6b�1z�������.B�I0%�̄i1�X!c��c��̷B�C�	�@�R��GhN�A���NW2B�	8K�(   ܁=���avd׬|JB��
�p��r�G�E���X��u.�#?a���?���?Y��e86!0b "? >ѣ�ע"q�]Be�i�R�'��'���'Q��'T��'�B`�"��J�,ڎ@ߌQI��q�8�d�O����O���O ���O<���O�$s���U]Q���[�`P8㦡�����	ǟ���ӟ��	۟��ߟ82"�'��)�g��)���w�K�M����?���?���?Y��?���?���j�����<O�49�.Ai��'�2�'�b�'���'|B�'OR��5B^�����k^���)Z)SX�6-�O����O��D�O���O���OZ���+o:`�BE��2��i��DP,|X�lmʟ�������֟���ٟH���x��L�t���,��]�FA���@�gG�yH۴�?y���?����?���?Q���?��-�L��E/��YŮ=#A^��Td�T�i�b�'#"�'���'���')�'�蝡PN9|�2� 1��(:�e��r����O���O4�d�O��$�O���O�ɋ��_G@H���G�|ʊQ��Lަ��IȟT�	���	����	ҟl��ޟ�k!`�?�v}`�ět3l�b�.�$�M���?A��?A��?)���?����?ydBE�V�0����N"aڜ"ֈ'|'����l�	cy"�x)`-�� L�&3bd2�Se�Dl�%�b�X�Sl�Ӫ�M��w�V�{�<@Z����̽$J�o��Mk�'B�Iy�_�m�h?i�ꊲ`�|���I�*Y���.�ڟ�v$�9�DE����|����6O��PRÀ�(�����J��L��P �'4�	k�I��M���v̓�� ���mW;i.��� �/�>!s��$�s}Aw�ܝoZ�<i.��<���$5�P�#�F��=%���'�P��P#A�^�I�O�)ܣC�l�]��y�끸~l�AC��mE�� ���D�<���h��dO�������W<J�.ܢ� �N2lx�������X�4����$�7��M҆ �0IZ�e�!��zd�fxӐo�ӟ(
T
Ц9�'e��- N�i$R㺻a�^�1/��8G/*G0ZA��S�'N�\�4�|���'����i��H��B�$Sy��b�\E���(�����|#!Fϡg�v��ā��>���X�O�8oZ)�Mۛ'i�>�{sI�>��htO����!T�T�~.T0#Q�;?AB��\�HHQ^w�6�=���	EJ�"��t����B��?�)Op���W�&(��~r�²w���.Uc�eH�ɂ1lP����6�Ms���y�y�doZ�<I7�$@�b@;9�޸���%s�9n�<Y%��KZ"��.0WO��s�뎗�������bX��`O#'�����OؘyRB���O�ʓ���Ӟ[�Z債 �(C�����$P-�O��o�I�R�j�����z�ПS���p����b{�D�>�r�i͘6��O`�p�l�6�ɢ&V���@�LMa��@�e$�=���Ey>J���[u��Ol����T���4O^0�p`¿Rx�c�*�7g���Ic�ɱ�M����J̓���EW�Ѹ���?�����`I�I7�����%��4�yb���O�u"�I]41�r�ar-��.vf���F^�������~Cϯ�uw �2qZ8�<���BX�Ƅ\3~u�e�/gS�)DV����uyR���O�l+g���$��rӎ �M
c0ų�"+?��iQ�O�9Ob\mZ�;�z�	�Q�|0đ2��b��۴�?�,D��Mc�O���u�Q<�DAJ|�i/iI@�H�lU����������'���'��'b��'��#;����'�8p�B�	�OR��~�n�}��I�h��h�韘��4�y�C�S�(ip3F�b<0���. �v�y����d}��Tޖ8b�v�Ot!	���y����1N�f��Ġ��'z}�B[{��a6�|��'�"�'�"�"9�<�@b�ĀWޜ]�ohe��'���'�剸�M�ub�<���ik�O�h�Y��՝l���w�=lcџ�ߴ����~�&�O���D�d��,�%F�;z����?Q�,	������!������H�r5�b�A��z�U�a�̮3�8��Q�J�%��:B���$��*Y`8���>&� Y���,2p+��v���y��W�iQ�8�DN��<�<��+��;Wf��R�L�j�O�;���2��L�}y�L����h�B�1-�64z�` %})�(q�ˑ7�L�J���1�z�r֡�I�d���HҧBU2!�c)/i��7��>�]��8�^�"V�8e~�c3� "�!�`I=S�z1
��
�U��8�n��=�PK�kܼ�Z䞠���  s�$�ƅ�"�
�Pw��_V� �D�8oh����ڢhU, �p�6��i2QFZƝ�G�Cf����,G8� g�ѴD�������A����k��U�1.�l�0P��d��[�(XU蠃�MS
	�x9�盹��59�
� ��u9sK�-=Hi4ΐH��!*c��1�Z��M��v4�D���b�	����IK�Izyr��F���C���
`��m&f5� ���|"�'��'��I=~)�uk�4M2�I��FM4I�H���h���X.O ���O��O"�-|8��=��J��[�,(�����A�'�R�'��'�"L����6-�O4����0��H� �\c�k�� |6���i"�'��Ɵ�k��c>Y�I�<��$�����ܺ
k������՟��	ğ��Iʟ,�Θ,�M3��?	���Rrj��M�`Thd���a@flx����?������O����5���$�<ͧM��`B�A�x���!�����D����?���|:��{W�iG�'���O�d�'��zh��>ۀE{�!�,*V�A0�S�h��1Vx\�	̟�I�.���U�4�
�9��Z�F���K���%�?���W.dn�v�'"2�')��Or�')�C#T.��$�X-a�kG�@B�ӂ_@��'��i>%?���M�P��Să'J��J���4�?Y���?	Ѯ�������?���?i�;�m�hވY�*`4� XN:�/Ob˓v�����'h"�'���R�m�$#�,�����y��:s�'�R��XQ�6��Ob�d�Oh�$�_��4O4T@+^��n�T��>q� B@�'KH�w.�y�W�4�����Iޟ��	��"���cu���$�� ��d9�Ɠ��M����?���?��S?��'9Bˑ-ud\���	tnxa�f�>=��yb�'.��'���'��L�COq������o�N !���p��a���O���O��$�O����<��{o
�ͧ}U6	X�.�����r!ş`r�Y���?I��?Q����酳=4bQl�H�	�:;r��U�	4I�UAAΎ�=/"��	� �	՟T�'�b-�����'p�d�+Czt9���g���C�=[Wr�'sb�'5�M�,�|6�O����O�iJ�T~�2!���Z *�_<}�����O~ʓ�?a����|���?1�@�|��`��q��]Bvo'�X)���ߤ�?���?���@��Ϥ�?Q���?����b�d���Ђ�wXfi���B�{���*.O���v����3}R�K� ��P�fܤo|�P��י�?���&]m�&�'���'X�$�O�B�'F���Yx�1�k��9����vN@�/�c�]��Iyy���4�@�d	�m^3 GԢ|���$Y�ʽo��������B�\�?��	ן8�	��4��x�? \d��C�(IAXy&�ۚ�v����';�'�V� �����'�b�'<���p�Hb��X���r�6�H1�'?2 ֯xH�6��O����O���[��8O6�+��PźL�ք�2w�� Z��a�	q����`��ԟ\����I�5+��a��h���r Dq%��[$艑�M���?a���?�2R?��'�r��.&�d����H$$?��w@��EX�'���'�z����'��'<¡�}a�7M�tɐ$z�L� GN4j� Y�%�����Of���O����O�ʓ�?D���|"l����h��k�%q|� �Ǎ���D�O��$�O���O�`��I�ߦ��	� p�듾�RHk���/y�.�X&��l������py��'�1�O��I������	�J6��jp N.I+��CNF� �	���		Iz0�ܴ�?A��?�'ZVԤ���ι% �䠘�S�t8��?A.OL��[���I�O*��|�!��
_?�〬�^N����?����?	��:'��f�'�R�'��d�O'DP����tF�2~~0�CIK��ٟ�1�L�x$��Se�$N)��X20��L�4���bD�?�-Z&U@���'�r�'7�$e(��O����b��{�P��b�)������Oz�S`-5�)§�?!c��N�
��a�f�;W��or����4�?9��?�	ؕ��'��'�*or*� �o�<��tٵ�ݒA�r�|rL�G?�O��'�2GA4@7�і[�x*��u�E|�2�'m0=��"���O�D=��F�B�RTST�ч<���c!OV6xʓ-
�ϓ���O��d�Ol˓H�1� U/^.���� Y3�3��?
�'�r�'n�'�b�'bґz6��.�ꅸ�-#�P�i4��y�^���Iϟ��I{yB	]4A�����4p�zѯ �!�d�)�k��
������Ij������ɨ%���	�	��+�@� ����\�V��'+��'t�[�(�C�ӆ��'b�J� ��A�Q�QzD�۞Y�	H���?�M>A��?�,F%�?q�O@h���p�6��5Fɜ{�Pu�v�'LR�'b�%0�0e2I|���
�'ϳJ��L�퓢ZX�"Ə�����?)�uư�Γ����TMT�"�0��$) ��­H!�?!*O*��*�����O��OY��@��d�s�	?͂u�qŁ$GHH�	Ɵ��Ʌ��L�Ie�)��%QT�!)Ǝj�XL�R�q����'��p�g�f���O����� �$���I+g��T&�ݖ8E� ��'/��4���O�e��K�)§�?q��=�Lp�D�H jub˄
���'�R�'������1���O�����h�뉩P[��BA�/��T3���O��O�h��?���OD�$�O���M�5Nb�s� S�6L-:���'�R���o$�d�O���=�DÔ��eRe9 � �:W�ۮJ��˓Ť	
������OR�D�O��>��c���k��cp��dt��PO3z��'���'��'���'^$�8d#����8� ��*[�R�����y��x"��(�d�b�@��$*�+0Ҩ)���5|����Ga4>��s�Y(Gq�8�.^+r"�d�O����O�O��D�O`��iP���q�.R�65�U��N�Ot���O$�O �'����'!���kd9�e,�<U�x�B6��y���'��'�r@پd��,���3S�B�)��v���[%OG$��E�FMگ$�,��1�<D����@N#eS�O��^�()	�A:�1s�48��[y���:����x��pF��Pr�%��
��ldܽZ%�Q�!��I�dD]���xjG߮[�$���H��|*Eh��X��\���h�̪z�1���u%��s��	�m�\��K�P{�i�7��:�ɑ��"[Z��V@�EDdHS��"d�ku���!Y6� vFt����N#�qke)џ4���tJ#�w���R�j�)��0���?�=i�
�|��qI���+N^"�ㆌ�,o�d���&I��V@�d�,�q+��j�����S��d�w[!	�����F�
��@p1�$�H����$?il�%*񰗬�h܂����Ep��i��������� !�fiطM�Z�l�aUԺ�p>I��>��'��'�]��j, W^����z?���
�]
���'w�S>-2��֟��	Ǧ�ڕ�d/$	����c,�l!��ޫUH��D�3LDO�S~��%�2a6V<�L���=el�X�H~ӆ�˅-�O��E'�"~nw����# �	^���'�ƥ3x�7�μY��i�L��j��i�,0�'�(��Tb�X2D���C�'b��'�F42�h9St �s`�Ѯ;UF�C��B�'��p�&]PU���f7p3���Ed&����?� -�.O�$�b��?Q��?�����dt�D)�e�_�i(��b�e=��W��� f�,�f��"�'�̹5��K^<;"Oӵ�x��OFt9a$�i�l!�ϓI�� !��\,�AR�ȁ�F9��'|�������(?��OL�D�>IԎ�q��y��K�)�f����US�<I��(�F��CF��#�F�1S��$�n"=�)�L��r�x��M)�t�F��[*=�2�<B�؄���?���?iD)�?a�����')��CF�.�e���Z��tbG�J :����q��� cۣ6�L���#L��X�v珎�1h�H� hp�ZW+	ԨO����'�fON�B��4�=U
T1#�^#P�,��O�˓�?A�*��	���U���+R��=N��%"O�  �I���&k9��"郄a>VHc �OȤ�'��	�=k��A�4�?����i[<���r���.+��p�őwA��3�kL����ٟ\IE�V!c�P�G�4���XR'KE/tuz4͜�{VX0�l�@�B�y�hQ��	�/�]�Z)��L� I�_��p��BE:K��C�-��N*l<X�lރo�:�K)b�'� ���?�H~ٴtwf�f���2q�#��]��H��'��O?�R�;A�A�1a�&��Q�*���hO�)Sq�Đ?=�2�[%b�6�na�EDݺ]O��S�1 $�oZ��D�It�Do��Y���'��6a�	G�0��ץ��}��A��PV�	.2J}�p��o"@pD
e��p��9�4�%�s�9 �b^�g��2�2M	4`k�Fp��pJa�_R�� ���X��#�I'��QP��\c��H@"��8/d<T��ĞMε�ش
K���	˟T��'��&AlM�7DK��!+5�ʺJ^��jt��!�o�0M1�A!�	�7)\N@�=���Qؑ��Sݦ�b�6=Аm�1�^�����G�+�?���CL�X�U0�?���?�����ͦ�1F���`I�m@�	op��r�J���	�+@/�
���Fٕeh�'loh���F!���4� U`#�Ů}�T��-�1n(<�@
l�
G�Įj����Q?�#ۤØ'��$�T��o;�|3a*F� $\���k�O��#�O����O�Y��	P}"�!yZ��Ү �~��	+�)W#�Px�i�(��G���4�~4��
�>T�fi�t�'
���'L�	�ʱg�E?Ԃ@���ʿ{@�$��Ȓ�x4�0��'<��'���_��'|�Z>)� )X2��^�����!�%0�h=yv�"v����lӝYu����rS��`���+����$F�:l
"��6A(�� ��;㨙��l�P��	18v"P@&ŝ�#e��@!>vx�''�MK�����O��ʧd�*�;t�$�x�v�Ȕ1�f0�ȓ~��p�+�8v��5��G%����.F���[yb��W�֝�T�ID���7]	����f;a���q�[����`�O����O������	J`.XQ�f a�hy�"&�l����$}nx@f/
z�M:6�8O�Q������M���e�
ZB�ke	J!x�(��T�\]tp8�#��K9@����H�Q�̈d��O�xlZ�M+���)�,��MaV�ݘu��a�O�(�D�IX�S��?���>*�� 	A�N"'�E`�l	\�D*��|���>ᡍ�<j�,! d�OH,
���.W?��#H�l~�f�',�Y>�Y���ɟ����%T'��o���j��-��{�b]I2|)مNB�A������PO��ا�?��|�1��8�⃍g޸����H���oچ#�|��.��	P<�Ґ���~X��0�����P1�F4D��d��G�d6�ab�i-�ܨ�vSɧ���C_�	�ց�B�N7���)r픠�y��9���M.Y�$z�L���(O*�Dz�O6�FC?r(��s��S�\=L�0�L
 4���O��Q��4�Z���O(�$�Oh����?��5�R�P'+��p� X{�D!v���ȡh�N�:裇�I�k[J�K��~�7g�h .�OfMa ��C� ��s(���l��IZ�?R4(*5�P0�8��n�h���n�:$8�|R�Ө/�xr�k�"_��+W�<l�$�D
�g�X�����ه]?��?�Oh��Nb�4�b.Tˈ-��
O�7�cV�%�s�d��1Ja��c��ʉ�D⟐�D�<	�l�=(Ǭ�kpf�#>f($�"� 8<�r�OG:�?���?A���;��?�O8�8���MSp��>��*�Q:2^���u�\MX�<Pdm�>qF�L:m�]P�d4X����IX��7��O2�Ig�, ��ɻ"�U.�p��&��y�%��J��i逭)7�����y��Ł5�X�$*A�y��Eq����~2M'���*Z0��4�?�������0�HU8�gB�D�
T{��W?9J��0�ǟ��Iퟄ�h�0/�{�8C���6D�]�p���>��);�Ê�М	��+���+բ2�qB�:��89���˶�ݦ�l=_�$��`@�`P č�&b�ڐ�3h�i�'�n����raQ>5�,�	q��R��
�j �y�%4D�0GN\.�=�ސL>Nԓ�	&}��i>�	N���ʒ�:�
M�cA�3H
�駟��ʕ��M#���?(��ͩ%E�O���k�e�夓�HK�!�".�Z��"1�P"v&�a*�����S���iu��p�N�R�(��ӂ؋w�Hy�41�J	HW�>��S��MdA[>Y*�'�#f]�h;4H�a*`��O<�$�O�D"�禑KQ�4��Ő*{��Y�c���t��ZX������Bw>tJ�h��`�R��`"ʓu���'=�؅A$�K 8<a��OK
�Ӄ�'�"��E:4�1P�'o"�'���o�%��ئUCw�-7C~��@�����5(tp�àƗ�vH.P!����La���d
�G'����mAp�Z�+�"� 3!�Ѱ�V8�$ʳc��f!�n& j���~:�]`"В�Nݸ�~���?Of��A$_(jj$��l�?P�\�$D���Ҧ��Z?˓�?I�O�P`R�T�sC
� �D2q"
�P
O$6m\�z"`��
|B�ɑ�àt��YS���F=2��<9Q�ݣ�D� ��;�M՚�V�M�8~�%�§������ߟh�I3���	ȟx̧tEA�%��p�ȅ��ܜE�^+�ϒ�s*�1��1X�u`I�,���qT$1ʓd*ʡ���*k��d1��G[n[���f������C��@�E,wrl�(uh"�Q�&����B�!�e��,-Aզ�1K����2"O�U��#X�A���?j�p���'v���	� P��
a�F�|��￟|!�4���M�i�1O���ʮ%�m��l�rQ�{d���'�ў��s��7��dQ���;7���	� �@E+����B4��ch��v���˥Xs.���lB)_�xl��(��={!�ՓH����0(�/@�&�g�� �!�$ûv���6h��p`���܉\!�
M�@��C�7�~�����/S!��6J�̙I�����U�x!��R9��HA�C�<1#'X�S!��1^���P�^�Sʼ�1���p�!�$���baJDL�d����G�0�!�"f���p�
A�#�4�	�%��C*!�dҊ��������{=�*�D^�@	!�$Ʀ``��wݩ�Lɒ"R��!��D�&�M����2z����gO
F�!�*�ԁG-��lYy���(5�!�L�T�>m1��N�H�6� �"!�t�P�`��&dGH��4D�]!�$��U��]�DO�%���> �ج��{����ϟ1�X�S�8~��m��=ZBT�1�����@ ��?e�Q�ȓM6����Ż>�o04 d�ȓEk(�;EA����\��GJ$P�a��ɐ'.�ͩ0m�I�&`�>�ڐ�0b�	5�}�2�&T�2؄�4�h!�6*@�_�fq����/�<T�'���FK�w\u�������>��+NM���в�X�:���p�,D�L��m
c.T�ro
�{�$i"��ԥ(�~�(��+!���+R&p�D��qO�l2�HO9$��T*!KS�c��`B�"O$��1�0j��v+(@nx
�"O^h�d�	'��!y	�D��TO���TM�8 1��Ʋ����v*,D��DF�6l�v�Q�"G�i���a�m�lG{��\b�OB��Tg>i���Nf0�!�"O*81�D�{���� �H}�ES���4&Z�<�}�q+
�G�:}سN^�H���$�Ubx��,OV�dd�&� �'JJ�@�s�d^���<A��C�]B�A��1s�iS�u�'6�)F��J$�6�S׆A:>��8qj�//)�IZ	�'�X�� ��fa΅j!C�B��ĊشP���S21�@㞀(#�Ptn^ಗ%ݞm蘿��d!D��@ �N? ��!��]�J�Ju�rN�>	�'��\b�����-1��hS���yӦ\�EH�#!�!�䑲CD
`E!G��:� �ș8��O)��'��c�o]�wU�5�k��$��(��'	z�@"B-tr�0� �U�M�%{�)G+�Px�-E�4`0)M)6���a��0��<IpI�i�w�z0A���c��O\���ȓ80���R��&� ��͆PU��&��05�-�S�'tw���uǕ�m>�P�(�<)*\�ȓi�����Yq�n�8 h�	�L(�?�p�I8��{�lI1S�J����$F04��'[='�qO����<qbJۊr�~,#��+t� (A>v�����	�s�����C:L��U)ʳ��9�&��9<��P�鉃�T��˲b�8dp��m�\5���&/O���D6K�xŠ��>y2���H��L�t*�^6�e󳏖T�	 _4�#<�}�%JE^�xZt!�H"vP�3L�K~���(�H��؟��@E��S�P5)�P)ۍ[g���! �1��'2h:�"V�[��&P@��aPWx�`2����X��[�f���!�3�d]�����#!�� �2��Ԇ\���'B*l�� ��c�K|hV�aԨ��X���p�:C�0t��ƕG��Oذ��}��0#���u̙N�(�����O���j�3b �
0H�6��+b�xYt�&*����{�O��������X�qQ#G%>7>�y�*:��������F�e�����f�Ou 8���($DS4nж!#�ڎD$<Ob�aG(��5`��/Z[�����s��d��'�H�5�H�	 �Ϙ'��m��/@�f��bFM;%4�=��',�y�o��k7R�%�Wr��� CS�x��Ҧ��TzrQ8�'	",����u�ހ�3��M H���F	q��*��&R5>,�Ah>a2��*:�	���S7X$�� �:D��+�	M�D����E�?Tdd�&�<YӇԒ�x�1%��[�qJ���Z
f�	d%T�jX������ִ���v 
�в��J��R�/T��:�!wb��,��D�}�h��w)�;Vl�O��;u��y7cȯd.��׆X9a�vP��#R�x"#�f�J|��یC�.� p���E*�P����l���y�(��
��@Â6��UJ�{�)_�0"�	t�؝��A��p<)��!�%K7.O��yrg��� �k�'!6��k�$�0�V��0�R�56bh"CڼO���$�-f�6t�Ĥ�����I]�����Q e�p���ɇLH�c�-OVމ)�,d�X��
��Ki2l��&��%S����(4�08�j9�P�Bˈ5�-����c���
r^H���n�I�
8��݅p,t��O
�l��w"pHrd��7T6l�b�.���2�'a.����C�eN�
�A���c��C�~�*���E.b@�I�(A��OBO\�y�,V�O�٠�iƏ!�rOX�I��W9d��+�KM�e��� !iI�`�1BQ���u���M�n�Є<,Ofi"4�ܱ���M]5t���I0r�~�����r�*�q��\���G �;��¥'Knpq��C:\}!�%*[i�+�B�-�&)�^���կ��Nxu�ǩ�;s�6m�� ��_��U�$������C�O����3�l#��38$R�2�'sĜ{�ˀ��٠E ��գŧ:`�T(�
�KR � ��_w̐c�;��Հd��"��۝w���J�s�.�c�&ʟ�Q�w����"13rA���:8��a+ck��pnej�CV)�
���Y57�x0 ���58h}�� �?��O�|!��ϯ^�:��dO
�/�,a���#)[Dy�S��1�&���
;FB�be���p�ߞR�Y�%���FM�W�؁D&���A4YA�����9"2\�g��+S�XX���<<H�&'D���)��Y�M��,�w�Ȼ3xRL���	�T�����-M�}p��sg�9"�04쁞 �"��dL�1�DB�,�L�+�`@�hjP<��	�R'n�:`k�T��&�?�	5bV��\��  +kbD�� �U(p��$%j�ճ�i?'�\lh��]�<D��D��Q j��t�L�!�|������"48C��?4�� 2���i��9�� 5I����&�b��vK�8 �<�Ō�?|� )���|�zZR�E�'�$�ZV�^=y��A%�=W2т+�a�q#�aQ׮�:����}.��ֵg Aɀ)u��D��0LOj�qT)A*�D�4���]p�aE�i쪙�(O�X(��A�-0����+U�N��	�<s���>ꦙb��I�0<{�+ܚ`VX$a�@ D����_��0�kۏbr���&�f�d-��N!(����a���<q�֐\��(���ml�l�ü�i�TE*y��JB�|�ekPfX��ٔ+�"I:>����
K0��3O�-����K �C��DQ�<+�H�R��>�b�OB�L?���%��'�������w�ڄJE��(��"��]���3��fb\�Z�蚗�j��%��8j�E�F�e3&�:�]T���s&��j+�m �C+�}��	K�0M��3阺k�ک2�i�@����w8!+���rN��8Q����F��s0)ϓsJ��p�Nh,��/U�Pע8�T�4>g�B�I�4D���Ŗ.A�냫��A�~����Z�LH�rI�?�R@����ʵ��$G�ɹ%��b0��L�y����OA�u)�!�)J�a}r��+P�A;"c�HK �GP�Q#����^*�.��'��R��Y�`�L���i�'"����H*J1Ob�����PB�dZ�q֢�٢"ʓ,�(ܠ� Ƣ1�Nm:B��wݰ��b�n�qcC8m,���ʘ1W�q��G�< �'&�.��C�@:LO� �ET"�,4PP��5��lP7�βVJz�k���� C�̅pJ������6�*nӬ��ش9�~H)��F(CE֕����H֨X�V�N�<����Vl {!���o��T�pA�4-�n�	��2�8�V�J����M�)7��@`'�4\^4@�P�{�ڒ�^�|�z�냘<�8`��<�O���A���Q1��R�m�̹���
b�(8Hu^�,,��%O\�4�^��������P#�n�K[�$ێy��+�� ���aA�ճ����O�����ʺ:X��9��H.͜�ӗ�X�+�����E�/hN�d�#��!7�|�eD�s����č5=�)*�k@6SXaz2J�&n��3�j[�,9e#��4�u�v��t���`� S�V9\�0ê�i��)'�����O���h��]+l|�`.�^u��pb"O�r��Q7�~�I#��5mF`�mʢp&8�+ל�MӖ�iZ*7-Q9���e��~0����
&�y� �� �̓��F�ѷ�� Q�����'n��Dp�D$�f�@�9̨Т�A�)u�f��g��7�
�o�XR,�kuΚ�7�0x*&{|�mٵ%B�T��j#/�g}B��"T~�@0.Y�s$|2$ŋ�O��HA��C�������1s�V�X��	�- T
�s��i���L�s��yP�[3U�Hg,��{�Ҡa�_���%se�����O�|S��)\�qj�lԹK��IA��6F	̼���[$ �\���\�#�@+ ̪[�]2";�M�2$��l����J�r���8T�-E.�k��
J�(� �=�O^���ώ3vV �g
$P@�D�ybI�6|^�$� Z�`D�$���0c��Oy慸���n����a�A)�lQ�q��BU�a�a|�S���8#G��tt����j�j$ZB"�B��l#�H�b��p���Ƣ$&`0Dȋ�cz��Pv�ɕo�|�B@�G��p��i��r��	�)�t�H,*x��S��I~�0�a$�]�`;�]_椉7�RG�Е�d��k_h���K:=�<H�N�H�*W );�5�teQ�0��&`��tGz⏆�:4�+Ǭ$�& #Gh�(T�n��Ã9w���8r�C�t�<�"U��9>=��l��'�04[�8O~��c��)���1��?i��lFp� )1�OlD��j[�o��h��"��m��Ѡ�,�9��%�f�K&o,I�fL��Ě,-���p�!ڱs9vϻ<3�+q�W=)�K
��l���6�OZ��E��]rp�{G	�%�e匰o�.y��J�Z����'f�u+FI)R[����&B�ڢ�4e���z%e��Mo���#ȲT� �ā�)D:�rb)�i�'�HY�ad��/v�A��NU�i�dU'J�i*��ɨAz��עS&Mm�Hc�%Uޞ�bT'ϊ{"$Y�F@	3I*u��*Dv�"<If+��#k�H�ӏL"1tM�bg	�T#�FK�8��J��-y�,2�� 6$f�l�/�#5~��.�Z�!�f���D����WI�`!G��%` �y�N�RH��䗼3��ذT�Y6SA�m�7�� A�f�S��̎M:�]K�Y�~\d�NerdnZ�VJ�a��#G�|��� ��x�c�oSLu@pJ�Ia�~�&RX\�����"�Pb`�N��As�I��~r�y��J�1������H�t4����I��)y	I�8X�dYUH�u.x�����lE8���z�'��[��L\ɶDc"�H�zʑB/<�&P�aU�	���R�&�r��;�lӂNi�`*I�CgHlYw��=� 	`�aV�����YM��� �����'_2�J�D'DndCȆ�E�"�2F�Ӯ$6F�%6�h8k�H�P�B9�1�� �d㐂-���q��U��`�@�,|O�D�p�He�vq�#FH%Q�Rܐ@��%p��8&�V�:k�H"�'w�d��<�w+ʜ7N2��%b�:aG� 5i9�d�+b��s��y��2Iď�1SS�x��P��?yAN�@� Uō8Y�E%D�:Q9T�²U^�T؃�P�X\L X`�U�DQ�EBRLf��bO���=A���\|ȑEe�(��a#�c�V��=�!�ն���vC5w38�Q�
��$Ru���-i>�u;���\������?10z�`ً�0��5+X�Od	��!�{kr�B3*�v�<(ے���px��_�N<Ta�-��hW:�rp'A6[��M�D�#�O]��eU�U��9��f,O���i�JP�+[Z�b�l\�Ii����'��Y�Jիe�IJS��ZMܼh�w�&��O�,�)x���	P��\H�'����`*��AwR4aԃϖIX�O� ��I�~�L� h �C��	�%�v��r�a��j�r$���	�*��"�g����>1���z��u9�+Ŋ1L�Ѫ��!=7f�jCÍ%�V�Ӕ>a��J r�>O��,D'�R ("�êb\�a��	�5�����1�'=+B �`�K��Q��,$��ȓ8O6�J`A�/Y�#݉C�.�ȓdH�jǯh��D���I|����8򖨀Ԡ��s@��U�ʋC� �ȓ9���j��ҳc%T����!��Y�ȓ Ԫ `U�pm�Y2�	�"���yȐA��
#8�6���KK�9}���ȓ3��!�ESr��U�	�4Y�ȓ_Π��b��-2i�A� ɉ��ybBX�5�t�ul�.�@��`ĝ�y��Yr8:XA �]�r4���y��X!*�P\"�g�<6"Np�`b�;�yF�d�ֽ�T��,�dx�0dO��y�d�4l��GN�"H���D8�y��͕.;��ȷ�Q'4p� �BX��y�JQ�k���&�I����{���:�y��V�3KxB�#
�`��z6,���y�d��,�����6X�d��@`8�yB��??\I�G��(��I��Q��y��MGV�	�+�(|S���"�y㐛+��� �ئ _�9��E�y� =��1�®11���f�Y�yҮ��!�N40f�6�0�&μ�ybH��7����3��|(���%G�y
� ��P^�2����b,e('"O��;��	~�E�a��m�9��"O��� ȇW�$Ui��D�pz��"O�8d��$j}8���CTz5{�"O�[㫆��y��dݪv�M)u"O.�2%�/�qh��%a5���%"O����%��ʠ՝Y�f���"O�8�'A�8�yXwK
e���rg"O�Y�,�p��M #4�i+"O��z7��$[��RG�ѐsP� "O8��A�@�{`�����~�)�"O�<��G�4eJް)g�IE�PP�	0v�t+V�u����{�H�I�P�dȸ
MfV��2�'j#B�	��.ثl��S��!G.��B�I =�̑���dˢ�9�@�;x|�C�I'��d���j=�nT�-��B䉾7�Jh�f�^9E���V"�Y�<C�ɦZ<��a3��
4��ź��'	�rB�	�s����a�0L�	�$j��k�FB�� @���(�-Wvmz"�NV��C��6�P��a!ZZ^��E�=
F�C��z��R�˷s�e�(�,}�C䉛ZN�ٰ7eL1z����8.�C�	" �nɠtct��$^��X ""O�ɪPHȎ�	�$�N$��"O���$�=R�pjf��
F@�V"O�%K�N�l�Nt+d�O�5��V�J�<	s���
m�p�M�'״BrJ�K�<��ѐ>S����n_9*�!��H�<1��Wssz�{smB6��큒�M�<y�KE�(�$�F]0dp]�4��P�<1a�_i� 6�I.C�4��$ȁL�<Y�/�3=� ��%R�$UP�i%�D�<�6�W0V����刼ќ@����e�<a�WA,9�<Ot޴w�_`�<UB�5�pyk7/F�sD�s%h�_�<��m�g���G�5wl����H^�<iĮ6a(��R��4(F��0�^A�<�p��)"zL�4��\��X�ۗ"Ox͈�i��p�I2��Ab�`;"Ox��w�H7O,��R�iީpB�1�"O:��f��5- %2&���"OP��P��+���!��-�p"O���EH|A��D�V@��R"O`K��;3�29e�+}��Xs"O��S�LT
~��"q�B!Aj	[B�'��	0]� Y�UB_��m����ͅ�s�^A�ע�PF;�
+;�q����'玙!�����5+���+��= ���/����	�'0��Ge	*{��	P���R�U)0+>܆��7�.��O\��l:��O�d�$e�C�{�`��>���J�';<ջ�G�2E���׍�����;NX��I0�M��ˁ>#�Q�r���p=��O\;)  ��g>��rk�`��~�Z`���6�AF+�9E��}��ƪ���G*�̹R!�T�f�L!���y�J��6���@V�c�*��¦�A$����aS�h�d�9Ҥn�Y�B�[J~�w�&�K���i֪��e��6"�����y���a�>ź��O�������;�N �O�Z#Y�7��4dȇ�^��1�Ğ�U���Q��8Ă�X#��6�1O�[%��������M�0� �������<aC�0˥E� �($8�('*.`bG�@ˡM�5@(%:� G����@�˼+a�,�P
љ"�LucoI�kT�͹nقO%�+f�D��������i~B%Ծ(F������'s�9haĚ���x�$,�|YȔB�l��Jԣ�NH�ϟ�li��Dz��)v��!��/��`�s$Ҩvf�x�K�t/��{��>��<y�C�,� �x��d�"�hC��/������ �fhy��Ș'gfi{��6��0��$��a� 	�y
� �E���s ���c�W�d	mQ4�|b�G�ɔlR2�F$z�^3(�>�M�$��m
�ԉF+T�+�� �4뀌eV�@K��$Vy�7�3 f��4|P����']�#?����|3J��rJR�0i(�i�l�X� ��1���K'$	���6�����<�J���O,2�'3p��a���q�>*FJη1��`�Y���	]f���͡3��b�-&z��g"پK/^�2��~��T����
�¥�i��Z�ȈV�pĉ���T��'V�hHa�	^X��XU��f>V� %�'s�(���d7p�B��<�����:t�oZWp$���7R�f���w�p��k��V TH����C��{�Љa��ٱIGL�s��).˒��TJ��дf@9�uo�3\|��A��N$��c�hY#M�VX3�4w?"��ױisX0X�@��u��7�G�V}��*V3f	��"��}�Js�c͇h+b4a��ɀo
��ůL yV|��|�'k�i�8T�5aI&#����֩t�|���S����b6�'�:��DD�#���b�n�3*�f��b�\;DĴ9 �B=Vo�<��aN~r�O��-2m�.��c��k%�Fg����`E�R�xҬ�2�\XƏG�y6I���+��3A��P���F�y��<���V�96m�;|�B`"�
:�����+pe�%@��@��M׍<�=���)�DϽ\�h<���i��� �I;H��踕��'���&\����`B�`8hWI�)aBRi�1�i�lA�D�,Gm*H1!DX�?������_�j�꓁l�M��Mܞw̨Y�۴ mR|0���	�����%?��O*�x\�����Y�[��B�_���/\�����<�}��Xy��R�L�'� Y+����>����Y
`���y��զ��O�T$>��e ���Ԩ9U��?и��s  9=M�����Q8��u,}M��X�B��f����k�B !��� $��[`Έ�\<�	�,=�!�n���ݴI�pH?�	Z��Ak��O%R��|*�(*�ғO�}(�$ez� n�(����'�@�H�?1x�h>4�Yu�]���Ż@ �w��"�.��s�L�g̓�^�`�ɮ���kٮl��7�������/�Mۑ-J�Q�&��|ڑ%Z�<Y�D���,A�K79�=�p���V�H%+ta=�O
����ئe�ȣ��׶_t���N�Y�m[t�O���7�F�B���'r���Y��nn4YC �8[}�iCgF]�j`�鉍^54�0���N}b�ҟՊaP5*K���3��.r�(�+U�&#���a<v��O�B��?�I��2r��r*bı� ʣe\1Oİ�$ڃ%���;P`�QO�h*'OV=pR����E��9y�l(kћ�>���M� �D�Q���y"V1��D����QbJ�CU�dB`�4�O�W�/�^�? ��'eN��[Yx�jDo��]��=z��-Ht,���W�t6����Z*� �0�ȝ,���G&�y�'ِ�I.��	�D�*q��$+��ց
O����D�2V��RϓJϠ���L�C֛�`�$ET|� ��jy�󡚟@�*c�A�7Q�">a�I/�>U��D����I�RL>тb��_���@4�%�'?P�`?z�1�W���Lѣ�}ҁ
�XHV�+��ޯ~�6�iQ�\58����le�4�����&w�
���3��Qi��[�A�iNt�I�d�|F��n��Jř�L׾��=��[�Z���ioӛ-�n��Q� 3z���	���Y3s
[�}ݼ����9�:pԉ�77��u�W�Jd��oZj�*q�}�U��Y1w��G�5�ᄘ���<�tЄ#����m��{���I��@P�>*�`�톫A��Pk�Y7C���àCB�~�Z��R��Us���0z�:�"`嗉a�q)a�HU~�ģm$�KrK
�Q�Hͻ@Ó���l#r��s��u'v�zШ��?�~h��"�=�xY�b�����*��.w���F�<P�t 
���#^/��v�,���QA��p<��Kߛ#(�΍���Xb�?>��+4���<i̩�"�'�@`�cCιF�	��4q�Bd���i�A�6��A��%�x�LL�!��a����W=�p��h������|:lE�	U�&Y�0�nӐ��O�|b����)C�fY>2�Á-�6c��5BA�= ₨+�e��0=!��01���6�,�8��N�3J��	1kΆrt* �6)�
-�4�d�P���Lhǧ�m�"6��#�(�jǾIm�uB�eC$U�rNee����S�`	�dB֘'��a�lR9g�ARR�Z,.�.#h�d�6�#�F&!�¨�6FFΡ��T ]�<���*�����@�T1���#��]�X��e2ړxcJm3L�w:���I)�\��3��S1�Ez���)?��b��ԛ<�ZLq�]��MseBs���9��HK�ps�����lC�ά1�������2 �v��t�!�(L�����%R!�A�H�7M�M� �'���`�6h��NϰAb�A9�ρC�V="��{�ؘ��-V<&��=;ؘ�#.���� �	���H5��bAg��]c��4� x��U\%0F��Ǧu��� A�t�(��ԠBFp�$��OJL�c�6>[ڑ��D,n������|��T. ����Ԥ86.@�7�;k�\堂➫-wZm�烃�$Z`��F�/��Q+�'J��(�Ȧ��N�o�P)�/Z�PR(�	�6ړ|�&eXe*	�"	�1��ę�����bB�&�)��ŌXQh�8&6D�"��Mc���S�	Q<$��{S@ȫM�Y�r�J�M+�AV���w�a}Zc���b B��p�@14�ԛj�r�i�*O,*D�H-G+���Z,0��OF�:��Jp%D���h��K�8d��Ùm>�rVEY�V��x���L�L���I5%�Z����	b���R#�E  ��b�B3�9c���.1�N$B�H�R#���o�&8����Td�- 1�'�I�\�'�T^��Q$���
�(�Z<4��@#A�XP.��	��FO�^4$�A&@!E�Hp*0��b�? �t�cW������ּ\���X�mX�y6p�S��/�h���د]ax�֐9�j�#nҦ#�d�B�`�
Z�`�W�V2`6Lx�I(0&��Uǲ}z�a���O�]���ȓ!�"m ��і1�1�P`��_�a}R9�Zh
3�U�a�-���@����4�p ��$D��6-�,�&�>�;�64Zi7$���� `���tLZ8c���sџ�a`��%r��0k��7������'(�$�%-©(R�F�ӵ� �1�J0[�2�ʲ!ԩe,(}�S<c����%Ӌl�B�X�W~2,�G@�<�u��$;��q��LK����ơ2�ŁÉm=~�C��g�|<j��_<�� �V�֒<L�
���h��U8���+ �=�%����^h�� H�I� g�#x��֛�\}��V���Mh��ߠV�`�+t��'y`�u�ކb��-*�
ǹFL\�7 gӞb>�+�K��9�r�@Ҡ�HE��Hכ"<-��I�&� 灕�\�x$#�O�9`�E2%a�,vH��U�F�iô�L�4L����тa:�yǀ»G�̐��XY�R�:����p>I��D�s@r1�t�>1�F%C����Nܣ��p�V�S#kU0`���	d��?^* ACa�u2V���@���!�ry�!2~s�7A���3%�
*�(O��`�)'M�~q�Y��1!Q��1�	]��F\��	,r��`o�2�)TkȨ+bP|#�M�![A�g�		r�@�gj�/4yZLJ��J<4� s �=&��@��Մ${걢�Ki�'�(�SGF��C����%�/�E)D�B5�ȇ��,�T���a��F�iq�g�L�6G���p=�B�ɕ�y�C�2�:4���]�y���k�[���>Y���d�t)QBJ�F����텨Wư�d���E>��,�%KSp��JĪk��i0�L�>��e��+{
x��];M�}"P/�T�'�������ܴ�p��Bu�L���^*�R-�'Gp��#π,Ί��᭒ mU�yp �ѯ~�������O���t��3ܡ�%�Yq�`��_��r�b��8Pf��V�b?$�)1���X	�B��HИ[�}���_���?)!g�����yK��v&Z<�BݎR�=�� ۸0T�nZ�g|R��>1�O����^�x!��W�{<�A�$�"*�!�dѼ2�0�蓠��t�-b����)G��S+���IW�D���f�%d�ɬ�6Ij��؉O* �ӕ����DP%3Je�.^=�a �9~����nY��M��
�=w�%1�GN`�,)w.L\�'P�<��D�!3@(�� +Ϊ]P���كi�T�5������?�-͋~��H��,�-0O8��d��{Pҽ��'��h �g�]v�T�������c�'(��:�	���K�ӕ!�p�%D��5���A)F48jC�	k��@�閭u%�	ڳA��A��k�&`�&A�ɧ������%n҄�vH�`:��o��yBAV�
�Nq�\7[���!\�&	��;� E�Y�%�ҭRPʔ�+z&��\�r�����t��r5�ś8 ���� -��K�_%6�R�FO�1@,�ȓm}D89�� Z���J�#�����/!N���i�Q�����Au�-�ȓ��Phs,;E��a��>W5|���q����D��")���9�m�/��	��)$�qZ�j�0=�8� 
#L���S�^$ȧ��D,� Wm
I���8�
��&�)a�t��n� 6��)�ȓ\bl�!#�NĬ�K�����ȓ(%^YÄ8WD��*�CA�~���ȓ�@t!ޘ1sޑ:ԆV���ȓs�+Ԏo�4�V
�PA�Q��Z6>9فO���rݑ�N�T!�@�ȓJ?ɱ�aM
�~E�"��F�n��?�e9���?@*��d�I,E*H��W=�S7F̵Yp��C��+R����t�YF��?z͘VͲ)Q\I��~�������!m���$�u}�u��L'6��A#Ѥ����!.&s�Ʉ�nf�`�ؑؠ�@)�#;��h��n�Ŋ��{k���V��~�\��ȓ@8�"WA\�}��&��Fԇ�?Z�X� �N�R�F�	2Z�lŇ�x�$L��d�2zx�y6�ɵ�,���S�����쐝v�	c󉈗bԔц�(Μ��Js�� �&�!��9��S�? �$!�ľJl�̚�j��0�ځA�"O E�!G5-�(pw��_�����"O�=ɥn�D�
1���.Z*U�"O��V�A$Iʆ�#��bD��"O.��RAh�hH�B�l��"O��QU��
m��QE� p5���'���UM�A��Y�>��*�'[0�pU�՗b������d
����'՜���
F�_������6�)��'"DkB"�����e���\T��'V�@���߰$��$N�[^���'i�ԃ���9� C�-�;@��b�'���: ĺ���P�(�:@&���'��4�$�C<8�N��A�6����'	2)���#>���f�ʰ/q����'$T��#U�B��j���%-�] �'�.��5��}���j��+��1��' 	y��̡8���!Uż8��l��'���1��?���L��@.��s�'<��c���sh�A�jۅ:1�P
�'&ޡ0a���o���C	5V��'D��AS�U/"��`�%8&&���'��Tx��� �`�At���9�'���
��g�0y����;_M��'0�J1'Ï-m�1��	I*�Єʓ?<Xl�*� �2��[�bi�ȓoV�	i2$�6�)���F���U�ȓg�ཱt	�}��]:�������ȓ�B�j�'L�<�q)ѭ�/VL�ȓ ���[�F]2Y)�P*ݯ
p��ȓ/%ʸXw� =xۦ8���٫(���ȓQ> �x�oL,��,a�!V��X�ȓ8��5r���g
@���"�RQ<��.����k{�Llx�1*�̇ȓ}DD��G-)�,�A��	.6d��5�f�0'$��j�LA�*J*��l�<IP�­R\�[�B�
g.�33E�P�<�N֥h�ک�w$�F0A�%�g�<�s*Q����&N�:v6k�]m�<�g���)��T{#kK������j�<Tţ3���'��	>��K�<���>;89�ǩ�����L]]�<�w�@�#�r�+g�O��p!�^�<���0[�ztꐈF䠰���W�<��N�`�  �WB�/�6!C!�K�<�� ǨE_��飍H�Vrj!�� J�<�Cl&vS�����f��u����l�<iׂ�9AO���E��+����j�<�qGO=s�L(Р���Mq6g@P�<ad���0�"7a_P�K%	3b=!��M�aG
_J�H�MOvI!�$݃}�^�A��^�|1�$a- ;!�ԑ-��`���7mCJ�{'ȊC�!�ĖwKܝi�X�7��Zo�a�!�]����BNV�\ȳq�C:�!��D���w!�L��z�F�Wx!�D�]"mk$��n�R�EԗY[!��`��]�ϗ5/��,Y��S$,U!�$_t���(�`�_r� $�<!��s>bkЃ^
��Y��U	19!��J�akM����{��8�6�L�e�!�DP̘�㛛��@�!�"j�!�$T��2<s$^�5�4�QE�~�!�D�h��cN,0�^��ǠB9	q!�� b-s�� +�ԝ��!"�咑"O�	�'�K��0
g��/��9b%"O
��g�� �؄�!�*�~�J"O~��b��,�T9��ǂ�)�le�"O��Q�Q�U���2M!'��SS"O�;F+@!�nų�lǬy���"O��#1�C0�zy�"�^�<X�"O"���_i��U[��ڠJ�"OX�A��be�K�Cΐ���"O\53�� pѐ|2���#� ��"OF YT�_�'x���H��D/䄠7"O<�$Y�5^m+g�'7���t"O,����ޠ^�x�����"Od�p�oFd�[2.�����	��0<�G��*,�*p���5ip�m�Uh d�<Y I[9-�!�"�g���E��E�<i��7c��$���U�Zp�y�D�<�����RD��)4�����@�<!��@�&���	/�,{�ZE9���S�<�O�4j�8�yAG�zP:L���W�<��"�$� q�'I�#s�	)�m�S�<��(̍3F�c⫝���UKŃ�i�<a�	�8���ੀ�F�Rc��K�<Q�C��7+�p�CW�O~�dJ�AK�<!��-@��A%��5�,`R��r�<���%WU��{Ei��A�
�Pa�h�<�3,�5�)��!�te.IЖ�d�<����ȍ��I��+����%�Zg�<�"j�����2Pm��y�|!��l�<�gYȴ��!�^0^V� �w�[g�<Q!I��n"#���:�ʴpa�_`�<�2AËc��i�瘎BHP�J�b�<!R�Ϡ�a�E��,���MXc�<� /i��\�� �)C�`P�kN`�<ق�כ����)I�Jxεxv
�_�<q�GE�J؂(�rb�-~���c�^�<�T�;B��LȒb[�O����'�RY�<���l���r�(C�vT��R^�<y�n�]h�< ѣ̅5@h2��V�<5/r��,ZcO��)|,²o�K�<!ToJ8X�B�hm��;�A��	�J�<�b���v�B�ǔ5�j�җ�Vo�<��H�7���#�320����j�<���T�Z��U+scʲ=���h4�K^�<A	�=��P���,���c����y�����d�)�PE��3B:�y�N�Wئ)��E��VIt<��	��yB�ɝ.P05�w�!��j����yb�@�g�H8��ӈچ�PHH��yb �$%�6��,.��ر�]+�y��}A*��۫v�����y"�J5�� Hf�#ma44P#�8�yRoX#"�H,���I��1W���y��%����$MS<�T 3F��y�a#5�UrRh��4���!W+��yR J�G򕋤�E:��F��2�y�IΒ/z�%1��+IK�1C� ��b�ySSNO�SN��#GE�N���ȓJ���eܧ>���R����L�ȓ,L���-Zb��5��Lݴ7u�q�ȓ�^���Gm����W�`wJ ��Eܒ�#�\~C$p8� ؀ʒņȓ9�r)�B#E�2�x=P,��q&���mѶX��kā'J��bDmQ�F���S�? �R�#E�A	�g��"O� �&*ӷg���p��W�@�A"O�i��ʒ�&S"��4��-h� �"O������t�ZC�<��8�"O�y��H %��=qG��%,���y2� .p�ZL���e8��,��y҅�0N����ϼH���FǍ��y���f{��#@0/D0��R��y�j_���9 cې)k����)�y2�V#^(���1W;�qX�Bˑ�yr�ν	��i�%n܈+������yrK���`�WJU�I��A*�f��yB��#_��z�ᘿ>0A�)C5�y�hP��.!�)]>0WT '�"�y���c�$00 �w3^PxVf�:�yN/	HP��tIă;0B��ɮ�y�M��	>�E�s	 /�����E�y�a	�eCج��c�-�̈Ӱ���yb/;�ň�h�/'e0uQ�$��yB-^*�� ��*L�����{�B��,
H��M+>P^��G@ ��B�ɂ̞|�a'�=&�<���^�P�C�5���4'^49����@|K�C�Ɋ�*�Þ���p���^/�pC�QLe�ŉF����ȅ-�b��C�	�\�(�K��-�<%���Y�Aj�C�I�'ƚia#bX+V.J@��+^"�C��0:��`A��ټ �be�gN�'4�C�ɑ>@x��"T
�2�rҠ���'m��h��W�D��U�E@���'���R��WSl!��
�C�����'��������n��$h���6Z��x
�'H|c�A'�D��82�\Q�'`llؠ��1)��Ec��N YUȭj�'��Ql�!iQ�i�Cg��XŸ�+�'�,� �
&
��1����Hr�
�'g:,ڦ�QOfSEǚ)~���a
�'+�|hb����Xt$�|�ȵ��'��1�(���]b��9?$Y��'�r�3��H�r]��R��=���a�'�]��ꐡ�*
��<��	�'k�r`���<j4��A�2�I�'�H�k牎�v��j��	�:��)�'�.(��
^�@t8��E+@����'�B���'M8NS$�r���9�N��'��h	aɉ.X ǃ�30H�{�'zvԡ2+��BB.���E�^�xd(�'���E�rDZ ��іX�t�'ֱ+��Mp�4-�eR-I�@0
�'7����ͪN)J��&���t��	�'6���
_C ᨃ,M����'ۈ�y�n�-[��9�S�؄q`F���'{��գH�z���D�׿n
B���'10a�@���c�
��j�fȊ#�'�a����R��N^�X�L Y�'e"�c��ȧ� �����J���'��L�	��,�s�K4D�PC�'�=r���t�"��f��e�P�'�� *ai�7sz98���"�@�#�'�ʐ 6�G�L9���+K�v�P�'� ����A���pI+EY�� 	�'V��2AE�9��0��[�1}����'�|�s�%\�*��y�O�'RR���'�ܱ�EQ�:���1�˽SԠ���S�? ��!v�Z6l���I�BF�e�~���"O*a�uĆO�*<#R�^#!Y�U��"OX��B厼D۶U���HX����"OF1(6�Þ<<���ـ^��Y�"Ot1��΄,��4K �� n���!�"O���g� srl2�!�
�zw"Ov䲢*|٬|2����|h��Ҕ"Oj�C�)܁��1 �?_Q`1%"O�X�G�Y�"0�PS�(,�6"O�ms��ʓ�ބ3���j��͢�"OX�SƂߖY��N��.�Q�"O��J�E��4vD�8"�\&#����"O�d��G�2+��٣,�
�&5��"O
�r��?�)D,�9Q���Ж"O0q��M<��ɋVA����U"O��#�+=�\L�*!V�`E�`"OҼ�ׁ}�\#/A; P�D�u"O�#�BK�Z3m��CE��hU"O�P`�ɒ�F�xcΤS-��D"OhH��Y!g"��v��(~m؈y$"O���Vm�9� R�IZ4B�,�7"Oj�c�La�$����W,5dHa��"O>��英X��ɢ��� d؈�F"O�M[�*=�0��$ _����"O]SUl�����X�nݕFd�e�"O ��T�&� �&.-�H��"O��� �A�����ٺ��P"O�5�ǡY8$�@�C��>�b|��"O����fE���l 6 �Ji�w�<�蒸&!&h�c	4 i���$�q�<Q��Jx�=S��O�Lȓ�$w�<Q�nʽ�1A!��'R0Ru#�t�<	��E�F�p���:yK^Y��gg�<�a�9&_���tb�<.]@įOK�<��cT!\����UB[H~l����H�<�#�I�\c�r!eP�)\Y�<��ږÊ���a��5�������_�<��^zN�)�ʚW�"8��W�<)g'�<S��pg��+I�0`f�[�<�dҬ)��[�/S9U�&��v/]Y�<Y7a� /�J�A���4[�&q�OU�<�E�/Q�f��u%�(�@�	�\�<���)�!��h$�`�����Y�<�6E�r�:�ӣFt�&�H�lJM�<i�C(s��@��dQ?]L6A�&�H�<�!��	8�^0!֡>/Դ ��WB�<�N�-L�qSKX :�@����t�<1�S����LM�)!��1W�y�<a��^%m f�q�ߺ*�����'�x�(�d�@C$p��X(�'�xX3�U�H62��G~2� ��':4<�L�#}�DY#��p)|-X	�'�,e��	��80�w��6K�I�<	�cޘA���b�@�q]L��r�B�<��M�s%,d���yb��4�BI�<��CǑ�<��G�=Wl%��G�<�rΝ� E��c�	[�9�4T!uO@H�<�ů��X�Hb0�J�#ke	�DLj�<�IL:W���9D��Bn(�z�ƄO�<q��,����!#ִ:��8��S�<��C��N͎�9plM�C��\�!��J�<�1�'K����M^�)(�� � q�<��J�=����c�[H�J=
�u�<���A�V�N�S��H��QR�\�<� ���]z,��%�mD��9�"O�|2�&̈^.�x3�F����!	�"O(��F�4�m�� ��!�l�#�"OF��$�/! �Cm
.vv��X�"O��(SI�z�y��,JE\U��"O�R�É [����C1WȖ�"O0b�f�J`���bύ4z���P"O�%9� �9x�\piҷZ��@"O`�q����l��H�*�<B5"O.��r�΅$09A$�
{�dPH4"O~T�dA^��=�^y����"O������L$�$`ڢbF��"O|1��f�
�$���iŗol�@��O��=E��&_�|�: ��t�ՊBkԚ�y�É3촙jR-��TTPX�`��yb�#�|ݒ B�Qz��Cp�R��y�D�v|�jq������N��yB̉~�b�� �$8[���y"��=��pd��! �D�j���y��0,�ޅ(U� �i|b혐����=!�{"m�*vv�4j�n\�/�L���!M��y��va�a��ÇU4:���9�y�J�R�~a��SM
���k��y�R�n����mI�
Y�`o̬�yR�_�
#5��H��:����y�CADqPۀ#�?<MF�uA>�yRj�!*�=:0 ��J��
冁5�ybƉ�]u"����Ps.�Weэ�yr��2Z5��᳋�
I�D��pK�,�O��=�O}�`�5�r�d���Ѿ��Qp
�''�}8��'.DĤQ�ɂ\|��	�',tM[S'�8E�L�j`-7W�	�'z֐C��W��f������0sb\ �'�!�p�@2\l��w���q؞T�	�':N�˥  �:��IQ �Ãgw��x�''vM��͉O1� ����=e@���'��ER�$Y-��M��4G�H��
�'�����/2TQ�6(��-���X���*O��C�!A�����Q�/;6�	�"Oޱ��d�Z݋g�څ{ �лiء��HIhD@�0�)A�V� w
��ȓ,P�!�2iܛM�	�v�	r|��aX2���L&(u0A��)Ԍ���s�����»�̃�aϊD��Ȇȓ*�.���E�1M.P���?(�f=��|�򁺥,�$+��0d�ǲ.`~Ї�h���A��/�~���F6$Mbu��k���FJ �|Fa��@�1��%��Fy2���/7����ޖ04rA9")X:/X!�$�6>G&�:���64����#ʛ9+d!�DK C�����7ZX����9[!�D°%y��a�GD�?$�!P	� L!�A�;��*�	D�^mB��Q�/h!��)4�y��D��I�X颇E�c!�dJ����o��^� $��^P!�$��,���C���=R�nG����!�dV�G�Vm�1���/��ISDT�#%f�E{���'��aY�n<���,G�h��0��'�� �C��nTc��M�� �'�T�؂kT��ڷ��n�2C�	"<��Pd'�z��C	M�m�B�	�"�l�Y��G� �J ���P�	B��P�b ����{��� �>���-D��{�C8!����o��yr4i�1D�� XD10GJ�I�z���lWʩ��"O��[+�3)9̩˥m
5<�0S"O���tK?yp�`i���e#$Mт�'��'ڤ�c��"�h)����d���'x�j�����z���۽_VF�Q�'��A�f�?m�0��jT],H�
�'�6�3M&��A��+НS���'1�\�@EÛ2�x�J��~]8�'����G��:\zB� v�$y��d�'h�(�N A���H�,�/=���
��~�KY	.�P���*n�(	����y�E{XVt�wˏgܬpH�,�y�'�\�rM�'���ŏǶ��'�Q:H��m�P5"d�� 0��'�'��)�<��a�"�Zͣ��X�"��o�u�<QPhWf2��H3��M#h1+��H�<)�cO�r�$0хi��Ȳ!��E�<��(�Rx�����-t ��aKk�<�f����[&�̓*�	��BMf�<�

�:�RB��"�H�����i�<�a�TX_���"��<D��Thp�q�<q�`\�,.r�"�NW�gdD����j�<�A 1I��H����g�4 �Jj�<��O�7yڭ���B�}{�]}�'�Q?ɫG%G�`.��@��H���[�j9D�3�j^��p"H�.� �.<D�x����|#�T���*d"�x��7D��j��rI��b���W�t��7D���2'K��8q�a/C�pk�k6D�ԋҏ�48Z�8VI�v��: �>D��q���s�@9U� \PD˒�;D�H[�� 3/��S�*��$(<A��e;D�� ����L�����o��̘6�4D���%��%�^)c�jW�s���3D��Kҥ�a�z��*� ��1ʓ�hO�,Z�,4����2�~����gC�	a�������:�6���ϓ:PB�	Q��S �� C�ɱe�&7�2B�I�qİ�`��Ñ"�8�j��
dT\C�	�V�V��V�>p�pPk��7r�rC�I�~X¡`�c˧,+(�l��PKB��*	u^T���ñ��QB"G84B䉕)�8�B�a\�}�
�f-�A��C䉻��;]�D�C��,$�f4�$"Odi*�£
w���V�L?�*��A"O��Ѵ��X\��K�I� ØEr�"O�}kb ��*��x8�G�&�z|�2"O�4�G�S�>Wrms�l�r�lir7"O����C?=�lQUm�:ce�Au"O�`T�l-�6��7S��;�"O ���a]+q�ƴKö~��EL�`�<QD �vv�-c�/�a����rcY�<��#H�?���
�nBi[�c�W�<�� �9 d��r��m�D��"�T�<�wAQ�?�F���'�=��A�r��Q�<Qɖ,s@��J(��F��K�<a��6�^�`gP�8��T�M�<I�iJ-	���+�.�	7˞��J�<Y���(z�,���T�M��B��F�<aW�B�2tZ(��m��@%J�x�<iF��N�
��l߅ZFΨ2��\�<�FZ%(�\%9��܁)��h�k�m�<	UFW�L�d� V��X\2Ӫ)T��W�J:TX���˂7!$%xd�/D�� ��ĥ0.�P�� �0z��d�D"O� ��M�[�
0��O�I��i�"O^�����\*���9���+�"O6xB6��H�4��a�I&i��6"O0�c%�9 ��!2�H��t�$u�R"O�@�m�\/�Pʇ��x��$2"O��P�ܕ$�|����<K�lh�"Of!7�Q)VUfhAAiD�)iv"O�  Ð
6(���7EE3!�X��"Ony���).�) ���6�Х�"O2Q/	�T���Z��Pς��yBhB��$scJS"aC
��y" �����1@LM3S]4Ջ�Z��y"͜,�R�FkG/O�ԩ�G�yBـX^�h��CG��H��*�y�� 
���Q�
:@�y�Ǻ�yBg�U���!�D�'��)2	�y����`��%	Q�v��֮U!�yB��3tv8�#�$��$�p��ၩ�yr
*,�\�C d�?%���,+�y�NQ!S~x�ȡ���N��+���yR!�0>����F<t�Uqs�J��yb �(`8��S8  4qYC�ڮ�y���U���8�P)	S���y��]�S.�؛�땉z)�Ҭ��y�%��@� �ы	�u�Z\w��"�y��%�Te�D�C*8�i ���y"K�5f�t�0
I�~-2�*�� �y��[;
����²?ܶ�/ݬ�y�Ü.���c�#�!0?F�*��(�y�kϤ8�aɅ���7���;Չ��ybOE���st���44��r�
�1�y�'�
��e��)Y�m<-��-ѽ�y��6lPD��@Ѫe���;fj9�y2Jf��A��׿O>����F��y�/
Z����$�=^�Hmkʱ�y(ϴ,�v���M]^X�;$����y�!"Z�zD� >,x�r���y�9��8R�ɬ0��\�4�\)�yR��T8��c����n��E����'lZ�2��TN�,��ւA��U�'%�����PR,�Q/6e`8��'g�tK�"�+(�8���W�Fi�	�'���q���7[��@���SZ���''�(�E��e¨eiu��;�)��'`�엂#��	"e�+s$��'�Tq�A�d]������*�֤R�'A�TQ�g��G_�ź���/!u��x�'�pM0vc�7 A��u�Y(�TP�'����`# ^�/�6�\�i�'Q��A=S� ���+Z���'��!˃M����*�1XPM�	�'���:FT`H�S��.m����'�!j�b�
�H��<%�-q�' Z�b�i�(������-f�N���'���͕hl�(�J*\���0�'Y�xf��|���e��a�:Ղ�'D�	0p T�g���H�\�d��'H���E&[7A-f��g�|�R��'s���VBK*(��)W��$&�LQ�'���xEo�.������*:8*�'�|l���>{�8��J��ޡa�'��-h���@�A��B�4���
�'H�!�t情w�;R�����
��� .t��C٩6t�<�g�	�F���"Od��c�h��k��2}�\r�"O\�3��n|��'���?�da0"O:X��z)�ʠ��vn"�9E"O$"�P�F��`�'̗S�;p"O!���*����'�		>d��"O<���aM?
 ��'ݲy�� 9�"O|D[���҅����[L�%@g"O@�9�/�4�ҙ�o�6$��sv"O����߯�z��t$
�iʽ��"O1��f��:e�(1����C�Ĉ�w"Oꄈ��Cp�:ȃaO�δ2"O�t�@�B|��5��0�pQ "O��8���0{/b	YS ~��ԓ�"O<9cwF2���I#�x��"Oԕ�.�����R� B��`�"O�L�fǈ0j�|@i &J+4�!�"O��@)6����jGj! 82"O�A�eK�`s� �+i @1R"O�i�n��v�1E蔮@8"1+"O���H�:~��2ҧ��m2f�$"O� �G�:�y��'�W0�I��"O�=J�P�,��@�3�H0��"Ot���Eg�=���((B�P�"Ob�p���.H|jD0c��l6�R"O�0ȵ��
a��@��ҥ��MjP"O�H˷K�t$��"���FRJ�<馎���J��̕(��}����<��cW����#�H&s�jU��]{�<�0�ה+�N(؃�Ӌ{(����z�<����:|S�R���d�RW��o�<�F�ǢZ|�\
3��)?��B�Ok�<a��V4]�
���&c���D��k�<Q�`��K�4�ϒ���]�BL�n�<V��B�� $Q� �b�2��j�<��J�/B�<�A&߁�:���bW\�<9�����R'���|�,��cXV�<�FCK4f)�K��Х!��9�ĎL�<1�ϝ)0a���dC{�(�Y��s�<�Ղ�6}4yCb䄅`�h���!�l�<��oIB�̐�1JU�I��\�d�g�<�t�ԙnQ=P�#�Ԓe)TC�`�<�a�k>b���(�����MG�<��@ԏ+��[3�Z �ck�~�<�&B�)"�Ľz��S���̸��H|�<A�C�(*n��@1�
sN1��w�<�'	��l����K�*Z��B��H�<yt�:�Z�o
 1����p�<�b-��&E�� �M���8@��l�<�!.A%B�x�S��P��ҍj�<	�0���J��I7Q�4���n�<�BnK�I�$q��=h��)`�,i�<a6�^:>yaGgH�$�:YPG�^�<A6��-iجk���Tj��#�Ma�<A�R�;7��	��DbEl@a�)Rv�<a���d�[m����m���Fo�<����e�0��ǔ#5l	���h�<Q�'�a��$#��'o�4���Ae�<I�k� �(⅂)j8�t�`�<!�K��7=Z}Qf�^(�l�0��e�<�c���
�­�sC'���Z���F�<1�@R�6���XulN,�L(B��j�<1�k���R�	w��<�0�7f2D�@���ņ	* d�mO:�B!#2D�� .�3�ʆ?5�b��g҉̍k�"O,������z�l��e��/�(qp�"O������{�����N38�b"O��%mMN�nY�kقw$�T[C"O�ْ1�P�\��rSIL�5-̱�"O�$h�k�o!ܱ)��� O r"OE�T���s����"�*x"���"O�,S3�6���(7��a���"O����M!�z,2���8D��A"O4� ��.0�@��3���_
dѦ"O��Z?WE�T��I'N
4�$"O ���� R���b&-�Q�0HȄ"O���v�]��v`�2l�'���s"O��lD�z1T�7+�-0��=�P"O�Ra�0{�*LbCOX��"O�l��o�_j��%d��H�rP"O�#d �59?��1"�D�-^�i�"O2��P���T��<���߂:8�"O���Wq�N 4�2 �TkB"Op����M44[�-�FĄ���y!"O�
���Zܸf�DzR��"O�-�1�M"&���栗69�z��X�<9#���z݀�wŞ�PL���k�<Q`>'�Xt�VHT��n%�6�f�<�$�/^���s�LŚTC�T�f�|�<9S
B�f�}�bn���5k�)E`�<��o]��Bm�V�W�),*Cb�f�<9@ퟄM��ST���%�U,�F�<�#��6||�� �$V�D�ٵ��B�<!Q$��U����BO7ྍ	�#�A�<9&��6v�P���Ŏ3TH���o�v�<�n�{�R��h�� V Aaq��q�<a�m +�����-�((l�<��oY����W 
15�l|�'fq�<�@A�-Wd� ڑ�)=	�qk �o�<�[�70�a`�(4�Z���F�u�<�e�%|�!7/V�0�.9fC�|�<�s�92����L�=4�R� ��p�<qIC��&< $E72�~e8�ENl�<�S
���<eC`��	p��5�T�<Q���5�D��fi���Xh�<�!��L��jצ� ]7����I�<T㘌+2��WG#s��xp҃�B�<�T-186L�f�,�E�#JV~�<�T��� ��Q��� �X�a�Ta�<y��kDN0�`�יp�*�z�fYh�<�Uk�sL>�"���8y2��t�Gz�<)�JП	~���P� �Bl2�JeE��<	ʗ�Y֭K�FX�b�D�@�c�<��E�O<����fQ*�� ʆM�a�<y�F0p��I��o�9k��q��_�<�1����%IF ͢�l��!�X[�<y�
K�V��k��z|��v�M�<����V�����Kd����!m��<��
�8R|ژ��K}7�)F�Q|�<�	�$˲�K%a��uu0a�j�c�<A�nQ��\@"6a�C�H0AmDX�<Y�m�/<��"MR��楈F�HR�<��nI�N.�v��S�
YXjy�<1SL�M�ldq��R��ne@�\u�<	P�H�Q��f��c�,`�"`�t�<A�ۻ���#�(:=0�O�t�<97��=u��X�u�Ϟ!"�eA��o�<��#U&�"�� ���$�s��j�<� .9�P���S�J�ZQ�
"V��d"OP�џcb�D�eɜ�^d�(t"O��A&�Ӎ*�j�vL '0D9�"O��CA٤r���	梑'3�qr�"O(�r��K#��`�����`s"O�XE�C
4����Хs1�H(�"O��e�ʕg��0��ss��X�"O��REmQk�5��J��dRI[ "OX�b瑂 �ؕ3��� \�ܙ�"OvM��d��W��H�ʷ!Xx�G"O�4��B�&�A#7$V�09�t[�"O���aNwS��{�#��q/�]C"O�ѱNE�y&�I��Ȗ4�8��"O��� &�P��Q�C�o(O!�A�M��"d�4,�A�s��#Z�!�d4`�v�1�)U�9JX���C=+�!�䁰<{��C�#������Z��!��_F��� ^��Ժc2�!��ςd��T �&(�T���׋Dm!��&C�Zd	�FU5�i�� �!�ēf�5P"-\
%+,P�ʌ�M�!�D�7刭rQɔ�K5�uj�2m|!�dЛ<�0h+�-��a*����@i!���P��YC)�* �D�@�5M!�$��[�Xlr�'�=}6/�$mA!��� 8�&����G�\�;�N��s�!�0?�&��-�q>� �-2j�!�D��g�h��@����<A�}�!��;yL=� "^1y��h�2d!�$K�+����CͶșReU3M!�$�Y����F�j�p$J#ҢG�!��E�Q��2q�ݨl�Xs �	�w�!�H� Q!ǭA�*�R�k@@�<z!�ā�M<����k�eж�X�mB�0�!�d�w��H!J	Q�yR!�@;6�!��T� K�m� ~����+I�!��J�`�����=Ou8=j�d��\]!�@�C�(ä/�`�U:��*pR!�$�d��0��*W�CW U�W�$c>!��#�`�n�99*��;�.E�+!�� p�X��+�d"�� Kx�!�dĊ@8�w�Q)F����?�!�F&N�B� l�N��8���[�y�!��R�r��XXr%�*3���C"4�!��)_E�Y92�	�Z����͑
�!�Ą7�0����x��i�i��0f"O�%#phW�r������\:UW���Q"O4u��&�ZB���U�ь	S�{�"O�x��cƆ8G�8�3F�>V3�)b"O�i��%�Fx0��K,0��B"O�ؠ��l	��&��z���"O���919�U`��\�b��a�p"OXt#ի��u�[�eE�S�T��5"O&Uz��U�`T��d4V��Px"O$l�f�̔a�V�Æßn��IYG"O�m#2�3�=�w�� 9���p!"O����H�mu,��r�cs�ia"O:��	�%)�,��#E��ggL*�"O��Xc�[/4n�FÙAg�I"�"O#�IÂ8��z6�ܓM]ȝ�w"O�E��-��AMԤѣ������"O�i����n�\�3��.t��!"O�i[�@��f�����I*�n��g"O�M�6 �%Π,r#oմa�vI*S"O� �D��L�#a�:��4m�W@z���"O��ʢY�Sly�U.�&7&���"O&=��?[fl�r�
,m� ��`"O$�Ps��
s>K�i7&����"O<����q6Ø�lp��"O��y��
Pq����>�\�!4"O�<J��;��8�4,��z��b�"OD�!�!�r�diW�J�E�0$��"OZ�2��3@�`� �9-Ǽ	YR"O��R��Cb��8$@ ��a@5"O�h�AN��-w($so�0r�]!U"O>h:��u[��2PN�.پ@��"O>Mr4�P�yi�m2u�H�Xw"O��@�� A$b5fK�Ef ���*O�0Q��c�l	#bF2�3�'�V�F� g�D��1-��;**���'}�|[��Ź���`��j��Q��'ɀ���(D�L�mh�e�d��
�'���pnP+7�P�5̓h��|��'�PiF���|z�,����/s�$\Z�'f��4���Q캕��db	��'�~\kd.W4/lB٢�n����x�'�6�@A�S�u~�,�J_����Y�'�}�GGÌw� a�b��zHx��'}.ԡ�ţT��IS�X�6��*�'���Al�=0`P��Ӭ6��	[
�'�h@��G�N |�k�ݐ*�y��'(�-��ɀ"���kwn��Vfm��'��@Äɣ{Q�d��A�\��J�'kni;�/�lbHI#���J�Е�ʓlL��ؕ��'x�4���ə;
f�ȓ2#��g�L��d��<R
)��n��:�	�,v}J��e;���ȓ&�)�'ڲ<f�1�d��.BY��tJtأ�O�	�2�˴��D�ȓz�H"&��/G�Y��K�?4���6�,�����fn��I��X�cU����/�Z8��*�
K,���ó�`,�ȓ8�ay��/�f�Q6+<Є��^.��1lE���uq�E+�<܅�I� -1�ڞ�$��B/��N�������@��ɓ����3?¦̈́ȓtW�l��ۭC��hAN�<Շ����Pn�.�*�X2*��Q�hl�ȓ2L���v/H�<�E���˥<���U�"����.N&�M��McK~Іȓ�D� J�$�x�6��D���`ʌB@H?�$%*��e�`!�ȓ?�� �O>A�|�c�I:c7P(��hQ��Q�'\��6E�歁�sz ��r�`s��8�);q5o
&]��m�X���(n\^�"��0|�`D�ȓ,�$��p������K*l��y��?���f��g�,̓��A_����ȓ&��
�D����d(�x;F��S����&
;��6� �o�VB剘2c����5vj�,8���YutB�3K�}��"����(N�%�xB�-K]�D�ǌ�%��hD��!HqRB䉏'��̣��"�b�yAj��*�B�	�7\J��3�	N���5ن`�C�	$s Z��F�+$�`��$3vB�*L"�ȩB�8GN���W W;KB�I I��y0�jтHG�1��U�]U�C�)� ��i�j��*%vAi�p�9�"O�<aS	Q5r0t���)0^�r�"OZ��d�N]3���EFF�+r��r�"O&5z�Iޑ=<J�i�e�7J
-h�"OL��j�5�e�j�'
F��"O����4����k��T�x��"O�t�d��i1`q�h�A0"OZ�9t�?]�������R"OܤH���84�����28p���&"O`�#L8:[�D�1� ���x�"Op�Jc�2[(�9d&ˢ|��]��"O�KC�C�iI�bE�@�U�xa	t"O\��B�/[?��@׫�s���b"Ol�Hs��}��a��F�"O�9�^#1��q+2��/k�
"O��x�dݣi���s
0 ��0S"O"��A ؃p��I6�����8"O}����<cF��<��P@�"O(Z��³ᬅ�P��uU\i�"Ox0��OD=U1J���,K#8�pyR"O�Т����C1*�{T��	5��"O�-�J�"F��i�E��%O��T"OP(��gƐI�ac�	\�xe~UR"O�="#�}�~��iDl���A"O�-k�L�_��]���wX��"OL��t's�4� w�]�lT�i"O^�b�/����qQ�|B\EjW"OmQ�%��KDl���,F�,&H1e"O2E�O��F����s�Μ*E09��"O�
���Ґ�ג8��l�����`�!��3�t�I��3.��hQ��1!� �x�3�Z�(��AIp��1	?!�D_%t��ǄW �����ՎO[!�$2o�=�c/֙-�-����&R!�dL�Z�(�*�"D*bdj���t�!�d�+v��3��\8U�1Gѫ.�!�$��>U0��W+�U$J�8!�D\z�^<1D��6K*��3�L�q(!򄈁t��A�����r\y�PKX�]3!�M�&�X�1�,��9 ��qR�D.;&!�:��U( ^���a&[6!!�D�=E�r��@DE�,�
CO�z!�ÓD���S�\�zz訸�cͧ{!�ҍE@�M��$Q�Q`���W��d!�d��d8�o׸CCd�B����C�!���f���q4'�YKؤ�B	�'J!���w��e�'r4h���GA��!���4�@�!U?L�b�-�2,�!�$H�*d��ن@:��m�;�!����(��/@K�L�}�!�W��R8�` ��&�\JEaQ��!�DL�[�:�9"�Ţ~
,�+�Ꮍq�!�D�E��G�]	f�ta8�m�'$�!�d�%\��Qr̃�! D���fa!򤏐NDL=���\�.�4
'�M�T0!��܆μ�#2!6(�h:S+MT!�D�l��1�w@N�"R���_�!�d��[i��r��h���+�(�!��X6n�J � ��B�B��G�|�!�f�k؁=8T�[`O�k"t�V"O�!rg�U6QH8��`[�|�&	"Ov|0�ÄN+�8`5
�M�Qx�"O��uϜ'~�R�S�o�>-B�"O��c�XNPĬPr�ܔ
u��s�"O� �<J�LL:;*� Ĝ_F82v"O�� �,��9A*!q�� >�rY�""O2p0�k��g��!Bn׏Y+�"O�P�4dQ��JMBfMA�%�M�@"OH]+��˚rV�9�1��t��S2"OT-�d�ű[���[rO���D���"O��)��!p�Y�D_ ��x��"O�����>0�)��|z
չ�"Od�2/	a�t����8���9�"O����Z�q�QZu�E=&�z4[$"O��#�S���r�o�#"O���u�P�2�5%G�lb���'"O<l�1^t|��H4/��"s>�
"O�(ө�=�d�j�MV5G�x�"ON��d�r���ҐC��o`@���"O�T����)D`D�s��sy�|� "O���U���8'����A"|Q�g"O�� �@�#�Q¢*O%X@�"ON`R��2Fy��#& V�$т|8�"O \�#�^�!�|9U�]8 ��x�"O�a�rO@"����O�v��! �"OֽC�Ͼ7;L���+u]i%"O*)hեF�JJJ� -��A�,��ybE�o��]���W4&�j�˓�=�y�m҃Ekp�ZB��	�y+@d��y���9���;sO��P�
��y��Ŵ����ƈ~�� �F��yBH@�|X�P2N�>,��ŋ�Nj�<YR�P���`!��C?T|K���A�<����,j	��q�	��&P��A�<�b��7R���oݑ���8��PW�<�E��<��53�e�NK��Y	R�<��AU�C�"�����z��;d2D�P���ʕ_�ٸ��^�YP��=D���NQ;b-~��%´t�h����=D�4Ȧ Ÿ�6���Fݾ]bm��L:D�Ԙ%��)#��c��w&�0�*O攙Š�d�<� '�޹V��� "O�9�fA�;������ J�b�"O��zbF	�Ht\dC��/J��QX"O�0p%GA���s��PE޹H��'�Oz�Ė�a�q+L	9�P�S"Op��@�o�VJ?`���Hb"O����$,P�U�A�΁;B6D�Q"O�p��!�plpĈVD�$~V
\�B"O�%y,_	�ƅ�6dD+{78���"O�Q$M��9�9�r���8!:�R"O�L��Q�^A*��g�üt�%hc"O�I#��9 ��Ȳ�23a���D"O����H
}WL��3�C{ᚘ�"OT(OQ����3�2q{�p��"O��q2K�	CwR��6�әW�8`A"O��3Q�7i����$,Ҕ/k\�P"O��	SM�/@����̏#%��"O0⎟y�,0���Z6�N��1"O�L���N��LX�L��9�]�""O�TQ!P�=>\���߻�6T�"O�!V �XȘ��J֯Q��9I�"Ov���a�> �X�B�1��\��"O��A7�:��&��7�t�yg"OK����wE��y��2�ဧ�y�CD�O1^�ۅ��up�T�eL6�y��ϱ��!4f��v���G���yb�Ԏ ��dp�	���Ȧ%C��y
� �(:C�Q�Sp�C4���M��dBG"O�)t�K���C�.ȨE��K�"OH���h� ;��)��,Ӊ����"O��"*pﮙ��,�"1�:ݐ�"O6A ��'	�4K�HU�nq��"O�+Cƕ�pP�!6eԑOz|���"O���D��C�&��d�4���s"O��9V?������7�a "OtȈw��e���h\*<p�P�"O���U���JsBX6'�Q`5"O�]bB��
EڮH�B�,g�`��"O��r&��&��I�E>јR"O P���އ �Z��@ �/F��Yۑ"OH�y���w�,0�6�Սe���A"O����сǺ�WJ�*|��mI"O|`�pg�:A�Zt+�#EU��I �"O��,�1���#�C��.uc"O�`kr�92089;e�[��R�"O�͹���j�B��#��Wإ�"Ob�A!gC! nH��*g��"O�@���:����I<^�ȃ"O4�Q�@�
���	pa��b�j�"O�5��\n�
�g/M3;1F�P�"O��GË�]�Tч'Q�M	,��"O<Lk�L/^��]����9N5S�"O����L�.��#@���4"O�+�#è�veѢ� �Y�	��"Ob��!FD�z~���E�KN5R�"Or���f�ol�iSG��9��#�"O�3�W�V�V�)�$̻}��B "O�I�Փa����	�MO��"V"O� ����F"��'��Ya��"O5�k��A�!&�_�&h�0"O��� �J.2H�KSd�1���!"O�����#ER�%�W�P3��]Q"OE��^g��L¢*{xz�rP"O2H�Q'�.��@!��&"��9"O|)+@�c�li���ղ�X�"O�H�7��<6��-
�$^�)�"O���b%_#u<Rl�c��Y$�U�e"O��(����u<6�Q�a�H4ZQb6"O����K	u~� U��(:���f"OS�jBjc���7�E�I�>�"�"O�$3Cj�P�D�PN4F(��)u"O����,�^#�%��,Z�>��1"O�9�rg@�YG@s`�ڶ��"O��pFQ3R1&(��e�%���5"O���Sh�Y*N8�$>B�bu�"O�U���!�֙�tm 'Q�rp�"O��HG��>f�r��)P�0���"O,� �m� jWgC)�J��"O��H,G�p0c�U{���"O|�aA��֑
�����a	1"O��$h�.$�\��M�,�.�ٱ"O�iۦ@�j�s
֌-�Y-X!�T�jx��ž)�:�Y�o�87!�D�<	rh����3A����N#{!�G�j�RH�!I�7Q�pc3N�7@!�D�K�n�HGDC*h�P��_�!�d[�1� �c�?tx�l�7fb!��.�*��A�
h�p	�@�);!�֢r�q��-OVb���N�{!��^�	<�8���P:V4`�*!��
��� B񭘛u�C%m��,W!�� v�i�$�`]f��E�ʱ�VŃ@"O��	�C��M�������p�xI@ "Oa	2��9n0D��%�ɾ?��"Of�`�?I�̌�@]��
%�""OH����x/z������)B$"O�h�n� >]�Ȑ� �f��"O�����v��T��G�*��1"O^=��\-���'D�\o�*"OL�#' ����K�l��^��i��"Ob��`k��L�2L���RѼ��"O�)k&�ɾ�\D0�/M,��t�"O�����B�޲����h��S�"OV
(^}��c��Q�u�􌋧"OT���fY-oO�hRfӮ+���"OP�����M�-���X�p�#�"Orar����DLV���:��Zs"O�MxuEY�m�ȴz-�!��Y�"O��Ӣ��mJġF+�����[#"O�hI���Qx4-�`�:��h�$"OZa�֡D q�vβ��i["OD��fQ�j۞]��L��n�Δ�"O`���Lń>X �RFE��V�4P�"O(=J�C�gx x �ƳD�
Ta�"O�<��m�3gf��a+��2,���"O`л����r�R�! �;8Iڂ"O���pٝq�x/߈DKZ�:r"O$ �#G���-	�m��غE��"O0�(��m�����X�'�<P"O>�Zp��8A���l\SjnH�6"O*��b�D��r�kا:��d��"O@��͒'mp`iZum�0E�:%��"O�1a-�"GVt�-��b���h�"O�b��=]z���nC'{�JQ�"O�ep��̢k�0��J�%�"O�|1s��q!j���m�*!���"O�� �g�G��`�.K3Hz`\j�"O�t�`�_�Ne��Ҁe`$!1"O^�A5B� _���%ػ0m(`"O���`Ɨ�p/��YC�Ua�t�"O��K$�$[��1�l�UF��p"O.p�=#����ɽKBh��W"O��{�ã%�Y ��]	nYh���"Om$�ͷjѼ$��) |U,�7"O���H5�"���jF�U�"OF�8'œ26�6؊Հ�	z>�%�S"O�A;�A����/EN*p�)C"O�]�(:��Y0o�r�
�x�"O �4���Z^�u�A�3O��uX�"O
(RځY�q���6,K�"O��BרT� ಃ��6b�
�"O���'�I�V����$�Z�Vl�""O���"뒲BAR����� �2��"OdT����m��9���k�轡#"O���oϘ"� �+ ,��S���h�"O��sR�ӊO��xD@��+����t"Ot��d���x�ɂ7���Kc�(�"O�� ���a'�ѸTހ8G"O"�WH�� Hi��|���b"O����Y%M z�1�&��nߠ�I�"O2�[�	-ZL�i� +�F���"O� )W�(�Hy��6�M��"O|�PD���f�wʋ��Q"OAP�E<PDIʳɡ�(ڀ"Otѻѯ���`[r��mH�91"O� �(r��Y�2��CB��4�b#"O&�!��A$iu>��4�J%-�P��2"O�Q��\�HG��{�<�3�"O앲��	�>��{tʖ�zMX���"O?�v�C���$\�,\[��L9i�!��X���A3�7�J%���,l!�$ �o��	���ю��j�A��	m!�;Vz�٠m��MҾ�Q� �*i!��8D'*E�^%/�V�q䊟�gm!�]�N�!FΗi�P�)Q7vi!�DO%k���A�E�TT�1
��t`!�d��D�2��&H��]�.��q�U6Z!���47x�L���:�0��K"c�!��AG&M�q��6jӂE�e$Δ@�!�	[xf �S�DǄua��x�!�$ʹ^S���գ�D�V����D�!�]�uBGm,?���� �0cF!�DQ��QsAE��A�>DK@@�&8!�X�XLP�cL0B�R屰�%V�!�dI*����7O �[��(���O�!���/bz�[�K$�h�����.�!�����b�T8=�x٣��){�!��ߩ�|��'�O���G�ēlj!�Ĝ�P�x!��"ζj����
=g!��
S������\��x�d��2�!�$іˈxz�"C7,��+���N�!�d�Y�7�8�i@Ԣڜ7�!�D�&���І�L�ށ��⎫/�!��41�X�ٱ��lT�܃0��4K�!�P
D��T-�?LXYhA��'�!�ݼ(���ƀ�"4�4�ti�q�!�8$�z!����(;�G�*�!򄂈:�Ba��F�$�k3ǈ�B�!�ċ�$�"M�ׂ�5_�r]���T3	�!���}h�h!�e��*��Q�dB�<�!���#DЕZ.���a���_�!��D;F��Y��c�?l������ `�!�d�.�Qrף��&��s2��-*!��q�BS�@x܉`.��Lj!��A�&��#�G�Zs����GP�~Q!�D�w�`�AaH��D^$�C�m
,4�I`����52�
/>w���'���q��"Oyr���'U-4��B�X�("Oz�b�!�3yhĹ���
���§"O��P@�[�>��c�6x��a��"O���C�ٍR�
h��;G�4u�"OB�1�� 3��`A��Y�A�Q"O�ĺ�W����V��Q�Di�"O����	í|o�����5!.t �"On@ۣnɄԄ�A_�E�y�"O4�`С�
-<B�j��M�V#""O�e�"Y�(4��A#1�&I�@"O��hʘ�N��qE�Q \�$�
1"O����Սq��=�p�Քo!�i�`"O��@R狿~���#��U�hIP"O�,RPZ`(��A8J��Y�b"OY�DCX�c�l��᠜�U��Ap"OB}�7c�FNb���^�5w��"O�M:�̃ ' <�/��a�Ѻ�"O�Ԫ��D,��V��9Q�<|9"O���@I8J"[+�^���"Onm𡨍�t�����i��fEd�I`"O*�ֈ�1T0xG�d�R"O�	@���	n��0Q�y�"O� x�J��'.��{�j�i1(�)�"O�p��#�Fz�R$��:��9p�"OYQ�+�-u_V�QE�G�@���"O�+��%'������P�Gjp%+&"O12f��m���4΅�6[�L��"O��h�]x���@df@�y;�Mڵ"O�+t
�
rS�hUf���@�"O�ر4��67B$B%�^�}�"O�Ɂ���.���#�;�Lp("O�!iw��=w��󒢋7d:��&"O,0��fވK��}8E@K^	�"O����Ľ6b�����bT.�
�"O�=��c2����;J�!%"O�I�`kو�
�Q��U��)��"Of��(���Ҵ�!F�G��d{�"O��XT��9v�����ʡo���"O^\�5�9�~�[�
�9��<��"O�]�� ��`�1�f����"O��%�K��pQg��xB:��"O�hQ�aJ9}�8��e�C�\�0�qb"O�x�ȋ��E5��HG��x "O� :'(�m���4&T8=0��X�"O�d����,y4�hC3%#�I��"O�}!��6;|1�-��6!¬0U"OD*�D�?��t葍F5���X�"O�	b'ʍ�m^�[@������"O���ъߞz���!������:�"Oh��v�����H����0Y��"O�kў �`� @�&Y�z��1"O�:PT"�����l�B@ g"O��3�_�@��06.����0�s"OTP׈�X�4Tybꍔ|�\��"O� �Ѧ@7%��f�	H�
0:5"O�a�F�H5��Z���s�hF"O�;��3"��ۃ(�)��"O��Y�#�_��P2Fh�j�� �"O�� &�P�H�\@�(�
Jl���"O�邕l�>7�`tc2�9i5�(f"O�q�D�ʱ"�H{\ �"O�\*%��%���u���/�Ds�"O �:w��&~p੒���^����"O�)Ȁ������I�'�>���"Or��Ni-��Ӭ�W��+"O��H�n�;4���נ!�&��"O�88ѦZ.]�^�b��Q�O� ��"O�캑��a@�T�2#ѳ	��(�1"O��4��se��쏉&ӌ��"O0U&�_$^*��1K	C���"O�\C$�Ǆ5���2�^8D�JH��"O��I��&y��h֕�)*�"O��� f=I�N�5J`v�9"O�D�dR	ِ�XbM�,VdP�rv"O��)�Q�ؙ�ׁI�1�Z4["O��j�
���!���/:��K�"O�1R�x�ƠKԯҫn����"O�� L"hGT���,C2}����"O�C)Bq�L�G��n`4�*�"O�GZ +�N墷�U!A�hp"O(�!�jP�rP�A��K�j%����"OZY�j«_ўa�	1���"O$�v%ј���QpkK�F���ʵ"O�<Xg�׃=bu��,�V�
�"O��a���%DgBqC� ��*"OnqQc �_���e�P�k���"O� �@q��ӆ���2J�&JB�Mx""O����lŮR̼�A�4Y9��е"O�X�@�� IB�� ō�?2II&"O&x��.D�t�\��F��|�$�	A"O���&իEJ�*%C]�w�HӢ"O�lY��ƖS�2s#T�P�H0 "Opxy�I-!dh3�,S�k�L�1�"OM�b��*�L��䗈)�mI4"O��dT/)<5З�W	{ܨyx "O��4�|s�I0�,����W"O��JҠC����ŁB�pi�"O����V?9�D�c�P�T+L��3"O�!�Q���׃%T)����"O��yp�ї/*�Kb�):���3"OpQ��b�2*�� աQ#�^���"O��K4��r�,�P� ��$ ���"O<���+8	\ iB�M�w�^�"O�� ʐ�'����ͻT+DH�"O�@8�l�_�f5�$E�~m,D�"O���Ό�nό� e��!3�qð"Oj��Q�M�-�J��Ed�"%E �A�"Oԙ�P �Vj1;�m�#><�C�"OX���0��\�3�^7��X�"O��s+�2&Ϟ�:��=6Є"e"O@鲡H�P�$p[$
�	���Җ"Opr��ґ0��$A@gRa��%�"O��reȓbVv�����8-n����"O�%���x`����*$q~��"On�y��$�� X����`}����"O��8chX�(��oǮ6N:�ɠ"O���E��h�YR�ـw�^��"Oꔃr�Y#lT�:F�6l��@S"OzQ"��F�Q	�-���G�nc"��"OX�� �:DE��*�@�[Ir���"O̼cR��.Fz�y��(VH�x��"O���� �q�5낍�2A`��V"O<ܺ4a��OO���P-��T"O�(2_f�8� o�`����y2l��|_�}�ׂK�80�]��"O4�y���hP�З�H6�L���Ǭ�y�c�.|à��9?�RE[!����yr'	 ��)h⬙�i��!D���y�_�)M���S5`�z�bΜ3�y��˱@��2'm_,AtF��Hγ�y.-/��'��$+0��D	�y� >FP2$Ct��`d��&��y���v!AڙB�=�%d��y�1d#TZ��. .j�����y⠎('k ��� �{ߖl�A���y�uY��m� |;�)�y�H�6���
�9I���Q���y���W�L���>!��01�� �y2*�]�u��G/|yK�# �y�oC�zxɒ0��y�X��`U-�yR��'`o��3 Ǉ�r>v\2-��y"Œ6S!>�%�6x�����"S��y��k Q��	S7oq^�����y⦅�
@�`Q�j�
�@����yR͙l\L'��
P�����/Ď�yb
��Gx�A�m In���� ��y��Jv'2�@Te��2kt,�w���y�G�^�M�4�C/7��0wĄ�ybޑJ�܍a`�_%F�n܊�-�,�y���\�����oP9GU@����ʒ�y
� �a����Y'-(P�S5.�F$8"O�t��a]�&�FC~���) "O�4[���8+c��$G&ZZ���"O���_]���r��:kI�1"OL����edD�vN	+h\�2�"Oa�B.q�X���G#�v�� "O<Lz� �3��D	�N8�~I9"O���[�n���c�ӡ@���b"O�p�A�P�1N���C�4�H��"O�4K��Oj��R��� �x ��"O4�!�O[���ݫw��.�"OT����V�@f�P�S��DQ�"O\y�	K�{��Q��Ax��!"O.@SqD�7j����͑*=�i�"OT�K�BH��>;n�!�,��"O"�J��:]g�����'F��#D"O�%#ǮιG�XH(-�R]7"O�a�5�@%2@�Ye(�11�$ ��"O�(�7kfexX�B�L1M�U�<��g�8�4<����#-q�� S�<�A��9��i:L�X��g�M�<1��6=���0J�3o�<4x�OM�<��Aƃ\��fl��#�Yp��p�<a�@A�JDb0�U�ٵq����Al�<�(��9(���g ^51�Q��*�k�<�T�զŔx���21%&Y�E�n�<��ރ� �" 	[2VtX�$Tl�<9	�01r)aJF-dm���FdKq�<�A�L-mR(�0a��Y�*��qXk�<�LWh��9�*��/�v����Lf�<1��ͼRo�UKq+	�|�����Ea�<�_�D����Q(V�jʚ��]�<�r�^L��p��Үs������`�<���U<����k݄�R�	JB�<p��?e���@fgC�5���H~�<ʆf�Fi�2K� xj�`�d�@�<��D� (5�ŧ�1�&���G�<YG��OP&�[�L��F����F�<�$߃Y��d�֌J�r�2�ҧa�@�<��̕���`1IÐ�T�I�{�<Y�o*V���e��1��+��y�<�BᏇ7��!� ��I�|Az�͟v�<���^�d�r��0��M��	׊�\�<��E'I�.��*Qt��t��$�Y�<�`�ڏGR�pq����d8�iR�<qQHY�U��D�!!ЇJ�����Q�<IRf����H9"!ց>�$)c�LJ�<�#ę(AA.��NZ;/_�=�s�m�<Q�	I�s( ؃��P9M-(I���j�<��@�~� f��6q��$a��NM�<��K�\��h��mM���qK���K�<��珒2�P� ��ÖmK�GP�<9�A�9�ؙ0fҹ\πAӅOE�<	���j��E��5j�9�&B�e�<�G �v^@18��ܪ$��i@�@�e�<�W큾W����m�5�h$�ө�_�<�� �;Uv�!	�
�U���D����Yg���v#Д~U1:���� �dą�@4u��� �[L4R�I�|@2��ȓD"�ɱ��:�h}(r�Ç#ٶ��&!�MBFl��d�, ���9�T��ȓB��5&۫F���3$�`����Ll*4�6�Y\bEX�X�.��ȓ<I6	۲Ɏ�f�,��#JN���S�? ��acI+]�F���	�8�@Iɥ"O6��V�G:`\6�K��[��Lp"OZi��:�	)�fW	�`x�1"O, q�F[�v��!������p6m�<Y��S�9ᔪ�-#���3e�e�<)@%ۦ1$��u%��Hp`g�k�<��aXu"��QĀV)RR�3��HL�<9bB2b�4��֋S������,[J�<�e�@&~�����J��I ͒�y�K;S69y�2���&�
�y*�B"�QE\2cy��Ԍ-�y��Υj��x�%��"oN�1qg͗�y�M�_2t@SA]483R��1l��y�ɿ2{:t{��C0`�vU� ���y��P�\"(���NU*/����y��W�#pLp�Ϻ ���rd��y����b�d�rk� 	� ��(���y�)��PY�t)e��rM\���X�yG W��i.��h 6���j	�y2�QV�!R��Vbt 􂜯�yrM ƄЛc�LH_P��4)[-��QX��X����Xb������;g�U���,D��	�-�3�ҵ
�\�b����Ī������13< U&�`X���Ŗ֘B�I�s� hgo��k���@N��cZB�ɋ�@P[���(0�X[aD}vC�I^�~͈f�/ܪ�P�޼9��B�	&#_ޠB � �3�F�Z��_r`2���4�,x&�C�L�t�^�:Eɟ�6K�Ԅ�IQ�I[�D	��3�X��r� �FB�	�o��! ��,iL�;�D�:X��C�	6PʥA��Px��2��e��C䉵Gb̐)�+[n8�s��||hB�ɽc����sH-P0��
Ѓ^8PB�Ib���p�	+9��#��άg��C�I'۠�+�-�- ���`�O ":�fC��s<�T��쀤��@�g>LC�I+'�<�I�T�7��������<C�	�.I�ƍ^��
qC�B�C䉡q�0ѐ���p���
ǈX�_2C�ɵY���3j��?3�� �D��B�I�s� �QR-P�C���S�&�*^i�B�I�g�DqV�J�dWx��lQ�urC�	������J�e��CȈ#��㟀�鉥,�.�S�e��T-�R�K�~��C�	a�4��5A�xp\�"	�"I�C䉂Hh 	7�p��D�.[�����5|O�b�LyU�� =����f!B�6c��)#�1D���kũM'��"��_��x�Fd3D��aF�9ن�s�Z�l\h1��=D�+&dm��mX�&T�T|�d�%9D�4���"1�z��K� ]���f�6D��QG��g>��n�<:��H3D� �'� ��`;5I�U�6���`2O#=Q`�:n��h+�bRpt�+3�c�<I5'*m�~Y�ɗuH�5�`̓�hO1��(s ����F�`�L�D"Ov8�v��\����)� �h�¦�Mx�HPnØpQ�Ӧ,�
o�!;��&��<��.������4u�2�A�%A���
O����8�E/G�FR]��"O�[`dK^��ʑ�� [ YQ�"O�]9��׎��AT)q1��T����4��'��?�e�Mu��4���a�JLeM'D�� R�G#JT�[�D�`$��p"O�I!6��m���E�H4�0���	q?��Ɋ�i �Zΐe^���g�MP��B�&Y��ٳ*�o�~�ªS$DI���'��	N�O�H$C�JF�63��Ba"Ev
L�
ד�~���t��K�9b���Ç��^�� ���O��3�kh �%W�'
�>��!F7����c�h�B�i��x8��#�O���u�T�G9(,C��&���B�\��D�Lx���U(^�Ef�Mj�L�H��X�
?LO����,I�S�p1"��U�`��`�dK>D�\��m�.:!���),;���f}��n�G~��O���&�F�����<�zS���B(,��ȓUYى6F_=	~1`���^����hO�>��v�buq���%�>Aa�F.D���`�L�0"����	�s�޵��g�<�
���TX�l�`��xI�:�L��IZ~r��
@�؝���y��
r��y",�n uH��'uԵZ`��(Ox�=�O�0���	�irJ��6$�8y�ђ
ߓۘ'�a"3'P�LB8���vr�B�l�O��"~�	�EO������
-��P'�ě��=�)O��	G� ���v�N��a��#o:��	�'��;q����q�#eF`ě�}�̕�I��D0�	i��+r>�@ZU똼@b�� ��%�jC�I#k�ʡ��b� _=U�4 A6P􆸰6��IG�t��P�X�E�O����N �+_h��$�O>b��"θX��9����;q�܊�O2���ns�6b��E|����{�ܤk�M�X�$X���p?��ON�
�yq��YՊ2plP�QP�X��N�S8��#�E�OV�,��Tk�Hp�a=�O��W�l�j��D$e���Ï�TJ���M����Z�J�Z�HϬQ����@���D%��<��� �5�6lb�%�$����	n~b8O����1Z>���E�7wQ*��"O���щ z�n���">��[U��7�S��҇S1Na��m���M���
&]!�ď</�底�ɬUx	�#oK\Q�D���ʑY_�a�"��P�hhG(^n!�]e��	�Ά햔�1GG?h\�'ў�>���DB�l��\1vlF�|$��(D��Q�o�IO�@�A�2*� ��-3D��+���y*bkߔ,����1D�qW��){�h���h��w�o��C�$����D*H��!P� L�E��B�	��X� ��.^�mY��go�B�I�:üQ:��as�a�2�J�m���� ʓ'���Hq�D�#J���� u��u�ȓ��,F�g�\i��y�]��nf�)���X�2$A�Ⱥ!�Y�ȓHGʁPР�~�0AS�\4�(4E{��'1��S��;*�z(�+��c^|ͨ˓�(O0W�Q�p���6k��W[�-A�"Ol��T�C�8��j�J@���r"O�`%.�$��S��+%\���"O"���YG�͘�@�8�~p�"��Bg���Ә*��u#�c���
5��l�*B��`PCA�U/2���J �S�a$B��7�ʽ���ˊ<"6���K_��C�	�� ���U������ޣ{%�7�%���r�C������}T(�R�K#D�0�+�H����$�<��D7D�Pqs$�=#dt��晪m���f	5D���K��B��sda�q�M�6	>D�p
���cZ�e��9G�Q��;D�� �p��gJ�1�6�����UFP٘�"O&��'DF�$"b�	�	�N<R-@"O�%��X�2�P�r�����q�"O��Q&!�+w�<0s+�H�\�� "Oi���9}b���SQ�|蜐T"O��G��DtI���9�j�"O��h�&� ���Ѯ�1�\űp"O�t�����o��# �>eJB"ODӦ	I�AjdDKrL����0"OFa"q�F�\�F�p�ͅ�i�F�A"O�){B#J<>C���\:�}�"O�4�Q���&(T����~6:���"O*5�"�S�ja��X�FH@=s�"O�Mx∛'�Rd��B׮E�@p3"O�5�7%�6h2�e��2;�>8��"O���
�2=Y@�cb�A�<!u"O�-2@焩/Ⱌ8���.V�%9"O��{[�*Ң����ƈGT �a�"O9���1(Xb�%8D�ͣ6"O(ї�4�t- S*�-{�ܼ��"O��S�fC/\��Yi��$�pc"O����Ʊ#,�0�-�&B���ɧ"Ob�h�ہ`RZ��ݪq�4��d"O\����Y�"`�Ӡ�M��TQ"O���(AI��q�K�W�ZE��"O��'� .BH���0T���qq"OH�٧�H�j�U�@�E�"��t�r"OڅHR��6:�.X� �S�k���e"OY�ąͼnTm�AQ�Sv���"O
dS�g�2��n��F�V�ڗ"O��z���L�� ��Ña�~Q�"ORՃoE�~��b�jŤ��Z"O��Y�HەY�˙;TyY�"O*�0��ζ�bmq�I&r���"O�E��a�q
I���ܲ^� q�"O��b\�cGDi�KM09�hA1a"Of�j��T����N}8��"O���Ȑ>�ڤ�GM:0|2�i'"O|���G� e�y���w�А��"O�AiTLk���5��UeU a"O�x��ⅦQY
��ԫ77V���"Ol�(B�Q�8f@E��c!�b!"O�a1�
n���
�n���"O.lA��	g�B�B��d����"O��QD.�m?&Ȋ���nFj� u"Or�Stf��N���B0�8�����L�<I�]/}���
ֽ%��a�OPP�<	��wBR�����*�cH�r�<I�f�����ʑ��y +�u�<�EҾ^�9�#�]	��,aA)o�<�q�A[�z2k͈I$.)�D�R�<���9y�����<9���@ C]O�<� 鉸h@����5�\�PDS�<�&V�!^f!��g���` �VL�<�׍Զ> �Ãړ`���f��K�<����%^�� KWo���LE�<9CM�on�D�[;� ��DfD�<���
�ꘋ �H$�� �~�<�vn�2p���LHF\��9���d�<��Ԫr��[NT�6�f���A\l�<au�Z	'�}�Aʑ�m�|Q1�]q�<��%)db���Ѣ&ؖ�S��Q�<qG��]�|�:�\�D�X���Q�<���'P�n<{&�L�&�lbb�t�<� ��92%V?C����.i�4q"O��xp�����FX�op�9#"O 1cnЍ|�RX;D��La�ds�"Ox���צ��e��ጽ^�*��S"O4�3�+D�N���A���"Ox�*�L%[}�����R�\�p5"O�á?U��d��ǕF��0e"Ov�a�Ց�����b�$e�2R"O�!��O_*~Y4<c��֒3Y�ݣ"O����f]�o���WB�&opy�"O��R�A&g^�e��BS�oZ�H�"Ol���T��D���I:.u"OhE�bK�b ���"�[�tȒ"O�����I-!�H�⁖[x Qv"O4�$��G��K�
*S;����"OL8Y��K���}aR�E�S�(a!"OZe�th�9SH�JέJ�Z�Q"O����&�ZSj��6�>e�"OD���D�,}�:��H�hpv(�D"Ol|y$�PJe�@K�QN$�2"Ox��1&�5��SK
�Q�uh��IR�O	&�8aB�+G��i��;"�P�C�'/p�dM�T��:�GA�-�bݐ�'��d:����?�y��5D|ڳmq���:��)D��{s�Yy�@�Z���<}QZ	c�E&}r�'�~���^	B�6p���&^��J�HO/[/�}�>OQm����Dj`��'@۰�p7��4���?��S���dê8��d+!0��%��,kfa}r�>i���-�x���
Z,� ��RVo�<�#�q4�U�"��H>j�g���<����tվ��Я�"���9VI�JiNB�4gxIB��	|>�eC:6/�C�I.Ӱ�Q�O��o�x�0D_��&B�	�ӆ��G�N}��I�W�B�I:.�ά����h_(��n\<R�#?I����$Mb\H�fK�su����S�!���Mځ�eB��+��y�M��!�:9�� ���t��4Ɠ�!�ZG�@�1P��d��Đ ^!!�$�Z����e!�, ��ٹ0#�)>!��.0¶I�Q m��j���}	��=E��'�8���#� �%���,�p�K��;�S�$d�#8��t �b��u06XZ�Ļ�?Q��'�h�qH���( WC�dI������%c��ϢW�FdSc�-HV(��ȓ}Y��"�D�4>0 �sN�7<����2h��x2�]n�= �� $<2h��	Dy��K�6J�Z��RxQ��q�l��yb��a�]��l�xbi�n��yB�R0j^`���B�v	��j�I1�y�-V!V�"�HqDz���b�͜3�yLH & ;��=c��,��$V��y򦜥`���:�H�er���G�y�dL]F�EaD�]�d�"�	@��y�g z�&ɂ�g� 3ͱ&Nݴ�yZx"G�6	��XF�C)`C\5)�'��u��u�r0q�\瘥��'�-������*��Q���"+���'k(�qP��<�1pf҇�>Dr�'a4��P"ʁ��)�� ��`�y
�'�b|z ��$6t��b�`ӾDa��'*8�Qm�C��y��>'7����'ӚD�q	�1��S�KJ"��0�'ؠ1R���8�Ĕ���?	 �d���� �}����^�����	���a"O�P�vo�Q%8I!�(T	
M�s"O:�P�ȑ	P�d�t(۹�>%C�"O�l� ���@�X��tI�5�����"O`��W�D�F�P�Q���=u�D�"O� �/�91��T1FQ�odj�i��'���,	nՖnHȑ#�K*^��̸�&D�|Qa��$	��ŀ���rP�3�$�d.�O A�� �"<��Җt����e"O~��a���q���r��^,c��"O����C��d=ty�F�ŸeW�<H�"O�0J���P_&��dnG�4V��"c"O�}Q3H�03�4�LU�r�T�7"Ov4����	M�$ *��P(��3B"O��@V��(lQ��:]	�@S7"O��ڤ�$jy�Th��Q����"O���0��gWf����d�jȓ"O�C���E����Q��7"Oxi�.� �E�Rzs@"O�� �薼A������5���R�"OH\3���(� %�S��7D�0̘�"O���'��!X �H���v,<S�"O`EQf�'.I�p�S�۶z.���"O|�C �&:��dqv,�>]*j4xP"O��1Co��u�J���m
큄"O6�i���.J1�D��L5_�a
V"O���Aj�8RϲAb��B2`��7"O�	��ɝ}D�+B�̲UW���"OpQ'Y2>�$n�x1B�m"D����#�ݤM1� Ue׎�� 0D�4��斳O`��aE(&f���*-D��1@�����
0�I��j��*D��an�#HpI��ā!<-n��Q"=D� Zdo�er��A�*�1d]�&0��0<�$e���N8�q�N�2ьa
���s�<�R腇 �|���7cj�,rQ�YG8��Fz�@�0�v����d�ta�'�<�y�)�^�NB0�����BaG��y��ǏS����%�K^V����	���hOf���U�|�D��=�T�Z�Bڔ0N!��ؒ-��y`bP�^���ӗ�N�)!�	�7 ����l���! \�!��q�-���;�����̰I�ȓn
��37'X\��Ν�H%��ȓI�,�C� �aH�@�BG�7�݆�ENTd0�c�.f ��q��-2( ��M�҇@a|%�E؂i�b|j%��<����9S�Ld��y;��F" t�]G��Ob�O�0|�$�^�|䰄+1�N	<����'ܮ�Bq���Sql��a�;��Z-O��=E�D�ֺ4�FCQ��V�"D���7�y��!g�<������q��ۨ��'��{rm^�)��e1U;0[���s�ն�y�N�B��x���Y&I��E׃�y��W�z>���^�MrEx��Z(�y�`�+�f����E,J�v�����7�y�k̓XyN�� A2�T�p� ?�y �Y���b�>
�}������yB�И-"�y24��7����V�U��y���sl�*��w�$����y�GK�S��+'C�F���5�b�C�I(H�r(��N�V�T8s X�L�RC�I�&4�A0AU�� ����.N��C�	Jz�&�/�DT�Rf5FtC�)� ��름�5Q��X�Ï.Rv����"O����A���ft1�რM[� "O�U�
�b�QE�S9E$(�s"O>��g��Q��PA/c-�q �"O�-
Re�q�4��NڵX)�}��"O���E׎q�Ƶ�0,�^��"O�� q&Ԣj7@�pT-:�h�T"On�C�D�>@fd\�j`�@"Or�C�K��1�	�S�
�7~)�"Op�����d� V�-�t|zP"Ò#3�ВŰ*6 _�fP��"O���4/�{�ܹ�MB"�u[�"O< a쑽?����Yw���y���x���hI�H�Y�e� �y���=t�r)���O�9t�Hw�)�y�+\�(4��!�_oP�Yv�θ�yr͇qAD	����jy���B�ݧ�yҥTI;=8��5o�4�' ��yB
Ciج�
�n�,�Iu����yҫU0�9[fnS�c�NM�n��y�##�}QA
ڗ`d��W�6�yB��L�V����)lJ-�g���y��
� M�@�y�|� g��0�y�N�k��LC�)H�j�af�W��y��_�A#��Y��<k�0%;��
�y���qP�����	O�Miŉ��y"�䮱�A��<�"�Q�ș��y���+{���"����(kX)���Y��y�
=~Y��̵,����D��y��1i (��%���yS�[��y�E8Fd�
Exf"��i���yrÈ�%sX�;v+ش{3�ٛC"�yM]�2@���'e� ��<PÎ7�y�Ɗ�A>f�:�
2tlh2�؆�y��@2U|tr��&L�!y���	�y�*��(�TX�e ˂[�t��[�y�'L�!��<���<"�uD��y�k�7�l�Go��ac�Qat��7�y��d��u���� V�Z�h�$Ђ�y".G�����֡Jߎ���S��y�I���v|��
O;�h�b� ���yR�0H ��	�NZ�e
�ؖ���y�m�8�i�#B���z���I
��yB��+.>��%fK�v�*�*ra��y�M[�Ox���n¸ >��(BJQ��y�hY^{���v�(�T��fH��yB��ufԵ�.�'����vI+�y� ���Ӄ�24$Ȣvg���O��yB�ɛ72&Y��C�mx(���'�b�c�J�]��k��2f���x�'8�uH$�Ձ|�����X�-��'�x��e�(ax|8W�ЀW֞��'"��U�
04M>U�vl�F����'~��@�韌(�`�lK�=�F!��'i$�9�# @�*M�Pj�!-X���'P�#�!0Mw ��#�8!�R�J�'ov�aV��?Gj$��ꃫo$f���'�T��d';F/�i�˖�`󌝘�'/��FֺX�%:�/�*]n�)y�'��œr�� �D�B�f>���'D��6
Պ��(K��6��tC�'���c�O�$��`�(5�v�S�'bm����.��<�'�� *T8��'�\	 !Fʗa.Psfc	�*��ٚ
�'g>q������F��&ΐ]���� *U�2d�+2Mx�K���74�b!"O�R��s��tД��+/�t"O���q@ʹ>�9PB
�S:�I$"O�t1��Z=KW: � (�4�~xs0�'��p��*h8�����O�9�f-0~T���!��!W����"OT��W�Ad�)`e-��&L8��� [���$7�A�@h*3>��F�aC�"���� K%b�x �NX��y��"0,�j�&D?4ӲI�6��z�8"󠒬'o@�Kmo��a;H~�=A��H�o�,Q@�VL�肢�D�<٥�'��|J��I(Q��¦���<�#*��+����kZ�_��<�F��`h<9���3HqN�a"F
<lZMB ���y2�-|>�8��Ʌ2�6l�����y��韊e�?yCd�8e�8��jU�B���f�Y�<����Y?8�b�ך7�Q; gURyR�e��̰���I� DO\Ay��[�ԃ'mM�l�}2-�<9�Ζn� Xr�
)IC��R|�a�z��	2 T��Ϙ:$���B�]1�����ӈl�����[5UE�!R6�Ǵ1�(ۖ�=�h:R�)#�f����ۊW��i�3�v�h�Dz�O7|Uh�{"��;v�l��
	�^q��ƍ5�y�H��P����aO�������$v�8`�/�S�'U޶= �"�rK����ʕ7 4BɄ�m>��F�_,\��쪧���M�?�"V`8�4�SoJ�~� �s�*�mb�cb,4�X9��WSޭBe)F�;���&�L�qDC�Md�����ܬg��- ";V���D�-f�qO�L���7Pi�5���ɑ@��s"OZYxU���]�\��qΗ�)��ѻ��|"NW��Oq�H��hJ�n��4�2G69bF�[�"OH 3������	1oT|	���$��@�x�Ɣoǀ��M�g��S�U�PnbH�=����h���D	<OƉ�P��\~j���ص/*�����'L��"W(�zލ�Cנ�:�����s��l򀧝x�'�́҉{���oJ"�`��I'����4BϦ�p<��ㅗ$t�$:��S���Dzװ� Q��f/��PD��?l�'+��X�����$hF��m &C�b�F�Y8O�� M��� m��s�$����6,^�1�����hw�y����p##�<O^��k�10�B=*����+�`�J���K�>�'��MivKW���Y ^fµGd$\�R)[%V%�&�@��d����)�\A!1+�S�4q&����l��⏔�B��	S��b������D$4y�g�6W�(�Jao3�v�T�@���HE�ċE=��� Ϳ��HA!fA��X4dV5����<�}r'JDBv�CŢNB���BmYXy�nU
9I$�s�˷`iҝ
��sq�p/�7��x�aY�'z2���Fx���T�է8�cI�<���
pЮHLa"���O�Kqˌ�*��1O^E�uLZ�POR9PC��4��IP8�O�I�L�u��A���N���6ϰM8h��X7]�>�)��-�Oֱ��bۖR��E�\K~����Il^F�R�@ws>�AW�O�|��C�|�(��bZ�(���CE|�<)uIQ!�.9Z�͜= 4ISzy�(ݶqA�T�pdh�@MBD���4�Y)ҟW�
Qs��,"Z`�'�
�ߓ	���XQ��R����*����0]�����'Q�0�8�T�|�j����>�ꥁ�t���D�����6bv����P�0�!�$�#E��M3�� t�x��Co�-�e���[�RZ
xI�4y�d�#-�Ri��K -�D�8��$3�L	��p�jT���{i�x2��|%ʹ�Eֲf{���j��f� �%
n��]�i��rm���1͐Y�Vx���&N��
��P9+d�h��E�lOT�B���pѰ�'��ׂE�J�]�ѨW(J���4�<�+�+	-3��IH�H����xb�@��D�H�"M�Z}SwO&��@�q*U�ڸ��y� �={�x�]?�ۦ�i�%�7�_���A��o�\l�A9D� 3W�)c��ҋ�}���9��԰v~xMȂf+��7����^c>��O<�Pj����a�!��a^�My'n�\<���)�H%�r���)H���/ի3�����
+*1A"�L�\�3��� �)K�W(Pţ�%� �T��%��_u��/�a��*�G�l����"T�pR��0af��i��!�ğ w���L[>_��!��j�,u��	�g���
un��R$x����=c��Q�m߯S��B�"�:����W-:.*%�ǭ�5d=d�[�e�ybaJ������&^p�\�	���(��
-gW�|�%g�-���" ኈ��&\v�@�"iY-�y�C٘Q�|��acP�_���<�0?QD͞�ԨB�
L�b��io�t��!˻cd��i`�ժ'&|�f��6-��&�˞ R�b��$Zm�j�8#A\�d���ў�V�ۯ^9�`���3��<�W�G=m��2C� } �J� Z�u� E��07�1��(g�؀:\O`<�R+�/:�2P�M6-4�p�2�iVlu��B�]
0��veG�	^�����[!f���hSz\�����ETh�Um��V�p�VFZI�>���G'D�'��k��ё��+C8$*�oD�v�ָ��ʙ����b$C�@�N4I���i��ũq��.N&RT�e�u�'8K����H@�eSZ�E�%�O���C�Y�:��sBFI&;>�!8W�I�b����ĭ&f�l�ӣ�v���Cv���@R�
����<1�P�J|̓R夀FͶ-TX�+��[Z��qFz��(q[V9{S��-#�)�M�.^�&�Rץ��X�P<��K��x@���6#	)y����ul� ?�����)h7���DY�8����f��D �ι�6'ܗ|I��y ��/��Aa\1~�Y���	�re�u�5�P�+r9"��U�ފ)�zI�֍H.a��C��;B�Gd�Aݪ�ua��|k��[d���vI�U[�-�![~�ΓD�	!'��6BԼ!څ�F,{d���p͒�m�4%�"]��e�
�����˃7��+�.� _�q�bɊm�v��1!xD��'䘴�&  9g�� kR'��X�M��	j
��<Ip�0]F�(�&O���Hæ! v�'�=�qk٭$a�]��΅Zn�]�������Z��( ����Fo��-)�X+C�Փϐ���	��az����G�v)��S5fܘ�Z��M���Az�I�6LC���h3&L h���*��$o�0�	6a��%��H��F��Q����6�
�9aQ!�E��\���X#��!P��S�G&�84I�6���1���:�I�Kp���LQN��8I	��y'��n<;�Lŗ,趤i H$��>Y���L}���'-�>V��D���9����iّQ
��	��9`,IĔ�
`��(m{8Р��͟Ҙ'!���`���sM�ȶ�0���l'��VZ1g��4���K
DO� ��l��m��#�H���RGD�&�!���Y1\}�4�.rH��ӓ�r�
lB�_�t��'K�jСѨ�)#�4�U�Ƹ~�ؔ�G�j�b��!Y�b��ߴ��7M������ɍ�@��= 2Ä�֪L�!��D+"� �R�J[�V�"����8/1R�z�L�*A��1H�k�l�4�dL-Z%m�)X��L�w�]�y�K��-�����'T�DhhwaC��0>!e��:"�U�o4�Ё�p0����մF�6P��'جۑ�^�(��	Zg!S0	�L��2�z���y�l̾3����L��-rdS��O�|���{h6 �c���Z#�	%kv����&�Q.#���=e��Y�U�K~�1i��%� ��h�^waz�!�*J�x#n�#%�����Z:��dI��e�B��΂~�M���M�D'���ÇW�Jh�K8_����C<�X�X"O*�(B�]?(6��W�4α��JC
%����cN�M�²i.&6m����I���I<���؁n���y�op�*4�r�͖>9���Q'W�a|��Ѝl�,��7�q�ŀ �Ƨ6���3 <U��(i��_	R���^�9s��w*�"�������Hb�!�S����6q)"\�l����'?t�0s�ƅ�S�ft�f�>/� ����Hs�	�L�
����->*:��w��8��3�d�	d�V���|)��`��TC��xv�U	l��ا�<�B������%T߶�Y�A�2q�M0���<#�a:%͊HP��E����s➦QԠ�P `����0�۝\n$\�e�æ=,*���ȤW��Ɂ�BXC4`��V��(�.	>?��%!�'O3�b8 ne���s�pz���.Q�� �	>8��aWG�4�x�;�����l%O���8�&�Mr�p��I5��L�SfJ	_Lĵ���R��T\����	%���K:~+$�K 
�N�وpBJ�/1���g��9�Bp�4��.���rC��Mӳ�.-�	�ˆgҪ�RG�P�'��0!2�	QDC⬅ĲyI�%sD��!��|j^9�զ65�St*���� \b0�9�c�@�4���cH#=a4��0
�ݲb�lR��B-�F�P�H��-��|���@�*٘:��D
4���OȕhY���'�B�`'k�	�IR��I�O�H��T P�p��!� `��'�#cȑ2�,4Kbf�:H����==8� As��3%mF��c�Hy�͸˞�y�φ.���.�
X9�錠0g�̺+�D���\�1�0B��6�P� !�L�A/j�١�$'����UN}BcL4v()!O�y�l�h�F�#8��8�gӑg�ڑ�w��
j��ӂ���S���x%	,G^�DzҢ�6��Mj�*ueb��bf�$ R�8����	�'U8G[�2���/�VQ��_3>~L�D�H�e� �� ����-�Ӈ4�h1���֤ѿ8���`��W1�J��ɏoI�����s"hxSL��o>�ɘĐ=;��� 7R���'�fI��SX[�a�Qk��7(|�3��
�.Q�Ņ'��{�B 6�hhgkU�[�jR�	6 �cn�q�J��Ekע2 Z��r	*6�^�lJ�B
2-�+�7#b��ȋYK@-�5$Ĳ�p?�l�/W��|��瞒=:L�A"˨FHU�G�w?ّ��M{d�'rZD�t'�6,`���
+@ZI���6Iq�aT�D�2��,�ED��8�օs_�"?�u"�_W�9����܈L�j	� �,�%V8H�����O�
��id� Px��4��&��`��(�A��4:��ֹK����ŏ��V��XF�E8P�$��Ъ�<)��H�pn�*Y<T�[�8g9�Ap!�'�<���Cսw=�,y�Z�A��X���P�@��C���
��{J�\�Ra� +N{���F��g�X�OT�����	��<avJD"X�@E����}�頷�Ag�7�U&P"YJɣtҌ��#��y�lA�_���A2]�x\hrG���?���X$��� �&&|��6���_���y�a\3~DD:r���o����O�<X��#�=w:�DN���=����� ��A���^�|�!��n=Y����1����s�.�`��@��F���#SIK�:^5���x���o&lG\M���
�BS�PCd���O� uf��99��ң(��DQݦ�����7:�����+�.�1b�Yq��s�Y�S+� ���_��A�끰/6�۰� #t8����U��r�C?� Z��O��� 
�u�@�;qP�P5��!
� �= ���ՁSwa����"O:��D�L�H���� N��̔�V�L�7��s��xf&4��;|�9"cQ���i�Y~��Nۼ?����G��N�}�' �J��5A�V� �&�e�Q��]��@pe+}2+X�7 ��}&�tK��'_VtЕ'\�D $��H0�nh�����N�O�H�"��=
��y�"���X	R�'�f�Λ��Ɛ3��Ϧ�;�'*��i�� sr%��EM�
�'+Zu�`Z��N��GO�=*����'�.�Zr� O��ȹ6�:?�|��'�|�b�_:h.��j����]��'�yA�nq�Ӆ	Ǭ���0�'�h�`lԐu��	��?6}I��'%l����G��`���S�h���'	|�y�LāO(�(���"KN�
�'����"�,�`1&
��H��'�>���ظ(S(�+���"��'8.t㶡��i���ܘ���{�'>T�%��s�͋�%Fz4�L�
�'v<4H!�'쀝c��6$�k
�'��h41TXYR�U<G��	�'��×C�W���/u  	�'�~0�N�:���:���	hgd��'�VY�dCþP�� ɋx]����'� hb�L`0�js�ǥz���'�荐��L�}�u��eK?$�2p�'���ɦ�r�@ya-�(NIS	�'$j�SNGa�<zsm>[�
aR	�'jz�r�#�*~:$�{���,y�<�h	�'�}٧U�x� ��c_`���'�^�c6�U=�=ywfP"l�+
�'f¡�ƩT�@}h4�Q�}Y@��	�'	4Yq4���|b�X�x�`R
�'�<	AgK����\���V`�<���А��=�a��8FEt��wK_]�<I�Oi@qaE�X9X������]�<��场W��ih���U%�H�n^S�<���
�'J�Y����lЀ#��[O�<9G�S�����M�5^��" �H�<9�O�N�l��M�"�ND;�LG�<	��!����#B#O�hX�a�JH�<'
�V����b�1#rh��D�<y`C�6H�h���%oʰ�sVc^D�<���_|���"I�s���`����<��ZN��lR)5�H �`�<wj�[�	+s�H'Eݜ@bRt�<��Յ}�
�a��4�p��Gk�<1��_�G�Pp�U�VG����*�k�<�č�tq��Eĕ�rw(�� Cd�<���3@��	c��3v����d��k�<I�nӿ6<����H�����fM}�<��H)/@a*��U�a� в�}�<1�M��Yw����:���"A�}�<� \I(�ჽ$&��k�H��=^Jiʆ"OPZa��Q�h�k���[冁�"O
Y:���)2��-Ȱ�J�^�� �"O
9�C�-o]p`��s��m�`"O������ʜ�A�Շf��C"O��@�׊[v08�PΘ����"O�ˤ�T6T���"�_R�RHC�"O� �#������
�h)H3"O�p g��B:��y��8;�0���"O�,��O�fJ1�p�@&���"O�В�G�e�
�hp�ø� �"O��#s��f���0`~@ܒ@"O�#��D����L��*D��"O������8Hr�ɢUOO^M9"O��چ"��N��1sP�׵ָ@y�"Ox�a/� ��h��� �F�1�"Ob�����r���-ch�s�"OD]�5��<��Y A�3u?�hYF"O���
�6����a]o��tó"Oč	�C��b�B@qro˺=�X�s&"OZ�������"t��G(����"O� B�ʻ2c�5�'�K�;�N�#"O�`�Ы�]>�墅��.���{"O�QR#�+<8R�`�:��1@"O�=K�G�1jjf�
6�=ߎ��"O0���)X>a� ���]L^ ���"OH:w��X�6i���Qh�~3�"O`���-�(Rh���G�W�o�ܱ@4"O�(X�g�;a �� �D)T�V	z3"O�9i���)E��BG.ەxƦ�"OF����R\0PQ"��[<Z�0���"O�U�$���W:�q��mGi�J1b`"O�ub� ì.��]{1�L�tC"OL|{�j;U�T �R��(?Pd�:�"O�QHq��>��,���(�x��g"O����`ˆ}L��-ܡW��a��"Ot�h�@�BeR�h	. �h���"OT��%Ǖ`����tq��(�"O8}�Q
݆�Ag�3��9w"O�a���Y&	�aj�G�>aդ�!t"OR�+�@M��j��� ��_˴q�d"OʡP2*�&�}�'Dفf�(�"O,R���B�0��س-
�O�!� + �l�'HD�J�H�+�01�!�DM-��gh��Nl������I	!��H�G'���dً6B2a�uK��!�޺�6,�F
+,epA�H��!����Ґ�wM��� 맊��8e!�$��F U�PM�8~����ʅ8W!��ΓN�
r��;|���I�o!�V�rx �wL�J3�\� �ȜK!��ܛ$�q��Gܙ_:~��*V� �!�d�������"l��0i@�t!򤑌	F��p�xX�Zg�A�p!��I�c�tP�%�A0^��--9!�dYL�
�	�c�=��1`�ؔEZ!�D̂$�p]zU	T�5� L[0*׳L1OHKjW�N�$X"*�e�O��j��M�v�P�?~��c	�'�L,��(R�	���Хͭk�ҩHQKă�*Ż��<��H�K���I/�r�en�$ ��Ögž(`C�I2/@�@`�|-�UץߗF��H
���
J���B�$rX�qy�Yc���%K�\�YS���?�Ƽ��	�D�~h���$ �(#��V�-�\t
4m��l)��[7e��b�%4�����=X��5��0=D��ؤ�#?٣��&br��s!iB=$��w���<���� $|��Gv응���M�J%[G"O ��ʅ�93,-�%L�2�ȼIe�.�J4���Ӑ|]��C�M![1���%��S��H	`��1͈��1�)� �3T���s�"p����di6`����H�=��j��H�kO$,O����Ƙ�gl��D\Ϭ�W�ɚb�J���&Ӳll�F�
e%b���g�f�6=�0
3}�2�
ģ*}!��:r�i�0� �W�+���B���'������3��kRE�s����Z K��up�J? [��S�k�9���]�h��x����te�B�ɤq�p��J�N� � �$~�qb ΄j������sJxp�ڥs�x�'O�#����s��ݛZ�8����F��܉ĩ�xɸ��μf����U)O�mh����@.A?�Ђ`.~�찓A��Nv�j$cL�K|��w	�:bv��$'�m�bw��`��! ��Ը1��3w�QG{b�؜d,��h��7:p����h؞�A�҂���*��@>�1����l1�J�1�S	ד �RXQ�Z ���4M,e���n�*']Y�k�~��}�U[0�蒂Q����Iۦ\�L��u ��+ؘ|AF�kU��%�^D(��'t���
K"�̀�l*;GY��"n��9��
�H� ��3d��S�5ʖ��J'���Q�<Heb�w����1��<)^����GG�U{�^���F�S5}7�ӊ?�ʰ�fg����:1�<��!�͉l���ٰ_3^ �{#jҼ�Є�����(��KJ�~�9��Y�S�����d��rC
l���æK��  L*[I��	�V���[����3t�,�&�]�V�8��;Rw�5r3Gσ�0=!�h��H�X��F�O�z/�oZ2,;��@��?0������dk�"��
Gh�#�<OD({6��3/>��u��,.hءc2��%?����';��B� �[�>�bZf
�P���:n�@Y���fn!F,��y¦��q ���f��(rf��;���l�KG��������CvX��f�Oi*���W��(k�@I(u�� )�=����P��D��Q�8$�ra�_�f0Y�J�l�^uP�JC���'	 �kWEx�\	eOEW��䠌�d�Й����?!���W�E(JCll2�����r��V���?/|���CP%?@8�C�J�i
��#��m;]�鉔U�Ա�c��6b��#�P�7�;5p>��'�M{mm��˺.���'Ө`����'��V��A*��	|�,$�aQ%
jx S�$D���2�\��@`����=F�L�c��*>�Qp�lE�Oi��s4H�x?���C�c&�@2CF� D)܍+r1��9z䅐�U�*M�P��,k.�y{��'�T��f���@����IL��X�	��^6��ą�l}�B��Ԭȡ�O�+o|Ͳ��@'�����B-��!Q�!�4 Y@��d�$9RQ�@�c%����)"�A�'TZ���%G&?_4���(�U�����I=���Fă�{A�� ukH�>O��k�KA?nFaz�W�r�X����H�j�����&mv�w��u]ֵ��O�"u!RfV>t�B�`�]M���#�⦭�� c�p�KT�7z5C�bK,l�B��M���w�1-!*��bn�7e����
��{��R"�*/�>q�'��3W��HMIG)�5S�B:�̬"890���C�M��I e��9b��S	{��yvŝR�d�2�&���Z���Y?�gkU3dZz�Ʈ�	�� ��M*{�X-c��䎀5t�t�<}�ȪVM��j������f����w���M[�d2��i@&���� KdL�;���(�˕+	���p��3Cɚ�����Q�X���Z�G�p�0$�wV��8��h{��IdO�L��	���	$����F'�@�L�H<i�Mn�,�7�H�s�D"5��jx���]�y�
њ���"ۖr�Ḳ| ��2e�n�t�S�-kӤ�l���M�r��g1�fEݠ.? �{ �m��P$b�����Q�Q�K!�3�+�O�|hR(�Svz� ��a���Q�]����XlbQ޴6;f�Ð�G|L%�k��l���C8->`�����aq�#�+u
���/L�V�t0@��D�O���L�Q�(��M�7���p$`a��H3{��l�uG]$��@�iY�[K�ˇ��5[x�� ��E��$	���O^�pwNK�LZX Y5��ȀZ��t��TeDS�2xAo�+B�@���� KWN,��Á�MkH*���CT��,Mzr ٰ�
f;nXӠ�>GD��g'�O���Ǎ_)tl����A#��1U�ܜ~���GF�^s(P)tSG���W-��tp����D-��Y�4�8���G`@��&�Y����8 �'�R�(�e����<*C�^j�}"t�<�B�D"â#0����'C���@k�J&,("�c��a�Qz�n��T$��"# 9�7M�Mwx��p�
~ћ��
�k;�P��Ǆ1��� G�(����H�dL#�O"ZV�hP�22�H���07�n,�%E���KS��)d�,+��G�\X�0����nM$0�.�^�xP�|&�M��D�V����H�D���XjD6,p�Κ�]�!�di�l�Ğ;!e��L&c�Hqp�a�L���{�� �r��h��Ip�%9�ٿF��y��b����x׉А7��sT�X%	$��{�[� (vO�a�<�з�D��y�H�eIll�q`�+m��V�.�p>!"l�\�������bv46�Z-�x�rt�Z)F��	�W�l	�V�y�Bt9�n�CC�3.ۘ\a� ~�TPr%�284��z�����Cx�ܩ6+���HO iV
Y��FĚ��Ϣ:W�h�e���d���@a�7��Ը:��B�L&98ᘀcA�o^��pc�󲒆��~T��`$���)���-C��P�Ņ�^����C���r��P� SJ��%͏	���QD���@�� U��gGS�&��ؙp��^:�%���ѱ$o*������ȕ�;|O� d�3�C"LD�i2+
�%P�u�$��] Z0��!��(2�EG?�"�P¦�1��ˡ$S�M�e��8�y®�8d�bJ�2]L����'!�t���:F+�,:4���@���W%6)jyi�'٨��'�i:vE2#�WA+�r���6�Z�jT��5/biY��J c�0  H]�3t��V�'Y��hE~R��B����h7.7*�R��J�qL
<����h�i�SO��[��9k�O�!\0<�V�Q�<���%�01�J ��a��k�M�?� �/�jdQ�N�y<MY#�_y�e�18�~��D�M�{*���%PN�3�O� �q�B:�h�� ��5f��t 1'B3;8ȗ�0�d\�[�ji4��3�'\"ak1�#a���b��5Lh\!â�7�Hj�����Aϓ-[2E#��ġd���
`i�HcT)���wF�us3��
ԠGO�9���P
�'f\k�h׼n�ab7e��?���u�p����uU����nDk��W=|g�Q
��\?;��a�5wj6)��,z��F�Ze���cٌ,+#�MY{�@��B2C�F�g��},�x���ñW2cT�ԡ~ft���l�.83� �B��._���'��D� 2U�ȺQĞA�4D��R�j4�Y6ɸEc���e�'�.7-C�0ĺ�QQ�G�-=<�)��N���-���vH�#C�*|����k]㷫�:��cU�-`��C�&�}�tP�3���~m]�4���󵣊�EƐ��E�yw�Q��2$�Yؼ�a�V��ybf�1F�����JB���{Q�����ĕW��H�o�q� !)\�\8⢙�s+��Of�,P��Y�Z+@)y��F+z�<��{�,�$��D�Q��4=�Vl�'K�3oF8	cDD�%�g߈x��(�3��&8�#��3(��ÌY�]h����'~�4"|
�H�1K8�Z��Y�m��Ț�iBU�<�C#��f�{�L�n�J�M�R�<��)H��E3�*��-� �`�\J�<1ӠD�4�&�[�!��a�8�ĭM�<ٴ�,Y��-9�炾Y�hR�YP�<�v��
fz��-�5=�B� J�M�<�� Ց@���8�̄,L�d	�D�|�<1�ϴ�4mh�
�)�Q�3��}�<���R�8	��̄&B�*o�\�<��"�^}�P/��L�bQR�@�<���K		ptx�%�$V�r�c�|�<�uiP>j�6�ңϟ�a�]Eg�`�<)D'��Y��ȣ��r��;��c�<)Р�	H:�`��Zg�����O�\�<��M�*y�Z��ǔP�I��b�<��%?h�I���],�>���e�]�<)��[BND� &�S��A�D��G�<a�/�?g���^�\����E�<��E�b�f��g���_bu�@�G�<ɴ��/j$�P� �)���1�Q|�<A6n@��R�A�T�0q��\a�<�Љk/���E�c���0��A�<�t�K�x�nЙE�X��I��+�D�<iՌY�<ᔅ�t)ț%����ME�<I#�ذ"II�F��M�N�t�<Ѧ�+0�B�u�0L��: #Tu�<F�^?b��Ѣ���	 `�����^�<1��X)�(H���;WO�YC5@�a�<+�/��	����~xj� "��b�<��H�6',��f"cp� p�<�ѯM�L�6��#Ɏd��(@e�<qGM�&P�D�bK�JZ��U��`�<��WfW(݀�	��	�0�'�HG�<�D�}a�Lw  �H�y6
�z�<��!זO'�<"ǏG+un�I�"�~�<��E��� �O��HS�lq��m�'T*2�Aڂ�������@�`����i�*��V��p�f���A;v��Fz�%�t�O�t��D�>�, JB�Il��e�p9OB���B $��0���Z6�H���S�_h���cպ�lr���Fi4��&٭o1T��A^�0B��O���iό �ZDK�ċ�fV�h$ �1����'_N1�R c>=:WB�1�p|)�C2|#��04�#s$��P� �'�يC"R��iU�J��pR���	��m8q`��K��x�-�fk�)��	�0q�m6~m��rDeJ=ۈ���l��c۴GU�����		-��\B��_�ňd���s��vCQ�yb�|���U?� }���$a�PpbC��H4rABL�W?�2O�6��$��N��h�N`qg
� F�<�  �n8���R�Dw��$�  Zp�A�O�u�^>Y$?7m��
@>A ���-V�:��䁓�Z��	�[��q�C���	V�m?���Zh�v,����H��9��������L���툤+:?E��CK%0*�zR)QXX�9� �~�� Y��)'��M<E�$�Lo��;�M�"nB��BfV�W#�<���Y�,�a��ݓZ�<�3��HIY $��/G�@QܓO" ��*@P1O�O
D�B�,@vh��3L� @ld��O���Gؐ�O#|�w����p�#��$h���$̔؟���,�"@
L�6�>E���W|n�zQ��O��^q�h�*��U[�\�"t擲�~R�O�ʈ�5G'���!X��"�̈]r��a��Q?Q�E�P>�C�I�h"vY�L�P���D�d���6BѦ�AJ��#�����T�}ӉO��5�#�!ȲC�i�H@*QJ3QA�<���H�T"I�T�S�	� Xqq�7f5f]F�U�P��Y�4�![��H?��)��s����#��O D�Z��B�4��Ё�`Z�zЭ��=D�����<hdX�4�R85��� wn D��sp���	�du���4*�%�$L?D�����q'�)
�g�+ FqQR�=D���-�*@�.���a0x\zѐ�<D�$S�	�Y�8b(X�#�"=0�E9D�$ ��
|@�HR�21J�R�8D���p�لrD�c���`��qQ��7D�8���$#��u�i�-t�6��a0D�,�s�h���1�ɇ dQСh#/D�Tن�O3R&D�{S�J�&|x;FD,D����-��z 2f`� h���*+D��$)�P��je��7��9(qm*D�,���D�[
P�n�*�Z#�/&D�X!���5����BIW$3����(0D��`Bƙ=1YP�1��V15��Q�B.D�< �$Q�*9Ԡ��̉ʀ�*D�t�q�L		���Jf!��`��U:O'D�x�F� J� �h�h֬^�t�z��*D�(`3�L�����l�p<U#�5D���uZ����X*�N�hѣ3D��:T	�(.�����07nD`�e0D��2���tr����c�lt���8D�i���;ai�4+Ӯ�N��z�I7D�$�7��(� ��ꒇo<�!�)D��k�Νq#h�s7�3g	�X�`3D����܏/QIT!Z~-� "4D�L� G�)&f�	�`(�

����
2D���Z�8�fm!��A7,�\4sWM#D�|0�K	�_��P�mKyD�A�l-D��hL�$�`���^\���,D�ܫ��ָ6²Q�v�R�/NL�D�7D�BAO�M?b�g��[� hY�*D�Ă���5u� ���"�+'@�D�(D�4�3AJ�����bc�%P��
S,#D���E���֔��gDB����m D��r�&H����x5
�o D����K���H;2��5�4�=D���+��Z����/d�61X"`6D��uk\:f�0�[!����G�3D��sbf�,����rhɤ3�0��.D��`�͠:����5��<WC� ���+D�l"#��f��V!��{�t5�f(D�����B�W@� @��݆=��	��L4D��:ܘ{�@)@aF��.o��G$�X�<����2&���c
}y΄S�b�{�<�D9%b@��u�V�V���k�P�<�d�݀_�� X�+�a�f�"DI@L�<�ۡ1��6&YG����G�<� �E�cF��=��
�'�/{�M�g"O6 s%Aly�t�W��xHd*�"Ob��R�	0[(L�.X4>c�5�t"O���닜n�as0�5`���0"O*]y��� @:�,FhۄUM~L��"OB@ �/OAZ��g�7�̱�"OL\If*F)p�����F+b ����"O�r��T�<7��h�A��ݹ�"Od�� F\�zLv�#4M���:�s"OB�-�E(�x�F��*?\4�T"OH��$}�B�J�x�KE"OȄQ�"�Z\5�ā�G�>��"O�%P&��B0�E�G��
Tz�a�"OHqieȜ�Yp����V�{N0��E"O��٠'��t1Z9�+ʽGU�"Op���oo�I����7��t"O��y'��3p�����F?�L��"O�u���!aB���朚�E��"OD��倕gt�e�-n�@��"O��u"�4/�ʡ�A�J�XT3�"O�Ū���2)��|�Ҡ�)y�p�c"O�QI3�_�!�Ԁ2���p���$"O�<ɲ���RpX��M	3W�!#V"O��U��$p���a��ح?��"O$������J J_&�Yc�"O����Eu��#�G( ��@��"O$8�d-��Z���`F�̂�y""O�tJ�):tH�lX"W� �@"O�m���6��SL��%����"Ō+勍mg���#�Y$B���"O����&Ҿ��S��$jq��"O�9�e�
�@cV�k�.�G[�]A5"Ob������|t�QjG� G�J`"OpeJtcV�Wy�l+�)�0i!�"O�����7�h�&B�`��"Ov�k�	8a8�5i���c=� "OPD�ǀ� (�3b�ԣPR��"O��q��.*L[��E(@��"Ot<ppmCg#��B5戡x*�k�"O**�AT�6��q�-
�T<s@"O&�!E��>�.q(��<9���C�"O�Ia���4|D��g��)j�d"Op�K���'*���&��o����"O�D��%ǧjpM抾42"OV,3��ٶh`Փ��	.vt���"O<S�Α'<j�0@�dR�Od���"O�������
&��jG�i��"O�!(�s�\dDQ_9V�;�"O�œ�N"iZ�a GAP"10ձ""O @��(��Ua���p�����"Oʼ	fM��+�0Dq/G�uh}HR"O.�I�L���B��,%�Uۗ"O�����B�}u�_�XȈ "O0y	���_e]����~��� T"O�$���W+v���a	ѕ<���4"O��R�#� �����!��O�x�G"O��A���a�"U��嗠1��
�"O��XA��H`ABХ��*	
qz�"O!��ąNx:���D�<P�X(�"O.�XA�x����C�����"O��$ٜ^*�[-��d�V��"Oh�9�����E@�W��,�'"O��c_�m�*�ɲʟ/�N���"Of؁�=/���A�V;�y�"O� 줹�\:5�h����$p~9XF"O��Rl��r��4C��:n�~�r�"O|�(�ȕ�d�4���Y�g�ti"O�dЖ�N�TT�-��B�Tb�Ir"O�Q8�� 6Uv)#� Z/;��f"O��(7 Ĳ0Ҋ�(49�0��"O����+My΂8�B��41�Ib"O)��.�u��HX��Տ$��iw"OP�B�Fˢ=�6�K��	1�����"O�p�w ��,Sp��o�$�j8�0"ONꆉ��5�̜"����L��"Ox�����eX� $�\�o���[�<Q�B�j��+3�ʑR�Ge�<�&$����PA��Aoq�%
^�<��ir��41��D%t�eBa�Z�<!��?��x@�Q��t����U�<�Q*2X:�LIE�8�y��nm�<���ض;ȰyŢN�!{(�*TC�]�<	��2v�V��m�L?��
��p�<q"a��G�~`�Ċ�.&�J�b�H�F�<qӭZ
\��9��ϒ*73�2�a�f�<�!+�����,�$�YA�Z�<�smڱR1�$���Yp摩�A�<�4E�%@{�� 	Ъ`=���B��<Q��!,���&��)���Z�{�<1�J�<K�=��@�-B�rab�A�<)Č�.���'㒎3�pQ�i�}�<�R*E+_�h��5(N�&$}�OUw�<�h/P�-k�ށi����D�L�<��y��Py�B�?$4�1���K�<Y�E��@��$)��=,��T.�D�<y�*�U���(�U�0f��ƚk�<AA	�)��Y;B��9w�8�Ȱ��e�<�g�:y�p	�g�5S�,��c�<i�O)!])Ȳ"�)�|2�+�i�<	q.޼^���bV	�AIG��M�<� �Z�?�
qA���vKd��%d�<1&��q��p��ESW�pxD��[�<����'�:)�n[;O��ĞQ�<Y7F�.eA*]xcM��I���*���I�<Y���z,����"T)�I��]��y�N�f��T` M"D�	U�Չ�y�+�!2�
-�q�K�p�P��Wo�yBA��O㺔��ռc�nd+���y�a֜,��Ļ���3M���Z�k���y�l�pr4cc,�=��$[��y�%��y��k�
 /��
󣞯�y"�Ɩp ����
�v�D��`K��yR�;$�q�g#�>�2P�R��/�yB�� j,�]�g��
"���eb���y"��&�db�'U%~�����iK$�y$��`����sBo�:��L��y�Z!~�81w��d���a����yr#ͼ��t{��p3�3�]��y���(x��j��8��M��B�y���<)Y�o��x3w�Q'�yB�M8#��Q�%�u�D��V���ybcȚ^�Y����k#&(5�y���of�4�)G�k�V�G&�4�y���sb�U`ũ��`�����yb�)}M\5Ӳ��S��\������yB钣?$��0�S#ZD��$����yF`����0ƏO�Ψ��A��y2 H9h~����]�������)�y
� >���hِ�"&+�Hr0�"O�	zծ��U����2IQ�*����"O䵠D��9>ɔ��,(lP�"O�J��Z�*�"X�D��W"O$�(��l�2	�E�=>1(�ش"O�̹2���5|@�E!Y�x��0�"OX!�DO3P8a1��ǎo�Y��"O���F�Ϣ���B�˸MR�%�'Q���ٵH2�C��P:����'�ڕ��2|� 7ENc0Ջ�'QB,����s ���Ɔ��XD^T	�'�J���#�K����v��,QG6��'�\,���T�i6^؉wc�+Fy��
�',̲��79~t2w!��
�Ιi
�'�`9�g�ܛ�<��"�7WՖ)H	�'>z R&xDJ�!�Q��r�'�@@3�)�.R�V�C��JX�'\�	�	�̈́�� -͜�����'���Ϣ�tl` &�6��i��'# DH�,�<K�9x���!)讴��'�,E*�
�16�X���	�5��\ ��?a֧@��7�>��H]qh�+ae�������N�w�'��&""�)#��R�� |���$@�� �ՔA2iKW�Z�P>��葂R^���d
2��jT�P	`J*̀���Tң�l?�}+�%�'���ЀG"\0���4���I�R�a@Z?1��T�K���*�<2��(
y?Y���?�K>Q���5�������K8�P���&F���B�Q��E���M�0iD�$Oޣˈ�`���Ԧ��'�(�d�f���d�Ol�'>D���4Q�<��#78Ҥ90bԦ�dt��'_�BG9G�����a��U�ږ� G6��e��(�OI���D���to�:�^	f�x���`�u	��W \@{� �*���a܋���a���Z� !2�%�c0��`!$l���V� ;�7m��GB�v�He���I|��V�?���$�ݏ:�a*�}��?)�R�xB!�*N̘�z�Z+]R �
1Σ=ͧ"����k�X���o��s��bS�H�ȑBq#��77��h7�i��Z���A���?yFz���"'�]��ću��l��Ζ"C���P��Ɣ�Y.�	_�`]J�?��$��g:�P��ğ�|!�A��,�WK^��b�,>0��T�,�Xy[d�<-_��>�#���L����;^����(	�3����N�[��7-��1�Ɏ{��(�)�<�۴Tz9:���s�`ca��dX1�'cў�}�$ z�t0�)�3R}��Bi�B����[�4��\����'������E�0�%���QՎ�YL���h�ae�t�	ҟ��I��<�XwR�'U�/ȸ��<KWH�+d�a�e��b��ɚ"K��S�<�t�U+bC�e��)���J��17��=�p��;H���j3�KCuP)�CN���9&�ײ&v��ס�:��i�0��#1�,RD�~�8�@��6�ɨ�K�OP�l���HO�c��Aa��_�����	�~\a$�Ҙ�?��&�����h�D,ٱ%i4rF�8�mO�+�$mCT�'ڀ7M�O��m��M[,��	�Eڦ��	զ�#s���s閒]R�Qʰ��`D����Of����O��D�O�ݻ0nK[�����V-�0��Ab�8�1�cբ]�	1`BN��hQE
M�dWQ�T)e㛻Mtp���� x��P��~����]R�Ը�#�5?J@���.j�Z2Aj݃N�'*b����'��f���<��MP#'�^"`P��36�	Z?���?����d��$]M�)v�>�>pk�+���(OnEz�'��§#$A|$
��љk8i��U)|�`7�<	]�h0�i�R�'6�>#��n��f ��61T�<��\5{�nI����?�s@Q5�]�dl�.����;H< �Ѯ����s��h�7�H826ص��ڴHH�'&�lj�[�2�Cs�
���DD0	_	8�k�4|;�I~X@"��*5�) ��F�:'�\�A��O��o�2�M�����OȊtiEI�6#w*��gb]�%*j��{b�'��	V�'Ƅ�8����42�pR��4-��xz���f�.Ov-9��K:��@�)�/��7jיc��p�	k�IU�'��l� ��      Ĵ���	��Zd�i��,O���dC}"�ײK*<ac�ʄ��iZ�pW��lZ8 �m�7� ��N�I��3��J�J�"�\J���ٴ?ڛ�S�V��֝A�����������?	�E�CLE�q��'7���`O՗��C�<�]�{@2iyd�>!�f�=�9��� (v����uR4��ᱤ��D�p����#�D�U!��M&~��"�G�l.��	�h��R*M>�r�(�/w-^P�2�'�8��x��V-i >ErD�>)�W�P՚�s���)�|�`��ۇj�2�{�����4٫w!���ɹ@�����ʡ�� �럴_���"���;_F��u����U��c�J��J�4�6�T��*�O���vKS"E�H�둢��,��˟� @�L>�u'1�  ���$�?���aa�,C�l�Z�'X"m��,6w�кK<�p�A<w}�%�t;���re�ʓ�p-�cgB���"���GgN���iJl�:��-���"���@&́��$�: �+1��D����� J�=�. f�7��\2�	�f���y2!}�X1siVk�����y�y0q��25��2���M��K�O�}���=WD�I%�r��=Ԕ�m����	�-���c�-^j |u����<
�J�1%Z�q���(�"�J�4�>� �]�d	1&&�3#T}B�F�Rj�9�f��/bD���<�V��"
dT���S*s�i��'��|	� �Tƴ�8�E	]\�� �O���H\%|�J�OB�06��F��'��1k1��a�<p8p���<�n��I���k��$�&@��ȇ[`��A״E�bycaTA�dT��f�*[���/�7$\�'4XJY�EL�"�u�4!ީ�� 	�d���ļD4X �'�h�2t��!���ڡ�c�]t�ɠ�0!qn��c�B���(�6 �e��S���OP�c��F�_�1O6�U�g�z��=:,�+'aZ�^#��+b"O���C�  �PV�X$|y9�"O�T��`0w���E.B�n֨�"Or���.b30$�t���=^�wj,D���qAT�p�f�9dg��)
ת*D��Xb��4`�8�CJ�5�tE*�D%D��X�@�y?�P����69
��>D�H�W��K�:VH�*[��<Sk/D����� x�dc�n\�Sj�C6�,D��ڷ��u���/ܴ<�0�*tF*D��y��T�,�aB��[�3��¡!-D���6�   �  �  U  �  �+  �6  �>  �J  �T  ![  za  �g  n  ]t  �z  �  &�  g�  ��  �  7�  ~�  ¬  �  I�  ǿ  -�  ��  d�  $�  ��  }�  �  � & h � �  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p �<y���/m@*�y4��"m>2������&�!�-F�H�+�暶m:(��T��V��I}����	�q�P#��P����5.�Y�s"O��B�ڋI.�:�B��&�jE"OĄ�#k�L�Pb�6.��!"O����D��1:%�rFʔx��9"O��s$/Q�gn�{q��<gX�Yb�3O֢=Y��D�z�Lh�#��I�,!�f��r(!���$��c���+^���v�͟@,�'�a|���;�$Z�c��c��V���y�Cv�~]�IZY�
Ƣ��y��=C���@Ɔ	(D�4��P����y��"�Z�`�Df�2H�CKJ��y�,rGjqSIF�b��!����y����S;D�QţT<W/>�3�aB0�y��ϟ\`���o��G��HsQ�y��$*d��&�B���&E��y2!/j�܈2�-�Gc��e��?�y���y �;0FD0l#�e��.��y
� ��5퀀���z�LB�x�Nt�6"OԠ� �(/�꬙�jMH��j�"O�$ �	*Vv�j�JP�Z�>��&"O�L�%٫��[�N�C�����d����	�8=Ё}�&`�vϘ�S�!�Z3V�\E8�Ί�*���O��0y!��L�W|,��)�R��PꔏB5Bn!�$9��	s,8T�\��BnL�m�'��|��=��k�ʘm�� I���y2E��$ʡC�Wl6tQ��� �y2d�����P��Q�vU�t �$�y��@�qA�۳�ƨCS{��D��yn +}�z$ssD�N�m�q���y"J$�p��*�U��@:�"�y�.˶���F��+bƜ�y��'��1�u�Ӳ%'ܗ�y8�U��Bx���'�̨��.\�TL��*� KtK�yp�'��=�##�g�К傜�q���D;��(�o0�:Ar�I�� ���r>�Y�K[?ê{gk��#�履�F{��ɒ��~  c	�7�(4[#OP�0$!�.;�uy�O��w/` 7J�k!�D�>!~T�W&;a�Yr�[&G�'2����[�Dހ"��m����X��+�E�%!�4H`������	N��bEN�	�!��=$`�+��� 7�N���
n��ĀFl��҅]�#�Yb�B	�`ѐ���<�(Ol">y�
 �`��x#'��:w`F�2p!�m�	u���O���0TAC��;��K&	�L��AX����I1$��ys�%o����C���?94h�>1�'�T�ɉp���'i㸡�p	���s��
Y
2���"O�jU�ni��#4Ș�M� �"��!���\�Q��)�3�	 p� ����d��AJ��d��C�I#��5��]�`���t��4;�˓�0?9�#��,�z$��Z����KFy��iV�b>�͓'x�8�@$�c�t�J�JH>��{�O�s��nD��K��07�K��0=�R��0̜x�5D�@Lr&���y��u�h[ԯnv�Y�"���ē�hO�����6Gʠ!-60�����q!"O.�':�@!
���l�l�%�d+\O�"Cs#�@p�Ɋ�$�]�1O���n�"��
0i��D� �m!��I~Z<�5)�!Mt�q�%kھg�'�qO8�D$�I�o��BB�#m��P��+�/Z�B�I5j�0p��+\ք���K�O���p<i��������A��}�s��P�'��� [w(�N�b{�$�'�0��ո��Ž�M�K>�דx0)��
2�&��`Ǚ����ɻb�Q���C�'٘��f�ȿ!_Z|��`��^yB���x�]�!DN9!`�C5P��4n�����Q@n7�9�I�?M�}r���b� b�F�20X=���f�<)�ҿT����E�3y��wMCJ�d�$87�3�|�'i���@שL!����t�R��'+�Z�]�[��!	��q �c��d0<O�T�1Q)9�1�tÜ-;�J�9��1�S�Og�I�`��A�b
EV�h�N�F�TY��oJR-����w|p8PL��P��ĦO���p<� �;b8�؂��u�D�0w��s؟���]�4����1\���FM�9����S����N@��R!1 Ō.y�9�ȓ9o�iJ2�	(_e0��7g�/{��X��O~�J�I�qX�s�Q�<U�is�'��l��$�䁹m�28��h�^g�,��S�? ��9A�Ȱ
`��V�ıl� |��"O�y!bM�	L�`֮K��*�"OL ��nءN��D�J�p茑h�OȢ=E��F�fU�PoT<\idI���ϭ�yo�?z�m�B��!H��4����?�y�-լb�� [JU��-�&���yr��.o�j�iqD�,|�T�(����~�'V�z7��q��2L8O���
�'�T!�G�_��:�#�L0iv�S
�'{�G�S2�"�� ��!t`ny���D"�.5Z�J�,[�MD�p@��8p!��J�H�2!�݅zL,��*�v���ذ?1�C�
疵p�3I��9�̙T�<9�e�  V��Jܡ(��Q�<�S��*�
X1�̛�K����`h؟d�'� ��)�g�D%2"��	��	��'0髧
�E�&��v�R7 �����'t	�w!�<2V���·|�� ��'�IY��.� �ǐx�ԩ)�'�ў�}"b(�#/�
ȹ7���<X{���E�<y%@�p�6�P`��W�h�	���j�<�U�ۅS���t���)f���"\�<����dJ�ȟo����m�<�paY1'�D���(�W�-:��DQ�<)����#�*_�%���`�MO�<�gdۀg�Q%���dt��2v �M�<IfgP�u@� 0��OՀ��SG�<E���e�ڑ����US� r�Y�<A�η�td;�$�? �����j�<��nX�}�]ӗ�T!} �Qs��i�<��Eݻ<ʑ@"nݴD����,e�<�vo
� �w�
�]H�Y�1jv�<!���)'`d�K�$/��we�t�<qE�SNU�e��N��B��cUn�<�p䖞v������%2�R�q!Om�<)qǘ�Ivx�{�a]�S�ęA7��h�<yc���"|
�s���IC]�gHK�<a2E�0b���l#T��bFG�<1�>*8�Z1�G�9N�#�c�A�<	���Jܨ�k���{[� Ф�u�<�dN!:ݎ 	������[�NMn�<a5*�5~�8H��X %)D��P_�<i0M���p�-�>Zf����c�]�<y֣$Ho�h:���?W*��s� �o�<�s`�*����' �MB��s�Ka�<���V�o�ak*�枵�v�YC�<�%	��X1�1�A��հqI�y�<�B��HE���v�͏<f�1�5�Rt�<i0�֨K`�AdLńbnb���U�<�f�U	Dɪ	��$@�5vr�z�ϙu�<�q��!Ἴyv����E$m�M�<�'�N���Mv�2��5��H�<�b�U�\C�S˟#>L�5�f��A�<�S���oB���]j�P�@ C�<A��ތN�NX E� h��v�Z�<)gF1o���!d�@���P�%�U�<I�A�-���!ّ*y����Z�<dۋ5�$���'ʒXHr�Uq�<�@�]//��Q�݂5�& ��E�<��  �R)c	�vw��#3�J~�<i݌g�0|� 'Q�*x���A�|�<��ޑ�8�Rp Ʉu��K5%�x�<�Pf�rhҥyf�Vep���"s�<٧�ٽx��\"p���c�Ѡ�En�<� Јp���?a�ܻ�EA�R����"O�`F��9,O�Y�E)b�p5Rg"Odl;բ���wJ�e1�Г2"O� �s�˴D� �+��'V��PQ&"OliBg-F�%��5jP���Q7�?����?q��?����?!���?����?�da3*��	�B��]��Zr�$�?����?����?q���?���?����?�@X�&ʂ�u� 'ixV��3��6�?���?A���?���?I���?���?9C%ڦS���(H�! ��L�*�?���?���?���?���?����?QGaX'�$=�P�[�:i$h�#�7�?A��?���?Q��?���?i��?I��B7q�2ms$�^�#2�!�O��?����?����?Q��?1��?���?)�	�D�q+�>+��rR��?����?����?	��?1���?���?y#�ǿ6` �j#(�/����� �?���?!���?���?����?Q��?�/&}C���O� 7��Pz���?)���?���?���?���?)���?Y`J���W`R�A ��X�	�?����?���?����?Q���?	��?����(ېٱ��Zl�f��?9���?)��?9��?��?���?I�Ai
�����_¹��?����?9��?����?1��?���?�T�ҽ�b��g'�J����B��?���?���?����?Q�OK��'X"h��L)}ӄ�K�4S�g��4�Tʓ�?(O1��I��M�W���,�Re!�/��0K�킞cE���'.7�O��O�9Om��0+d��T	��쁒��7>��۴�?Ad���M+�O�|�NˆB�XAI?��%4�ޡH��E�X�Q�M3��͟��'y�>%�!G�9p�HaÇ/Z� <=�����M�.h���O�6=�(�b��]���C��.6k��z���즹 ܴ�y�[�b>9��ۦϓ0v�[��T~����B���͓ Yp���F�y[��)��4�����<����!�^'����WkO'gc�D�<N>�&�i�:��y���2e6>p�"�s'��P%(�:%��O���'�<6����̓���4BR`Pb����0{��U�I��/Z���PC���c>��{F�'B�`�%
Mp�!&#8(��a�Q�0�'���9O,0 �"����$D��L���ہ;Ol�l�Ԍ�*[�v�4���� ��B�j�P�➮���a9O��lZ�M��Jh0��4����/�h�1�@���!�46q�c6 M�`���u�;��|�)OҒ� (
u��#| q��\E����Й�X �4kE���<	��t����5Iw!ƻe"ް���3v���k0�&�m�*��]��?I��$<h>����@���a�%Y�y�
xA�2���/Ɇ̣��O��E���O�(�'�)	1��6�B� 	,Z�	��'2�IBy��|�Am���C@>O�U���Ro�����j�px�33O�%l~��|�T����sӄ��F:x]�kVj��)��БH�Y��%zSgu��扲2�6W�p�J(��ٟ��	�]�j��10N�����n�ƕ��mħs�!̓�?�.O��S�OE҈R��ۣ9'Τ�FMG�N=�i��y2,c�|�0��й�4��p��x��ٟ<�@x��@�V��࢟'K���M#�i��M�#Q�V<O��:�kY�t�a����'���p���w3,t��ꖔ<v�(�J+�5?�'����O2ŢC�ǆ~�5�)._��!9O~�O�lZ�X>@b���O풑�������yG�C�N�.���OF��'2,7��a���Om� ���g�D,p�dͥ?���!p�ީ'ˬ�������4�dq9��y��CJ>1� Q�J���	�(O�Y( hJ���?�?	���?Y���?�|�/O��lړK{<<	�!�0���[���0*�*ܺ�ӟ��ɩ�M#�Bo�>�׻i���Iv��+h���Į�B������jӮ��ۥv��6�+?9��Y81ђeѷ !��$E!Ny{O�)�00�։ݐ ��O��$�O���O�D�Op���|B�G���9V�KfMT�a��?^���Q��y�c�D�$-���|λԵ��틹Y�*8QCd�3Jb�g�i�7�W���1�O����
�i��'��6m�Lk�jR=��!re��b�=0i��<�W�Io�9A�Aĝ]�����۸W��·��*|�y%O��jC�7Ap��ֿ���!���|�<�šH��	�w �	h��I�zy�M^�~.|�꒤ �dIP��!~��Ex!f��W���̓35�2eCWk�M+E%��B� ���']"\��q Яd �9�׏O�?�X�s�DX,(���#��v��4Z�1qzlѲ��
��*��W�й� �gJ*^��y���oe�U���=BަI�"4_��c�iJR�'SD �����e{��H�N,���z�`��5�$�<�P��b?�d�_�
P�3�)�/T/�du�����O2�L�0r��i�S˟(�s��&�D�yp���Q%]�tk/9�D�<�3FDu�O��I.(5�V-����Rq��/��v�'��B�Q�H7��OX�d�O��I៌�$�>�
�a#`@�}���s��]�`�$]�'bI�j�R�'�i>����pH��)>i�t*�M�t'lQ���i���BUJm���$�O��柺�I�O.��O��X���)yD9c��/���I�'��[p��蟰�	~y�O��O�RE�w�DQ���}-*�7N���7-�O���O�v�B�������������i���-��L(�a�[���+vH�I��')���) �*����럪���O��� ��`��.&�%���I�Kt��3�i�d�#�:7��O&�d�OZ��_g���O��a��rP���<u��CW��qD�t���I���˟��_��_�g�A��Y�5{�8��-M��� �.k�����O����O�e�Or����	��c����� �$���7���X��?����?���?I�� �Rĳi�����N3J7LHcq�	 g�eӖ���O��$�O����<��3Z���{a&�:c��Y(W�{�R�ڰ$EN}���?���'(��'T���b�P��O�����M���k��	�4-�	���㦙�I��<�ICyr�'O������E� O�4�`K���	P,���n�ܟX�	ӟ���% �d�b�4�?!���?���(O\�����I��	CEU�`��u�B�i��V� �I�!���ڟ�����4B��5"��Mh`UA�&ġmHnZ�����%���#ܴ�?1��?Q�'�R��	�T	Q�A�|�J�@6�1tm�a��V����7h����ܟ������~j�aȞ\�4�5�#gM�=��¦�1��!�M;��?i�����'�?9���?���]�#�]2�D��x�����6$I�zg�'��-@��t����OFP��HO���'֏k:q��{Ӏ�D�O����WloZ�����|��ş֝���u ��ɼS!q���0�<b�PJ��*�	Ɵ����s'���v�Y�6�x�+��׾�M��b:K�i���'�R�'Y��'�~2���m�TQ���$5�BPI3G5����9�����<��ɟx�I՟\����MCs�X�8��bF��:H�94 H���':��'���~*.O����nư)R�o���.�3�CR��AP�=O�ʓ�?��?a��?����9��M�?\�mh%�gz��j`���L06M�O��d�OL�$�O���?TC��|�2��t*��{aB��_B�Y�����M���?���?���?���*t��v�'6b��Ԝ�@�ԑ5�xY��Y� �6�O���O`ʓ�?)��|����?�Ti�'!��z$a��H�4�7��<k7X����?����?Yp��U����'���'��$��W�vL��^�2������L/B6��O���?��F�|�N>��E+i��r=���f��W� �J��b�"���O��������I�����?U������L��b3P��8�N�j�/�����O�5���OTʓ���̧��S�+p�qr(��^*��%�?	I�6��ZL��o�̟d�IП����?���� �	vM�}�Q`E�J1�1�&�_�'6��R�40�� ��?�+O�0���OV����N���� �o�+3�hB�Ǧ�	��,�I!�^���4�?���?!��?���z�2Ȗ�"�}�C�	����l�O�'>��)"��?Y��:��w@�8v'��H�9A��Eғ�i����:O��$�O8�Ok��$j<Y9w'I[��	�������I����&�l���	Ey�C���5q���-ʹy���(;��
�F>��O`��/���Ob�$ܣF�$��+	%��(��!��L�����'t�	՟��Iԟԕ'u���7o>Ij�'��.�F�Ӡ l��򦯬>���?�M>����?i3I�<��loH�g�x��`9b��a_�Iϟx�I؟�'r��4�Iۛ���I�o�f$�rA)$Q���l�l$�h�I�\�A�f���O���� !���ʰ 	!c�Ig�i���'�I03E]AM|"���z��Ѻ9���pH?f� ���S�}A�'1"�'��<�'�'�ɧ��Q6�N8z���  B�PDn�q?��V�| 2A��M+�S?����?"�ORy@ɵj=F}1�o��q-�=(��iB�'�B��'�'�ɧ�O�B᪐i����h �Ҥ}����ߴLUV���i�"�'/��OVOT��WW�BI9�/؞O�<���A�K}J�o�8v�4��G�	h�'�?�%��=B��%���� N�z5 + �v�'�"�'�h��=��O������C��qU&yT����0ԧ}�t�O�E�O{������؟�В��+T�b�h�
Рx�(2rHڪ�MC�M<�#�x��'{��|Zc���	���$�R���A�#J�	�OYx���O�ʓ�?���?�+Ovrb�R�*D����*BJjh�"#r���&���Iğ�%���	ğ��� �,p�l��� �
���=���	Wy�'K��']剾!+�1O�<ق�M$3���F��;}k�aӫO&�D�O��O$�d�Otl�U(�OhAi����|{hE1ǋ4}_py����W}2�'0��'�	TfћN|:����.H(g��
r�hl��L �yE�f�'��'�r�'O6���'��k+�A��o�)vv~K��εHJ ��唊5��h�!�-:�nZ?�H��ɗ�\�C�+C٬� E�]�ZNC�	�U~n�"��>_n���D�5�2�x�'.f�D|�#%�>4^0͙P�ьYgZ���ƒ.~*Y㢆Ց�b=84%��phW�X	 ��Q��{�S4���`f�ZWح�۴PŠS���JN �4ۇ;���;��Ԛ}gԡ��BZ'�|�C�Mc���a��S\J�O)% \�u����a`���?I��?٧���5�E�> F,)t)
�K����+�h���	�B�N���H� 0�c>M����^x�;I~<��k��$,|�/!(������8��L9�ǂ*�쥰dOܧ]���-�y2�H-PuA����`��Z��ēLl���hy���Oq�B�'d���}��r��`o�@�f.R����(�`�JS�[�4zA�b&I��	�HO��OV˓MTݓE㒀N�����ŞU�D-
�c]4A�����?y���?1U��*���O�瓛C������a;<Lc�nå5����!8^��Xq�XЦ� r��Q�܏^�(X��I�O�3����
(Y��P 	���?i�ՁV	D,H�@O_şp�4��''��'i�O�E����e;Ԋͯi8���"O��2L�KI�i	J-�\��c�@��O0�MkF��q�i���'��a�Fפ)�<����oxe�v�'{2�ê= b�'��)ݸJ�|���Җ����6��hp��sfp�#�>��x��϶Z�&���o~��� �j$��C��'�����Z��p<���N�p��4%��	�T��*&D�0\2<��hV��N�	�D��s�S�O58�a0S�0&�,��Ͳ<�� 
�'��7M�<���`E!�:I	s�ӊ��d�<a���=S*���'A�V>Ap�d���(����m=��䀿(�b¦�џ���84)�0*�ź��S�DX>���ǆo���b�L	�+�a���.}�T	M��eh�N�(A�-��ct��|��\�;vj�j�b/�y��[C�D��	���'�b�'��P��&��1�� ���2v&�`Q�D�O���F)l��l9�h9
�����
q�axr�4ғ?+�)r`�FGU^P��n1�UZ��i	��'Qҫ�>T�j�r4�'	R�'��wB�uXwJ��������Y.��"VG�Lȹ��W*jz�D�e�9{C1� ��&�U"�y��ՎG@,c�(ӍZ��� �,CƄ�ا��:b���֍�-\�Qj��t�V�0���ϓ�)��L�1s�U��#C4R��MK����Dǆh������?���t�a�N_�X���d��{Gd	S�'7��g-�x<�!'�سN�����'�2 ғ������$�
8d�ذa� S�މ`$�)��U��3*���O����O��;�?1����T�ˆI*x(v��:'HD�>SN�sD�UA�Zc	x��5��b�(}m��Dy҃� ��\"�L�D�y��D;?����ЈM�D��b'I��P�J`B I�4��Fy2��@daJ��'y�bM�&���\OD�	���?��8�I:v���;�o)���C�Ф~X����.�DҴ^�\���<l���D�T	1Oo�ɟ(�'(֍Q��>�A
���ɜ6#1j�*�٥�.!���?�TN_��?�����퐭|�&y3�̗�+�.� B⍕~� Qt㚡��(���07�XDFA^p�Gy�!!.�r����9t�Qg!O\�f���d̢p�*rNڞn��(�V�/< "=�a������ɟd���<i�G�Y��(�ĥP9�'7����`�เ�nʢ��$�e��'8��"<���4���l& 8�a烾@0�<�f�< J���I_y��U��6��O*�ĸ|BR�@��?��/ׇ���3�@΁8��	��?y�3�`���R)J�X��(���7]>��O���6���6�(���	�4h�i�J�\��ݝPs8��aAYq���򉏹m䞴3���7?��p�!�
�Z]�n��I�M#A�iL��ɀ(�XX3c��������.iU1O��D!<Ojm!�C�S���@[3CJ�U���'�6#=1�PJ����,l�~U8g�&m�@(��?a��3��X�m�?���?���/l���~`��*慑�[d<	���ڍf��p��b~����YV�=�S-���a�8O�b�.աJS��y�烒��t�d��7똭�4�F�B��q���Jq�: 駦���y2�W0HS`�8ab��n�\l��d]�5K|7m�̦��ɬ�"��)�<��{=4�`���7S��y���sD�!�'���OA�V�e
5b�k�fES�'��J"������'F����F�9z�K�>:@"�(��Z�<�r���O�$�O��;�?!����dG�!T��+&��%CQI[: ,�`f(�0r�(�I(#�u��?�`�^i@Aҕ^Ed�P_O&�%я�� zd��VF'9�"M�g��&����#kAb1�=�R�^.�xD�*�R�D�c؟�dIQ7I�8hׁy��0�5D��ы��j~Ľ��+Y+��䀥�'扔�M�I>��F, ̛��'��-X3.�hI`Je��"��=E���'��p��'r>���`�	��G�����=U�H�J�I�6]�b��'��^�P�1�9����V
K2�(O>�7��~ښ^C69���R-W���/]�D�!�k��eYDDцJ`�"��E��@�'��X��P��!jӘ�č8jk ��ug_>Rͣ%��$e�ʓ�?���[T�d���ߞ������M�0���E{�O"�7�ػhL�񍜽a�Ј�ለA����<��j�=������4��	��f���]8:�D=���{����p(�f���D�O����M�O�b��g~B,J�I���"�9T�9Y#DF���D��"<�2Ch�L5��֧;�b�\a���Os�3��	��C��ua���! ��ju��i !�P�G����"µ=��(�b��V�ax��(��!��D�)NU�M��-�'t�l#ѰiW�'M�Ą�H���bb�'���'Y�w�t����Փd�@��ef�?~�8�b�h�� �舛`�����N�!�1�hA�Ċ���y�)�.��Q�Ǫݕ)�Ex��� �P�.��L��fB�)�0U���i��q�x���� 6����f��%E�!6�Z|@��Ma�I 4�R���|��6)����B�({x�% ��y�i��e'b��
E�	��M�Ѫ�&�y�'_�#=�'��8RX���$ܓMbb8��D_if�ȷ�ЗA.\-����?i���?9���2�D�O��
w0���b��4~���3�٤J�"�� >�`����4
�p�rcƀQ�9�V#�#h�Zi1E8u�Ѕ���8u�]J0K�2j�H3���򬅁��O��d�O~�D�<�����'�
��oM-w"0(7��#�2 ��'G^�"P�,>^�ڦkƢ���yR��>i.O��H��J�M�Iß��c�]�9�r�ۋ�hp��FP����������I�d�'{|85����-��Ě�^�<8�10@@54/l9��8,��}�����AoƄ
 +ʓ�u✫X�X ����	zȽQ�iV�Cep}+��E��Wǀ�v��7@:�l����]�Q�'�n�+��%��Np����\�%R�@��M�*}�D��bB5dR���?����I<wT�`�6hݻnf¤���Gr6��D{�O56-�(]"����z�����ݣ�`�ĳ<y�*߄q�6����?9,��죂k�Ob�"e�Ը�� ��02{�H�o�O����!o�S�E=1��0C�M��������ʧhX.!�GN��i�2��%��4ŧOV�I M�0zB���E+Ǿ�)�W*��v�͟X�,XU�P<(dD߷O��)g�>AȈ�� J>�"���H|L�2*M�U�歀2
_k�<��ݶe�����RL���scc��hO�]�'C@�Jo/���d���gڅ)�'��R!�9C0|8�L=6�60PEaŊ�y�JƉHC$�J��ّ'�lu��L��y��[#X%0�Rf 2VU�e�ԅ�y�hXyT͙���O �TS���y2N����0���9K~N�����ybʀ�9t*�!�l��4x�=`���y"�P�R�dˁF�,v0����_�y�K܃-�68X��K�vܐe[�,
>�yrU� _ �7��"n"h���G_��y2C�8D�բ��\S�]H�O4�y2M�	(��U��E�`m۠���y�,��0j�T�$�h�� �y�m]w'�PDf�>W��P�S��%�yA�.ˆXS1��;j�m�"ƚ�y"%�M�<����$�I9�-F�ybi�4�8�`f��E ��h0���y��@ ���`$��=G�d�
���y��ރ$2��8 �ѽG�Z���_��y2m�[�<4e
.>��x0����y�g˴=�`��_�8�\ة��[��yB��87�4��$$E�+o��P䊼�y���N~^e��ʕ ,�9R����yB��m��(!e�#�@!�',ء�yR�,Vp�R���P*�j�` ��y��B(_b���!��|��7���!�dO 6H�g&"�M"�φ�!�D	�+M��ӫȜ7Ѯ%@�dȉC!��i# �" ��Z���	>�!�;*��𰵩������
A�:�!�$f�$E��D��f�2�醻[�!�D_/�t(p�m�!��!��?A�!��[�+zՠ k�=�Ô7c!��=x�x$����i�!�+aS!�D��m1H�І��}���Q�̬A��'{ўb?ͪ��b�Bq��ʆ �� Aթ1�O
��d�Љj�ZL���®M�&�9Qn�\㞜*3�1<O�C�iX�L��E4������e	"��<�f�S�v�*��R�P:t�
�SP��1�i%�����Y�&�oo��hTLV
�򤋦K���Ӓ�A��քѿ>�U��I�צ�><�q	� 5:B��fl�*YW"O�@Z18;��h+`�ݒM�ά�Q�U� ���&��N��4�'��O���6aĹU��٠%�J@@D���X2�!��(�a���,@;����8�93���4X]�U�Oxi�G"�s�hMA�����A9��)� �!sc�}�P����6!4%+���<qg�0=lP�� ��v�4$)ҦM���A�08� �rf;{�ҽi���Y�U
��'%�d)%�Y%E^M3�D�$�D�R�i%�9��ON�'˲7�)}�̂(!��.ؖP=b`A�������2o�a}"��%^���W�V5P�	G'*i+�Ʈe.�O�wQvY�HI\����LZ;�����ȣG�-�
����TL<Gzb�I(<��� �d�6�H��E���D��m��I7(>���9!쑟}8"�40Ұ�@�SB�ۃK����O�Uy���4�L���Vi@H��0�i����Ί�b���&	u����'L��{r-E�I@Rm��L� *�͡ �i����2X��p?a�!R�6z�(��Y���!1Ý���"a�O��Ct��IB?�Gj�ۦ��ؐB*��e��4�*�k��S��}��C'{4*�V���SOD��C��;Wp1O��G�'�	�p��`�@<Oظq��P�{r���J����XC"���C�	�g/�`b�JD�5:Rˀ(d��z���M��\�է$����H�L�NY$����X��?�P��5�Z�B6� �I��i�7�]�.Lƭ*'�4*T���4SZ��hĚ2��Jg�R�Z��h�3�M�n�Ƭ$�����!	DA��I�9���;va���M3 �� �0�6Ϗv��0�"�b4���Íad&Bw�3+�Ҁh��>?y\�Db���=?�皟�S�:���� ��O��I� �vo����N8c��x�!]�#j�(Ra�t�'�&e(��C�'q �*O��2�O��^'�h�I�}�)'���\�R�ɞF��lQ�o�??���g�LW�
�����e��ۦ"�?�XDp���*��x��pWB��
�]�'��؈c��*w�]y������j�T>��<��`��ֹ�g���"b.�a`�#g4V��a��H�C%\�3Dg��=F��g}�X�jB�db��0`���7��om�D�"�Z�`fh	��K��0=������{Q�^��4̎�m>���T�ioJتB�j�.�'��1O��OU2%Y��HN^��m��i����)���S)k�T*�´f��z�*�bG�0���Q�R*M��N~��9�����<ڈ��\?U�LJz�\AT�-p�p�BA'�]U(�Պ��5��p�O��M��x�tQ� ;���+�	��w�ܥx�i��b���M�e�M7��ԝ?�ˈy���l��d(�`�~�(��d;�M#���L��{�']1%є�c�Z�K4�~R���l�����ƔZ-�� dѬJ
Z�ِ��[�jM�ъ��@�̄뉽Pu"����C�EM:l�B��	Q/�<�%��M{�P?��oA��]#��ܴ���r��8��ck^)K��ԇ�ɜl��3�U){�S�[�J���H<U��A�4%O�`(w�'���cH1�3}G��I׊&;N@���X/8����1�F�����cU�]� a�;NT�w+�>���P7���K�( ��8hu'�䟄r��٘��I�	5^��'5���iW��t��#�����qv�{4�Q���צZ��������L8��P	;�ٶ/�>}=zU�ɤ#���'	߻-{a{���L-�8��K�6E�$:0��n:Z��Ъ�s�d�+V]t�L�U%��l�H�uEB�e��B���Y���䅩]2�{���me
��G�]Be��+N���m�R�-/iz��!A�K:�ċP����yǍN�%�T-p1�P�i	��:`�[��HO:��B�ϲ*��ɔD`J��U����$^� R	XE�8H�̹��"ʓ+�.���,N�`�RZ�}�N��X��sƫ^�P2�0�A��M���2Nx�	�i��%C�%B��Y���5A��,Fq�&�2�
 !!'@�49�fL �a�b,��'hVPs��^!�����ɨ=
�"�n�p7��p�{�wh4���lFx�)�`P�c�L���G��b�L��IӬB27@�pb'뇑o-L\�N�t������}ie�J�4��kR)i�yd�)6�=b�K��DAX�	�"b���И`��&<D��D5�8�;��ĢA��Q�g��P���_5a�\Z�('x~L�- �-_�T��Հ�p���I(~ 
��IJ���F��.7sD��s)� {��Ɍ,D��0�OU
:�H0�-�¤{��
�'A��Q�ߠ#�vY�"K��x�F]@���[��8fc'�O&�� �Y;d\�``K�cz�BbC�L���F%�	��Aɰ�%,�	�S�'a��n K씪q葡eJB���"q�a}2�Ufb(L�lٜ����� T\h��o.V�y�p� Y �
�c�Ĩ9��! � ��E �1bT��	qVL��w*�D��`��D±q�@�+��qDz2��)b�X2��baؙ $��7k(�b�n��vM�D��f���+&ܚk ��AhֆNP�)���"����"��X�fl��	��"jqO���FfM
�� "d�>vW�P�'�֥"�Y!`��asm@:Dm���n\(V)�5B�l�2ߛ��X[��8c�.4�"I��o �yk���s���@� �z��vh(LO
��Vb܌o�,�zb��F�e:D��)���"�S�#(F�)t�P�GL���ԘY_q�
�oڇ��cѪ�0g.*���N%a�~��d��
Bt��4*H#i.�B�j��_��QmH�h �q�f�⦍Rv��6+�-���3���t�nT��iU�eղ rBE�+/ �e�R�{s��g��<u������/	��a�B�;s��c��1=���`+P( '�՟6��@��@�^"�r� u:L�)��֦I �cS� p�F��{���v)1�Ɂ?��ܚ��5���X���P?�7K���#��;��y��V�G������
96����5H�զ�Js��� �x�W��5;�^����"LG|y�ǝ�;�X���ՠI{8(�p�'�L�Q���w�^ͩ��5�ejǦضY�N�;��Ԟx�/A��M����K�S��#Ӽi��q
��|�hTz��"Q�Z�"��80�!4��T�*.����b�$J]�B�	Om�FE�yJL��C�/HD�S-PT�����<���L�W�=��̶%�paQ&�1+\ʭ�[�Q��/o� :��U�d�X����6��QHq�
�w�������i�\�C��R�0��	n���������1��(��A���"��>-Lb�(�ӡ	�q$]�C��"|S�2~��C���y$n���!�5u��	�W��5�|���<H27���|��Z=IA脒O-,��4�p Ǜ8�ԑ�N�?�ߓ!��^(�k��S�(>�a��فe	���*��R�.E���Bbǌ=l�c�O���41����0� �(�   ��C#a{"h�Q���q`�?)�r�ԋ�� �3I'O�@�A闻D�H6� s� �$��L;8��'Zw�6o�
���ð��3z�D���7��!7�6 �U��n�M@j�a� x�a2�KϨW�E���G30�G���"#�%R�M�	�M���L<z�h��Z q�$��t��.�l1�����f��3�I���8�e�SZ�U�t�\��*��Ą��\�F8��M'Δ8ĬC�LD���m���t���m����H�h�H�7��`��߬d&�� 'J�&q�5x��'|ji!��H� l0Iw��:x�4B@��fў�I���p�����K!�MG���ƴ�Vn6KN��S��d8�[�NGf��8�D�ÛEmte�Rf)�$h��J���C�ee4�ЂH�Ħ}�w��e�lc l���TcƷ>���SF�FBI%�$M"�Ube푝+Ě((rh	�+�]{�d^TaKZUy:�0C��^@d��&�J�t�r��7�Ѫ��@�m��}��F��aW:�qǈ	��EEx� ͏^�l	U䋛?��D	A��%����7w����� ��5�ڿi)�]3w��l��f"t�vy�#��.lwpH���
�~*���N�y���r�$<˪���Ȳ-�*��f朅-��P�ԅcV�-٦��<,��X�v�����"��/3"(�V+*u(�U���{<��*�4J�vD1'K�Z[���CnO�a�D�剠w4�;��̾RC4��F�Ϯh���@��Q�  ��Ak�)�I�Fd�ăw���2���:�쉷��n�	JF՝(��}e*$�
�{��<��D�}q���%I�OΐH�n��!�H��ܴyFn8�#�>����)s��r�O�9R��,�4LNc��lx��/�7-g\5*�_��l�Ö7R}�v�E���=�!�\Q?���v*	�e�~Y�'�^Yʴ��8)'�qXb��E��2�R�g���X�ȧ�P�o�C�6Q������6:�I�d�+x?�i���G��H�ӵlX2f{^�����,�� �|�
%i�/A7'y\�yR�W��tq�'X�MM�����B_�@Qd��m̈�j�a����\[�1���T"�FxRFڤ`O <�!Ƈ-����Ծ��O�<��8_�T��v,�;{��2!�;v���%2v��@��U%��r�kW�yؒ�#g�?�O~jV�U�LA�/�?JA�ݣg�$�
��ܡc�W�F`�X��}��?��U�bX���Fj_-3fL(�Ë5D��iu(Y �:�� �
$�f4PB!���R� �3�>%?5RF)rޝ �3ʀQ#�[�**\���.D�|��#�!7��h��Z�%�F�[V�>�5�xR�7|�2����O��)w�Ѥ[8 iю��6�2��u�'|�'�ܠ����}���p��,p��)�:����.a|Bo	�P�T��Iԇa�"5�MV�y�M�s:|0lW�Wdz-F_��y�G��#[`�&h�9�B�S5���y�H�:Z�VEZ�E3��$����&�yB��w:�u;���'�2�3a	D<�yr��"~dɵ(Ƒm	�1&!�y�ٱ|nxC%̑>b2d!��C���y�!
�dm
�����\l&�0@��4�yRn _��4jE�MY&�j�ҡ�y�dC�u�����f�-�zX��]��y��S%i0��Ӎ��
����y�NAk`H�d�?5F�E���y�V�Wt��Q�0�����/��y���<u����dB������K��y�E>1�,�H�d�6X�������yB�K1XE���(�H1 ��=�y�V�z���Z���>~�iu��6�y��υ8R�|�n�;vF�9ŮF��yr�"O�H����:�\�{���<�y�F�Z.�#���-eO0@5� �yb��9p�d�N\9�-���y
� ���˘(��Ӌ+]lj�Ic"O��K�oX��BUQ�L�Cd�Z�"O`1y@F%>�6���m�LY��d�<��B�8��a+�Ƽ�$	�^�<ELK�t[B���ѨW�V��QoZ�<�b�ףLNM�A�H#��,�5e�U�<9��3"��թ	 �b���&�\�<�%fȇ$�T���W�I|�l!��MX�<Y��E}�-� ��C=L91�ɞH�<��+G
V����#�/~�ІM�F�<9�ǅ�M�z��+�ș` �]g�<i�6Zb ����/��Y`n�`�<�l�U&ƨ��%7P�&[�<I�*��;&%+��V	9]$9KoZX�<�T�˂v"tZ��Or�B6��h�<Iv��7�9�Tϑ�&����\�<��������J�
��ǏVV�<�6	���hV����LA�䨋M�<���ԉt6�<��J3z*��u�H�<�"f�9w�
��פI,F�����F�<1D�G&�Х�B��9�^��э�}�<�g�ʣ|X���,H
?R�@�q��c�<Y��1vJ.aQFae�X�!�F�<Qš�\�`V
��yڌ����C�<���X��.!A����EB�<1��{�<k��
�H��%{�-v�<����/`h���у� ��$[���Z�<���	����7�W�r��X��[Y�<�f�SC�
( �O�v�0�R�Nq�<y!	�e�1�b��57\�Z�)�S�<�f�
L�0��&ʢ�BU�S/^t�<��� Ck��c� �!nOT	��,�l�<�!��]�UZ�)��@)��yCFQB�<�aN�<]�v��=��	Ɗ}�<�%�ü"$p` A�q��A|�<�@��8
�B'�>Ƃ��#�R�<i ��;]y�)	�
�<#&���L�Q�<!�Ȇ�s�N-aA*H�SL��B'��J�<9&�۾u�ڸ�v`�@�� ��
N�<�'j�kڂQ�s(�%�b��GoRO�<�K_&<2��@� �~��VK�q�<Ѱ�P�l���`6��;`��%�W��c�<�#�5/T���(T�/ٶ��`��i�<�':���fM�2�<5���z�<y�O�%%�R� q��L�����&s�<ٱH�yM
}rC����%e�ȓo�ni�����*���@�6K�`�ȓn� @u�<�"�pR�"�)���j���E8_�����J՛{�VU��O�y�V�Ŀn1��{�5Lr��ȓh��'^%��Q��k�dd^���P%�\($�ϭvz*�x&KΣJ���ȓ��Y���+�f�y���:r5��kR,=ck�/Hxqb�S[�0�ȓq8��Cđ0Ϭ�#�A�?u�(�� "��P���@m� K��>	��̈́ȓG���!��
>�R��ǹ)V)���Tx����:+FQ�R�C�%�4@��D��ƉQ�5�0UR���"M��?��p�w��M�l�b���e$���&pXT�Fm c\�r�Y+
���ȓU�~@�#��/,�QAE��s� d��EŞP����K#H0A���]����p�ƅ� �6,n��d�Z�U�X���S�? �����-7������7^�*3"O:�0��Ԥ�誶� �����"O��0$�)�l ��/��S�L��"O��ҕ$)E���M6P��-�W"O�`k#ΐ1KK�!�'B�6Gv\�P�"O��hd��xL���q�]c�h��"O����Wb�!�1ǔ4 ;�zS"O�$�S���	����Xn �V"OTՒF�̹DЄ������HM	�"O���s�^,b1cwJф7�t��g"O��3"���y�恻5�
\VRg"OP$3�̎��@p�͜q��}"O��A)�8��)l�v8��"O�,����� !�w��X���"O����
h׊�R���Ar�c"O:�е�<Cв0T'�2:���1"O,�I��=yS�L{���u&�r"O��	RG����uڼ+Fڌ��c64���ЎE��7�ǏG�Z ��&D��Q3F:t[`<1�?4��՛3C#D�6OHMfR�!5�\�nV:���Z�<���T)��J>�yk@ɖT�<A�-�v�Q��e�N�h@��VX�<遁�&L�0��c"N��He���\�<�eZ3
��{䢈3$Rج���	W?ы��,�B��4O�_��q�ɗ	k�B�	�_�n-x �V\dHD�ɂ�^�2C�	�N8����b�`�8�#���fC䉌'��e��o�}�
)CD�Q�x���y��RaK�)L��Q�Km�$��C�ZUV&�:|>9AgSņ�&��Xs�<a�
 qb���a��X��BqI��A�]�$�@G�\��P��:=��1)��(��99�K8'�|$�؄�I;T&����+�@:@a	�
B�	2QAP�p��9�.a4�H-w�B�I�D%��"�N%�DĒ����hB�<O�����)�m�2��B�r�`B�I�@Ί�
6H��>��J����B�	�� C�#4s�M�5�?`��C�ɺ(��0Pq��D���g����B�8>�Z&˂C��q[u���2*������ ���n̼����{:� �3D�4�7�\'	�>!�p`̈́/6h�B�.��ȟꀁ�U�o��Y�eظ)X���"O����?u�C*��,w��c"O�"��I��,ɣK���I&"O��xQ��66��K��[ ^�Hd"O�1H��_1/r�!�	��(�i"O�i3U#	'(&�u��I>sp9��"O����g9�R����#�"O�=Y�'v5�e ���=k��$"Oj�釡K�J"dト��f�Z�;V?Od�:��+��� ˦C�%3�H� j�6s�݅ȓ5�$��B��'��i��u��U��dK�#ЧU�r̻ ��y\Np�ȓ��M�%��+m=4|#r�S�0+ ��ȓ��y�3GP<����i^�R^`��8}��X����u!�y u�[�od~P��-�f�qA�P	X:�2����M��?hc��C�L�puBB'�@~����?9Q�p�b���"̃����ȓ"�=�7�^ܘ\ֆW� �Y�ȓ(�TDJq�H��x̹R�Żh���S�? ���S����l��+Q.a�~�S"O���tL�)���r *�+�����	l�O�|�b`�'1�r���Gh����'R`(0&���l���y-�IOЕ��'�r0�Q3cT��2d��?rzP��'eE�3j͢GZ��!�4�&5��'�B�sWC�	r�4@��6&�.Y�'ۨ���K�@�&�{�l]��4�X�OB�=E�	��/T��)�
�~���&�y�!�=S0�K�#��}OR�	6�yrcɦQA�#t��w�n��!H��yr ��Rtji�;uhv8�/�=�y�H�0��Q��	4g��a����y2�,6�8����^���C���y�, E6dD�Tf�=mWl�Z���2��'Xў�����s)�!M�H�r3�\�/��St��{�O^����N�S'��i��Q�
�'C$$��N�)���xT�ݫ:�b�����Q���*r��:^px�vf�4"�C�	�d�@@4l
�Z%�6Lɓ��C��<v/| �@Z�5o�}X����z��C䉯@V\4#��0f�.�qE@���C�	�=��Sie4�wM^(+�C�ə&TU�΋-�ܬ����"	�^C��=m6�0��t��P�'�*JC�{�ĐE�+[�]�c�>m��C�I�*qș����P���J�qe�C�ɐO0���ˎP9F�TKš̸C��,`>�� P� �*��ǫya��<)˓8[pMH@S�_����J���ȓK�L�#��-��i��E�3��X��2�Q�����(ԯ�-�DɅ�z��
�遟D��L�0�

_�$�ȓx]��0F
N�K�� y�L���M�ȓ(f�R�*_�Vm���ԹE
(�ȓ$�n*��),�r��`�!=b���ȓ=�x�d�8Ta��	%q�ȓrx&�p���x��xCUr�����{Ԫ�H��F� ث`�I�f�u�<��a�%�`�DƷ>����'Ɍb���=1���'G4Q�So�P]��1�Bb�<a�O��0sů\��X�p	�a�<Q�́+p�ڱ�0]�Z��@(�^�<)�
�o��MPʝWj�zn�F�<�B�:	��u����9�(TC�<i���� �,��4��a6���ևS�<@���E �1���f�%��q�<1V��IJ�p��$$j �hE�<��P�B�z]�u� s
E��L^~�<��@�=�h�`�бļ�&��N�<��Z�~�Pp�WG$��0p�b�_�<��`�
 �F�R��N�>ކ�Sv�_�<��L-[f�x͛t�z��`*LX�<��kI����S��6oA&]S��R�<�;^��Tb�d��6���A�\P�<9&`N,7��yBE��%R޵B���w�<����&s�:�ǌ��t���ckHr�<�1)P%Z24��#7�h�� �S�<y�@Le��j��P6��Bm�D�<1�璡&���H���3#v�I bZ}�<1�ϖ=�� 
��Y->V�����y�<Yi�j��)�KR&=Y模C@[a�<y֩W
m�Ը6F£v<m�3j�^�<!s�0����)��)�Z�Ad�Z^�<� P���
�c�"=K��kd���"O�͛vb]�ĝ8�aҘ4aL�	A"O \��B㨴��`�062�1"O�i�S�c��(SeRrI���+�D�<�����u�P�J����=/���� �x�<)�NH(\ �a�"c� ���p��w�<�4A�T��)ֈ�%)(���ƅZ�<1�G��#�L��k����`�[�<i o�" Ĩ=�p�"@� q�BY�<Ѷˎ��aTlM j~�c�IQM�<�f�.�hի$Ĝ�&7��A5��G�<٧ ]4R�p9�5N�GH,��"�n�<q�l8mZ�Q��
�0l���Wg�<�Sb�-+���	������IK�<�0�X�x��+�����'GL�<��gb'��S!S!s}d����K�<q���p���cR�O<�Xы��MD�<�t��1t�X��X$9��UU�< �5$Җ`:��^P�֍X�#N�<$M7���%J�F�V�BNH�<�#j�$)����	��H�@|��c[�<�d	�{k~�n�<Ǧ�Q�iS�<��D�Q���3�CA�
����L�<C�R Q7Bȓ��\\���H�<��4{SФ��f�;-o*-�w��F�<a��ތT�xRm�5S�!�uhXF�<���X_�8ؠ���$(:��F�<��>s�h�� 9P�vT]�<����%���U	^�@Ī���\�<��㙐g�h���� �>��m�Z�<	��B�a�D� ��bA`R�Y�<y"�_x� +�OL�$^.8@��U�<���EҴ�!�C'�քa�S�<��bK�~�̭B��y
�|[Ҧ�N�<A��@u�Q�!/Ɨ�,��ԢL�<�&��gu �5n�3�|�
��N�<Q�ӗ6I����ЊC�l���`I�<a�nFwC�d�&m#t�xuO�A�<�0	�6�p���N��HA��p'��C�<��+o�@�jB/b�n�H`,@g�<Q��^�o�>��ݬ(�IX`Me�<4於��tI��\*f��`���`�<�B�(dm��L��*R��ɷEKg�<�'eڎ�*�9s��-FIx��"Gz�<Y �A7C����N��x]�W��z�<�w�P��M����M�f�9'�o�<�#�x��x (?���C�l�<Ywl�$c��T��;EDЭ�C�_r�<�B�g�(���4:�,���Mp�<��K��V>ԩ��A��w�0$ـp�<its�N�"�dE�W9�!�7 C�<q���"r�]�&�hta�҈�T�<�C�M:���r@F�3-a*��P�<��Æ5r&i[u-&*p�1�4�KT�<ٲ+Y�(��t1����5)BnPL�<�P� <Q�1�Ʊ3���� J�<)i������d��L4;!�DA�4^��[�bR�$��ذ%"[6<S!�J3�M�ŏ��=}zm�U��-;!���7�6��桗�%d!# �ϐ]9!�Ĕ�,����)���d�)!�_�x�R�w&���,�� ��!�$g*P���֘\�a��띙cN!���< ��cFɓ�p���2����!�� �p��U�r@��h@�Z��p�"O:(�T#��@ �+��H���2�"O�XȒj�5Sl(��'̃c���"O�$��q0�{Gh��H�0�ұ"OF����f�J9�@9k�"O���"/~�UE�y�  �"O���*��x_F�C!�B&/䪨в"O���)�����g��?��mRq"O��ґb�<j��\8h��{C"O.���J�;-L"���l�AT�H"OP��bo9k,jŻ �L�&�J8Ic"O�u���1:t�m��%�'���a6"O�����?-���h��X�@.��"O�ɨ%�ƳI�0� ���8v��"�"O���Q)5������R�G�N�e"O岆&^h�hp�N×d�P1�"O��F��@#�{SطD%��1�"O<��HՀD���UV�Y��Kp"O�(cv'Δe��t:�� �c2֬��"O��{�◱h�:dsc��V$�I�"O��ha����͛W/À��A`"O&�)��קV]hࢦ�\T�!�e"O�5�G�^� l%�I֫H�� ��"Od����}�1��#��
�"O�jfF]1d�Ĩ�b�5@&u�"O¼���N�u= U��=?zh�f"OxzR�q. �q�@�1�a�"ODZ��*�y��ȕ5���a "O��N.$���A`G���r0J�"Ob("��;��8C���$RpP��"O��I�LD�D�����%�Q=8��"O P�2nC���Dc�$ƐwJ�Lʶ"OhȪ��X4��B��J�,@����"O�y���$T^��z�ك)>6�s"O$Xi����B��D�`n ����"O$!�ӏ�E�V�0��ڪ�x�6"Ohv�і"�ĵ����q��	�E"O:a��H� $݋�E��\�� �"O���!��P��b�#�Nٌ��%"O q���$Q��
�s�b�U"Oh�3g��_�j�	���I�.԰�"O�PõC����H:O{̌A&"O�)T�	x[���3OAB��%�D"O~ hD�Y��i1��Ɛ=�:D�v"O@|��G" �X,lIȁsG"O���	��F��U4y�z���"O��SN�>���1i�{���
�"O�i"ř��r�@�Q� yF@��"Oh�r���9XM9�Hǧ1r8(8�"OF��ʓ�`�(����f$5�'"O�Y"f��!s� ���h�fd����"OpH� Bi�՛F��x�X �"O`�4��iwVX�=ؚd""OFY��ߑ��)��, �����"O�#!��X=hu�UJŦ��ܻt"Oԝ �)��'x����ьU�����"ONi��� 2Yi,���'F�,�J(�"OH�[FF6~|4��&�$�
���"Oz\�^0tE4щb���v�4���"ODHB���,/L��=~��ES"OI)�G2}l�DKȼ~��:7"O��� <O��<ȃJ�bS�5��"O�����S	t[R��i�d�8�"OiH�k@?8�4��E�>JU"�"O� F	;$/�6V֡R��lY,�J""O�V�:j���
�Gx��q"O@`CT�N�(���ʒ�?R 0�x�"O&��#�h�4E��&��R�|C�"O�i��^�0�S�&�+2*Z���"O my�V �l��ň*�	H`"O�ݐ�

ά�ic�Y�t����"O|xK��
2JJ���"���ų�"O"��b)ȩ!2J�3��	�"O��W��lf���)���b0"Od��Q��X^F5���V-4�����"OhqH���S��pY��8��̉�"O:H��`ɭY`С�R�@:Q�����"O69�h@Ԩ�Dʽs�p��p"Ox�����Q޸��	�K��8�7"O���a* ~�:pF�0���s "O����'ZU�Fy����:��1��"O��;FM� rP��b@$��"OԈsmԆsɠi�W��-=�8�G"Oꤸ2�R�ST���"&��I�"O�1�^�-�J	�$ԂV��}1�"O�ٲj�9D�|���F�y�$) �"Otxj�/�t	&x�'�ڀ2����""O�x0����k(��ZCP�nԼD�w"O����J�|Q��b�*j�	�P"O� ��/��!���!ŅQ�&� �"O�J��CW��ay�/�@�@�p1"O����DrW�U��N��e���Q"ObP�k�!��1@��#��`�q"OJeрa-I�D�cY�R����D"O�8�*��ua��S" �2c��� �"O�82D��7�̪w�8�ԥr�"O2eY�'�!#
�H҈׋L��p"O���� g�]Z�hY2���a"O�1@wH�#)�<�8�m��!t�z�"O�MiW'��Rٛ�G2"X�|K"OV�k�h��z��EE��&�`���"O0�f�	,��@��x� �"O*����M�#^� T$Q�:.qk�"O�p"ɛ�8�AXGJ2e�6-I�"O�T�@�"C`�d)�$:h��"O�p�V�F��u�RBE"|�� "O���H�j���96�ыt��#�"O�)z����>��0x@�L�?�~TV"O�EqB��Yq��1����a,��"O|�����'G�������'���"O�� u�D�/w�r��Y8�x�q"O�pv�ǈ�p}:gUZ� 	S"O6�� 
��i�e#teA)I�\��"OL�C���0}�����6��r"O�-)F7D��X'.�%:�Zq"O�ti0N��8^e�r� �i
p�RV"O4�X�ӈ[j�� EC":P.��"O6(B��Oo�Dar�	=&�����"Ofmq��J+o�X��P#ޫ �\��"O\��$����	Yg *S�� w"OJY��� V<�׀�����"O�q�՜X�*4C��8,�^�5"O �r����,�$��-� <+��9�"O�@��'_�P��,U�"���a"O��`+	[,uƋ�4L�:�"O��KK+@cD�FK\�#��e"O@��	%��XP,>8�W"O��hv/���}v��5B,a�"O� �	1�(�
U9��n�[a�d"O���M��80��,�%�(�"O�X��EG�^I�G&��`"O�ܒ�[6$�����T�v����"ON�Z��҂vD�t�K�i�p�"O��01ǚ�/T��׏<"u�"O� ����Bm�� ."9�"O�Py�HΥqu��f��d"�$�"O $�/�g����)�%����s"Od1Y��P�u��#CѾ��"ON@���u���3F@����ju"O����+P\ZC��[�Bu�@"O�q{����M2��3dL x�"O�}��坏"��cǂh&d��"O�31D���R���N-!�8i�@"O��8�L�?^ �Q`�!�M����"O>�x�F��P\Qe�� &Nqa"O≀���Sv�D���VN��"O��bdDJ  ��m�7)BH��dA�"O6����QIL�� �ަ,xH��"O�P�ċ�H���i�oʾCs�!#""O�;A�՛V����NR=wv�"O�]��� �@��f'>
ޅ�!"O��{d�����2f�@� �|�"O8Ȑ 2KS8���Cߒ:�Ht"O��C&�U8`K��֫�/
i��"O�	c1��A���f��ԩ�"O���mԏ�"�`�
�k�B���"O���!���p]f,@V�*&�{�"O�)2 ��Ep�q���%
DP�f"O�)q�H�;hNNt�H�-qҥq"Oڡ��+�y>M��'�#6X2"OH�b�E��1�6D���$K�Q3�"O�ͫrʗw�����ʤkK	�"Op��v'� ��cDa�7
|�"Ob�Y�!Ր���Kc�ѱ| T�"O�����\&�|\;�����&%0""O�m��@�9X��Q�Z���Q"O����t�h�UFj�FH��"O���-�d�ν1��\=#����"O �J��8R^���W� 
	��4"O���FD�"� �9G��T��4"�"O�q��I�b�X�A�..�{"OT b@@��Y.d�q�gG�~�&A�"O��q��Q��AhS'�����!�E$D��B`'S�؁
f���]^\�0a�%D�Ի�s����E��	S-����%D�8�Cƙ_SΥ�e�*"�d�.$D�L���=U��lm�?Q�"I��Y�<'aĽa�R��d�4�:Q�aHS�<�3iL�/j�c�4P����A�	Q�<�fkU+R�Vihv�ߊO�(	[�k�F�<q6��%�Fy@R
V�C�N��Ǣ��<�C�$g�	�gN�y}Y��AC�<1������t2�E�%ff�2�z�<�QUV���"��aQ{�iv�<�Bh�`5�t"`Y (��8�t�n�<aƯǢI܈��+�2Ę �#JOB�<��#P��M8B��8�,�2B��y�ɛ�/����d�^��msrBC��y"�̣Fh^����W�P����P��y� ­Z�F}3pe%C�.��⥅��y��9z;��
_�g���Ҏ�7�y�C�:e]�I�IW�Jt\L�RIH��y
� 9��!�./ ɰa�/_@:Q�B"Ol���a�3d?ր� �?\Qx2�"ORP&@Ӗ�|���	'xE���5"O���C��hv�p�+qCT�0"O}:��Q�]�n!�/%����"ODԈ�g��,Ҥ�@b�U�6&\E��"O8}�!�M�`��hR��_h� P"O�4���nE�����KR%�a"O-��������E΀"O������*`�<�ф�)B~}*�"O����iӓd����'��V"�� �"O�!ky���pЃ�+��"O�p��	.q��y�����)�"OJh��<8%H�R�.�7<mZ�"O,dx��4������{ZIp�"OH\Z�/U�G�+����fhb"O�EsCזX�c�]�l�Y�"O���f����"���a���Rx{�"O�u��]f���Da������"O&��k��_��� 7��)q�"O�9%o��pU�G�;	�Ip�"O䨀�On��= q%�.��F"O$�-��V��*�T��hb "O���m
488�`�闝�����"O��k�!bvtܑ�\�2sj���y��ҨNnl���Y)>~�å'�y�H�jSX���'�$/d�%�5��y2
�g�>�� a��#���ꔧT��y"E�D�0�s��� �T�݁�yrH	�3����Z�`���3�yB�T0k�{�n�55EsD'F6�y�j�gfH1u���}5�أ��/�y��V�Vd��2�d_�$<��s�Q5�y���mb�������Q�$�RnS��ybϔ�R���M�4��=�@��y䖥~��P���%��j�,G!�y�E�"k{^�!���g���*�A��y�:Pɲ��c�˶�F��yB��.�`sJΈ%sDh�թ��yR�0s���@�\�?t5�����yb��?w�4x�J��J���Ϙ��y§w9^��E	��A�'A6�y�D?``�C�H�ZD��`�ď�yi�?.@��n�Q
~�+�)���yR	b�ҥ��M�@5嘼�y҅ ��Bȣ��I���0@���yR�\SW��!3W�H�m�w;�y�H�%���dm��A�����Ǝ��y2ɛA�����=�(��3�B:�y�f�#Њ�3M92��j�l�'�y2D�+���
�,�*�f��@
N�yRښ?0:a��Ǎ9H&�cm];�y�� �o�|Ţ !��Am�؉�G�<�yR	�����Y����8ubhAcÇ6�y�޷�ĥ1�͜�7`�#3B�y��S>�T����3��3���y���ŘC�q`�P�a�ȓ@�H1��(Z�O5q�����Sg<����ſ'Ǻ����y�0�ȓj��ģB����h5@�'Y���ȓH��L���9H���ck�&Wa>T��Q0���v�@4�1�ǈ[�E���ȓfb@��V��]O��u��>S���ȓ��W`�"}hH��F��l,��S�? d��C��j����V�@��a"O�4hwc�!?���H$W��I�"O�����:,ٴ���C!R��D"Ot����͵5 �W�0P�����*O
Л��]�hlZ%���T����'�DK�	��q8�g{�yi�'���E��#��$���7zЌpk�'<hQ�o�B�biy�æk2A���Z�I !	�T>J`� �3l�����{���ΝX�B��v�ٲ~�|�ȓi�e�$��:�L�R�ܤ��P��3��Ȑ/���%I�ȗ%he`�ȓ�:$��mȧIbN�P��,C��d��o�R� �ěR���x�F\�y4le��C3p��3G-��Y��$A+?�p]�ȓ8������UOXyRe[=>����ȓKٜɹ�J.���5l�7H��܄�u�i�7*��in�ѩ�lX��z���ּA�'acԸ	ug�'P4��ȓSʘ��w�=X����`�'lzԅȓi�X�Yv����dE�l�F��ȓK�D ��MջH�x ���8�"���m4�y!��Y(E�1�_�y߈݄���\��ŪY5������,���fF�q�4FN)�Xq�'Fخ>�N�ȓ+1ZTۇ#L��E��+�,Xk0��ȓ>z�u�'-Ήe؞�B�,It�-�ȓn>��ѕE�2Kΰ]��Y�X^Նȓ6;�x���%a_��"0�0E~Նȓ7p�7G$lu�vd̢^-z��W�L,P��1�D���߉(<�!��N��9�-�3K��1�5C�G6Їȓ,�Px�PD)�~�� �O�$�x���fH��2E�r�^�@3��"@Y�ȓ@�bi"�,�/�|}�����v%�ȓx��M0�fCT7칢�χ�`M�ȓ8*�4aט`*���eW<c>i�ȓ��u ާT��@fb�:Zh�Ň�eA������ r�6I��������ʓw�:�Y�o�.��y����C�I�
�Np06K�8C�q�#*4��C�-:�r�N�"��QIJ���C䉑�&�;S�]�P(�Y��[B|C�	�s���,ǡT���J�K� �XC�	=!j���EƁ1�P���S$+��B�I&D3���%LY ($�Ċ��CB�B�ɗW� tDi�=��D�D~bC�I�5B����+��{��O�XC�	?�6����^�0)��̩g�C�I	e���ؔ�7�{g��sR�C�G]r���L@)��
`�J�zH�C�I�&�D�GLjB�[	�C�	��"�)��Щ(��G��w�nC�	:h22ɹ�&U�`wZd2��H-FC�	)ኩp�`�+�:�C��Y#f.B�I�-Q���5@՞��25o�58��C䉭Ҩ��K�7�&1�R(ڂ�lC�	'B�z����=V�=a�]+y�dC�I�b��	��%T<!�*�'+Lx�B�	�v!�pc@f^�O.�T�Viث��B�I�0|T����?�`�3�e%nA�B�	J���J;|vVh/�%�nC�Z�|T�U#\�$�H�ص
c�jC�	�����`)���DP���=9C�)� B�`#��o|��ja��VR�T"O�@y�B��*ԁaN"g4~<�f"O���V�`��v7"����"O1��k��'��U�aW;��Zg"O6�񒄙�"�
�f/E�N1�c"OpQ8`8&.�3(G1���� "OT$���(團v!��Q:q��"O�����q����oJ/.H U�F"O�H[�+N�sTĥ��hG
X/ ��"O~q�q �&(��ɇG��.,�"""O�Ax@��,CN��'��l+�Q�W"O"-������m��F�0%��c�"Oք	��]4�����gS&e�V<�"O<`���'z���b�S�Y�4��"O����$��t���a��-�p�h�"ORh��E��M��	J�Ĉ�#�"�q�"OR����-P7|�WB�j� )��"O��q��G.�i��@�F����E"O��q��1:q���P��fuV���y�+Ȟ�CN�~ �iق�׍�y�ǐ,?ܵ�Mܨ_6tZ�����y"�<\?�D���1)��Pҗ"[	�y�A�˚�PG��k�F���*���y�Ǒ&b^�Z��0e}<Yk`�
��y"*�B$"��,`�T)C#���yn�[_J�p�fP�X�vȳ2�A+�y"CD�A�B$#v��XA0��BF�!�y҉��o|f����]��ibE�ՠ�y"H��T�R�!���]z�Q�̀$�y"O��Z�I�cT!XN���jǱ�y2J&~�p(C�Weʒ�����yb��]� �6�>-�2�V���y2�|��9d �D���c/�y���H� ��@��V�"�O���y2gN<�@X��?/f ����yr�E�cenpׁ̜	JE����1�y�ГF�zQ���Hk�lq����"�yri�93�ֹY�b�Qf�Cӌ���y�� +�� o��HP�(;֠��y���!h�Щ�D(��@U#M)�y�Ŋ6u��Aq	��d��k<�yȁ�}d�p3��~����$!��yR�\������MH�Pŉ��>�y�M� �^Țw�M8Q� �9�=�y2�&*>����\}%rm�����y�l�l3�DْG�v�T�+����?ٌ��S6 m"D���N�Х�A��X�ޅ��}��=IwKE�'w<Q��ڿq Ʉ�D�eL�	��5Kt�'3q>��L��)��+��$����J�+�,��c*�A�4�A�U� `��/�\�U�ȓ:<�5���)��1�ʖ:(2�m��"������I�Y�cI�sQ�y��P��yi҄��`�΁����؅ȓ��z�f]�2zHuHa@ն�D!����H:SJO�.��'�B��}�ȓ,u�3HF�g�n1!")�#>®ԅ�ON��KF-�2g�|Ѹ�ᑝ}�|��ȓpt�x9q-W����� ��b�ְ����(X#း-Ήȧh����pp�����^�n-�#�F=kI ݇ȓ��BS)X"x��}���0O5Z���A��`��8ҙ�u���6�����8@�JR~�L�kE�4ZQ��S�? EaCoŮˠ-�POV�a�͡�"O��Y'��\'�)�R��a�"O|�b���gM�$�2�"O�]b6����!*[���0��"O�x����8P����g�(q����"O*��VN߯�����J =�Б�"O����'��\:Z� ���^��A"OT�*R�J >hy�'�e"O�ek5���m��MJf��U�@�"�"O�9��f�@���ɦiH�W�\��!"O4�q�)V�L�����S!DZe "OZ@g#�� �\$ࢭ"O�5����1)<�0�;9�b��"Ol���Y7Kg�}�d&�%�^M1"OB�eA�%%T���9}���;�"O�8�'M9z� ɡ�"%�.��"O��bW
��BDT�5J){t�M�"O2AcQG�N��舄ȃ�C?,+P"OP=��pu%����[����"O,%kv��dD2i󒄌Q��� "O�٧d�'1�B�B �·{X�=R%"O:%υ](|��@�ҹWߠ�SS"O��!֤a���i�l�  �"O�9�"ίG����q��(�#�"O@p��G|��|)0-��L��A"Of�(�K^7v��	86�©h�"���"O.40�H�|�����N�<�b��"O��Cv
g#��s O�g���A"OF,r�v�CC�&߲P��ѭEN!���(
)�����k��j��@�!��C�q>�a���
`�h9%$�+@�!��ڃt���;�͓3HB|��bל�!�^'�a�R�ܩ ,��KbG�;�!�$���-��U�|���˪d!��c�}�5�?j�3�@�gv!�dG"Ŏ�q�\��D0
G.�(j!�$�,�JUE8sI��@�k�.Q0!��m�X��G	S�>���gs!��4� �*x��� "��9Z:!�đ�av ��i��$���3�H{!��34�5JW�E p쉶�#!�D	ކ-s3�7O��I��4AS!����<ıQ�Fwx��!�$��54D=�`'Kt:��ҋ�7!�$̲n%9S���Je����EZ�|�!�Һjނ§��5N�и�Ù�V�!�$��+4\�&�P�Qh��	�C���!�d)k'*|��ϝ ?�@�"��y��'�f#�,P�c�,���A?5P%��'Z@Zu�PE�㇇+�Ƥ�
�'��$��R�}W&xJQ��>xY��'iTD�.��Q��t;bl��l3�� 
�'�	Ri�.WR|0��g�и`�'0j�`U��6*���j҇F5e���
�'�Lp�R�]�20�0V��R
�'�
�T
P�zj���� �5�
�'ڢ%[�
�>ov�HpC�Ʌ+	�'�v+�	O�*��l�B
6c�X�	�')84�ՠ�K�p�ұ≀X�BP3�'@�|1ӌ��DT�j1j�/Fj����'}���'p���� �ͻR���'����՜9Z��2�)L$� J�'˺�xb��|���gX�h��'C��1F��Z�0I��.�R6	���� ����F�n�a�H�#�2y"O��I�#� �&�?T����s"O��ـ�,jL�Q`���p)�"O �� ���i���AB��#Uq���s"OH����ܵv��]QdW5M>ep2"OH��%P�n<չ��GP֩�w"O�L1�ܪt� �p���5(��5"O�Բ��B �����BG��0"O�4�D
6U��C���A/����"O���靸-�.5��jL�f�Ta0"O�"�n�{�\Aqρ�U��� "O�Y2�`�~�@ Un�7�b�"O�Z�#]�/�*�#cL�\����4"OlQ@�lĹ>� �J�b�=��Q�"O�j�'bp�����1fl�w"O���ϖ#<\}C�@T�CT�"O��TD�H�j��۬M4~)�"O�U��En��r/	�O�X 5"O���@
/6�$���O�<�xr"O���k�����޺pN��#�"O��#��!�4TP�-�$m�"OL��D�Ž}�I�s��S(�xP"O�A:�+R/�<t2A@�-��3G"O~x�p�J#Ap��ギD�fB+1"O,1�'W.l9��#2��.&Y
�Y�"O~��I���(����!SQ2�"O��i@@�3r��b�6l���"O��#g�,���pк2�\E��"O��)��ˊ�ʔ�T�Xg�,��"OV�h��ہzY�v�@����B"Oء��k�$S�zHH��1H�H�C@"O��x"J�2��b`��|��-��"O d�D 8)���y5�ض^��"O$DA�k�(Q�ƴ@�`Y�=�"O>�Bd�
� ��.�)�(�(P"O�qA��W��)�.S�5�܌�"O �qL��K�"��QD�[�P��"O�QM5>־��s�طCҀ �#"O���L�r#�LP�a�m�<�"O 㳫و.n�jR�'
����"Od5��W�uk���Sc�6E�2p��"O���e-:��0#"xޮ��"OJ����L*OV���W8h�V�*q"O�E����37*�y2�_n�N�x�"O"�y�ΐnf�-SF-ϲ���"OHX{��=b�����<;���;�"O�(����,s���IA�`�0HJa"O�����pG������Up2���"O>JS`[w4��r`��Ec�J�"O�m�G��~,��X�tUL���"O�-��'���j�lٴaG�d �"O��H�/Z� �b��׊V�
% �P�"O��p�e�)��a`�HE�e	B��c"Ov	�t�X(��Ҵ�
�+��x�"ODL���*@~ [W���Zߨ�9�"O�d��ֳ��a#�q:��b%"O
��qEޞy�ڡbc�R	 �9"B"O� ���>n3@أGi�����v"OT����Ϳb�h�Ċ�W�("""OԀ�C,N:!���Q�IF�{�&]2�"O"`@pM�}�v\�EIG-5����p"O��J�@D���b�gR(x��i@"O\���΄d&\�EB �t�%"O��鲆S�b�TlA��W�@��"O� p��q"�)��eJTȕ�^�����"O(�E�#u�ԍ*Ԭ@�3�@Z�"O�5ied���x�P��N�<�+�"O�c@@12��l��mU3H~��""Ouq�Κ�034@�%�ܚU��*R"O����+�&qXt���M�9�P$��"O����k�?�H�{fMN
l��	"O�� d�=���Jr��fj*��"Op�
ы-|�A ���c,�}Se"O�]���s�f�h����r!�"O��I&���J争:ai�?1O� ��"OF�Ya�Ӱ	��a`�ԇojHPY�"O��S,O�>'�x �K��W����a"O��B�BJ�kB�I�k�7I���"O�P�6e�9;�0y�	Y�-���"O�whU.�8ɖ�ҴC\V��"OdQ�ݑ�v��!�XN���s"O�)��6S���A
<��0Ҳ"O�x��d�0J��!&�j�����"OFT�f.�<����ғ<��Mx�"O�����,dP(d����:J`�a�"OFM�S�מr�t�&��;��Q"O��aRhɳo^����Z�_V(�$"O��hA�:]�Na�Ԁ$=@���"O�5j֚i8r���>m*���w"O�eӱ�3T�x�aV�"<�a2"O��CB+�ޡ(!jBqr���"O�D�u�ܮy�Ωx�K-2�Y`3"ONE��B^�?z����#n���P�"O��2boI	=���k$���:&"OԹ�dO:�| ��en��< �"O6$c���3��h �B� �,k&"OB�0��L\�wAI��Dx6"O�-������*0k���X�@4Z�"O�\�&�0\$@#_
c��H"O�l�Ã�;K�n�cDB�r��9�"O� H���f	yFc�4iv<B�"O\9Pbk��=HvP��'$\2�*g"O��kۛD;nph����Iĕ9"O��eܑb���J�,->}��"Ov� ̛�o��UҊ«]�\Hz�"OT-���m��:f�	/.�d��"Ob�v`�!+�Dy��:{0Ta1"O��q�C�n��3т�t��"OбsjS�g��l��K�g~�"�"O��I��]�+�T�����)tH A�%�'�!�J=����M�z
�����O s	!�Y�C�z�9��K>uv8SL�*8�!�$N�K�)1`䊔L��a�݄f�!�D�96��#�"��� �A%	��>�!�dJ�!�t0��ǘ??��(:��ηN�!�d3q>�ͳB�T?4�H�(K�b�!�dR�i�fpy�z�,d�GϮ�!����P#^1?���{���;l!�$8Md�	�B�W,{�)0�O�!��U8@����\mpAJ�j�!��&Ts̅�G�QE�,�&*G0#�!�� 0.��u�v�����ᶯ֛F!�d��=F.Xp,M���'�T�	l!�Ĝa2�X�r��<*|����ڟsY!�V��h���>Sy�Jr���QY!�d��R���HR���x�q���ƹ h!��sݰ� ��ڤd@�P�U�NR!�䎂iRJ8Qn"y�(�cS	I�W�!�� � �`D�}�$��늗?[���"Ob���*/iP�JGcM=	W�	ʑ"O,Д`��#>L�E��TB�E��"O�Q�3O'L<�]���)!�hrw"Oz�X��E�VU"㡜	S��X��"O�	�2�ʃ+�Z��� ��\i�"O��j�(��F�Y�gǯm�
���"O6�H��El8hm�EW�C��u��"OЈ@�i �i���� g�hЛ"O�頄�:�p%�E`�9"4@��"Oܼs��T7rM�u	���O��"O��)�m\��VՀfKZ3�,H;�"O�@��H-4��5�V��7)�mJ�"Ol�kVI�M� m*67	Z0"OD�I�j����`ƈ�82��$�"O�X�� �4pMj�H�<hc@"OX8Ke�T)!��hW�\b��r�"OP�P��U63�P�'%ӑGT�$�u"O��{��j`��ɲ���j��"Oxɡï@�������Ƣ:-��"O��K���J� =��K�$!h"O�y����9����#**{4P}�"O�[r�اe@���[�3B���f"O��!�:lJ�p��B��"O�hp���@��L�u�N�rǄ
�"O�Z	�&t�nE�����3"O���F.��=����B�,��"O|��aS?9V��a^"v( <J�"O�q�%-�k~�hȰ F�?a��"O�*2���񷯓3���"O��hd�}�DL����7 ���"OP�ɢ\)_���Q�"_?8�J=w"O2�S1� "��brJ��R�ZC"O@� �]�z(iT�Vs�t9"O��rddød�P�sCK����"OY�UIʣF`�M��b�;d�v�q"O:�Bs(��z�sB�ms�X��"O\�6��aҠ B�T0dÒtK�"O��R"&`H��3����<$�"O`Ū��!��Y�C�Y.�p(S!"O`�Q*�!V|�I�㞗	R��"O������KZa;'�:UY�4�T"O �#���3�Xm`c��bXfQyP"Od�Q�N�O���5G� qJJ�;�"O�Г��J�C,��@��e��[�"O��b��v���� C�{jAI"Ot�����xґ��OƗ}�f� �"O�͡�J�<J�!��U�~�aˑ"O����F��n` �EA�4����2"O��`�O�7l�����fh"(�"OΙ0��m��y�ʆ�@4b䑔"OL 0u� p���S)T��fY�"O0��Mb`� #֧����{�"OJ�����aO�ī ���D��v"O�8jf�6H�Х�J�y~��
�"O�|y��ض3X���.�"^r���"O�8�S�U6j��`"�<_V&�K�"Oc�˞uq��x��S�g;$5��"Oj�k&�!9�d��Cʖ>5�$s�"O��!Gʏ4�reZ��D�4�a�@"O��&�3S�LZP��(.�Rm�v"OPۇ
���
,J'+��Z��) �"O�4q��O�V��:������3"O�(��Ɨ�P��9P�ƍ�.8�0��"O� nԉP�R�HW��ՏGv��"Ol�c�٣D��ӡL8p���"O�#�dկ,��+,����	�"O
H�j��8<d�JB�)p�b5"O�!����-|^�h�DM�g�q��"Oh��+'N�X�Ӳ��L�5"Op)���Dkh5��CN#s�����"O��6�٧&��ɦB��0�.A p"O�Q��kѨ�����~0\��"O�(ز��T��h�]`@)�"O�ID��D�
��%IҬq]h C�"O ���)V9XE��zNF��"O�ș����V2�*�͉�v��"O�L��D��)�41�,�s�"O���ƒ�Y����Ǽ[�F��"O����h�>�^!{Qʭs���`A"O�s�+� Db���a���g�\{s"O�E�.5i�9R�N7}�"Op�P��	��y#f>Y�<5�s"Oԥ�4��&,}hQ
�/�*���"O�=�0�\�I���"iQ*mF.��E"O=����2�6�5J�0]��"O"� D�k�Z��aɖ�/��U��"O���J�UF��bS�ЬO��5"O���"μ2�sV�'y�:�ڇ"O�tA�k�F���լ��+���$"O&���jӷx����I����T"O�"G�ߩg���Z���چ"O�AB���p�+fS�FV9b�I�<)&k� 6��4fF�9z����Z[�<�aL� ��H��c4-5���A,�M�<a��&\�N%�0&c{ZL`P��M�<I�A
�[�4T"B)@�o�ؘ�G�<1����;���r�ញSÒI	"��y�<��'V��P�ȅ�Ԉ$n~%����u�<	�㊅NǢUB�J�Y�V��6̞}�<���SDR1Ѡ��Y�"���#�q�<��R���F�C,e�t��!�j�<Y4�&F~��v$��l*Y��)�b�<�B���|���i�k��]K�K"D��2�@ҥm�XU0� G#~r�!�u  D�8q���/��=I�j�B2�1��:D����߄.y��g+04�	)� ;D��:���A����jЫX}~�2��#D�����8H���7FOmh�Ӄ�!D�h�!b�+r�5#r�N(�e#0�=D���bE_�f�RT�)�0O���g:D��xbb��RY.Ȫ'�6,@�c�i<D�@�$�-
6����jN�'�As��-D�H��H3#����7��.Z����P>D��cR��'����� `���Q��0D��CR�X0�j�p���7�y��h-D�<I�`ݺ<XM:D.U�aR���Bb/D��g�O�P�P2�'p͌�r��+D�����.��)35�C7:(��#�)D�đ�/S�<�>�C3� Nd|� 	=D�ܻ���x�:�b'��^���%g0D�0�%l]&3�L����c`r�)e�!D�Ppt�!/��� �,@��݉��>D��A�E�G�e��$�<h���qQ.>D���V�
��!�d
�;c��͓@,1D��Rm	��\�����)�L9D�����J|�2VËL�XH9R$5D��k"���p�0�HHL'D�� � �d�S��4����of�ɠ"OFh��O7-��E)A �Vyx��"O� S&�9j9,�R�N8}j��"O�	���2/-�8Bc ؁4k���"O���R�W�`�:����+��1W"O4��.14ݤ<����+����`"OL����Jw�(��Xwm�x�T"Oν���+��pZ#!ҙhV��2""O�(I�)ћ{Ͷ�Qf��|�H��"O�m�!`� �؈c@�:�꽛D"O���Ò�A��q׎H2g�%+E"O�q��C��XYޙ�C�yw�%��"O�q�EN1'��3�W�aT��e"O��I�eڪ�h|yv�F����"O4,����"⨋�eY45��ب7"O�t�t�ߩG���v��?��cD"OpL��Ǔ/7�*�����@"O�8�T���X�ԁ��1.���"O��r�D�C�L�:�cZ�f�\1�A"O���ê%8��XcrA2�lEHt"O6��'�کS����Oݫ2:M�F"O2�@�J��^��m	�.��|K�"O
HP�N�R�����ѡv��,"O�+�JK�#�TM&" 'w,^��"OP� (����	���8s�j��"OT�J㈤\��1�0e�0��q�"O�4�PfG������C�{�Y�6"O�h��&lq��.ۭmrr��"OZ豖��F���y��E�Ra�q�"O�A2Gg���!� �hC�Q�"O d"K�[p2�Za��%�Ty�"O��K��ۜ`�@�U��	T�R"O����n P)�t2Sk��VZ0��3"OJ�;�nnaJCq	[�Q����"O�5�BN�5�D�˰���b�x�(�"O�u��Jm�����O�i��d!�"O�C�kH*'X�<Rb�� �µ��"O$US�0B� I�r�<���q�"O�)	���{���3���v�axC"OL5#�&\Z̱��=b��Q�"O:\c1�Zw�dx�,�����C"O�:�(Ϣ�(Y���`;0"O���1�T�Ai��q�KN�bQZ]9q"Oh�k �MbR�@�&�׊Jf��"O@�/K�
!;EF�"FE.��D"On�j��%I��p��./���"O�r�EG�X]�؈)*��ab"O�l{A��Z��t�6�
2�)�"Or|�bgC�Ɗ��EH^��m�"OLi��Ĥ����!��?rશ"O�m���N>E咅����l�Y�"Ot<��ʙ�9���*���KYN���"O� H���I��iT��79v8""O���f�j�|����c��"O�Hr���WŪͩ�֌'O�D��"O���RF9C=kG I2L;bL��"O�a0Ӏg�$`�t�(��)CD"Oj0��ᎈ4��q�2A�J��H�"O�Ų��B�UX2a�?s�d��"O�#&���;SR�"�bC:O� H 2"O���Ð�\�k��P.F����"O^-�턍��� t ����I�0"O|D�@P�?��k�%) �C"O���0)��q�\8`d�8=�(c$"O� \(i�UX����"ɪ �>���"O��R!��t��(!�	�h��}3"O~4A@��:�~�pQ��?�Z}��"O�#w�ϡ#Q�P�GJK�/O��i�"O.�Z�NF�k{�u��I��x1��"O��*�BNh(f!��I�d��:#"O�Tk��� ~���*A�T�`x&�rc"O�qR͘xR=�G�!di��sG"O� 	����`�dAqY��"O�l��"ӝa�2A�@�O� Y�u�"O@a���W b2�鄨C�ͳ�"O�� Q�/n���@HS�'(6I#6"Odus#⃫����f�&}� �U"O�9��Z�2�4S�[�M[B�b"O$�CC�ݬpT�4Y�N'-g\(`3"O&e�U���y�6��g�̴`b<9�"O��)��LV@��s�.^�|���"O$و�n�)js�����<���G"O��!��a�.�����	���8T"OH� S'���1�%��
� ��2"O��#%�d��%Sb�Ġ#Bx�"O쵳+H� z�	B��9z
����X��2&/K�	St��mǱ5��B��$D�L�Af0jdEʬ�8	IGC�훦��f�'0��3�
GJX��{�E�<t�i��,LO,���a�	3;�Ȍ��QZG��:cC4A�B�F�~���7o���r���Ig�OZ�	Ӹ����Ol��x2tњV��x�P�t`\�[!�ֿODp�'
�B*
d��5�0�>)���	/<�H���ۃI}�8$�ۘ%��$�-xi� �ق]z���m�>�<B�ɞ;e�0�UY0S��TH%�ө� B�I�J�K6-[-^�h9v�Q9B�{Z�<�qG;��zD��i�
B䉌��9y�n��[��OY+d/�C�	�Ki�A#c)T����I5�#V/У<y���񳣅�������&qSX��t�Z��5'ʃA���3�M�mFp���X�h��	4P.:�+`��R��t���)/�J�Z�	?�h���v �[��T3I�ij���<�Ȅ��	�<���m�B�-q4M�r�+/��B�	�P��@����[��T�ec�ԥO�eDzZw0��A�Z=J��8AvC�O����'����K�C�P�sPd�IPi�,O��=E��`���0 J�=�A%�՝�yb+ϕ)��P[+Q d�8�㎷�yr�W�(k�0+�替|ܜͺ�FL����hOq�^�Y�J$&M>�K���7g�xUh�"O�@)�8����«��k�ƌY#"OFA"r��8\�Jѹ��U�B�"Aju"O\�BOʷO�m�� ���a"O��ƍF���� �H	k�F�I�"O����ӸT0����K|��X!@"O�	��#��Dp"���1dYP"O��SHP�,��*��A�0q(Q""O~�(Dd��4ND� �v܀s���y��<�\$�W�	�c��QÏY��y�d����H���>�@�pc	��y��={n� C��3��8��KŠ�y2B�6"f��Ԯ@*1�~8jF��yr-)ֶ��$�"^��� ��yb��u�u��+E���&��y�aO�[d��4D+k�����/���y
� ��Q�3Pz�a`��x#�4�"O�-�U�ˈs�$H��N#��X�e"O��f��e�j�ZDk�$*��e��"O��d @V�� ������V"O��	�F;�u�@G�z�:H�"O�����?~*�S2M�2O�I�"ON0���V�C�M9�KT�TD��'o)�S��yb	��`�܁�6N��&	��bag��p=��}R�ӧ$��z@ܰu�1`J\��y���~!�J̀C
p!P�5�ybJőF�x|��C0���
Х�8�y��NJX!�U�|�1�"'I��y��\�18UK��+�<�2� ��y��_�/��0���L>q����ď��y��!E0XI�$M�hC��ɧ����yr��">&��"�"_kd���F��yR�Y%@<�Q5f��^H��b'E �y�J��ԅC��Z>�)Z$(��y爨61L�1�iT�M�vd+dE��y��R6u8�`��?C�$p3�dƴ�yktb!�5��}h1�a/�y�+&/U�[��9��(S�`H��y �
��q��G�&6�2� �^��yR���N�K$h49��8�o�y�%��*��1%��b��;�y�jD�Q��`�c��+~��FE��y2̛���ƙ*�bQfȒ��y��W#@�L��V)�%�Q�!ܙ�y2$Y�EԄ�Ei
5A�B�M��yR瓁?���e��C�~�c����y��OO�ȊCC[�pNQ� ^
�y���R$B%�Ĥ6����b��y�@�2mUL�3A&K7}(`���y��Z�l��2���t��H����?��'���@��ВC����q�I,;���j
�'TЈ�,]4��y!dH6{څ�	�'��Z�L0:D�J����1%����)��<q��k  ��w��9)0P	BGD	D�<QV�S� *�嫕��1*X�̑w��~�<�3��@���)�A�-@��Ԙb� t쓘p=�6�/#h ��%=.����Do�<yf ��bjDı�DP�|��!�k�<!�G��H��U_�	'l]��fO�<!@'��t ���+Y� �
�ӁNJ�<yթ�Y�b ZDkG������C�<�s>�������|�@�f�<��@�U+�H��D*��P�Kb�'h��B�OH
����X+=I6�Qp�ϊS�M2	�'�h�c#͊!di����b��\X�	��H��	�(DhFA�O��8Rl�,[4B�	�_@�V%v���D�	p䈐�#�a�fB�I�v�xi� gJ/-MP����%A���D;��5m�(Ёg��Yh^D���A� �C���)����X� P��ԙ�y��'���x7j��"��'E£�y���Tܴ��@�
9��Z����y"nޗ,��y`�&�v���ǩ�yB,�<v��4	B�ҾW��x��-�$�y��!-#"�PC/O�W�^h�孟�y�(��i�F��e,.%p�d�`DN��y��ۡVY$��6�ŷ%����X3�y�)K�d8�����T-#���d"�y�/�.{�4k����\�g��y�)^��
��J�����W+�y
� �	��KT�W�,��g&�J@��"O���U�Y5�ċQ�C�'�Ȓ"OD������LI����r�m�"O�(Yp�X�@��r�̄M�йC"O���	�]�n�	4�#5>�[!"O�iR#L��n~<��v,��ufz��"O���a�ͫG�$0x+J<@>���"OF;�n�6rK\ ru)�<t&�E !"Ox���ӑP���Ӧ�!$ƥB�"O�4�ЎTEjveQT�̀x�+P"O: ��fΤ]؆�ܡ
���ç"O�fh/F�`;v,�J��a
P"O�l� F��viH�S3�գ"��ݱ#"OE��)ݿZ����b���\�z]�"O�]R�� DP͐�� gw�p!R"Od$�+�({,�9iB�'fW�U�'"O*D�l�z��i��X3I�- �"O�p��j��9�f��S�L�&����"O�B�mX�t��SG�+U�H�"O��c���&K����,;���"O�A�`�ڢ=��ʇ�5�n���"O�I`��o0qp#�)m��(��"O�!��S	��m1l^��ȹQ�"O"�# �4E��i�Vk��4��"O�ipևkQ��`�JM=Jwbu+w"O�	(ejˑ]�����ǹ bF�p�"O4��ؔ,2XТ��%Xi�"O*��lJ�z�ʴj���,G���4"O���k�8WL@i�D͐#7�l*!"OJ�@�h�/;���t#�e4Ȱ�"O�I��$\�,��z�a=��]�v"O��3�@�h=��*�C�,D|��"O޸REbZ�[�4ق5�8H�p�!�"O�A�D��3�2�K��Y�uEt�BA"O00�'�˱nX܈"�=i_v@c�"O�52� �V�� z��>m�<���"O��R�ΉT���i�8�-x�"O@�	�	��d��W��Z*p��!"O |9�GL_i��)��B���3 "O�]��nř�#]�g�F�F/�O�<�AG�-'���B#_*`�@��ETK�<�����_渥�a�#(s�0hq�<� ��J����	@'c�$�I(p�<i�Å5[�p��f�%q]rP�g�Al�<�ٞa�����k�	�>8:&��}�<	�JR&*��!$IT�i7�Hy�<�l�_*<�Fϛ|�.8�Q�Jw�<Y���*Xo �K�$߽mt^�z�Άq�<�b
ԍ�:|�"B;4���A��Φ.�^�aH4+M>�;�(�\��0a��A�rO|����{�� y��=D��:��9d�����ި :n��&�!D�(�"�Yg��mJ��T�x��!*D�l���*7
5³�δ�p�1�#-D�6��=|[h�)�-W8�X�X5�|�<��U#Xf`9�Ӛ �⠨V+�p�<����d-^	3"睔yJuЀ-As�<�C��� ڵ�4���`Mn�<����#�T [;`�P�kCp�<a�I�'8q҄��L��L}k���p�<q�J�,]��Ԣ��@?V':��Ţs�<���E1�$� ��;'�zk�Of�<�soп"
D�qD\�
\�Z���g�<Qe��
�¬�V��*��Z�<��Mt0�c�6ib:�i��|�<� ���V���X#�q��2�"Od�1!�O�tQZ%O�>-�0!�"O��	3�P'N6��щ�5f�d�k "O�5�0.�H����i��N��A"O�%������N	9�(�m"(�qL�(y�������(��JW���@hi��@�����yRaY:*u�L���؆k��C��?�BI�m�a��N�;��hÓ;B펎P�N�a��w�xЅ�	>.�����8%~( CQ�1��p��
<�xy�CQ�3-
��'2��97d?{�>�x&GG�6�b�'�� �KH>65е�����M��'1t!��h�,S�Z���B�OZ(�،�D&�S��͘8�@\�6+XN��+�����x�ւ
~����+X,d��[uÐ�~�v�/�S��M%ː�'2,�2�MO67/>a�U`RNX�\���ۛ�(E����H����O�1t�I~��}�Ӫ��D��ЪW��ȋ�D�'��U����S�iO�	hh|�f�>{�Feq���$|�B�IHSHp;�F�:!�������K�������i��܉��T?��u�H=� 8U��IYP%hAi*����g����`�H��T�g�R�A����ڼ�O?7��;�U	�A�5ʺ��)�*v<�xB�/*�0�@+E�Nv�b��B&wp��X*vp����I�X (O�4;T �L�#/�>�����F\��>��)�'i�:b�̱A���.{�^B䉭<K܉y���% �52Z{�"=����^�O(^tc#�*��N�
i�^��
�'��2�ςCy�p�Xdn9A�4_U��Ex���i��l��
p~�:S�O?]� YK
�'�\|�W3�r�ХK�P]�DˮOz���'�Q��cX�5o��begǱO��@{�a��]�'�LŁ&�O�g������O+�իߓJ��,���>��#էo5��M�#S>N�qfM�'n`l���}Z��%N"@�	Z�e�"�qO��%Q�X���ۊ�陆}Ԇ�iT��63ryEÕQ�����O?7M�]�t��I
�j*�$�AD6��u�A&>��ʓ�v�F��O
kE`öBS�9��G�L� X��^��r�1�O
��!�js�p�w���6�c���>:(X�F��tǋL�'�0�k�O�`@�[��E��Hޔ���	p�'��U��Hߖ{���90͉ƦE�'�ʕ	 nD��E�g�����=ғ��G��`&e��B����(�L��آ�ēKS���)��@�����_��(�b0 ¸
�HH`��X�<�j�!�i'�EDy���i��;F��i�!�E�@NB���c���j��=�	�(�!��L<�!RzM4 ���al��E\t}��AY8�L�o�Dz@}�O��)��Di��R�w��i���V�`�ҏ�T�'Q�*�H�B�%P�R`� �  ]�1�則K�������G��[)�r1ڣ)���N �a� �.���Í�d?�S�dg���@�c���i�|)�F�
���8�����Y�(8�D�Ģ��(�<��-�.�$0�"A�m�p"O�-�2oT$JN�A�%�9��I�E� +�Ra℄�$�?)�K%Z���'y^�:B�˸~<�C%AMH����'���@�c�/h�ˡ�� ��x�G�V=� P�׹� q���v�1O2��hT��`���Ip�M�#�'V��P���Mx�Q�c@S�QCR���N�t;�@�2r������Su}�[�y���G��v��O�$3O<�hP%%���.�"f��C0 �`�I�#e��s@�!B�YB�?!���@�C����zR��+� �/5�!����l�Q��;�OZ�B�-�����}�r�����$���n�<��'uH��'�96Ǫ����`۞w���ad�$g5�AS�M�%q�8�*�'Y:�4��!
��O�<�"��Cw@�@!Q������� _Y8����ȟ�D�2;�n�`t����0�ΎN��{�Lq���'��k�B�8������t��ԍ �gc�����|&x� kV��b&�/"}	4�&n ����	_s����Z�x��i��Q�$4���C�ʢ�̷�����3T���aa$hx�����"@�h�ʥ��ph@�T�8��*��5�e��C�D�*E�ؓ4���*�� Ұ؇J;m�P�gc4T�]#�"O�1�Tw(%U���%x��!���bV�	wa�Vz02g�0��|�1�Fp��L '! Q)�I�$#n܀"6"O�Ab���,��9HW��ZA��.��&�F���kY r����䎚��Y",/��0�����0.�@|���r#��k����D����f���OޘM�Bӏ$~\:����f��hv�V�E�*�����@]s� Z�d�fyA��'��#O2K�<�8G�[{i$�M>)w-۔xa  ��aJ�}>�˔.�vݴM�צ�Z��'�<*��(��ᜓpĔYBnE}�ٻb�'<�mk'H̏����]v�l�bc4s�����ρ�h��] 놡-:�qSW���ц�݆w�`�w;�L�� �
�U��b��K
�'���%�z�܁*�k�6wK��iÏY�|���o�`�zuCǄ�2�\x�U�F��ƵBv��pD��s寧��0�݁}~F5��9[�4��%O��1�,��1�v�#"�Z��<�G����q&�߬)r29xRm����r���%e���GR"ޢ����h�'�n�1r/��q���QIC�A�Б�O�uC��N�[A.=I�y9�n�U<0]h�hT���³��&Y�����D1�\��¥<��D�E�I�p?�[�
��d�F�M���Ƨ�,}N��A�JQ�JYt��Da̿jwH��d�F��	*H���g�yE��]�n�2-i�'��`V��v	��C�ɷ�YH���k�$��ce̘
qX1T.�+:��9O���ԡF�}a"�-l�:쩓�~Fz�'��!���"S��%��+\�=k��s�n�@Y�'��,w��і/�&sG�Zֈ�6[B��JH�7���W ^#`�&U�@�|��h �L�z�-"&�I�]kF�[7�%JB4#�HV"7���'(��P�H�/Ca@���8��T��a��"T�\�<��29��<R�F\�B@�1 4��J*�O�48e"ӗ;����n���Ǌ� T),A�#۬+g6���|��`�2O�݊�Ə�m�攳:���h��n�@t�4���/T�Q
OJ$y�D�Gb�*��X�Q�Z"M�RDxpQ�֯�yr�Ѡ!�B�S�d�H|�RS�V�)"ҭ�|?��À_ �@T_�W2���HJo8�� 3��y�@����_�.��� �>mq(�Sv�H�mO`�Y��&*�TȻ�g��b����&��tD�Ҋ���O.�BB�̔�8��#C9��q��>a2	�(yr���YG6��b��!�bX��g�:%�牜:&i�7+̳1" (�K��5u���c�~��~R��'T�8�[ׇ�,<d9WA՘��E:5l8sqEQP"v\���\��MGn����%��Qh`杶*m�� Ã��kʤe��*Dl�v��DG�(k��A�:z��y"X�:�4 `d#EB���l|�F��4
� �'ц��s�f���� �N?i��Y�J4p�����;B �*�R�'�,���W�=  K�G �;��� d��q�7��#Sv�4b�*ǉ$�,(f�߄yLPj�ǈ�Q�h��1�ʃ�O� 8a���\ĩSf�,a�.t��S��RqGH���� m<P�Q��|���ԫ�(���̓	l �0�E�(�z���N	#`6X�@��	�\����V�H��([��9���r��m�-F��g��'^X'�Xuϋ�1B�� c�Yc� �Hy����/G�|YȈQ:�O�IS� O�c'&(���0�.$�	�Yt�5+N<Y������b}��i���>��k����+R+*��1�ʪ*�tˢi!��I�L�@�gѷ-��`#�J%���tLP��J�s���/"�`m�h�|�q0�O�0���ZB��x� %����G�'�:p�F�T����2��H=e���)Ot���Ŭ$����fG>	���H偁�,�R�Zڴڛ�b�Ќ2ZZ~0��/\;	����XeP=Yrk��*�ƽ�@�'���rf�^'�r�A���6Gu¼�wϬa��I�@����HCgL��6M]��Y�!�#7��AC^"�5ft��t2o������Ӡ���?1'M�p�L�����U��-�f�$E�9Y���);O&E`5/}�H�$��#��b��&��#�-�N�$�B��*U}��� ��2�����~������I�VzX��C�/���Gҡ|��	���J�.���<CH��Fߙ��	�ď�N��M��dU�k恱�m]L�6<�T�\T̓K�L$���ӚC�Z�JԘL:V��'iyR��
�Vl,�05gӮ��ͩ��$SM��J�&RVw8�Ja�C�I�i���ǍL�Hٵ�J��&��n�oSn��$hD�_h���䂣
�d�F�@�R��E���ݨyZ0� ��hqUi�?Iޙ��"	�r%��'�O�q೤�z]>$���
-�2H���
y਻�㜷 ը���ڕX'8��C�К`
���R���:�4phs�Z(=8�A&��)*g�4���3#P�d��ʂ&�<�"T ��*9?�W��+F�6���;>�h�9�*���oS�,��������|�!�� ?ĒE�ȅ=C� �z�H�P�D9�S'�B�KԩA,�j�yE�U�=a�H>it�#b�9�'`٥^X0p�w~B/��H��H���ʫi��I4�M�a��kJ�m���fH{�&q��#ic�}:TNT�Q)�!cō�z<h�Ʀ$E�V�(�B�rX� ���R>h��̒ ��>��8jز	�2��&��=�1��O�U���Ь�<����ܦ�xE*X2�$u��E��H�`bAؿ��uzRd@Z��%;@|��K��"(AB���X���k$gX�c����'Nf7�\";��-�'���>0|���=�p�R �3o$�Ai\�8��4(��'m"�11i<��pA�@(��*��~������Sʰ1��[�-ؒ�T3X�� 2��X�`]�AS��*�Z�=�6�m~�)ħgV�s@`Ρ|o*(z���'m,8Jf`[�p�RT���� �'�� d�9����0_�j]!q�0r��P���o�1��N�X5K�j��,Y��S�? �]ɢj�L��$���E����YBKZ�/�ZQ�Hm�Hp��j�� ��M��:O��FM7���9��)������Q/Ek��M�$5���`�X�x�!���_���#I��d��A�A72�V��%k�<��F�r�i�(�Y��=��)�5a��y!X�5�k�W-�h�B�J)u%�����)��1|O�,�'�A����6C�)����;����HA&X����@�R�
��C�)�DZE	���Cu
�
9����q�!?�Ї�*v80��JҎ�h a�J�'�|r���'E�F}�1�\�&��	&Vqh%:�®V�̜s���O�}.U�y�!��Vmؕ���%	�8���	 ��}�����*+TEG Q����~אL��a�#/1��� ɀ�M��/��&�e�U�I@(ܺ���{�hK�1��B����%�]�Jl!�$HR��`T	솁��K�M�dE�@��?��iWr�c�+��Rn�)4�#3�� ?��}�H��ѻ"9�а7`�%-I����7��AUS �Ж���:w�\J)�X% �o�:Q�Q!s�͹�⁊VT�ȶ؟�[R�tR�Mv���ґ�#3�����,6qҭ�"�#~����T��T��_�`�:��[�gYH�ΓL~��%��QM�yj�{�`9�*�)(tN�
�/�P/�%��8%*_3:�X�3�����Q-���/֣M��� s,Hn5��Ąiv���ȓk���"��R�#�j9:�� ��k?�I���O�(&7��V�K:N��"Oұ+��M(.��I:��ӰBTv��r"On)�p�Z������X�/�=b�"O<��v� 2[�4�c��+t!���"O,u�@�W�(��x��*&��$"O��+�Ξq'�E�&ېB����"O�͹p�� �4��D���t���"O����i�P�~�ґ�ԇI��|�"OB����X^=��#�M��2��"O�HJB�>]���Nèjo����"O��sE/T ~�`-Q�HHW���"O"�qQ,��%�V� ���YA �x1"O��EҀW�V��S�	'T1��`�"O��a#�����l+!���A"O#Q��\i8�"p�ʗBz5+�"OZ�P��RUَp`C�2��"O�ԸS���$)3!�Hd)#"O�,��nP�y�TF�(�МhU"O��J��G\�)�d��?�D�x�"O,XCck	4_��]�G催7f�DR"O�d��E� XObyrEE�=EЁ:3"O@��0	�OuD-���Y�f�� "O4s��%��`z�F��xށ�'"O���"�O��B� n�Ne��"O�d���F7�4@C n�C�D�2"O� �@&�2�r�� �Y��-P�"O��BOI�Z:�d ��̋M�
!"O�� E��*��YǬ��Q#n!�b"Od�`��v|~	�f�V-6)��"O8�)��8FC@䈤�$%�p��"O>Ɋae� >��!ʚ=!���"Ov��šJ�]������Ż��yE"OP(CF_Ht����J�*^���r"O
XA�#� oں��!J�jL�x"O�ᢩ	����o܆1?��ʁ"O���E�^	�Ջ����z�A"O�� (�(��婀��
$��q;�"O� 
P���r	���M	�@YRt"O�M3E[�+k\)�oD (�Q7"O�pR�dU�=�fh9T�$qc*���"OԑI&�_*���7�%Kd��"O,Q{��I�j��(a‮}p��"OvUɰA'�4A�G�ߔ��\�"O�!h$
�8l�^a��O��4Kʤ��"O8,Y"�fxS�OΕK�x4"Od�H1��m~�!����~:4�Qf"O�	T7� �CЪN��,4["O� ��9����Io���4H�qD���"OV�X6�ؑj̘T�c�@c"Ov�!��ŝpG��cc�)	[���1"O��@*ޏofr|X�]�]��4�"O����G�6d��B,Y��̘�"O���hׅ<��@J�?)�&(I1"O��9��Bb�8�@�ʅh����"O�\rC�^;$l-��ׂ�d���"O
\��J��x�!�
Td9�"Of�"$ �9�0��� 4$Ѐ"O�l���S<s���@�&�5+�ؓ"O������e a�Q}���3"O�q�R��:Z9.P��Ϊ-0����"O$�����K�(B3�i2�"OΤ�B��J>V�@�HK1W� �"O`��D�C�Pq"C�ђW�`$K�"Oȩ����T��	�y�.<�d"O������z��"��Y�$��|�"O�XhŤ�>s���⅕��*�xG"O��嫜�,���Ғ�������"O�yZ�b�@�e�!b JqvE�"ObYS�`���h��h
�s�XD2"O�<��H	!)��Ѐ�̞]��A��"O����s��@֥X�M$80"O^�D�0T:\Ѷ��F�nՁ�"O~�S�%U�>��Z$��%=����A"O3���
n���	D�������"O����(�������.Y���"O�m@&Iޮka�dc���7���"OR 
�)U�c�������T"O$��/�\,3D�ڞi��"Ol�Q�C�H�e��Pa+�X;�"O�PQ�k��偲�J"6���"O.��V!�q���ڑGa�"�rg"O a�!ET�h�1��ác�E9�"O��A���f/���A�J,>P�1"O���PE�VX��JG�
0�ܗ�y�/�)
`���փ�"pD��ք�yb���\�T ���%�@N���y",/_��FA#u��3F�y�b��=�����M e'z��e��y��#P�r�h|c6�{tF�Z"!�d�"]]��Y����]�����;!�$	�$~҈�����hr�ʓ�,!���P�7�K���yC�I)z!�d*C��򁏞���\���ʅ�!�䅦�Ɗֆx��I���~�!�Fa�����¼f��$j�o�-5�!��A�P��� �Q�61K��<�!�DL4�8IR�5�s�jV��!��#��b�%�1IVXz�#Zu!�DC=g�pMh�!]6O܎��Z��/D�xX �B�n����%��L�� ,D���A20�R�j��(�҄ 0�-D�X�r�܋�	z2/O;Q���0�M+D��9�eʈb�:d1��U��I"%@-D��KU�[G�R��#��=.�����)D��y���$��n&)���UY}��߼t�4�X�V��Ȣ?�h��@s�@�Э�x񥧚lX��2��O4[��1`���z��yWk\�T6d���$J��P��;�O@��	����+��~E
�YS�I4�J����M	|��)ԫJ���* ����,Ǡ9�Vc�.�]��C�ɪo*X�Bʇ-MSc��yJ����B��-�r4���67໗D:��<�nW�D��@p	�&}Ɛ��U	^q�<� ����FQ,.�D��hD!T&С�Ɥho��B	�H�T0
�"\����&1ړyf"�U`Z�b}�D���I��謆�	�Hi�t�a�(|m4< %&�1'Dp����Ԭ��b�Wi�032$�7��>��@Ňd�T�0� ��FI���z�h�����		��	�2��-*䕲�Q>�b��:J[ SZ�VK$IvB䉴N$����	�n��$���Y�$aC:���`�vE$�1��t�O����7y�xX�aI
 �|����eC�ɫ�8�jͺ ڵh�h������@���s �q���bѭΫ��J8pĉg�>�cmV?�h@���rB���Te�V����L��"�@a�§ʞl���bv.����s�/=]�$�&!��a��� �ν�����ҙ`�����&�9��UP��B��%��'R���2�͝!��"(PD��0���)���y�M��%��=a2"�	�����C�*$���4*�$ f��D]9A0Ad�\�*(���!�u���;�dR�F����r˒~x$Y��ݸF>])��),�����v��5B[RHR��6J�T�C��K�\{���ڡ/�$pb���w+�jd�R�{м(�C�vSv�Y��I�E�&e�� L��*P*G��q&�0�m�'|Ɛ��+�P���mM�h�� S/�o�(=���64��}��b>_�������cR��6?r�1۔@C&+u�F�<#~�A��'�H"H8"Е:n�;���� �"����"�>�`���lv�@�aBq�V�d���(󀛇(���Ĝ$�b�j&MO�3�)`��L�#UN b�d��w䏁sH@���'�H�#A�N /X�+�GR P�1j���8�r�95u>)Z0��0�\�K�'U �Ç�!B�Y�wȽ:Yڄ]0��ؕA��u�6�U(<1�*D`�H̯hՄ���GVfD��?c���	�]th����z�k��,oښāe���i��Y�*D
ף� 3:�2D	
�x2��	���+Ѧs;6$���5^$P2����q�x�f�7$|�ɫ��æT�6�S���0g�@+rg_�Y:�>)ׄ4�lI��i��A���!S�c���7x��)�F�=@�l�pFS�n�"Q��(�3i���'門
Q��'P��($!�:{؈�BCH*��u��Ii\@#�*��ygm�5"��Z��(�g&ķ��U㇆�Z(�x���	�zbF��5|nu�U�K^����R]��I+t��$2�${lB�	E��`���M��A{Ɔ�&i�:�Ō�)�
!�t:OLx���R	F^�D��	�0J��}6fE��#)�c?�S��`���ӊ˭1� ��g+�P8�p����+��L{��^.+L��o�H�N蹁B�0�n��m��QH�L�EW:xPSלX��dP��ʅϨO��+��վ+�v@���Rު	A#�>�F/ݧ"��ikr���~J����E�n��]�*�$c^�!\ic0���W5���X�$y4���"7!�~�/
8F�IBs��*�*h�@���8�l����ܧ2��e�rIä�B�cOv�oZ�3��&�n8Q��"߼sЅ�+QX�)��<�����a�n���j�EL�Y��	ƥ�!�`�D��Q��U��%IaX�m�m����.k�.@!���5I~��Smғ�P��'GP��J��H�*#�w�>Xi����_R�z�
�;�邐E��Qcdt�L�0g������O	ZHau�E�1��[*dV�Ճd@ėSn>Yzd�	�
C���@��"�;���]�6�B)-Hl�SLݜ�(+A�V+�^����D=���	�n�ڡy����1��٠�Q�Κ7unVl��I�p�K`,��B�|�C�ǁ�M�q�o�3�<5QDkF�Pq��L<y�H�v��hg�Aü+cM�`��΂<>�d`�BG�B��$�G�J��RF�r��5ғ�O��򕋄�x��_�.P�S��1L��p�n�?Au��т��}?w�P��@Pu�_1H��P�\S�'OT��!�y~� XEo��uBޡB$��>�!�e�)9zv�%L�n�>��3��!_h��S��8W�Δ��-���Oԙ�`��%�	 �lQ�g/J�5V�$F��1@@��@�D�r�:��)�d #$�i*�6���i��쌥
��9B��V(f����M��@��#U(h���ə,���Z���.-X�b˓�VN��2��-#���""Գ*�0x@���M�e�i2��He�K�ItYAfk��k�����8{�@Vpx��'.�O��[ӂI�0S�E���>���B*NZ�E�5vѠٴ7�T�
Ui�8j���� �9AciD�S��$�ÆK<f6��3��b1
 ��*+/��G�N9q��Q4���L���7/؎x�Ȩ�q�?#- �0�-���%�܀�Ѯ�&!�`%MV
�|�.͙��Sb"�W�1O~�y��78��T.ߡe��cR���2d;y����C.�Y`���̌(N>�����>�֠�eH�Gf�"bc�6�x�/�$@���TA�.%+�y�N�$�:D
ϓft="�oD�9o�� ��#W�,�v��D�PX�C&��$G8bUJ�ezz���?QRd #W� �(�����"��M�p�@�4��gݠE 	�'*�eρ�T"2�1��J�cay�f�W����PN��
�'m�PA�W$"�iud-nQ!bF��S�
�"E��oXڡP��K�zh��E���O�mI碕�B4a�Q��r- u��'L.��U�\��B�>7��H�d�I�@%��͎�
'J�C��"G8��n�_��0&�$���9r b�0G-��� �c'.?�QڡB'&=�'�c҂�K���1rD� s���i�N}a�f�s^�`��V���Ђ	��Pc<qI��C؎�HE9,O���eK�yZB(�mIu�~(��^(X�.M�w�E�-ވ�0��V2����+�D}b�f�l5 ���*]�����7g�2�����7��a�b0��?��fB%:GIz�e�>P�����ϟ�:4`҃d�1^4�~�����"� ��b��B��`�/��	&�y
� N��Χx��I����H�qR7�'���yƅ�"L�U
�IŨ<
X�OL=��� 惝;��I�� 妁�gc���b�S�Gñ5�!�� �;Pu�a,�}6�S<�& ��jx�H7��%����<Y�+&�Ή	�A !i	��V�rH��jҋ��<y�G�(M�pzp�ҁvH�1%��3rv�����$ (0) G$A�P��4��g2T�ICjH�b��)���&�|@F�E7���`fi_0>~�]z � e1\手d����'Z��T�cD?o�e���)�1�DVW������1����	&��0���-OZ-�E�X���t�q��O�1�բ^��-� I���<�h�HH��y�}j��هdZ�U⤛�L��|
%���=��M�QQ���`��d�T�Fm���[�F
=a�oL�M��]1dF@�E���C$�����X��l��Ek��J�>���ǆwL&�2�gU<2w����չ'������Z���Fρ4>Z���'��dL�9Q�ī��hBEǘ�K���S��K�E�l<�1�L�Vw���d��&�����G���0�T��$�L5�\x�O�����
�̦���iFA�ɑ�#ҞP�D��!�5���KƗK7\s�c��b8�H�QOr���O3W8�<P�"$�C��p9���� ڴ6���b��W.F�(K�
$@�K�I_�5����%Q  i(7`�*r>V4i�KN�!�%S���$O8$�"��yx�2��I�����!C�$��Z��W.",���T��>,�g�$�0>���@"G-x9!��U�Y�xBcۃg��е@2��R}%�x�M�)q����놺`��d�6��2��P�j��dU.-�����\�A}~��&���	�'���"��d��>�����R�ڢ�w�謋fo�:9h�!�!��/L��|	
\G�NQJt��d��ʌyb���f��ܴ����B%]���f��kH���z��I )<T��@���\��ȓuߠ��[�ND��aC��n�T�ȓV�l<r&O�.e�A�q��*uX*���F.�C ��2�LL�W�B�B&0�ȓ.<��a�Ig�Qy���#=�\��2��!򲇑8��1��5;�y�ȓ ��|�i�!U�:K��PU��m�ȓy��!9�f�<|+�]�cl�<I�,Y��JB!�0���f����艿Ob
���F��q �; :����S�8v~y�ȓ'BRx��ؚ4%�i��˛�"ȅȓ�}�'��J���#�RM{���ȓ3\d���Μ
K��I��k�@�4�ȓe��KcGC�1�^	���:p���
��x���] ܴ�$�/(=��'>ڑ�3@Y�Z� �*S?	����r� 
7K�K��YZ�	۸J�.x��bv�`&ӄM.52g$W�,�ć�dS4��6LHo*�P�ӿg,\��ȓw����F��`B5h�c��-��H��h��;�@�"��Q�U�*� ���g�|�� ��d��]آ�?����ȓ���I�
�}�4�P#W0�фȓ�,�ׂ�+?��Ӓɓ�k��Y���7䚞D0&$ �LZ�:�$"�"O�0a����$ْ�(_�<Q���"O���FT�xPΜj#&A;��и3"O�A�̑/=l��{���p"O�= E�Ձx�}���J-m�����"O���@LO7��7 �-
l���"O>��Q�xt�T�D�9A�mBe"O" x�E���`�ҹM6���"O����C�}K���B�	w�����"O=x2d�-"��ko�ƀ��"O����U7Z�"Ժ��t�^ À��
w@Iۅȃ.\���0��'��C�.2J%�uEB�i�*�y�{2�t~�O�2K!�e�O�*�q�'?^��CA�X��M�3�^%Y�TY�Õ�@<��ň�4<��Q����g}�
 �����kڀ�k�����,yj/޽���-�>!v�+x��A���Td2���j�� �ř�ꑰ#eڥA�OV XT��V��!��O�N!*"�C�h :mH���5:��Ѱ1\�@�I�ǮՑ��x���Ⱥ|����M�:K�0�"�T �d�:ݶ���dLC�~n:�ӿl�4�[bk͋l��+V��4y<�öo����N<E���π X���Όf��ݸga?��'�u���'���ظ��$��h��?=c���ds$`�ǃTN��n}�nQ̓�M�0%��ƹSO?�&>9��
I�$�F��O{Ԑ�F<ufR�(�'%��IϚr�ʥ���<E��`��X�t2/50>01���M[KۮC'����C~��� 
`��t"SLE�r�m�'du���O�2�V�O���)�=g68���T����q`�b,@�{v�SX≦V�Z���^�/�E��fi,�3��b"�!&�\@1F ��F�'�b>e�W�O���Ј>(��U��g!?�g�Q�|Q��'��E��'�7.`@�OYHoz�d����M��E )�-��x��)ʑ+��B�j��G~z1�VQ��R��d�D�'��O���M~2�I�"�l!AsJ�`@P���Þ�3!��"�V��~�B���c?����ᣂ+ؓ^��AɅj܊<`���u�[�*��9��T�T�	�m�.���We�OQر�!�7m��X�a�-P���]+s}o��:zP�E�1�a�$*�g���4�N>/��Y� � �P�ϓN����2��5��8)�:�Y��s�F@J��9UHd����e"O�Q!�o�e�thC�@�a���u"OB�Jb쎈f/������p�6�3s"O�ŀ���WގH��%޶@LH�E"O`lۗ"GV��rEޑuz��"O9��F�($T�( Í� �C"O���L��u�n����߁e��Ձa"O�xre�*h�����ӹ�� ""O�����0"詵O��=�=�e"O0U�NӋ��HU��5z���"OT\�"CIl,9� U�g(�=x�"O�ѣ�)�h��!���%�$	 "ON����{Ef0RF�Q�^FD �"O�8pG���̎lꆇD�j���B"O�@�뉳6������u���"O:���uT�c�K"H��̓"O�}�T"�	,�a� L�Rgn�"O\mXD �Z��Ӧ�O�3V��cG"OU����f�=��	6ߢ��"O����!T"Q�����9s�:�I"Ox!A�H�4 P��L���p�"O¡�1��<W�ʝ�S�f�~�#&"O�u����F�����y]j9aw"O�Г�j	t2B��֯�WGep�"O���f��k��8b�0U"��6"O�ȋ�AL#��LX�g̓3Z�e"O6͛�G�/�xeB,�pH�G"O(-1���z�H�CF
�X�j"O����ۉq0���oU*V�D�ca"O�5q���w���0�O��os��A"O4�����3�
8�OI."c�("O
�ɤM#L}�M7n�\�\�E"Or�c=A��)��K)*B�0P"OX,��F;s��9&�<F0��"O� YAI��=b����-N9d�� "O��c"/�Щ�*��`;�J"O��r�G�N���85)��y%��"O@ec�ĚF��0c(�	pP���"O\��w��U�M�d�A���;d,&D��pX�M�~5�0�˥}*X8�D%D�Ă���}�F�r%@�3_�p�a$D��ɑ̟�r�ܼ��5$�(��B'/D����暤)zr��UGK ��-D�p9d�D?C���4.��>	q@*D�8ʶ��l%�ȑ�.̒W�h��E(<D�|����I�)�$J�q�Z�z��9D�����7�@A�Do�"'4A0UO7D�6'�����(��Y�E*�no�<I�kD1�R�r�lҺ&�|90!TF�<�����y�(�	v��6h.�t��@�D�<� ���$�|�aCRl�5sd)�"OH�(�j�[�Ը�.�L`�h8�"O�q4�R�cW���-�;Nܵ��"OV��$��jt
�X/H��0"O�p���4%<�`@g9n �)��"O��Ĭs�T��b��v�H�
c"O4D�ׅ\74�	(�Fsu�5�G"O��a�� ��4y$EW _��|x�"OJ��,��t;����*˻1W�$Z "O�I�ë�|s�KL�BPfe��"O �(7��&Z|�@�b=�#%"O�H#�* r�
�jE4X�X�ٰ"O\� kŭ�8XBf�ӱ?]��;3"OpŸeg� 7̎�Xf�r>��r"O
`��-]�:�L��f��N� xK�"O���� �u�(0��E�X�R��"OR �'&�v;�Q8�NG�����"O�@s���T�Z4�͒s`��2"Oht;Tٝ|�V�u�O�[��h��"O��䯝3%j�Փ�bGM��5�"O�SgM6��� Q��)���+�"O�����W�}ZbAN\����yrʊ� (�a�2��:�1��-��y�#Ǯ*����!��w�q��§�yb�F"D]������6ip	�@�ۃ�y�B�8e�˖��p�S�ď>�y�m�i���X�&:|���(0�@�y��<MSV�
��?\LPvb��6D��B��tќ0�+	`Xxd�A�6D��1�i��z(�v!��3�p$�n6D����P��E3Df��\d�`S�5D��'��% '4dвOO�W�2��k5D���R$"76	�D"��%�\��4D��/�n�Rts
�.Y\���2D�H+�ND(�.	K�aヅXK�!��;��5;Qc�#I�|��ē�K!�$S�Tg&�B���(`����G�!�D��bP��M�v=R�����:La!��3�J�L:*1�0���H�N&!��[$(�����v�����}!�;}���AA�B������Fz!��:x��A��x��01� S�K^!�$Tm�
�+�ɶduDq4�T�HK!�$I!QF�4�4U�kx�#@��
L.!��^5T�R!�6mN�0v��<!�Ė,F؋)�j�4cj�c\!�$AB����f#��}ghq���ȁ`J!����aGE�Ya���3C��]h!��Y|��,��l�b��=Wg!�	�-y���!b�Sjܸ�`A�z�!�D �(<p�0���1>49�T`�#�!�d�&
�ɈCc'���Pϒk!�D�)H)�Ä�-wVAQ�׃	!�	�Ac�l�v`ȟ�t�`Շ�1!�>U
X� k�"RҌ\��X��!�ֆb�n!��L+�������!�D�X���c^�W:�S՗�!�䟐I�$�ȁb�)�t�w��X�!��ʚ1	��e�
x����!��Y�!�$	t�J�ҧ�i��
�o�6*(!��_4�B��VET�	Ӫ�hp`A�.!�$Z�1�굡g��=}j3�eP�#Q!�$O�(��
�����'*�!���P���(	}9�Ò|!�� ������	 2�o!�T(0"O�"�ZI=µ`�k٬��]��"O�ɻ4�Ԋ]�Ƭ#�l^M}V�k"OXI��<WvTL����^�0U"O�$P��խEX��:�Mpl���"Of�c�D�ӵ�+f���"O�)�ET�+�*��ТҪ	���u"O����\�>0f�@��7t�d��s"O<��2�5W� �s�MI��>t)�"O�4�@E��O͘��C퓡��ɛ�"OH�s��Ɖ`n�ܸ�&�VԲ��"OJ�Ђ��#8b坈�4�H&"O6�۶��.<X�{QDL/D�L��a"OhQ�1��[�z,�#�8�:lʗ"Oz$B�k�5WT��D"�t��(�4"O,�ӂ��,m���PdB�~&j1��"O\��.�0��Aa�6`u�4 D"O�ɨ`�	,�N�۶�V
a$�"OV9  fV�5��� J��DG�$h!"OL%#F�1.�l�p�I�5@�$"O���'-�8!�ͦ_����"O���WKI�S�*�8�,p"O0|2U鐝{�aY�n ���X��"O����#���̸J6N��C�"�3S"O��H6i��L�`"� y�r�C#"O�b%�
{��PrAX�m6.yX�"O�Y��,3=0� B�/,X/�\B"O�<9�	XW�T�qF�BS��m�s"O8<�c���B�ɔ�ڴa�� a"O��X�g�����o">O�!�"O�`�vE�R���?o�,��3�y�l�	X"D1�gDL�4?��8A���y�\�m��%�IH�����]<�y��J='�$��� >�i��Ź�y��@	}���ɒ
��8��#��yB�K%��3��<�v�
d-��yB��	L���DmM#m�����Ǆ�y2�^(`4�]�EM	J	>�����y��N�|܅i䆒4m�9 wo�8�yr@3�T� GAD�����A�yB �Lufi�0�ǐ�T=cqF�=�y2 �c��$Ra�E�x�*\H`���y��j�x���v,��i'#F�y� ��f�Q�J�o�Ѝ���Щ�yk0���čk��)R��Ԅ�y�I�\�"X���Z7c�8Q)fAI2�yr&R>a;����>O,���UoӴ�y�ņ0j�̬!��)AF�E�4�$�y�-(P�I!��=C��`R���y`�"D	��B9qz�К "�yA3*b�:h�	q��e�Ǘ��y�+NC���4�5f5&����1�y�Ε�%^�u͕*[_*a�Vc��yB�:&�^������u(��y!�^�r�P5O�%L�-bX��y2-G�oO��	�,B�ı���Z��yrf*u���se�J�b�B��.���y�n� ~'�����'W��Ȳ(�5�y����)��DS���"	���2�я�y�ךN6 5H�Ȉ6K��l���H,�y�`�P�Ba�È�n�9�B@��y�@!9}�����D�3.
�1B@���y��]�w��R�݋0�~�k�ƛ��y�IC1[A(Yz�N%�̘KDB�y
� Vi;�Lʿl-r1��ӡJn�r"O���V�&�$�1`��?4���s"O� i3(�:���Q,ݢ-�=j�"O��Ig�R+]�vlB�+�2��b"O4�ЫPx|r�Pu儩E9� U"O���̈́kh�QÒ�R��@�"O`y� ^ gB}�1A�X�21"O~z�J��?���ul^�[��(K�"OPt����Z��$X����("O�u D��9�p���ŞmB�3�"O�])��\�58�"�!��,�A"O�T�%��u�9cg���s�[�"OQ�LU�o�l��A�rBX���"O.�K���&���P�C R*���"Oʸ[f��d�z�gŅ�2��4��"O�����KQN鳇Ô(�^]s�"O����Qg-�9q�bE=����"O>�y�蝙3��-�PA	
�B�0g"O�Y��~`� ��4,���a"O�YzѨA3Ab,Ԋ0�/���J"Oq`#�6�LP�#TP�Hh�"O!�$%[�i��=�2(2?��"OLy��   ��   �  y  �    	'  11  t7  �=  D  HJ  �P  �V  ]  Sc  �i  �o  v  `|  ��  �  (�  i�  ��  �  `�  ��  Y�  ��  ��  ?�  ��  S�  <�  �  ��  �   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6�F{��'O��V���&�;�+0:��x	�'%��"J�[�]�R�K2r��"
�'Oe#W烹�R}aC��z��
�'��;��7�������L	�'�:<*b&K"4����M����9	�'نx!c̓>�D �,ݻ2zX�R�'��@ �F�9<�m�7I�"+�a�'ր����>��Y�
�%&���'��0��3L�r5��M/� HJ�'U����J08fx����I$p:<���'6�D�)n�N]	0��K'~8K�㊵�yŬJ�Da3gǋD|H����פ�y"*@-0NPI�-@�=�D@f���y2-ݘ;������H����u�O���ޗd���)�S0L!��҇���Y�� 9b����2?qEԁ#�]1Ѕ�'?/�tzV��J̓��=iWɋ'Z��(���Z�:H�p��P�'a��G�ԧ��/:9��ƌM.��s�B<tK&��ƓK��8�NG�&�����!x8��2.�L	�I�ǐ�+��F�A����ȓGs(��4��>Z��$��\�~�<	�����.&̕Q�/B��nͺ6��bC!�˦Yҡ�'��h�T��^�!�J�8q,M	Q��d���Z6�D-!!�d���6�K��2Ĵta D@"-!�$�jU��j�����c6L!�� ���h�#]�3�l�.x�2xP"O`����3Xwr� c˔�=�(�"OLx�W�D�B|�̭5S�8*1"O� ��Ɇ����v 
=>�{�"O0��5��9)����C-<�#�"Oڤ�[�Y�Ȕ�A!͖yq�q��i���W�+�P� t�H-�<5��˅6s�a{��d�@�t���Og~�rt�ď{!��2\|���H%9���CT
O�<��!�O�@�7�=��4k�� �d���"O�=���_+L�(�Pd�͸L��uip"OR�8�Q�c��-(�%�
#!��"���[���)	>Y��t���M/L��`jV@ h��$<�O4����Ǆ[�PmA����q�詚v�')1O-Kq���q�g ��LL�"O�Q�(P<l���dK�iذ��"OzY���)}G��
�%V�$���{s�'Z�d�<�Tl��X 2dX
I�>P[��t�<����
	��0���	R� �BF��ph<�Rg�f�mz)A��L��I>�y�I	F����pI�}ܤ5��V:�0>�K>Qq ʽJS& � �۹)ך5GeUh�<�M�4�T �,\�h�~D�a�UN�Z���O�Z\�@���<�dnN�(�ZX�'�*�f��:m��`3�l�&Mp�8���=<O�9�d��>�\9�V�;o<�|�O�8hEj�#q0�)p�Z�D�P��6aEkh<!C�W�#����U����b�a�\�<���)��ӬY�L��u��T�<�3�[�u(��xRB��Z�� G%Q���'��O0Mj7
��I9N%c�@���(8� "O�I(&,�'��1��L�6{�
����$�OL��DO�K��ra��zP�|��fΩ^�Q�E{*�8�#T �h'�=
T���O��)b�"O� zD��9IQȤJיL�G�':qO�(�ӫM�P�4�
pJL�D�^ ��"O�Q����R��D�?��R�"OD��'A8w��F�\,���Rf"O4��
�(j��u��I�w����f7Od��$W��qf#:l�z��� :!���."=���3"�8v�\0�ڎ2!�䋜&��ԋ��܏	�(*0 .1!���M!.�۲�I6nd�)�AB�|!��:ʉ�p�TH� �@���!�$Aq�, ga.900qw/�<�!�_�X�2��D^$wI.������~�!��F'���y��鄈B��ǐi�!�dͻr�Xw���3�|�(��X��!���P�j�r���%��5�����!��G7o���J���je�KJ?m�!�$U,�0,�Qc��F!���L	{�!�d��C��U�"v��ra�9h~!�d־h�h���T����Ko!�Ƶ�Px�WbA�ry�勇Ìt�!�䖺a����?c|�ژ4o!��P��x��&JX3�t��A��r!�d@�����R�1p14�&!Q�F!�Ւz�$r��X�|�;�
�1�!�S5�֐WMƓy��䋵�T�!�!�]$U�Z�j���2I�p�5�ɻI!��W�Z�0@��j	d���S�!�:{|Dd�Q�0�֜��ǔ>A�!�-d䨔�`�Ś� �#��a�!���?�}�v�U�l���ibdM1|�!�� :��k	,nE��j���B�&��"OZ�Qj&t)2�b��0=��a2"Ox��%�N�=dIs��	�|>D���"OԵ��Jȋ�L	3����Q�|��P"O|�Hfߡm$�3sg��/"XA"Or�Ш�	&_���ү�l���"O����L���2��:F��|QD"O�l3V+2���TaV5'�
��"O��$L�hb<D���Ûo˺ �"Op�:�E[�"�0 ��(TN}�7"O���Ю2o��b�	�~��u0�"O�h�Pa^�z��UJ��	3_��AS"O�-e���
����R��=x��#�y2 G�9��+V�mpv��7�yR!�\�8!��͉���V�`�j�'�������#GM\�uSe�'����.�	�>���B��hXpU��'g�d�5.O�V�,���`�	sf���	�'1T}S#�H\�Nsw+Q�<d���	�'�.�(�	�8r�Ll���T�J�JM	�'�\�YV..�ܰ����YRM��',�ā�Ȉ���:��?{vT�	�'-����H=6���L"dJH	�'�`�gF7J{���L�p���'����T�����񱫍�?SD
	�'�n��i�Oa�aZa�Z5�l͊�'��Ue���"�PlJ�.�j}Z�'�$]8�I"��1���)^`h
�'�xmt���	����������-D�$GK�,��*u�H�H^�[4 <D��Kä���ҍ�����P�A5D���lR�_�:|j�a��1�I�ï=D��jQ*Z%0��з��4^A.|�G#9D��B�% 0OΨ�JC윎]�R%s�I:D���!�(Y���G��;,��[�i8D�Ps���-V`(LԦ�&@�T�z��5D���p"��=�j}@'/X�R+P� �!)T�܁ԦߌG \$8#k���:싥"O���J͙n�E{���C�~�"O��ʀ��-�(H�6�F���	�"O�Ԡ� ߂qk�,K�j՞_���ӡ"OP	a`�ì;$*��&I��RDBk�"OƘ�T!E�s� }p&�/5��0R"O��Hcǔ@�����#���"O* ''F�m�ȥ	�M���	cg"O\�95�T~+�= fLH%<G� C"O�S kC{��fK6D�%Q"Or0�����Z2��
�l
&G+V��b"O Ɂ�mG�[/,,#�#0&��3�"O���'�B?�թ�B��Z�"O$���Vd��˔��&G�f��"O�d;��X�~����s��4W����"O���%��EYFd���� 8(�"O�\)u_�P�4Q���l4��r�"O�-��.ԓ;��}{���%�	X�"O�Q�'D
^1Qsc��V�S"Od�c$Rf��rd�',���T"OT����j�p�� A&����"O�@��?qj�=	!`��Z��9��"O,hP@��$E�Y��	!H��\v*O��W@ׂ[+�Ո��&@48���'�� �Mĸ[/���mU8 d��'>^Y��NdCZ�u��?}����'�x�1$Ŗ�����1d.j�.@���  A��䕃 _�Ȅ"�L����"O��P�n*@5E�ۉ$���ic"O���e�_ n��O�;}AL��v"Or` ��I�|�MV60$Ґ"O�:aG�\����U��
5�d��'p�I���IƟ@�	�����̟X�ɝu�5�!�G*L���dl�t�zm���l����h�	�������0�	ǟL�	�cҠ󡫚B�FXB��ԀaH�a����\���������џ���ƟH�	6"{�@���0&;^�P��څMخ ���|�	̟H���(�	����Iǟ(�I M�"���gK�8�X����ȗH�&�������şh�I��\����l�I՟��	���@3�D� [�PH�	�<����x�IҟT����(�Iş��֟��I0!x�b F�� ��ҠVM��	���	ß�����ޟ�I�8��"��̩����C�(�K$����4A�	۟��I���������	���	�h������Pd��moJ�1���*=����՟h��㟼����L�I���	���	�>�@����?3�&)����m/���ڟ��I�H�	П��	��p�Iǟ4�Igo ��ŷ#Z�\��v܌������	۟��	ٟ��I�����ʟ��	<y;0�wbʗLp�I�1f<��	ޟ�	Ɵ�	����IҟT������%�\��D�g%: X��R�p1���	ʟ���ޟ`���������Rش�?��u��W
#�j��d�^%�4�3^����My���O��m�:>�4��RR&�I�=z�h�%.?q��i���|��y��o��Ჰ�E"!{�x4��7�	���F���	�B��8B??��H�

-� .�ԅ����̞�b�����)؎��'��Y�xD���X(P�~�S�fE���� �,<9�4R���<i���ce���3"(��	��^�%Le�dAX�J,4oZ%�M�'��)�4i|8AW)|�t���'J����fW-"���#c�Ԣ�KK4<g�9A�'Z�����'�(�
���#)�2�1`�՝O�);�'���i�	��MC�	�@̓+xt#�l�������d�=#,%��R�>!�i�P7Mh�(�'z�mY�� %u+>������wZD�s�O|@�'�8M���85�)E:H®��7d�O�h��Z;GPL�Ɂ6a��)"�<I)O���s����!Ф'��i2N��q��T�to��z۴;MH�'@�66�i>�sЉ\�Q,l�"NТ(�$e��lk�D�4;����'挸��A����V�'��d96�f�$��GY>X�h�H�4�\X���+Ϛ|��O�P0T�M�����8�.�P�*ܦr���q1�K!B̅�`�
�Xq�Z
%�����#���I��A	���r�·$�6P�B��n�4dPP�^�7�@�����7��a�7�F�un!�u���LM�r�g��FVt��`�`��B�/j�i	��F�"�Ah����`\2`e��n�Hc*I(A&�-{��Pc�i���}zå�.�)[t��#�P�o�������L���D
]:
�薦ʺF�X]�1/��/��	������VM��Γ�?٥#��+a��Z%�^��h1 '���.\ Zh6��O����O��	�@�i>	#-[O�\���I?Lx�5sd��5�M���C���'8��y"�'<���o��<����zt��#�eӪ��O���Lˊ�$��S�T�	y�x� ��r.�,@���)a����4�?����?qg�	U �SܟH�������G��������_	�PH�$��[.�i�ݴ�?��e�vJ�'mr�'�ɧ5v�äsp�a���4��K��M���>8���?���?�������O��q��](x|�Ӥ����1
ϊR�P5%�0�IƟ��IO�	Ɵ$�a�B	z=ĕ�-�(���ء �y�b���	��,�	Yy�I�s���E�Q��8�\����D�vw�O��5���O��L��I�Gj6 ��#��2�A ��;\�듵?���?�*O��x"b�f�Ӛ�������G @�&4�J���4�?1�����?�T��C����%<b\����5g8��Y6%r�����O��kv(�������'*��$�"�\��4nH�Q��cňF, O8���O5��C�O���O��Oô]����v�h������@�3�4�?1�<��9�iŌ��?���=���_���q�VD !F)E�5���?�#�^���'E�L<��̙/U[�0���ޟ9-X`�Φ�� ����Ms���?���RÔx�O�|v����"�rd
��T�:�07����҇��O���O������˧��)XJ&�����S�0t�3k�:US2mlڟ���|J�fyʟ��'�d�P����l��N�*���O<���(������'��d	:E7�]��nXA�V�iF��*���'��R2X�8٨�v�,���ȼ�P�#��Xn��#���M���BX���K>���?�����ă%LvTYDD���ڬ�C�M�%-ҙ��G�Q�ڟ��	�l�'k��'�p,c�ęv�]����%+�L�����S� ��ߟ4��Oy�N[����S,�졠�ɚa6ڌ��9���?���?�)O����O$�Q��OZ��ɽt����r���Z^}��'�R�'���s[�\�I|br/��
x��J��G|�I�Ȏ&n���'�bR�0��ߟ H��U��O|���b
�0K� ���#&��@���l�>���O��_°���T�'�\c��uɢ��6�b�Q��.�aJ<q/O$�3o�O�����3� Xt����>p �f�O�|��|R!��p=�m0O��(�Tr��f�<Y6�Ծr���(�m�hn�0r$�(`�P�S�O�+�>�!&�$I�dТ6�P6cΌm�h�|F��2��&|� 5�$�!Z���7؁M��̰�iY ?�����NW�Mx��e��e�0!�7v��I�݋Y��l�gj^�-�5�܋�6�y�jܜ(�Ѝ�acIu�8Q���\�fZň����?)���?i��&���tY��2��d34f̵�������`��!0@yS�Ǭ�p<�����K_�1�v%	`�]��`�Q?a�k��i�y0jƽ1��xr��XGp�q�<R�<�R!��u$�G:��'m���D�O�����;����x�yg,ɖh�@h�ȓ+���k A4!��W�T:4E��@�IQ��Q����Ȓ�M�%3%�b|Pʒ:�����	�?���?A�ct,����?�O�N:u@̀<��RĢ2�BL���ޮ��񹷡J��0>ѕ(��P�b��u���K�Y>f\P�)]'Ap$�I�`0�O<���'s.6m�ID��d,#��a���\���%�������?�O[P��+<).�{w� *`44��'NXpR���--f�w�5n�YK�'���^Px(n˟T�I]�t��O������<�0�1�Q�W[�D�$�'�B�'��i��B�]���vUf}*����� %s_شJ7��K����	5�2l�Y����`b�'Z����%-���(f�8D3�aDy"���?����?!���i�%89uY�'�5< �!����!�r��4�)��<���z�@D�P�Ź(���Qօ|���I<�slփ)�$蛵Α�M��H D&Lz~"�'�r�'���x �;���
��8/8(��'�L��P�G����Gܾ6�]��'���b���A(u`���an����'%��h"��}�н�P��+�H��'����3ȏ�bu1��Q�9GJ��
�'E8�'���x�.����H:*��1��'�h��s���B�Ħ��/���
�'� i��6Lzz���� �d�
�'��Uj�T95��x:��ԵnK`W@�<�w��\�B,i<x�RĠ��R�XC�#kF�cq�QK~T�#��6�HC�ɻ�t�І�8�H�;m�+tB�ɒD�l� �Z�1�,������T�"C�I+'�.pˑ��7��a��F��B�I��t�Z���	9���"�߮�dC�I6"��󱥇�L,�2�B]wzB�I�F���
R�E|f��ӑv$�C�I�t5z�jE���sr8Y֭��C�I80Efx�QdD/h�`d�6��
�VC�	�.]1cm��n��)/?@C�I�E�y�w�">4v��ԁ
��B�ɖ3�h G_�8?�P˷�;4�.C�4!�xp��)E����ys�C䉣�pȣ�c�e�DDp&�O�@�C�I�[�>%c!��\�`�O,xTC�I�DĖ@!�~-�H � PC�	&\6P�#fi[1
�H�P�
�/C�B�ɭ_p�YrC,	�C����Z�,C�ɰP�:���Y'6����dڬ2��B�	�w�j�0"����Ac.��{y�B�I�n[�᣶��0����Ö	��B�D��a2n��x���ԣW�~B�I��=B�E��C3iL��W [��y��E��J�I�$\�W�XMө�y�a�-?�����ۓU��(Ӄb��p?d�\��Mc�E(	c���!���$��|�<) "B7�:���X�%����k�y�'�@Eꢈ@g�OMH � �\bҜ��Oս0�2�P�'P9æBֱe�l����V���'�dyU��V�S�O`6��Ѡ�<	����O)@#HtP
�'>�pѲ��|���3!	P�2�O
�
� :�p=���G;�\0Bq�P!�F\�c'_J8��p� ����uɞ������ N��,T0NQ`���	��Q�m�1��NB�YX�p�a��hv.������zޭI��#?!Q[;-u(�Y�D�'.��yB��E�?��f�F8!���`��u�����=D���$�Wd��M#0H
\f��F˩R~�B`�bD�O�'T8�1�������5E	����nؤP�󕁇X<��ܕ>ɮ����-/��a鐦� 5�4�'����-U3A� j�/ɕP��Fy ֡:.mQ��L�3&����.���0<�ua��5�3�Dԧ!��cV�Ȋ0�J<��h�&vKS��'nFD��3m�Qj�i7�O���RLƜT�
܃��>aF<�r�����=�z6��V�
ț��4��<ڷ�Ѻ��!a4�[V|�p"O�t�VA'NvU؆�� N���Wk['-�q�mO������� >�� S3�:uq��:��ʶ�ք1��O:tu
ݟt}d�X�/��TP�a0�O�!L��Iwi ]�fʟ������Z�Q�,p�G�!�&D�$�C*$0��"O�+3)�q�R0�� �	5Ֆ;�c��JY�Â�] ��a�ְ\[���D���x���	� m�Tۄ������O�$[����'�$���珔	68+�խ
[P��=�'N�d#"��9 :=�&Q� U�H��WA�<#q�P�w�ԥ$h����s��3r7��zB%�) `��U����;�|d���\%�����*Dg2�8��GM|e����5e�bip�B��6�#��l~�b�*w�l9$O֜����OL�'s��E���)㪙8�bI�O�ɳ�*=DLS�ԁV˛�Lcu�B��5��c�@�4 ��py���0a��P7F�6�L&�'��WT	b��`�D���G/��ե#?������
�:���)�^�P��?��u���z��ɸ�h��A����b%D�pf���,Ө ;�����:uk�)��d�@�,��rӡK��91TL]v���	�,[�d�R�NX�	�u�P��%.a���6�䑁��%sA�:0��b�(�QIA>��Y0L��C#ɧ����֥Ӓ���[�s����B� ���O.ܚ����OY�4�E���D�^}�� #���O�%���ÿ/���䗂y���1'Ӵ��2sO��	�y��#��?�;�/��4?ͩ�_;J
|Y@��k-��b)��yR�4eܮE�ԞY�Ddp�	A4�?Q��J$1^@�I&wD�Q ��<�ӾD�?)kp�
+Pr��ef�D�pC�k؟�q���5h���q�O�"g�c��*, M�"ځ[���	�6T`�`�O�)]�s҂�$j2dk��u `�Ӽ�xM�U�.�aS�Yy!� �&�Ǥu�%h�4��%�D��9|���zgKc&���j�H�1���ol��dۊ%W�̈Q�q픜)�I�*w�I���i��\��P��eղk�f�I{?y�'Wf,3��R*&��5M��8~�@x "O|]�'H�zb`jva�u�̘���Ǖ=� �#nF?��'���OM.�#�F�9p0�ݐ��$b��� 4���%��Z�$�����a��У�o��K�8MSD΋mN2M��OG?�'��8�0�](�b�8ST ��{r"�!}&��C*KAL	�0����O��7��>j�PXfJX�y-�:��it���QaGx��+�/�	5�@*@�ʨ�vE��cJ�}�x��	<Q*`��:-P^��Ţ���(��h��J�V����B��I(���~��O<) ���$�\�S�e�+3D�Y M0D�H����p���hќ"�ȴ�S��P���#=�	��?�3O�i��bh����߼�@�ǴE�V���O�8R�xh���\<�D��W4�]��t�|�S����Y�`9sAۥ	0rŗU�����O��	���'�t��D�yxꁑ�dC7;jD��'�+�:��-�ԅԮZ(ŀ��fP����Y�8�2`@�?GN�b���P�-�A����=	�F��H������W5�&�d~"���K.j5:5D�	�ީ�� :ḧ�v������(� �S�c�_�<in�t�>��V��Y]	�Df_�VamB�瓎.�n��=�O2�1P�ܞ�yw(-H N[�.�=+���2� �xr .��C�Gt1b��q��cȘyM��bW�̍yF(�3��<�𩀇&6��<.tL�Q��#
0D����H�J
��d�
'P�%��-m�jTP4�>W�dɢ$ۑ�&E���KZ¥[�G�j��[$fB�Y�P��d��9(�	MH
A��� ��%[���TČ1��O&x��j� ��4<m���} ��qg��[��Tӷ�X~��ȓ6a ���h!�Q�%����I�<��X�S06��0�t9��. ���>��R (� M�z��s�C ��9D�d�@ T&6[8-�BF� {��$%?Y6ƕ�J����D����0ãE�
���n�3@�~��&]���Ƌ')W�q	��W�*#`M����3�y
� �dS/�ޕ+EB"T�V�qq"O�=q��;.b�(*]>�t��"O��H��/7��%��K�ߌ�B�"O�\pǌ�j\��e��3.���"O�u��K/G�$�q��ј����6"O����لUm���t�?��3a"OBQ��\�]�����G�V-j��D"O88�U��,b�\@�OF�JL`�"O�Ժ���[� 4r�A�5fH)U"O,,[sm͖.�� �k���͛"O.�9WE՞$3V�;C�Y?�4@��"On��c�"b�,�@E�۞-��� "OD�R���p��� �D�8;�P貣"O��v��� j�����K����b"O. �� ���`qB��J�`"O�d�3,Z
|J��5dr��R�"O�,��C*-\�$��dB�LL�೧"OJ4�6R\��B��-�@��"O�Ĉ���3W��<2!�ϙ��=��"O�u�Z�.�js!U�乐�"O ��W��2i#� {4[7��Eq"O|��f��&���J@C݅M�VT�u"O@X��S�R��t��+X�xӊ\��"OhP��#�A(�.bzE�"O���a x��H�M]�6R�D��'&��vJL
d>�=2W"J3(і 	
�'������!
�0r�dH�4wl�'0�B�Hܶ*>��C7��2��R�'#�tj�N�z�jl�3+P�$D�-k�'s�(�����bM>X�B#�5-�*@j�'��dC7&�3b�4t��I��8��x�'b�Pa5�L�D����=�%C�'�W`\ $P�I�QB]9Ė�c�'߰�s �5T0-���'z�d��'Nh�;c�Ǐ���7Ѧ���	�'G�-[�$�
�>I�r�|�a	�'F�iCЃ��8p}	�J����q�!D�l��k�X� dC�E!n�e�g�?D�Ts��J�l��*fAC�[���K+D�R�A��d�x�I�))��qk-D��Т�u�J2 � �o��`,D���e��C�N=q�,�-9��!/(D�䚀��w�L(ӷ+S!z{�`�Sh3D��K�a�RHFY�kͺ,߂t�D3D�l
��O>%��Y��"�Dԃ��0D� ��90=�����Z�p�A�0D� Y�Ξ�^��b�Țg䕃�.D��#po^���U �X"=>D`�m8D� )ä�h}�s6HQ�X8a�E6D��׈�61���aQ#I�QX�;v�3D���s� YL:̪w�3|x���0D������'`��HQ?��i�h,D�d��cZ�Q�YY7� *�Iw�'D�P$��*��L@���LR��벡$D�Ī�kpҼi	fOUT�F��n%D���6L�!������"�4��B@"D����/|�bUs���sX�	�#�3D�9%E����>4���d/D�JP/	A<\�O��̍��$/D��QTd8{�|��h*��y�`�+D�h��F.]]�eR��K�b�Ӑ�(D��)���L'@�8$�?��bAl%D��8TLۏK�>��r�F Ё���(D��:�M�p��}!���%`�ı��*D�� �0[6�*k����q�S�_2(��"O���2��ElT�Kį_��=Z"O��b�A!	��S���W����"O�m �d_nN��q`��ל��7"Ob���IW
P���vȓ�\%��9�"O����'�v�R���M
�B�"O�y����L+̚QQ&Q��"O���F�	@n���b�8[�}��"O(Љ@�\3��r��}C��3�"O>�ac	҂;W0$ �ߠ!����"O����'�B��g��3lҍ�a"O��B���<Z}B��e�'c8I�"O�U*���k�����ͽ)�d�C"O������0����]�n�Xs"O�u�V��\O,�E�_�}�"O�L	Y&	 �T��9J�F��"OFL���� :~q���O4g�$4�"O��(��F�@�`�a�#=
:DE"O:�i���2#�|�Y��K,L	0-��"Oޡ���)>jy� �85�
""O�I����:x�@�Զ;TS"O�S�]Q��agn� g�xm�"OԌ+dGi��Ò'���ڒ"O�����,m�s���^��"Op�*'��������Pd"Ot����!z���	E���q!"O�ua� Z�[��40�ȕ�y�ȉ�"O|L� (C�z)�g!�5>o�M9�"O���Z���o��i����"O(����ni*��ț!��As!"Ov(�s͡�7g�c�@(a�"O"�%D�c6pi0d��X�B1ȳ"O�I:����Ui5H@�V�dP"O�6KÊ��`�M�3z�]q"O�5���
�z�Jd�A������"O\d�F�6���ӧ�$�����"O�8i��J�?��M)#!ԋ'�@@��"O��� ���U�(�����~�6qs�"O���r��]t�`vɓ"~f�9�"O&�Y�)���iT�ƈ t\)C"O�m��B�>p',BU(кur�4�"O �c'����haG1(f�S�"O�`�&
�'�|h2@�OUap�"O���ܵ$�n�A��
�3�p��"O:��b�Y�p�v9	�.\=TLQ� "O�|�1�� xk49+D=�����"O�(�Ë߯1׀����K��v���"Od�ī��v��t���ĵ;�px""O�𳕅J5t��E)��T�C�}�"O~�j��w�l��H���u"OF]���Y�+�����'tt�u7"O�I��ƾ��u�R枻F���"O����&,��kQ �5��{�"O�!"�ڲ*n�Ђ�oC�a\��
�"O�S)��q|.i��EI7MEh9Q�"On5pV
�>Q����J�%,:`	�3"O�+�J �2�l �U�Y�$�@p"Oֈ��3Tܶh25��=�A;b"O�1#���A|�q�N׍p��"O�1c Dc�U@��6E���""O���� Ҡng�M� ���<N��"O>80�$�RKF�;B�T��Q"Oz�F�5F��]��nB�,Bt�R��`�O����P'k��1�Gl&~� ��� t0S�D
�[[̈����C�I�""O����ðzâU2�˜�J��  "O��(�JP
�����T��"O�i �$�c*�Lᖀ�2K�
*E"O�hQ�D�b�AQ�-Q�fV��6"O ��ѧҕ��
q״�95+ID�!��z�p�(�op�uJ]�?�!��7�����1Bl�p�QJ�Lk!�DJ7��Q�<Yġ�v�A!�V�{i��Z��^�yQL1��'_�'��|bnD9<�\�K%�(&N
�{�"ի�y�AG�J�y�w�8�ޡ�C���y�
�e�D�RF��7V-`F+Y��yr+[�+���t�U�D�hu茗�y�	K',4H���m� UB��t#I��yR�8Tjz)`�N8� �1
���y�ȓZ����(��v��y�O���M
�'J\#��*I�
�a�o�847����'��!�"�� K���W恈]�4Ej	�'fv�9����
�|��º � ���'��`�GP�S�nQ�#�J�z�'Ҝ\*׈��t�I�ςRi�	�'��y��C�-�t�ɑ�=\�&��	�'�n����&nJ�8�-�l���	�'�JI ���
�� �`M;Dt�'t�|���T���q0 Ht���'HF��с����g�[${>��j�'Wli�#"T�H��M
�I)�'j����F�<J����ڸo��Y�'U0 �!��Z���aZ�i3
,X�'�l@�4�D VH-bdL�9�zlJ�'��p�dh[�>��,d�- t5 �'�����H��>^>5s�8,
A��'�X�rCʔ�`�T��W�A�$�'�`�XS��D{\�BϚ��,p��'[h�1a+�� �
�Y��'�(HVfT
3�z���nF=�Z�s�'�`)��+	<j���*P#|�z@B�'%||!�a��B]���#ԍ`CF	�'&�=#W	7^mhI&�^�&D ���'�iS��L�^���aA�|�*�'?�R����J� u�4-������'�P�U뙪u7*y�`�R7f9�'=�����R�∁�n��(�"�'�����ϒ�5��8�[Л�'�@,I�O�N���Н.�m��'�X�
��M	B�v� r��Fm ��'�J4âm�c���a���Lz��	�'9���3 �����3 04s�'�F�!$��2e��T�q�R80qtl�
�'���fJ�2 �9��Ċ<��l�'�820FUQ�
x°m�b���'�*��s�֢z�"��Po��b�vaa�'��T�5���X����L �@�[�'!���`�@y"	j�o[{��)��'�J�����{��#��PW��#�!D�BbϏ1�4@�UD�k^�8i��3D�Xc��Y'cʰZ���5l �Qp�$D��bf�P�
m	R�-h�,�ô�-D���g֧S���0���� � �>D�@jV�.)�����Y*A��{�%)D�l !�K8+���rn��S/�)�U�<D�|q'���:�[t��	H������.D�h�'�²5M��t�@�1��-���+D�� �8XA�վN�.b��Ͻ���p�"O� j�m0G�X��END'�0���"O�Xp6bAl�l���������"O(� �)Η#C��#�3�$�5"O���%����˷b�6�pl�"ON��r�S�F�0=�E�ET�8%"O�1p6�'m���
D�?M<���"Ov�� Ę[4"a5ˊ CRB"O\083f��*����oH�a�D|1�"OX񢔨	�	eL ��%��2��iq0"OD�S���i7�EY���.k�P�A�"O��q&��}��Ԁ`����F\ѕ"OV���K]�,\<�6��q'��C�"O�ᰣ��)
�kDõ��̙a"O��a!PѲ���$V]ʠ��"O��R%�Qe��a�U)Y�3w"O�DJ���H�\�X��ѽ6�T�c"O��A�77t��G	�hxe"Op8��)�'R<CB-�7$��A"Oj�����c�ԡ1D���LM�"O<E���
�vx(q����f=""O�\��)P�H���ڿro�L��"O��ӧ�R��X���6LzA�!"O�}� �ev�AG pC�	�A"O�s��W�1�����%4�\�S"O�y��ӥ���'�� � PR"O0�+6%�O�.���0�F��"O��d�&*������w�&� �"O�ajQh�A�P�yǎ�vM�W"O�lT�P��>���Ǆ"h|���"Ou ���pT� *fƓqiN�(!"O��s �E�a�����$*`��Ku"O$�1#$�:k��:rj�< Q8蓗"O0��Ǡ>N���n�9>K���"O2%AC◨JF�,G��"MF�ap"O��s�B�h��<��N�t�T�Ȓ"O�q�@��O�8����ƿ,���#"Op���j*c����R�����"O�ݱ��ұ#y��&�&�L��""O:9RN zE�9�OE�!^�Xp�"Of�sb��h�I?AH4��0"O�{P�?�������%?-�$C�"O���eC
)'��� rڧ'ͻ6"O����N�8u`<!F'ٕQ%�d�"O|l[��c��I�.{>���"O�(�C��-d&��Nc�Q9�"O��#'�r�r �`�� ��d"O>w+X/��t{6H�4`���P!"OZ=�3�V�i�D@ae��:�6�3�"O���g�!����Qd�;v��I��"O�%I���%��ҵ ́#��*a!�$ʆT��
�} *�(p�Kh!�!�j(KFkPM�x`򫇣{M!��T)��H��-OJ�����NM!��>x�쑰Δ0&&�����!�Ĝ6w�[��'A����C�$�!���k�y�m8D�,e��*(a1!�_3�t��$8�~p)���s&!�dU�3I�u���9�x����Ӑ�!�$J�7���N	!��e����#A�!�^1Pz��	�2�݈��V+0!�$�+:�LY@��	�p�=��Q�2!���
����R�C��L*��V�h!򄀅� =���Z�t��I���I$P�!�� �ŀ���ҡZ�V�u�Tا"O:ő��ȨW>`Ȋt go<e��"O"Ѫ�]i����߻O}��9�"O���΀Do��9`��,�>�$"Ol|�oP���Ð��\0��"O���%��h*x��s �4���IE"O��*�J��I�,�B�ĉz�ڈ�'"O�E��!�R;�!B@,�x����"O<P�D;�Pp�-N��2�"O�Crj![��	����> �֩c�"O�M�q��2u��#ч�!Q��DI�"OH�2�F��
%D�;�eT��zX��"O�q3d���c��#s�.)[T"OZ�**א��`�,G&|C����"O�����[����KA=��=k�"O�T�Ў
����C��Ѓ5Ƹ��"O�u��C��^ Rm�hǑ@1�Q2"O^@��%�o.���%H��i���"O�����ݖx\(�,ݒ@:��`a"O�� �/ʀ����iS%$���"O  ����g�68C6���8��"O�����B�<a���w�Y9S����"O"����Qa%/?G�I�%"O(���)�dI�J0&2� S "O"����C���4TB*r!�`"O^��6.��W.Bq��՝E���i "O�%��F�Q��8�C[/OrZ)Z�"O��	v��EL	��Ť0ł81"O�ps�.�1'���6�
�j��c"Oj��1��T������܌]���"O�Ka�
@��AJ�E��˲"O ZA%K" 4`q�E]�Na�"OP"�@L�G�<�9SL؛o���%"O�f�I�ѡ@*�V��c"O.MqIÖ?J3G�
�N��"OT�h枦`��)Y��5h�H�Q"O$=`P�Kv)��t��+U. ���"O�`��@[�0m�����(Y����"O&���U��5
僗$FwN��D"Oi�F	��(��@���v_ ���"O����A������3R��D"Ot0���LB5v԰��G�eE��{�"OFp�e�Ԭ>�l��i�?�j�"ORP`�癔AMڍ �ЍW,��w"O.�Ы�D= r���4|��S"OZ0;CI	Xz\P����>$��Y"O�A�o�$j �8)���0#�B�"O�`���2&�]b5iWSl1�V"O�lRCLP0B ���BR�*��7"O�uЇ�Ʈ�z��U�o��"O"��c��<iZ�T
�R8���Z�"O�)��
�E�!$˯o�M�3"O1Z4P�W�2a�1)�7MBTu�"O]�D�������]�6y�t"O���%O<v���G�c�����"O���4��ƴ뱅V�M�E��"O�qy���>]z����Å>y\�c'"O B�M�J��� 'Z��"O\��eS��]���.i��"O�ʂ��>k���P�N�҂���"O(�CO�;�`����Q$-�|[0"O����	e�Y!D���lz$�`"O��p(�=���' �^�B�S�"O\t�<B~l�E3:�:�!�"O� �U���V:]S�$Ѧe��W�P� �"O����IƗ],�jU�ҾI���V"O�!�M�_�^�bH%4��a��"O�}�`	.��3p� - �)�"OndJ�ˈ�\�y$�Ǭ,	����"O^��"�U n���!�ֿ�,I��"O� c��[��@`邰F�N�w"O�S��˔f!���b�Ö��"O��XPA�H� P�"�́e�p��5"O��#��V� lN�"�K)iR.pR�"O�����\	m�L��W�רGؘ�"O�!y%�Ϡ%&�RҊ�N&T8�"O��D��"e�lj@[6_�AZQ"O\���)�0�3�!ԆX�����"O�U:
F"��Ig���
��R"O�����7����da�g�<%�"O�T� ��P����/�2�T=9�"O���̈́o�.9E�Q��D�i�"O�!�"e	R�����'Ā"O0� Ђ��K���x�����\�e�!�$��G0���`/նg*�ɚ2�09�!�иb�N���7@$�0���!�dW8>oR\�1&�#ʽ�&J���!��	C���w�D2x�Z�(!�!�D&�.�q�lQ����P��%�!������d���*�ft[�� �!��NA��xW.��s��`�H!��5,v䕩�N��y�d�0i�!�>=�"m 0.p���I�	$�!�DQ�m�>��nW�/sx4����h�!�Q�;������,��aÇE:o�!�ok*B�K+�j�3F�U !�D�D�����)=1��X[ƊNm�!�D�����zצ�O�f�c#J4�!�D�3{h�EH�/^��C�ƕBg!�$�=N�Du w�(Fc$�D�nP!�D¬h���t���M �3e�=@!�D����Da���*b�H�Qa
2A!�$��P��(m�:���j�@!�d��{x�(���#�<h���QG3!�Ė�L�|Mb�C׉^{e�l&!�d�
0�9u�gm �����
!�Ʈ#}��p �
Xh��`�D�!�$�������!�D��j��#�!�d�$l����2�ƃ/�x�ЊӲ-�!��Z_v��E)v۴]X�2w!�䙞Hd��C�ȓ=�l����&X!�dަ=I�J�K���, @�̋p�!�$�	I��ECAVE�&!� ��I!�P�^]6ܒ$
��P���-C �!�$��/+��p3�]�Lr�(����<�!��T3��4�a
b��`w�!�H;sԶe��*y��ۣN] i�!��@�E`(!#-��Uffm��D%yZ!��Q(��=��T�Y����l�lJ!�D�2_�ը��Z�.�rq��%O"4C!��iʅKg&^�f���;��C�94!�dX��(�D�%�8 8��	�2�!��(NA�<b�eP>=��B�\�!�dƤ��ᣤR�6Dܢ��W�T�!�$V�KD��"q|*] �k�0rF!��x*I3�f9��%#c��;s2!���RRI22�w�-R��"*"!�D�9�$���T~Ptr���'h!�� r,�$Ӗ^�@ :���@yf�÷"O�PbȌ(t��i%��K�h��a"O��R��'�� dU���r "O��x&C��|�������q�(�[�"OD0�Oֿ,WZ����6Fc.�b�"O.,�Z3����#��r����"OB�x ��\!0��qAD��~[�"O�Jq�آ.���q�-á��s"Oļ0a�!*B-�$�R-Z�U�"O�-k&�Av?�Q���5N��C"O����2���DO��03�%�"O\�[���nm6��d�L�z�:���"Of�HЯFKH$�P �3aqv��1"On���OI�{�@!#F��X��"Ov�u��p�֑ Ū̫,��x"O!p��E�FdD�2�I����[S"OR��嬝<R>���"��"O&�+銒|?�X)�K�7Y����"O愉�$=
6�{��%I��e��"O@�t�C��&h#eC�pޙ��"O�(�&N4�Rӧ푲Mk��#�"Ol�y�]#s�l�@PC<6&4B�"O��R�P7p��$;!�Ju5��v"O`гQ�L-���U	��9�aI�"Oz�Q#l��jDS�G��"�*I�6"O�tZd�dab��	tL��']R�!�D "��q�ĳyf@�qGM*J�!��w��ܢtK��S�� AR�:�!򤁁zV���+��U>��K�`Ԣ!��3<�42�}:�}�"��Ac!�D�^��'���;��y���S!�D�!Y4t�ycB�j�ր:�Q7& !�$�}�f�Pu�ҳa����J�1k!�$F�
���	p@��Z=bkEi�}!�؄'��a�nM�R4���e�!�䆓\��yB�Q�k�R�3���:&�!��{�p۵ჱd����CƴUM!򤄻R��	�Ư���@3b�3i!���վy`c�-8��5S�*�&%3!�$M$Y|�(t�؞i����ڻ3-!�$^�nު�r�3]~r���2!�$�*�rMc׋ɿS*P����1f�!�D��{��-1&�1yL��bFN"@!�dĵ9�8Y�L��20�����rE!�5a40�4��,��pH��!�ē�Dن�#`��v���#�!��	�A(�0b���1���D'xa!�$��?�aBs ȟ�����cNS!�X�_[@A�mCd
�I���3bV!�@	;�4X�W�|����U�&K!��).�:�hĬ�̔��M�I+!�䅀nPкv	޼��P���A4!�dG]=	��Q"xm[�P�>T!�d�N 5iD�̡�X2�.y�!�S��B���B -�~���!�D�5\p�!���+�"\�5�݊WX!��Z���Z��NޜZr���wG!�x���F�ҳ2ɾ5R��?_�!���#���ek�(D���Bu�.+�!�$]��avI��~nĚ�����'� @�NU�N�����)5N2\��'z^� ���u��j�b!��ȓz�$��líY�Qðe��-W�8�ȓ�5��܋�$L{f��cP�x��S�? |I��ΖGV�H��ׯ}�D�a"O.�x#"�2e:���"��)dp��"O�Q��䕙]F��+e�,�LB�"O��hT`�
��T#"wt�K3"O�uq�nc��Pp��/X�Z�"O���!}��� &o �"�"O�ly�śH����.A#v�:��"ORh�Č0$L�Kp���NXغ�"O� Ӷf�P⤜���ߑ&F����"OH�b�OK"8�G
X�R$�#�yR��L@�����D��8�����y���dX�C�ŀ4R�!��F���y�h �]�ʔ�$+�L�bv���yb#�8Q:؂���$���Fo�)�y���fΠ��e`�7 ���R2�)�y�IH�9�����Mٳc����O ��yB�KFl�ؘ�ꃇqg��C�?�y�*� Yd�\{	��@��ea"ꞿ�y�$�z[ܹ�ͅ;�`����ժ�yr._�4�~��P�O?/��-x6����y���O�⬁eQ�r?����D��y����E<�Hk�nB�p�5�4�M�y2gϢ2W� A˕�b�h��d�ޔ�yҊ�l?v���d�U�@h��E��y�C
	�T�3U�_�"X.]��ܜ�yRG�� �ȹ�p�����8����y���L����5�,a'�R��y�덒$���k�-X�ZPH�'N�yb��06PA�!�@ ���&˿�y����|g~iwcɔ��ѲV#��y��E�*0P��X+ ��l��DO0�yb����h$옎�%�ٜ2&��ȓ1m�q��<\�}R��]�B<T�ȓL�� D��"���ӱ��?�D4�ȓr�4��&�(c�)R��Zo�q�ȓ##(�	��@ jWYX�*߯|����m�X����R���'�6�)�ȓ,�,��G��Onř3�D�3&��ȓr�����cb�j�4�+B&���g��A�B� ZG�W#QN�)P�"OB�5틀WC���v����<��"O�#��߂������o8j�"OΉy�����ȊwP�z
L��"O:�8gf#9#��IAm�>[��4�0"O�]�fJ{��R%�С:��Xy"O֔�p��I/l�Y'f	X�@�H0"O�xɧ �t6н`Q�M #����"O�Ɂ�iQ�N��+F�Ӷ=侸Z�"O����+fx]�㈋$�豰�"O���d�==5�yX�a�k)�d�q"O|u�6(�5v�:���73�T��"O!�h�'b�zX1�%�-k���D"Ob�Q��lT�-�!ƞ���� "OB�"cE½W���1!Eǻ-����"O��.mŠ
R-L5@��F#�y2�b����!g�B-Б�&�$�y�BJ��RUO^/2;|�1�.ɗ�y�n�* �<�rb��-�<�!'���yR���)�Ű�CJ�wd`��_�yb��TO�sj��m���3���y�K@9N����*�Gx\���]��yrm�gf`,�/�Wo*�ӂ	��y��N1O4��A��1R˚}`�A��y"o�	O������_!{���h���y
� �`0B!sP���Y"?�@��$"OF:��Fm"L�6�R!#Ϣu�"O�;PԬl��ic#�&�x� ""O-:)�M�vE#�/�����"OL����DP�2���� ��8@T"ObAbG$X�Z�:"�.�A"O�UᑣBl�4s�L
��d��E"O�\P�n_�b� ��
Y){����"O�4(�%�u��1����Ow�9P�"O�Q�c ˓K��|0�'�fa��""O�2�iͳi��2�Fük�|��"O$�qs��+���+��/Z2��i"O��c��x��XIB��=9#0���"OV��ʚ�(� �&�F�;,0��"O�=�rŪDb�i`H�{_�H�"O~�`��{Xz%sW�z+-��"O�� �&�.:M�(���H$�kG"O�E9"�	)7��ip>���"O��xd��~��U3ץX�c^e�"O���!�[9Ly�$R3\8��"Obe9UBE�-B=�C�ّA��D9�"O~\��G�p��� �A�N��"O8��LZ�p#b��Җ}�����"O�8��Nl4`�0���W����4"O�$����o����LJGn��S�"O}�s�;`&�F%Z4TNε�"O���VO�E�bۧ䉣Gת|��"OnH2�L�&�! F(T��۠"OlE�[����;q�����+�yr�տ|t�`�5"�1�vZc�Q��y���e�\0�s�ՉS<�Q��_��y�#xڌ��)O�1�2��y����bC�,q�ve"J��y���j@G坁g�h�[� �,�y�.�j7����Y��5 T���y��؅\>��[��W�r0JVM>�y�؏>�i�@��
Q����ej���y2&�D5*EC���S-f�R��y��.�R��(� !X�@˔�y�u�dY'H	^V�����y2̈́�j&ht˧�9W~p�R2�y&��x7�,0�C�"{�i'&��yB�ȰGR�\�ӈ�^Ϣ���@��y��U6i�D)!-H�)�봀�yaG���d��*!�m���\(�y"��A���Q�S4���Pʈ��y���*HO8���̤�b����y���8$����m�{?�X 5#���y�D1\٤�!��ߝ���d���y�^�h�T0 ����Dp��M�9�y�F�Y줜P�.5�|� ��yB�"z��u(,ws���a���y��r��Ws�hPka���y"Zn��a�ÈqB8((!���y❼.��$*r-�kb*I�@����y�^"\����Qg$/�x��	L��yr�;*e�ʧ1Hh����yrn�g��M����$x���f�۲�yr�]�x*֭h��U1W���3��,�y�̑71�yX����X"�����PyBÊ;��5�r�޼F�e!B��q�<A�g۳9�|����Ҿp�U�Wj�<�Ѝ��D���BD 	�_��"!�Kd�<As��)D �E@��� F��I�C�y�<� U�EnƝV�F�i��oP�q�"O$H���i�T��U� �m���"OԠ#�!� �ӥS!��]K#"OR�2 &QA�nV/U�l�9T"O�҄������@5W\iA�"O&r���O�����8Q���kG"Ox,[R�2Y�:,�a����I�F"O�`�u ���SGBUk�j�s"O�C��� >5�zD�N�k��Lb&"O
��mH�{|�e��'&Q��"OLqHf˹E�81"Dӎ*�m�u"Oe)�a5�L:N~�x���"O����&Q_��:�j� %f��U"O�=(��Kz;Ă�� �$�d`�"O���FI�'=�<�Z7	�<g9����"O|Ayak��Rm.����֧)�}�"O��pMM>#�pDaF�����t"O�٠Ӥ�jպɡ�J�@'lu�"O����x9��K�M1�0`"OT{Ӕ\���M'l�q�"O�e���݄{FPYqF�H����P"O��ʴ����Τ`�Z��ͣ�"O�\�#��"iV�i�@Ҝ^��A�"O�P�2D�
԰��C�|����"O` 2q�:LP�p��ŏEj�	"O��bL ��eXr�������"OZ��0��q|��v
�
�d@+"O,� 0
̵+ތ@��K���p�"O��aץ �x�&�:�h����'"O���e)	 ꔡ�&�Q�$y
%"O���Å�p��D��掃#�� �"O�qz��K�[Ԑ4O���"O荓шX�,v�O|�Y w"O�W�ۻ|�,�Y0l�^v�� �"O�!j�EB�1@�e
�T���@"O�u��c�2m���A�)��I�
��"O6謨Xf(4K�샏6�T��1'�Y�<�5���~o8P4�Ge��P��W�<IQF�9;�����ʛT@ ���8T�lpwπ���h�%�M�:��$D�Zd	�t���Scѯ7oF���!D� ��+׿[q��@�(��2(y f#D�t��o��t��=��i3.�9��!D�РqJ�9&q֡���"w/fA�Pd4D��W�� �
�k��I1}@����0D�Y���${�i��D/��Y��*D��a��(�rè�ƙK N%D� ��ģX\��j
��|����.D�����~B�\</�HU���,D��(mߪs^�[�W2?���rpg*D�@��ĚxL`��C���t:�C(D��'ƕ*L��(�RCU3iP��&.1D�|�.�#|�1�C���h@�2D����k�{&�����
���IVd0D��J�N�x�Ε u��
AC��0�(D��2g��?j"4i6��P�|U w�(D�@���$M��Hk!ZdZ�!&D�����M�b΅��O�4o��E#7D����Vl�~P�� |��H��i4D��J֊�3_L����ˎ�I4���c�0D��H�_�PS��%��E"I1D����ƭ2��87���	��Mz+*D��P�F��2�I!"v���*D� A�[^����-]�$�䱑 *D�� ��Bc�%��Q��G�"X$��"OV����C��P<�4�EQ��u"O��z���G�L(�\�J��Y�$"O6���-M(y���@5nM�p�a�u"O�Yƥ��{���ق�//f���u"OqB�@�P�|�Cv��,N���"OzeqSj�&���C��Цt�� R�"Ol�A6�C��0�[��[3W�
AQ�"O��9��z�8]��݉Di�0�"O��s4�L�H��]�X�2�"O�@XV�q��Y!1��$�e�2"On��疔�Dm
������$@�"O:����.(};�� d��b�"O|���/�7Oh�2��)[q,`0�"O�=	F�<>{��P���K�03�"O��!dG 9;R�gCBR<�K�"O���0����0�u�@�x<���"O쌸�e�1��BhQ�5�q�!"O<	�-P�0@R�+4H6>1*!Q"O�x�	�l}nޜDcB<�W�2D�|ٴe��E��L�e�΢|B�P�O2D�@q�*���H&�˸_�x@p&m/D��kqh͓L��Ы����/m0�a�*D��wK$
�԰��"Z�nР@�)D���g��#y�!����P�0����1D�ԓc�,|�A`��/Ta+�F2D��`a�Fu@�y�"�3(�`�Q��3D�����
kπ�	t%��4`Y$m3D��'�.�l�˙/;���Y �3D��`gC$�~��3��q�j A1D�I�5>��x�rB� baH�j.D���b)q�`�GMڛ_0�U;�>D���[[f��pE��W��-;D�D��"Ĩ%�ԔkAa=%���f�9D�dX0�}������PmF��L;D����$V���Q��A3K�j��3/?D�`�V��)���q,�#};�lc��9D�p
�g:l�A�_>0^�T&3D��D`�a�x�"�NX�M`J��� 1D�<�#ͦk�p����#�.���/D��h�훩W�d�f@,p\��{��+D��Q@�Z�9�����޶���,D�������$�h�Sƛ�e�I�1i%D�T§���o������*��b�j$D��:E�	��P�2���MQ�	)5� D�0�0G�45c�HP'��  F��F�0D���e 2cl>`R��ܸ+
���,D��� ˢ|}��It�T��H��E*D�@�n��F�%�,�FL�	e�(D�\���[�����E�E:9 �*S+:D�`��FХ'z�5J�@�z���5�6D�@��쇩i���g��x�p��w`6D��&��$J!6,97��1X\�ӡ�5D�\��ON}&f	�6�\7*V8e��'5D�hH��(� =Q��l�@���(D����!�Gp���7��%T�t=��('D���㟃5fx��D�+O����I1D������XI�1󆝤m+H!�Wd.D����'�@-xZ4�Y
y V0�g"-D�T� hؠ ���Y5�ݛmG�R¯?D�I�ҟ$#�����/�T!��*D�Xف��2z��av�s6�R�2D��*sf�<c��*�O� 1� #D�Ȃ���@��� �,�J���C�*?D�� ����ݽ)j}YTJ�u\���4"O@�Xl��Q�8���B�l>�P��"O~u�cA.|l��;gB%|0��2"O�a�f���R+�
|�Ћ�"O|�B���"r�98�*@�s�B��"Ozm��`0�AҒN��1ʦ"OXEz�a >j�� z"%]s���6"Ob5W��9ov��箍;qXlR"O����e�3������8]rQ�4"O~�2�I�k��) ,�;:T ِ"O�t�v"��ŰDi�%E�V")�d"OL8&�8:s���vZ�9EҤc"OpUA��GX�Be�n��f�d�d"O�x���1	$�a�g]�-&,tP"O�T���Ծ�>4@��PKb ��"O�D��%W�M�rL��-k���"O8��
1���E�7.>]�R"O
�#*���%Q1˒"t�h"O��r�KyFQ�`�-���"O�I"ˋ�Q\|c��%\<�ȱ"O����#lEЀs1��%����"O�4I��~W�ٗR�5�p�2b"Oܠj�,@)Zx�ˤ��R��8@�"O\,I7@�8<ۊ����/�p�٥"O`�bFC�Q�Z,K�YC�!�q"O���GLF�귅Z�%�pH�"O�c�+�7�aDC�9j��Y�"O"��3�ѓFr�Tr`�?>�h�e"O�� $ʏ�CNiS%�$>�Jq�"O�@귫��cIԵZ��n��Ը�"O��Csj\"�@���H!��M+3"Od}H�O�<Ug }	5�Z��~m�U"On-W��/`~�"�P4aƚ,�d"O��w�=[�䒳H@,��[�"Ott�"�
�0�����åV���2"OX	�F)ŠF���$��LK�u��"O|�R�)ߟ*T��@*/��8ct"O�!@��G�o������8.���v"O�9P�GR� ��y`�^�4q�"O8	��L�D%��_
Q�mp�"O
:�"8Dޜ��#ܢm���"OD%*�)S X8x���P�7Pu�@"Oԁ!�G��>M�ѤB!��p�"O��D��y��#Qc��8��u"O޹ ��QAB��A�!|��P`"O<�;aKD� ff�	�b�G`Eb@"O���׋@�a��Ç"�4+4Ja��"ON���!A
�}��<r.b q"O����ʤ)0���# < "O��+�j�	��X
-�	����"O����+� ����L_"#��U�D"O�|Q1�T%,�X�Q�\\jvUs�"O���!�S�GA���H���V}�C�IN�~��$�A���5��*@vC�I,a�f�c��?���@q��D�C�I�5p��a�b��g��+:�PB�I�~�^d�sN�-U.�����W��B�ɒA��i�M�0y�4�����VB�I�pDY"�D� �.�Ұ`_D��B�	�Z������>w<,!q�(��'�B�l��J�=g��Ȁ��XX�B�I�I�� `e�Q�h�ؔ�Fƕh�dB��(�fH0s):Xu�`��ƅ�(��B�	w��6%�;�j��soŢQw^B�)� .�c�bY��
4�"�|��m��"O��;��!|M�����|�Q�"O�th��ġM��2��\�����b"O�m�r(�4d;(���~)�p"O
��4�`��9S��Ge���"O��4���Y���@L4)hŐ�"O�8xc�I&Ll�E�%�V>b��8�"O�ă3�ިRx.�PR[^# �q "O԰*bk�;/�p-q�K Lpe"OF� 2�'��T35���4�(9kF"O>�q�B6hk�0�b���L�@�"O�g -+�����ɳ_��$k0"O��AG�Pu���@G8}�Y��"O�m���N$Q4�`��S� a�"O.�j�A�@�B���ԿQ���7"O8Qpt���Y����aE�<[2�:�"O���G��.6\�$$@8*P���""O�4F P�tNܠ�����<7d�"O��JQ��7k`A�G��~� ��"O�K�̑�Nϰ��cE�n��X��"O�<	@���ˮu��a�@�Z|	�"O(��r���~Qs�@ZF��UP�"O,��C�ד�ޅ�UO;,W��"O����n�8i�X
�N��
#��x�"O����ńgi:-��M�+s0�ja"O�-��(ј}2�٨��h�Ȋ�"Oin�x��ez L����RE"O�@+S�����(X��ͣw:���"O̰:�jG� �.�c�6�
 �"Oj-C��#���!C@J�H�"Orq��D8�4�P'G�欰%"O(�r����6�!��Q�G�nl�%"O�A�H� PQ�#Y�����'"O���R$�4g�H���M�=��IH�"O�(9ԣƪnE�Uy��	�[�"O9)�&ƱX��a�m_�S�j!�F"Oz�ZEG.-=���l�̂�k"O���EZ%0�ҋ��"8z!"O(h����
9�LrF�
0%�ּЦ"O�uH֋��{��IzH.���@�"O��+���6&Vq`
F� �lH"O��{)�b�������)� Ӷ"O�@��もG��0����#0��9J4"O�p����6 xj���x|2<��"O�5s��J�`�i�u-�d��q"O�KC��.9x��ۨ3Fb�J�"Od��D��DvRa�%����t"O�Y���ܻTQA�����	6"O8d��aR�h��-��E��!U"O������p��ؐ+�[�fM�W"OxaA�9@�� �ԫ�>n�Ա"O�b�(A
(�5��
�A
��"O���խ�2[�Mb���|��H8�"O�����I<�0�` J�-X��a�@"O���!���k��h��/L�vy�@�c"O�e�/
m"q��ݷ:X*)z�"O����;`��B�Aat|�;Q"O2H+�jŖ	qLHzqLY�j���"O"�@֌�:}����J�i�,�a'"O|T!%	l��MӲfԄ����,D�l �/ȍ"1�ĠnY����>D�КA�$3,�3��B�]�U�@�(D��3�f�'�P�8��E�9cO(D�$���e��D��4AQ�1"ad(D�� X�1�_ [�,��ѫ��L� X��"O�]X� 7�~0MM�M���"OfE���-]��}@�����Q��"OBAr�,��9�2�ݦĄ�3�"O�i�b��8X�p�-~S�Y��"OB}r�)
������¯n���@"O&��5k
��租�Wy�P��"OX���f�P�΍�c�9r9jf"OP�׉L��0��3	ه(0�(�"O8-QC˝�B��T����u�>�i"OV�E��|[���H��0@�q"O��XgđWR��p��S�M���HS"O���"�y3nDI�J��/N�ܻ"O�-�FF��Y��࣯�3+����"O*��Łՠ� �{�gX�a0(���"O����^=x�JYд]-a��"O�UQ'l���b�d��dl	�A"OL�A�-�9�:��4$+X�F�0"OčRàE��^U1���:t����"O�I�f�
r�J��EA��߮���"O����i�X��E/�)!�8�"OR�+��"kVD�!.�?89��R"O���C{R\��E I�Y u"O�8� 1X�.��R�Of��"O�ɤ��<]�x�q�M�=UhT��"O���!B�0I�A�| �q*S�y�R�B-p�PT3]*��0a���y2���q-ʕ����P�\YR�3�y�ᔏZ�saB��Q%ڴv��y��D�B�������\}�"�'*H�1`�<g��0�5EViq�'[(��@J�yj�Ё֟'r���'�ne�ŊZDBP�#u��%~��'��-*�\
�m0��M+$r�8�
�'1�D�� P�s��ӧ(ǣg� ���'��=�D �]����f�I���'��m�Ee��hI*=	F��Jrڑ0�'/ ܻ�F�-�f9�r0�LC?�C�I>�<���Fs�~p�4ˀY�B�I�+y<�"�G�/�<|�	��h�C�	B[j��G�Y�V5T@ƁAA�B�I��d����9�1ٗE}/"B�ɂ5Pf��7IXӖ���ոX��B�	7&t�yq2I��� ��g��H��C�	�eFe��
E�&�m��Q�B�C��X]Hm���,"z���"R���B�ɏW��P�$,ӳ��z"��K �B�6w5Hu ���7 ?8I2q� �2k�C�I�l<�Xbn�����(3h�#C&ZB� /� 0��E���p�ƀsFhC�I�D�RL`�,X��) =s�ZC�g��Y@Bf	�/��#/�~�C�	XT�nS�cΚ@��0R��B�	6S�-�$m��`?�%���)/��B�I5$�p3��0xR�=���ǹ8�BC�ɟȖ%ړ��4�إ4�Ʒs"C�3U�5A%�. ��`E��1H�B�I/`3�	��L�'u���	8Wd�B�5<HԌӆ��+p�Tl:2$½K��B�I�R�Qf����"t�ҩ���B�ɗLm�p�
)g�Q�S�5s%pB�I�Tن��$ll��s@�� B�ɔ*��ª�3�! Ը3��C�I�jd&X� E�:�V=[��S�FW�C�)� ��k���1cO�|4\�JW"ON�5G�����F�(�#"O��3��[=pI��z��BBЍAp"O��'I���Li��)a#��;�"O��A��*FH)I�
#���"Oli� L.C���S EB���"O��
`G,.`P�w�V�<��D"O̅�6���j�T��s(�;Ҧ)�#"O�LѶ`���쨥����b�"O��1bY
?�����D.'�ґ�D"OحJ���^G�� uE�'T�zH�a"O~y9F�D��փ�%X�
墠"OP���*\�H$:�cȈl���"O8�8�"�$c���ĔAb��"O ���+*� �C��eS`}��"O�(�d^�m�|$�3HDu7�H�"Op��� �:���U.����*O����Z� �hJ4��v��'�f��&A�] Z�!����ʉ�
�'�|�b�Dnz�`�"/I�~��	�'���RB�p�2ݠ�ʶ{�PP	�'�z�H�h
0>�ұ$�*v�l��	�'����g3-�j����g�Zq"�'O"���ޚI|l��Ы��[�-��'
��� ݵ�vL� A�U<%3�'���8W�w ��@�,�wu��k	�'���v�^�m��婅d�h�	��'��T<Bz�h�D��J+ܝ!�'�����ΌS�}�amΤo����'���z@���:"�u��4aFj�a	�'����a	�1��U̅�[����'՜�I懚L� �l�-[Jn,��'\�ܡो�X7����*LEd���'x*y���+�*Fˋ�{�̍�
�'n��Z���&sn]��	�m"��	�'i���*Ui`Dȡ��)V>E��'�x���f[�a�v�0�c��?��!�
�'��8�iH�H@5i��0����'m���f�0�pi��*̌-�r�'�t�X�p#�uc� �nl.P��'D(\�� �=[�\V�i��� �'�����2���hfkL2Xe����':�2"..X�vlїLv�q�'ʢ���$r���(@(��GI���
�'�A�䇖�`�� fǺ9��=a
�'RP��� '.j��^�.R�Y
�'�Z�HǮY!d����M�,��X�
�'k�x�̉
?��5Ȧ�̤$#��A�'��Hة/� �[����ZBd��'p�fa�����''R5 7�՛�'�\e�3��`e�l!G�
gH�D��'BZ���`ɏ]Y����K^�d<���'.���X}�mh�%Nb�"�K
�'�:A�5E�Ta�ӞV���	�'̚!hA�l|u$��$+b���'`ڴ�5G@�U�$u���S#�<���'ʰ�S�. ��b6�W/�l�8
�'�Dl2&�`\+�	S�!�D\X�<��!��B��cT)�?��\Y���}�<�*�}:�aƆ��y��� �v�<��ꟶ*d4m���:�
Qs�s�<s��F�������� #������r�<�F�r��@���$e<��A�v�<��i�<6;Xm��-�$	 d���M�<� 0YlR.H��ܻP��&�|:V"Oд6C[�/K��ا,�*�,�G"O�ieLㄋ�Wf���"O�U����5nC��� �H� (["O���Rɐl�\8�I�.߾գ	�'�4P��G�8�`Ek'��X	�'�
�ȇM�:qF����O������'����M�!T���r.S����'����шr���)b�Э-�Ĝ��' ���aa��HfE˱:Μ�R�'�8��Ve��dղq�ڿ �ꙉ
�'��H��e�A%~d�ʊ�)�R,h�'vH!AV�7e����� �e��	�'	P���fĬi�dƆH��]B�'���V�����\�E�\�{�',�[p��&l��;ӆ��7y����'�lY;��R�jl��(�.�(�'l �k�!��&�ԣu��V�а3�'OT�� K(l�v��$��q�ī�'��8�7��t�:DkA�%E\��'In�)��t�D��p�Yd��3�'���s3M]��d�7�Kr�X�'��`�&@�#�T$V=Rh��'�� "�Ǩvd�ڳ��5Ӭ�"�'� �"Q�V��H���/rh���'0�� ��2$Drq@�	�8�C
�'���1���J~��e@Z(YpeX	�')�%�vmF�3Q|���o�}��'��d���BX�䬍��&(�al�b�<�5�B�M����K��.=�.s�<#l�K�:5 �+�em,;s'r�<Q�Uh��J	7/�H ���KH�<	�߻"�j�c�AL>v����\�<I!�)zS�A��(K�> �;���X�<�TMԔ��l@c� N��T�NS�<�� ¡%��� saZ1�b���e�<�����M��S�,D�q�x0��m�X�<�`@%i9��2��!qHԘ3S�^�<)B�	�$������U�{�b���W�<���5~�1�МY�������Q�<��㌄L��Q@c�^��T3�EBY�<�W��x�[�P�0�ZȚvNa�<�b^�8��̂`�R��1�Մ�Y�<񔂉�$p@�!�Y��%R�<��h�m jV�Y�ؔ1�a�5�!�d_�C���w��iݢ�c�ɲ)�!�DjK�T��Q���'n(b�[�!���΄2��z1�,��Eۢ7�!��×:
�d�2�W�g0b@+�Z-H"!�$ m�(̚��ɓA,�dP��L�!�#�0ai3�U�:{�ũq���Lv!��Q���q�!O	
�D��cҌt!����@d{�KĔ!�J��6o�!�~t��d�F��#7�/l!�D��:�|��� �I�
�![�wa!򤟨J1~b�\�0�x�H��՛0�!��L9N$����ňM� �f�(N!�ɍ4W��*@��T��(��)Y�t;!��� #��r��)mw�� �gP�,K!���9�Pp�A@<ZV,�镥�);!�D�4�$�i�/�\9Xã�<%.!�䇨o��(G�%}H|�c�"�$l,!���_�T�@���j>D`�C�Ǆr!�ɰ{�a�ʐ?&���M�j!�� ���P��	p� �m0(�2e"O��Je놏mp$�p֎��.x�A"O�ka�0I{`|��g��L)H�"O��:��� jP��b�^�Z��J�"O�x�
��3��ʱ�	;�L[�"O��#WF��5ѳ��3R)S"Ot9�!Z�^@쌻w"�;!.P�{s"O%�Q �"�d!���F�d�� 3�"O�kE�M���H�*ȗmL$�:w"O%B�fR�<�P+w�Z�+�@�"O��@R
�� ���*��Ӽ�x�"OPL�4�O�7%%JK�V�P@�0"O�k6拜J�����@���"O,���Y��� 1R����A"OtԐ2�B�~�V�� �?i<�!�"O������]�pD�!�V�#nD( "O�)���(p���2G��v�Υp�"Of�C���`�C�"qxw"O�ԸB`
�f.���P�&Q d�"O��SJ��I4������7"O����o�Ϩ�H3A��"���z5"O ��/*B�F�9֯�&\����$"OB��`NK�K'�S�!��aO^��3"O�XSe�Q�J���M�B*P�"O̹�P��GU������ghՃ"Ot�0��D� ��r��8a��"O@Q	%�ؔe^e�ۮ/���%"O�Q��O�R)X�ʿv�x��"O�l������-��ZM[�<�4"O$�FϦV�$I8��V�M���"O��YTj���-���������"Od�����ei2MX�o�D"Ol�bA�C'<�鬘�����Nl�<9�kS83�"�T/N&
h�KQ�<q���'icF\�%�� j����b�_b�<�4-A�I�&�{r&E	 A[�<y�������B������U�#>!�$�6����+8NU6�H"f�2y8!�Ď%z�L"UJID�m[��Q4!��M�w
zpD�I�K�l`�����,�!��O��2ԍ�����褢�%w!򤞒 �dl���$>�X��T�%zi!��׷C��WEC�b� @g���Y!�Đ+T{�ɢ�J>J
BdKr�۔�PybJ�"^K(T3�'�<z5��0	ƿ�yRǄ6��=;7$K�vL��ᜎ�y�A\��a���L6�����מ�y��T�H'�#�f\~�`�:	4�yZ�E��'XZ�b��'�,!��4p�'Ѭ=ɕiU"A�I�0lӰ`U�
�'�tи�!�b'Be���o
dH
�'�x����:[j֥��lp���	�'G@�Q"�Fn��v��8�@��'&�YƧ͖:r���Sa��a�'eHxQh�K��I�$gH$_*´��'���S#��x�����.Z&��
�'M��1��
C�B��@�e
1
�'�ژ*���sD�q��@���k	�'!$Qq�M�?oI� ��3�:ݛ�'��XRD�ҏG>2�����	�'��u1�]�v�2�w�����[�'��E���~��p2�lвrJ�9��'èh�F�Rw9����jX$�!
�' �b�'�{�t%#1H
�7�bً��� >ū��0_&Bp�G:&j��Z�"O��zŊ�W��ys��
?9�h�"O&@�gǋf�!P�d6|%�z"O�51B�Y�2䈍�2� Px�9D�DQ-�Ar�D9�+.��J��;D�$1c�ʄXH%I�)��jU����:D����!A�8����Ҕ�M��3D�Ȱ�Bb
 ���R��,#%C/D�H���֕v�p I�Ȕ~ٌ�c&m"D�$��膲lP �!��ŃI�0���?D��'L�(M[�Nª��r&�;D�p)BBL&�0��߸�{��:D�X(��_����B U o9t�4D����+�7X{<�S�$=5�� b3D���C��
}��!�J�Cԝڔ�0D��hsa��������
��-r�-2D�|j�G/:�H��օAmP�Q�h+D�$���˚)dnL� j�N���)D���CDi���7m�!i���B7L(D��Ҷ
��%�䐸!O�vr���!$4D�\���\&B���حkb�-D�4A'i�P1HX�t��Hs�u��H,D�(���֡j���J��\�^|d�	&5D��0�dj-*��6��7t��Da�0D��x'f�9l�&)�sh�:*B`�"u�.D�d9D�]���B�h�byb,�J,D��@�U�z?��:VH[w
��0�'D���2j��nwf���H�:S��y���<!��哈o̥�p$ϜR<pe�#J٧�hB䉫�8a3v�W1)�Lmit�ԩXA0B�I�F�����T;[��	K�d��y>�C�	�"�p26#
�gøII�M]�?�C�I�?AJ����hVZE(�n�/S����?����%ڗ�f2n��$[Z�xV��y��8ܸe��C^�~�u��(T��y�&Q:�b1��%�0`F��fA.�yҊ^
l:=��.���*��I��y�ș,���# �d�4�p��O�y�!��1t8$�g� s 䝩�B-�yZ�N�iG�͊X�r-��L�m�2C�	 JH�IS���G�lUh��	��B�S�t��rCA�^�P�AG�ܸE�B�(�n��A�v�D����B�zB��h��0����]ܱ�SF�j�\B�	$Wt�S�/V?a٢�ҷI�B&���f���Gb�?t��4��D�=Δ���+D�����?*T��U�ŧ2HlQ��@5D��qEM�KZ,��ˁ?#`U:Fl6D��h7��&a�z���M�(�:�y�2D�L��C�+RQ��`0b !j�n�)r�5D�p �ޓ���p(�$J�^L��C2D�yP�� {�Xhd

���Q�1O�=Qt䍄{��Ta�ǒF��Ё ͊\���=�p-AM�r� �)T�ɵ�W�<��O� � )`�
S�������J�<�g�(W�llsEї��)�1��l�<��F�c]4(p'��;<feB�i�<!��E����&��zw����_e�<Q׉�G����&�H����%��^�'NG�D&� �4K#��/h��-�W�C���Q�F��d��j�l�5O:���(H�`�O^�=%>��GY�Rt�%h��.xkԍ*D���u�ӱf�8|�� �m�`lz厵�زe�>�&�5�g}�`
�l��b2�=�"�`�B�:�y
� ����Q��;gA�#�L�cqȏr�������B9rlaB��*����y��_�M��㵋U
���E�W��y��C�?�	�h�gX�s�J�y��c}
�9���&؁x����y2�Hx4���Q�*� ��y�cR�}�b����U>s��pUmY0�y"m�e5���$�ע4~��	�y"UcU�ԇ��9��A���y��ζtØLP��r.m����yBc�.fi�v��z�J��  H��yb
�->����r�~�3��
�yB��Z�Г�b۷}����ݵ�y�؁m����͕#z_>��f�>�y#-%^�P�p��3p�8AT	�y�N�m=J�AÃĸTi�"�K
�y��N���A��)�`�'�W�y��W�>s�U��`	$F����P �y��F�����hOɉw�U��y[1[|N��q/0e\�C���y"m�1(�)2��Uyk.<�Ҁʤ�y��M�6���!p��*��y���yb��r�<<��
ri"Q�[��yO��JM�j��"|A˰ Ƹ�y��N50|��V�|"��g����yrÀ�:t���q-��|�V����R��y�ΓC���6�\ ��$��.�$��ȓ:ĪiP�!BG{J\Pd��襆�[�,� �D!E%���&�\8���gS\8K� R�4(*�����u�y��oA p"��vY��R�D�z74��,r>�P�h�
(N��p�?���ȓK?���r�ȅ`h��ò��;à�����5���lo�T���7�(�ȓ))X�@�&�lQ����ͅ�(-�ɒu��W� ��sFbOjx��Ql�M�F��5^�@�s��}����ȓ#d]!eh�d�j%���G7;kJ)��ph�� G�[��]9QE�	N�=�ȓMA�}��nT"]��S� I�ȓ���aԯ)|�a�b�K�I������d��-+l� +�5l^�0�ȓB��ن��PH�\B�֚p�@�ȓ<���K!�?)�l�#e�"�ȓ4������*�(Cv₼OflB�Ic���u��\z$E�ר�sR�C�}|F��~����,%jB�ɺQ�*l2�Az�� J���/dB��H��9Af����C	DZ�+"O��;$M�3O�B8�3.�&Rl5*�"O�Y7">�nD�FnY���i*"O�y�Ё�<m)~�8���y��-�"O0 A�f���͹����� "O�� �j�J&������-g�ޤhv"O걇�T� �@�E�.9r�c�"OvE�'E�B��}���t9��	�"OT�K 	 ��$qgnę"%��V"O2�+	"�����ߘ=��pE"O�D���5�x���l�Pp���"O&�s"c��q�t��^��Œ�"O�� ��� �8jR��P+�ib"O�u!��ȅ7~>l;��K.(t�T"O��b�!�~��	Z0 ��5�$"O�=��ʜ4Yd u���F��pi��"O� |��@Xsv���g��B���a�"O���i�n�
����I�yL,3e"O��p����o.ΌH�
�D
F�"O�Dq��߫#�v�ق,ӆ>K��)�"O� �E���D���ڒ�44�+�"Oڴ�4��-Q�"`3�)0��%"O�}���֝a�B�&�[H�1��"O��{1͋�S �0�e�'\A�0��"O���CH���`䋚8%f��f"O��{"m�X�8p�T���Q"O�+`�J$8�R�"L����qp"OĹ Яٓ�����B�����y�"OH�xRcJ:+�4X1�R�����"O��!ef	�-$ UӲ�@5^�B��"OJ���5� )��+�3᪐�"O6������ �x���6�"���y�$Ӥ#�J� ��C�'�*d��N��y�a�.
|�*��G�pBu��y"��	(ly(��U�)_���^��yr���YC.�2��� |���2MA��y��#W�6@ GB��ˎܢrcё�yҭٟY`f��/� oRJ�
2����y�(�6�>�	��R�o٪�a$\��y����ܡ�aN��OZ��.�y��2s���2���o�*P9�ꄷ�y�N4H��΀aјL�t�]��yR͡���j�aPaGrX۔��9�yR� /Z"T����UY�����y�A#_D|���J�$.<t��J���y�e� �X��錅i��÷)�y�Ȋ2?����oN;a��9�Eð�y��O*��zf�Z\�uy�j���y�� ��U��X�Pa����y"�ڇS%�({��4bx�m�3�C�yb�U���2�lN9^R����ս�yb��[�>q�'ƄDf輪$��y�dk]�X8��
�B݀q[
���yR >mZ�
%�A8j�2���F�y��͕"���Rc�Зg�@�r@Ǐ"�yr�Ё��1Au��$/���Dd��yR�N�F4٠��X�0�k��y���-]�H�k���I���H��y� �-ǔl���::��%�yR����}��'8�P1+��Z�yRaJ(Nv��E`%.�S�7�yb��0>.䑰ρ;� �ʁ�L:�y(Q P�G.�N��!�ظ�yb'S
E@D́�By���"�y�KV+�,�{��ӕ�((�u���yb���d�*�ꆃn�Y�hˮ�y¨G-U�p�v�Q�\���O���Oi��"�wCe��L��Ȁp"ODH�ըIq)��	G��i��)�7"O�u)s��l�N�k�Ku�l��"OPP��ӢU�����\5C� U�"O�y�Ň0j=2S-]#X�`$�G"O��)p�4#>��u��2�b(��"O�*�#������ѢT��<��"O��銖Gd�i�׊�usN���"O�,���M'a�2�	�����&"O ����A,�&���N�"O��s�ǅPZԠ"��3�8�ە"O�Z@�ÕC�6�"��w$��3�"O�L��	�k����Fh=�	�"O��Xqd��Ae~�@���r�z!h1"O� ��P�nȆH (B̓�bǐ]�"Ond�6F˒/��y`�c��yQ"Oh1�B�eךD;S�	��D��!"OPM���E9c�zDqC	�k�z��"O$�"#K�z(�p胫���h�"O�U� N�
XH@�����T�f"O�����M��9�NF�	ވ�k&"O,��&��3<�[�(��5�И!e"O�:kL����ĢE'�袕�RB�<�5��_b)�����C��hB��x�<�Va!�h�Je'Ղ
�݉��w�<aUd�j���"u/�w�����VX�<�ⅉ*'|t�1�9Cl\	e.�O�<!���$����E^�{�.q�b`I�<��	p�(�0i�3ZF앋q��s�<! B�	� 9��(;��m���y�G�/\D��/;�&���ύ�y2�^a(�����L9�q*��J3Rh�5��/N��(��<E���:��M���Ԫ,c<\����-�!��B?��+��Ae��E���_%����I:r��IV����] �X�(�(�n�|3&B9S,�S��1lOF 0G�"{�6(r֥��Jhz���2ţT VG�M�Ė ��?�'NE:����� 4ݦ<���Le�nQ�B0&R�s/�9�@�^���N|WnWu(��#������R�Yg�<����6L0~�#��I~@�Ѡ\�|�d#׾2�@I��dǄ:F�tG�b?�����xd�VU�F�
��^h<遫Ę9~B�s��T8<�D�cM��J����<4,B9����?�>1�����O�)�re�w@`hR5C�$Lv�] ��'�����ƧJ����p$�&U�X�V��w�=�1i����D�E��|��I�O���d߮@��hq�I-I�:U��f�3\�'�y��/M�d��̛�)Ɯ=�EIQ�H�ܨ�O�z�M

Xlȹ0@ǬH���'�Z�SÆ�$E8J�d�%F<�#L�91e��¤B� B��pZ�$�c�%�IZ$E(ӛw�P��ѭf��Eh�+��$
ԙ!�')N�pC��F{���S�]Y��3D�7�<hI$ǟ9��M�1��9K��QHC�Es��H���ӹޡaď2-��=�V�*O``�&��ϤzWě.�b���V�$�����'��|(��#�n�Y5�B+@	��+F���p�K'd�c ��:J�'ʨ9
��F4x2`�(���jI��[�a	nD�����|ʳeC�je�� (�6<|q�ԡ�@�<1�&���ł'�����c���8d漋�J�~_���Q�
�'�ȹkp��9����7�\=���K�m���1�
�1A�![�kt6<e�0�Bzx�`����p�P�������(R��R𪐀\-�M� ߼vxq
�W�[ ����� (��K�'Ч-rO����ߍ;�v��Gm��&�)��ɲ.��Ӱlߌ9�|��7m̨#��R��3	ĤC9�08��O>@`�`��47��/z���!3|���i�z�����-:�����ú
�x�ȇ�M-�ȊӮ���0��@5o�f��TB/?� �˱L;	�l�f���'���$ո��Żv��`I؏��?Q��x	��a�@	���@��!�j��g@�2#�� @��'�r��� 6
��X�jϱ��!�;)�Ҥ���E3��A�@�6x� ��	u
�y��k-�¸���/�,�2�AB�$+�m�˦�ृ�_(0���`-�AA#��\<6�	p偀 ���b�>��J&/�"�Q�J� ��ikF�A�lΠ���r&QA��N#V,ba�ڱ/��Q�eҢw��"��`���-#�\*� 
�0j<@���{ip�.:*�G~����mJ��e��B���:�` '�a�P���W��`���Pd)��	g^��@e]�A��5@��#�Q��#�tЪ���_�b?�@�,A2<�i7�ZL��0JD�Z�4�iprE�fΐ]����"GM��)�͐�&U\P16��l��D[0�
i`�eaĄy��Ip�����}��@X��&��i:���԰=i�D��N/FY�GJ�&����0$޹�-Xc#L�l�����O�N��3QH��75�D���
y���`�^8��#M�h����'��á̗�O��݃ i|	�pM[�B H�C�Ѹg6��C�1x*��a�:k�#�c;�xa��)S�O�ڴ#�D.�t��W�~�&	��N�8d���x������O>9��"�5羈RQ��/ְ�;�dӲz#�9�.�+�|�2�ۺI2!���6ᴜr��,ޤ�S $�0 P�XĂ΂w-���̙�$od� �C�	F)� p�[��rMˋ_S �b�c\��2��n)Դ����ì"5�Q��(C�_�$���J�_Q:�""#�Ղ�C�3RD�����I��Ć,�����F&`�a{�ŗ^���\�����(�o��06J[-�t`B1CҳP����V��d��ͨ��&2*9�+Z	l��v��/�~tbq�3�~��4+� �i��{�)��h����'9���h��lBz�$S�!�hJ�#�?��ɢVa�ոmJ�@ACJqɓ���wx���ڷO,�h�(�++p"H����O� ����0I�`2BAK�b�A�$(�]AD$'���`EO���ޔ1K�h:R�� n�Td�*ze��i׉"�ؼ���٤�h��c��r���� K����&�?!�M�&�Z�t�p��o�zg��S"Xnt�%sW�H����7f�>#�U��4d�B�̻A�yt��iV���O[9U�|��}�̹�C����H�D	{�mp߬̕ö��J���g�7�������P�IA��<�U�ݪ�@���e[�%��@�j�'�R��eBݫ�H���EP̧(����eUO��]q�H�5?���3��t�l��G&�� �0O�$�Gm��B�ލ����C��$05�'�$0D�HL�O1�`]YP
�%�����L^$qZz�P���9��
Q	���xR+	�@��)�GN �=�H����\��L*���O��C�4�~�$�|Ė��=�]�@8}"��C<=�@�Ԇ� 4�`C�35�dJ׎�-%�h�!p�D��(��&v�6�z��'���c�
ӣlm:�)�ɉP=�q�wOZ���(���(��)x�r��g��[����4D�p�VGٙg/��8V@#�E*�N0J��5�V-.�;Pn���8�ȸ���8s@�I�ȓ>x��`ꑪ2��ca
՚�����=��"~ΓFr��"e�ݚr���clN�6L��:޴��+�=�2-�bL��A�)͓����Sm3�O�|�)�1��4r���rb5��'�]��P�(��DH�vj�jƤ��^���p-4D�̫gě�(j]��OY��h[#I!D��0�GE$y�|q�a�˙4�ԓ6A(D����I J���8��	�F`���-D���pf�j��T,J9j�F�F�4D�DD/ӆa�h`�C'J�p���V�3D�,j��T&s�V��§=X��}b�*+D�4�A)ڔ@�Te�v�ݦ}K����'*D���a�jƌ@�&�2�@@���,D��*�VfT��LS��2���,D� �Q�ד~#��C�r�U�h$D���$�	0x����ƄɅR�f���d$D������c�bx����R�n�(��0D�4ѣ#Ƞ-FQ�$�JE����C2D��9�Ά%�4��p$�&p���,D��6朤"
`3�MZ�	s�ZÊ+D�XPM1\^,Y�yE�	��V��y�`�	a��4{T@5InX���!�yB��3���s�����0&ߜ�y�E{߆��F��j*0��a\�y�鎫�F;�R�xRDi�o^��yB���8~�(��Q),*�*f���yc�
y.���q�C�*��8�B���y���s��#�̞N�iZ���y�?<tl���I�L	L�Х�G��y�-ʅz ���,�
���*5��y��ڕ'T�h��ӡ�Ҵ�j��y��
Jˆm�CC��p��U��kܙ�y"�$og�B�&ܾv��sS�^��y�bD�&�B��ML^�6���ђ�y���)��Q0)Z"TҪ@�q�S��y����:���2P�1;y ��6��y���zƺ����;2�*q�5�y��9?uP<�#�@�(�(��Pi��y�k9%�.��'H�_�t��f��y�J��k�h���a��U��Tn�y�/w�,�[1L�?M�1�����yR�J?��{�V8|���P��!�y���-1b�3�EY`mƉ��\*�y¡[�Bq�Q��i@5f7�L�4'F<�y�@��bH��N�'[zl4De��yr�� f� ]& ��y"DV�x�2�3��(V �����M��y"���N����ę�J�!)B)D0�y
� r@�S�#��P	���,X D�@b"O�ɰ�f�	x����I�)�u�"O�9���Γ{;�1��ň�f��!"O���Ć̡W�D��E��z�J-�b"O�p%�ƳD�&�P���qD����"O���#�ޒfn��G�
\-�JQ"OF��#EQ�80�J�)c�>��"O�\a�l�v�Z�b��. Fe�"O�����;p���䂩B�f�F"O��1�� !L�}6��'R��!��"O�XX�Ɗ}14�"��K(E�"B�"OP�G��!5�����̸d���"O�⤫�?4{x0r�� @`� �"O1�GIg�����Q�WO4��"Om�&�	G�P�eB�$챃�"O ���W�4�F}C��S��U�"O��*���cu�D"�)6�N�#�"O�A��B�TsN��Q��1�x���"O(��* $X���{�4a*�ш�"OLIèL�W�t���0{����"O��j����m�4@+2c	�.X�Y� "O�X[#�v��y3�C��I���;"O��(v�E%_��}�e@�(�TD��"O�=��@�J?� �!���"O�!�ë�:bg�IIV��K��4p�"O�	R�f�-;�@�5mZvNE"O� �'�$ӄ,:�쀀U6a�Q"OB����x�y�ՋE�ET���g"Oݪ�fX_�N,Y /�;c5���c"Ot(%�_�k|��{!G�G� �he"O0!8v�׬2���je��9h��7"O����Y�8	��K6�#0��9Y�"O��R���B�̨�`@V6?�F�ʖ"ORI�C�҃ulZmȆO�t���b$"O���#�Z�Kv��u��"O�XRrB\�x��������l	��"OjU�AS�W��(��R#�&dk�"O�	���1=��MR�g�j�$���"O:��5�ؚ2ò䂷��$3�>� �"O����+#4�����π	�b5��"O-��:9l YRe>e��E"O$QS"���V�*�"4��̜��s"O�H1��(c|R�	� Μ<�S�"ON�[Ѓ�:$�6���͡�(�;R"O�`:�[�T"�`�DcU� ��@�"O����RM��(�c�9c����"O���>;��j7���̑"Ob�qӈ�
J��y���G�fd�"O��h�aJ�N�0��GX���YB�"Op��d�B��89�SI�5֕3"O��-��m����pͪ9( |�"O�A��ʍ������ôT����"Oȴ˷IF�l������B�j`�z3"O��� Λ��P���đd9y"O� p���L���F̘%~���k�"O4�0��_%I�x��N���� ��"O�����D�D�Y0}3�=��"O
�A@�Ҫs��30��W ��r"O 쁷&����*��<D��"O�;KY�{q��H�);@��"O���7�͘I���@'�7��)�"OyʷE���](�'Q1?��P�"O�x���'{ϊ萔'@/7�X�"O�@r�ɘ�q���}�v(�"O� �M����0�u�ȒXҒ��"O�\r�D�J��LKg�Ov�-�u"O�}�b���7ܪ���S�[I�t��"O$�#1�Q.rV�*���g&l��f"O�m��"�+�iPRC�05�X�"OH����^؄�ӂ�J�z�pt�V*O���AIQ��� 0ƈz� \(�'=6D�b��y�4А ȏ#{1`U�'$��x���]� ! A�M-�pe �'�P�R�^���� �Q��e!�'�L)$*d��,�G$�*��z
�'LH!��Q�����G�->�	�'�%�b�Dn��	�]1JL	�'u2�I��U��J}+�*�/^�`	�'m\}����Y�$i�&��>��'
�QQ��y��t �&	p�n���'QZ����5l0h(�f��b�'}����+�<N���;�%�L�0�P�<rƃ���� E�E�`!D�Jx�<����;z/�������I
�*�)[z�<���_��%L�8P����O^�<a7	֌?���\�G �bӧY�<q�IZ9<t,�RhǳBb���P�<���F�Bɰ���9���!&�V�<�և��w��pI����gE�W�<����'3�^�	'��/M`�w��L�<��d�$`QT�Ya� qR����D�<�*ٹaM�M�c-^,���xTI�N�<1�.0����AN�'��	p �B�<�@ĀZ��0�e�G�u��#0�}�<I�i��)Ȏ	�M�u��p�$k�v�<)q�>J��B�ܮ}��e�q�<���p��t�B�E� �����U�<QgM�i���'�H 27,U�GeP�<�ɿOR� q�"]�d�A1�v�<�f���{LQ�Թ3��Vh�<�f��F�ڦ��<MjD �@e�e�<�� �4e���8M�~!����h�<��'X�nK~	!$f�1NIdx��F�@�<IPǕ�X�������8�Zݸ��x�<�u�މu�$0�IQ�!^:��gǆt�<3��7gFH$a�'M�Y�d��l�<A�-]�v�d����'4h  �m�<��cՐTM̨�jҙ`CH�S��P�<q$n��@�T�� J��-/�`�@cL�<�AC;u�����/׺UGCp�<i����a�r�-y.)s��h�<q�O��P8>9�d��~�ȺPJGe�<��4uώi	��&��eKU]�<0��s��%�h�ZHY�<�p�	Su��P%.#.���'W�<g�Ǉ"nv19�>l���AS�<�ŭ̖'��1�sKD!�|���JI�<y$M�Ѩ�#)�8Sb6�p�̗~�<I��3G�uh;d��(*a#Tr�<HF�y0�� V���+���цLs�<�b�M�8��ֿ[�z�i �j�<	2CW',zι�<����Cg�<��׆G�Щ d�Ȓp�����V�<Q'�*m ����ߌs��i�$�Q�<ITm�L�l�e�[�R��+f-�Z�<�Ԇ\�:|r�����P��W�<A��ݐ(`�T�d,N5���Q�<�AQ���y�
��Z�"��N�<� ����aڣ%`j%z��ZE���@V"Onaz�A>4�<�h�ǌ`m"OL#A��&}AJ�BAE�v���"O�u ��N�"Y�}A0 �1%+`a��"O� �q�^�>�ӑNB�
0���"O��NCE؊���X!b%9�P"O2͢c�X�g0�\3�D���
�2"O�H3H]TX�EA�u�\9�"O���i-���x� ӱ/괼��"O��Ӡ*^�?�l\��/�8o1�8�"O&�
��aI���$�/6~��F"O쵪Tc�m��
u�� R'~���"Oj�x2�.c����ӆ�H/RIg"On]*�ŝ81 )%�Z�a1A"O��᪋!~����あ5�Le�"O`�	������I#���z�"On�`6/ɤd}P�x������!;�"O��i �)q <]xEhT�n�%"O���%d�
�n���.���}"O�l�f�Y';� ��,�P�d�0#"O0��7c՛pf��7���%���"O��R���T}�BfؑJ���Y�"Ot��d	ω.�P�q2x����"OZq"�f*	�Z�R'��#���z�"O�Eq�	ˠ'�dM��H�=�<	��"O&$B��Z' M�a;�lR���s"O��iU�X�e�A�J^v�>�s3"O�qe�]>< ��ĊD���b�"O�� ���1;&��!�*��k�$�2�"O�ȸ�C�<2蔘���P�x�ԭ��"OT�����1~4}`�υ�5��\K0"Oޠ&훯YT1 �i��~���2"OP!��(������,2���("OXm����f8R����&�&e� "O
 ;�@�0
��S ѝ%�vIpg"Ox���(�a-���Na�*�3R"O8 �5D�"�! �b�!U��"O��A�� �J�2aX�@ �7"O�0{�iE�7e���t`�$s�t�b&"O6���뇲@?b�	%��6��eؤ"O���6Cߣ~��ت6���p@Ӓ"O�0�m�� TSw�t��\�B"Ot���B�y�4	G�䕓s"OJ`hd��#3�9  �Q;=�li0�"O�9�1�_�|~���gF�0�؊�"O"�y�N֮ ����&3$,x�"O`�zbk�=K��� �F�g�,��"O�rGc^'*����ǟ
�6�y�"O������%'���I(Z0lb�"O�T�(C%t���ad,~�ppu"O���	3PHQ3&�_	)k�Y��"O0	��67�@ �Kֽ}]z�F"Ol�B#b���頄�53��X�"OR�BE4ry���cY�5�M2�"O:��&Z�1�`T����MK:!�'"O-��f0���a� %�B);"O��	вO�(,��B�)��ś�"Oe��R09o��넠�V����%"O�I�&�@�d��q������Qp"O�q+���t@����Jp*1"OH@�+O�i�h�Z��
�-�p�a "O� (ܽU<}K��C�N}�� "O�9������ n�/�:����b�<��T�t�v-�&G\n��-��� `�<� xX ��5Z 6Q���#{�tqD"O <�1E��wa��2p�G�Ljl5"OVܢ%��lL�3eŃt��%��"O�Ti��� ���9��P��蘷"O�9yb)��<ȸ��h�3$�Lӓ"Oz���G1,��is51?�Q(s"OܕǢ�6.�}��Ȓ�$��
�"OH0�2��Mh6)�*؃i��a"O�����}
�xJh�!
�d� "O��9�6��Q�Ǖ�8�Ա�"O�� 6k٦<�#��W�i�ڄ�V"O$@�^v<�aGY�l��2�"O��g�:b���c�.��͋�"O"�Zb)[M�\��M)a���A"O�2��=�zU�a�S65z	�P"O�idf�E�u��u�x=�`"O�D�@J�1=v�T����X�����"OX�����MN��I�W�@��$І"O&q�a�9>���2D�4*�ق�"Oș@�c�7'J|�j�ťz��l��"OZ�b�`�!i��Y+	��M�d"Oh�H��_;x<кWͷdT1��"O�yP2j�K׎A CL *�0�"O� AA�4w�M2q�
1E\A�"O����K�c�����wŵ�t�e�<q&@ hmz4L�<Ŏ�`*a�<�/�=of�;��	+��Љ�f�@�<����<O��RA�[
�z����W�<��	�c\�l�6�ؘv�V!U�x�<I�G#D]����X]3^����n�<ѣ��L��@!�i�O�4P��m�s�<YV��2�ND!�D@�+�Y�3eWi�<���6h�6Ų�o9cj�Pb��f�<���Պ�z C�&�r��r�C\�<��*#�P�š+�$����\�<�`�Y�:�+EҫT4:�d�W|�<�)[�g8��YR���o�z���'Wc�<��͔������T>,���K�@]�<�	G9G�ٓ�M]8֤32lX�<��B�-f�,�t#S;���6KW�<I��?W�<�tIOF�9�	�Q�<1��`���N�2x�Θ!"'�O�<���LHh��eB�o�`X�DSG�<i�B��g>����g)*�Z|�!���<�S'l���C��I+y���	�	�n�<����=�p����A�MA|���n�n�<��D�Ia5�B�&F@������s�<�Aݱ�q�*�&v嬑��΃P�<���#mL々�"EN�Q��l�Q�<��JH�!&8}b�f&>r.�Dn�V�<ф�y�A�D� 6�T|i�.P�<	�N�nC�|X�@���X��VM�<y`�O @Q��1c�� _�hRs�<G�YQR0ٔ�_�R(��`�ij�<6C��,��Թ�H���6�P�!f�<��
�'R�H|C�C��f��)[�E�^�<biM2 ��<��K���ڂE�Z�<�a*Y���� `����H���Y�<��N��h��K'.��)��ʘr�'� l����� �lI
�8Z,Or� (�)�'c�(���דі9��'I�&���;v�hP|9�M٣y�J�x>Q��E2E��EK��N�&_�\b`bZ�~X [�i4�?a⅍�'���i�,"�^9(��A�/\���2���M�d�*��ßp�҅
-�8��D�O��@P��7έ�� �q�.ɻ�O�O
�pC��:�)���<�0|�휞;t,��@��q��TȚ�A���S�½?��7 �1K��&�ӵ��� ��
 ���H�t�쐲vY�ۃ�o�P��|��03��E��dF�  �&B���тd#�=�7D��� �a� ԫ`�)@&��}BFQ -0������ C$�{��ݜQ�4�KR)I�ldX!d�<w����n�8$�a�40kА-JE��M�L0�C$�.b��-�"T5�,ؤ�D3<E U�
çY�D��#�A�^����I�0і��oԈ>� ���!)�@ My��?�Bu�kizh�-�*%�ȓ��K�T�ĸ��6߰�Z½i��t���N~����ʇ�<�Ӣ��d��)��Q�.,�xp �icX0��W�|n:ҧ\�,���~t\����g��u�?����?�0<Iԧ��K�������P��OUr�<)�c�5N0t��nB�.�$���Ηi�<9 �Ԕ�`�Åjz(����Y�<�S �)AK�AI�jX�e�T����V�<��ƜM˄%A1Ɖ^E�����i�<��c�sx��f�Gu] ���̞P�<�6"�!��X!
���I�<!U	 6,�#���g��:u��E�<I lQ8����@�a�t8r�A�~�<Q���P�tɃ�_.d���LQq�<�Îy5�(�
��a������U�<�c	�$1�-��e3 ��(ȥjAP�<)�N��CaNP�I,7�bxX���g�<!�'��Z�F�yr/&�L%H�`�<���&R��Z�#��=l�U©`�<��b�5$����K#(��u�ht�<�"��U�5�W���XJ�lE�<a��~��2�
E�aߒP���X�<� , 4g��8��V=4����MSl�<�A��,HU��@��:%��K�f�<i�ɩ��D�ѧ�*����Y�<I��{��=%���`��q�<YF54]�u�6L�89��!�@�w�<��K�,%����7&M�`e⡚fbOl�<��F�3Ut��a�,�vE~(z�͎g�<y �&F�u	s@�� ^4����`�<��M��T��xt@��a׺M��!Td�<a6��&(�6��%�Z�2%i燃Y�<q�/�T�Ȑ��Z�i	����_R�<1&�J		0ԛQ�A�%�P�A�K�<	���61
M�¬G�;���q��H�<IƈV�m� �G�̢mTJu��JG�<��Bºh[@�R7{Jt��F�<�v��+d�J�Bδ&����V*D�<�Ĩ�^%�)I�%]��i�B�<���׊x�l0Y�oR�A�n=���B�<q	
�h�l�B��_�&ʬX�! }�<�3mT�sA�\<
r��y�<Y�H��R���
8_�.� %��r�<�rd�9e�F5p��ʉ/ƈՈ��^k�<����3O���SE�v�ұ.Hg�<!EB˃����&��4��ق@��n�<A��+C+ȕ9��_�E��6�m�<�u��1qX��C�N	��z�ESP�<Y ��rb����T���K�<��L�N�&p*D�Ѭ�(�bkE�<�\�+ˎ!V�
%���h�!�dBr�ޝ�b�3:D�%�s��q�!�Ban#�&G����bI$;�!�DL�C��ӂ�('~`�r�D2k<!��1�tP���6����z!�67m�u��y�BH㲡��0!��EE��"�H�&��7o�Y�!�d��)!8�tF;��Q��M�0�!��T�����H(��P�Q>h�!�$�/�p��� j�l��@$J�_�!�� �xk0 �Bޘ��*��[Cr�!�"O ��;�<�ҕ��<ʵr�"O�S�.!n��ԃt�ρ@8���$"O�5������B%@E5T1�,�	�'���ۺ���G`͊ej<���'��
�B�><�"	��/
*bv@i�'��s"�7�м"�3�­�
�'���*`/�-\k���� 'KHDz�'1��Á�$u*5	�#'!(P!Y�'���aܭ}q@ع���� ⌽8�'%@��r&��9�����Z	ָy���y��P�}��;2����YPhA<�y�f� P����A� ����*�yr�J�(��I�E�,�� R@�Ҽ�y�.Ŕ���6D�)ZV����@/�yRfD�b3����.s|�8$ �0�y����13�@R�N!"`zd���y��F
k��␯� �����y�BD�_����ʇ��r=HP,K�y�՞U��a{F��t6RP1�M��y�!�1l�C�(x��ܑ�)G�i !�ă�4k��
X�<� d�W�2!���3"�!���P��=��.��rg!��W<��1�$��b���PpB%I!�� �J���gǦT�B��G '*!���88���2ǃ�:Mz5���2,!�$\�e1�O��i�a�&�Ɠp!���;�`1UE5T��)���^�!��R�&���9Aza2�K��D�!��_�>�r-s��<(��`�k� M�!�D�i�䡋](`BW$$��$"Or5�%�y�P�[��@�u�a�*O�< ��P�r0r�����i��'+�D��U�LB�1��D�-�*S�'#J��r�\�P|�,�CG	w�"Y��'L�q��mDY��@�*��Պ�"�'g�$�BaO/9h��K�
)��ѱ
�'^����c��E���B60ޑc	�'�<5I&�_�P��%p�!Q%+	�'�f]�m	 "��`��BO��t�'��1P�ē3d�����aɞ 0b���'� E�S�d�ൺ�M�Eb�ț
�'�\��&�ڀa�,��?��$;	�'��\adL]>T	yc��8ô���'��I���-x���#Cc*��Z�'$���L�&r�|aRG	�0:0��'9r�a���"�X��&��$i�'�����/��	 at��B���h�'
��Y���?g�8���.٬k�9r�'3`������b���鄌�M��	[�'b�qcU�׸f��J1�A���*�'1���X�~��0U�d�I�'. y�`Aڒ �I����H0D�'�v����*���&����2�'sД�0�<��<�ckû"5����'Έ��g$��/@\d3,ھ��q��'����Ç)
,tɑ�'O��R�H�'�V�sT�)r*erD��8����'
�D���?��8�b��(�|L3�'�����W7	�B���lh���'��=��A��f�����$7�-�'7z]�d*�-ꜼÓA\+Hi|�	�'���CD!����A��M�l�	�'t���¬�^R��͜ ���	��� P`�@-��fly7��#�*y2d"O��� jE��Ԩsp���>�l��"O(9�rnU�8���P�Ú
[���i�"OT�b',ݵ6z�<��ѩ.�ha�"O�����>)�������-�����"O��{qFR%~��+�c9�6�1"OZ�Yש\�&`*`�Ƨ/05�"�7D��B�ᓔ~�j�"�fq�;&*!D�����N )ީ��fex��`M$D�< T��I��i�ةWf:
��?D�<r�b0C���nַi�^���;D�0+C	�+�x!�)� w�zrƎ<D��ZU��x���j�y�f��&%D�0x�D[2`��Pc���bA<m��$%D���&�3���\6&(D\�#�0D�����8C�|u�q�Vh�f*Ox`RW)�8[���Q�ƅ!2��"O̬�@у~���2'�*=Zՙ�"O�d�͈'L�J���%��|Y��"OұC!�ڱMۘ���Y�9_��"Od�{�@g�hL��M�M]UPg"OJ�	&A�U,��"c�\<��H�c"OЉ�2�2z��|KV��;|�Ȣ�"O䭻��6v�M��JY�)<8�%"O��3o^�{z��Am����"O�<�Un9P�}��K-nؓ"O�M8���^9�e�@�f�МP"O�SM˨H<��@�@�5�N��3"ON}�b��n��I0�Ə*Â��b"O�3U(ݏx�ܵk��V�Z�xLS"O��;a�/�ґPG"ĨI�� �G"Oh��qBD�o+ĕ����0�!�"O�1;�j0�VD��`F�z��a`�"O�xG�E-D���)yv]`"O��i��
D�j#���2Z@^��"O��FM�.�6��W�c.��""O�9�VE�.������cz�%�C"O>�φ�bA��K�f��6e�(c�"O�iRF�=���]��衶"O��W�'VU�����i�(8"O�|�7#̰q�`  �ϊwtN1pt"Ođ+5� Q
�S��TZp�s"O��[��=[�|!!�F�+Cl�;P"O��s�N(q�s��}���P"OZ�;Â�o��I�@�Q��L#�"O"I��%J�������g����"O��8�K�3�taz$��:�2�#F"O�䮇d����փb�!���9�y<'M.�	�C������$ԫ�y���$Z�.p�v/�vu�4��O���y���C��+fH�y�t�A&T�yI�|� �u��&y�4T9��	%�yr�e�,�m����B�y2*_G�Q�tb�6^�����yBc�7$���1O���Ī���yMߡy�����`ܗ�2(��)N�yr��Z	�p�&Մ���c����y�
(*��|r�+U�v@%���@��y���,�&pPwO$u�x�R����y�N��'�����M�$}���ӐC��y�E:db�:tͲ���K.�y#��x��u�fK$�43m7�y�%�O��!jQBݷ��]���ە�y���{��z���1:�#���y
� �*��$V�|a��)�![`"O4l{� wʔ�r��փV�dh��"O���@Íl�ъE�Oކy��"OF ;�O�/�̤��ϝN΂��d"Oȵ��a 0�̌�OM(|���"O��b��:|t�!c�T;)��\b"O4���/��s�H5�`n��'�Z9+'"OTTr˘����Iu��$p��i�"Od��1�
kq"� D�+B�6�;u"O���4J�:�̥�ӂE�A�=;b"O��­H�|X t!u!\���p؄"O�mi@R�	��b��Đ7|%�P"O�-#�P.{b��
A���t�:e��"O��P��Y	���s�N�8RƱ�c"O�Er!c�*GGF܈7�1�*t��"O�q��	D�(���:]s>��"O�-�ь�[p=)lQ7&���"OB�'�L &^�S� #A�x8h�"O��S �@|�2αt� �G"Op$a���?Q��
D6}J`+�"O� �D.4|� a` ��Ii2"O�q��ÝT5�Ѭ�@R09�"Oա��ҾhP��K�>[\b(��'u��{  ���     �  �#  �.  :  HE  CQ  *\  c  �i  %q  :x  !�  ��  �  5�  |�  ��  �  ~�  ��  �  G�  ��  ��  �  S�  ��  ��  �  b�  ��  � �  Y � �% D, �2 M: �@ �F (M �S �Z �` 4g Cp  `� u�	����Zv)A�'ld\�0"Jz+�D�/g�2T����OĴ�7Bڭ�?Y����?�`�҅w+�ؘw�[�r���f�;BX8��D:QgH�kD�Y|$�Y䀝���<<�8��7���S�@�9oM�~=����� *�"]��arjJ �B��p-�-V�l$�_wj:�C�O�26M��i^-p@)�,4,�ȰUB��:�4-�+�^�-�4�տ$��5S��L�nE�!�ݴ�?���?9��?��EA�]
��E�@_�	A���Uz���?1v�i�2V�����/
��؟��	4��\⥠����4���R�z���Iş���ҟ�����X�I`~<��N��w/ǡ<v��G�M�@�~Q���"Y?r�i2'Gk}����!�'�j�'�N�jTc�-*
�,P��&E`j�j��Z�>���<�I>Y�'��ц�Б[0��'v� ��D��=(���֠��b�ON�$�O����O��oZğL��_�$;�$�dA�Du��h��9BM[6�'�V7�����;޴,����M�a��W盦��f�� %�� �p@�e_4CbQ`�J*b�x��?Y(O����Z)���F�Jn7����ם���x��̂!]j�Թ�K���{�H��t�|2sf^�%�`����I��4��O4�Դ�l��D!�6���`��e�)��``�>���D̦N?�����3*��	(&�Y�iB$h�#����{޴}��a�	^�hK�h�& bu����Eh�"�T�PGbӾ�mڙ�M���{��Uh1!�w�� @Y,
�^e��I�*.^��'�X0����V�*�ځi��+�fjx�h�nZ�N�t`1l�0	6���/�_�2� ,�W�ؙ�C�U.kKj�8�m��Mk�E8CzZ��bM�F���  	)�?1���!8-�I� �>`U�l���qr����O����O��m�џ$�I�"u>)���0n�H�ug�g"����֟��H�ǟ$�	՟ )��1��� 7��Q"� �A�P�δ��/h�@�gW?A?n� �@�Ԣ<aci�4(����&w?.�	�m�U����2�]�UZ�KT�ƅ!�"Hx�����<��KYy�B�<q����EU�� tcU$X:L�Pg������	���&� ��͟(�'�⬕��6�:A�
b�,�"�y�2�'hU���=R'�'������A�O� 8(�nJvB�a� (�"�'��ɿ>�"�(ش�?����?��'""�h���F��T��˓�2`�U�b�4
���?� &2b%<��C��2*� ���ޕ7W�������I�� �ĥɷ�:��1C$'7��UH��B��a'�x�B�����+T���M��dyyTj�$����ݼE�Iyv��D!�c�O��o�/�H���t��aF�!.�[%�/ؒO���O���O2#|�W�N��H�W��9/��%`A��W�'=7mO���ϓ�M��O����D�h\�A0'�A�>l ��i��T�4k�	��?Y�	ҟ�	wy�����J�Q�@ڼ�����h]J�+	�zt��*���*��W>���6F�����涟� ,��o���*�Z�PƬe!�@��B���铵5�F�3��b>B�*V�5i��ʬ\3�U ��F��j�;���8:�6m�cyc�9�?1�'���|2�ɲk��`D(�a��뱂ɒB��)�@uK�@ڵ�C���;�Ȭb�j������M�U�i�ɧ�4�O<�I.B?ޡ�V6�@�����ų埤R�rA���$�I���B^wA��'��NE�
M�$�>L&� dC��h�8@�'(~�|lS6�{S�)�i�/|������$��s���QT�߇����怀�.�LyZ"Yb�0��r��\m଒���uU@9P���TU���XeH��mc��M++ѐ���'6�7�i�'��4�7cW�|u��$�gb�͡��<��,R�!I�%�5�'/�7��%��ߴ`H��_�� d���M��?I�b��{4�%K!g�o���ȝ(�?9��F������?I�{x�RwÔ�%O�$R�4A������ i�c/?k��p�.-���,]�(OHQiS��Y�V̨��7
A<����)^D,&�ײ
���{䏟�Q$F8��G�Rʒ��L%��R���e�\mZɟ�Y�j��8 ^���f�LA���U�py�i�D�D0��O�q�X11S�¢ �6<��K��E�| ��:���Od�'	���/7w����Ce��<�ԏ\�F �7��O��n��B�x9c����#"��'���|���
ch��jV���Rߔ�D�̜*P2�d�O�!��:�@}P�B"��$d�	�}R���h����n�*ʠ�Ȣ�T����T�m<\�rCW�~n�e ��#��C$��+YtEӷ����LA%&X�怂�n�%T< 9 ����G�O�Ln�ħ��O���H��x���gj��^�,�9N>y���䓅?Q���$�>W�=b��� 3D��Pj����G~��O6�O��m����d��ݞ$9A@W�W��v����M����?��bo҅�t�?y���?����y���`(��E�Y�Ao`�5.ׅO��1!5߄jS��j�{��٣�_>�����N3�I����	%K�L1�!�> ��0F�T(` �Ay�$��gt�Hc��xӞU�範����6���
U=�Z)���]�Z@Z�a���I�0���w�~1�'�TM���ܘ�?����?9��J�h�H	���m�0@�Ę
���0>�S�Jj9j�0D��nh<щ�CƟ|�I��M�ǽi}�'��t�O7�I�9'�̢̛��|{���&Tf�k!�B�F�=�	��(�	���[w���'j��O42�:����14z���.V,>���SC�G��IQ�$������W��x
��DD�I���ac�_�x&0�s��D"a�3��
I4��%���
���3���1�)ʓ� �+>y㐬"�V�y�@�{pj]�p����p�?y��IL�TV�D�@�;J6�[���!��I���V���o�<e�G�:R��'V�6-�O��x�\��it�'-�؋' 0�~ȁ��G�T�4���'a�)C�.���'�gH:�2�3��,c�4��u�=,� �|`�5:�Jqٷg��m�j�!c��VUr�҈�ď5;�
9�T��_�a"��dub4 ����0�{uN��C��T������ {`�+c�Z�O,{��'a\6�Wy� �2!N�����%c^�Y�P�����3�S.�VY��G�:[�a�Fi��Oi��D{�O�6��)�v ��L�0A��tbpLRzh6��<q��W�la��'�R]>m�p�ݟ�+@�Ż1x��8�e�-M�Vށ`p��':��x�Cˈ!}��8T ��H��D�+f�h �?���Q:�AJǫ<dc��s7	.?�fZx����ZV^�����I�z���t�!�d�E�j5Leq4� ��G��9���G��"��:Pvq�%I�â�Kd���B�ɘQ��=��D � g���*دs~�?� � ( ���E�2�N����M�`lZC��,1���ßl��񟈖'��i�H�qH�������,s���l.`\�ķc�����N2@�S�?��`�����	�� �#�Dǃw��"�K�v�i��&Qi��Q�l��f?�Q$,�6��H�OX5�f\��yw+�0T%����N�Sp�pC�,j���C�<����؟��Sl�L>AUǐ.M���㲂!P-Xܮ�?����$�O��?��'Qԑ��jյ��a���.�U���?Aa�i��7��Ob�m�W�4�O��B}6ibŊ?;g=�$܀Q$������M���?����D�|�O�Hz�_(n��	@f�)�^<S��+3熍���G&�0��..��=���Us�'܊��7�N��A���� Q��ƀ#R��FL%~�qҩr���2�^�� �|bb�XL~L�䄖�
rU��D�q�����:M�F%-ғ�O8MP��Ɣ��Ҵm��Ւ\�`�'��y��Dº}Pʤ�₡)T�e��N�O&�'��7��ަ�'/z�iS�}Ӑ�d�O�xzp��-.�2�T��nPV�+��O���ϩ}�$���O2��Y��4��&i��\<��#0�n��چ�	�y
��|⤊� O0<�)ދ%��9�`!U�R�7�Xi@��Ș6�r�I��4?j�b�mٟ͈O���'f<7OYy��P4	r�$�}���������0>I�jDx��!�DB3BH.}���ty��'��6��&��� 	��E���B�ɇ�ruo�EyO\kR<6m�Ob�d�|��&%�?!�뚫T�a3QF�)u:���A����?I�"�-s�����>��q��Ȳ�3,L�P�@Jg~�$�O>}i�*�OI
9��fXk��9:��1?Iv�M��L>E���8�XȲ��`�Y�ҳ�y��J�}a�Gʌ`d��O��x���8�F���7iJ��(��o�5��Ɋ?�Ms���?	��Q���1T��<���?���y���Q,��3�)�q�w�ݦM���Sc�ܘA��BWL�0m�/���i�P�I�*�ܜS�f�1w�r����ݵs��T��hâWv�B��ɂ��-K��!擘2��'��`��o	��"ADR��z��U�i$��!��`���?����v����@��Q~�K�O�x��Ґ� D{����>2�����$�ʕ#�*����A�ݴ�?A�iw�S�?��O���.�}��!z��;?� C�,;^�P듞?�����D�|��O�%ۤ�ÇL�t�4̑$7�0�"�a�-w��ɕ.����H1�eᚦwk>�<qe@M��J���c4X񤏊�->�[�jM�"���h3DΌ�b�p���!!�
�<!� �slz`�U(�E,�AH�j�V}�A�	��MӖ�	p�S�xmq�EP�W�'+V���K��?	���hO�c� ��G$E�<�D4���0�/�D���ݴ���Ra٨��O�����_�B�@7)��2����߃g���$�O�ʀ��O���`>�9�/��5�u�E�S�H�:np��Jcd��.=�ŀƥRՒ��2(Q�4JC䒡]��։f�����ڠ�@	 �!����1�a#�v�"�;ÉښgrQ��Y&��O�|'����%�,׊)���F���a"D���$\4K��QǁR �ó�-�A���I�ҟ����Nm�d��t�=��,��ǔ<D�9oZ�	K���'v���� �I/���GÏ[��}�@�'l���M4@��?�n�����sI�L��`����M'i0����l�<d�2١���:L��P�L����WR�sg*
.,�tU�d*U��.�O��NXqE��o@�;~�+�O&4���'�>6�Sc�O��I�|ny*u�����"H�#��'���'�B� %zI"S�s�~�Ð�V�v?��F{��'B7�ɦ�'��2rm�(p����h\��fM��� �M���?Q��(�~u;q@��?A���?	���yW���k;���fԾrm�D�a�v��au�R5GS�9��! *�����F9-i�1��]�.��Wk�&ͮ��K�6a��1��/ I�v�AqJD7T��#��՘g��m�,��Y35��`c�zTƝc��7p��̀�+�@�6�Axy�4�?I�����|B%\%_@ �a�۱{x��a�JƏ<D�h@��.w
�����W�Q6��*�O`��e�����'��IL�4蓴H�op� ��0$l��	"��I���	蟈�	ݟ��^w��'��)ޓ"�8H@gT����R���M��uZ��+K�Ј�g���(OFL�q�  4P5�9K���K_~��� r�l��5M��}�z�X&FK�!�ތQ�J1h�*�OЀQԨM	*]r�G�7Ts��`4�Fy}R`w�~�Fz��ɸ`nD�%�΋U2�X���|w����+�I�w�͹V�ƈ5\V�A��S&
���O�0n��Ȕ'�\t㠥�~���L�p`M�+�F��bk׽@��x���?���ļ�?�������h�L+mS,r�>�QP�M],��[^<�>٠�Ҕ>2�k��_�>}Fy�޺.��Y�b�V^r���BY�d�����_�<� ����G9���zĭ��'6&=Ey��?a²i*8�J���"�$]pl�a�fɗ* ��&����	}�@d���kxе���MZ��F{�O�V����<Ά�[GG��iz�B��8A�Y����Zyb�'K�&�4��0iP��I���S�Х�g��=1���ş#7/�L	���a�8\%Z�9"�*d��)�|��#� k  ӵ��($� I���T����%h<,ɫ'@�=e����]�A:��y�,}�Nh�t�K/^n>l���yz�^��x�ɝ�M�7�i&2�~گ�he�ɛ�L�l��c� �b@�E�'���Ɵ(�	^�3�I0o��`$H�3����/��?i��ib�7�O.�n���zeFO1Ujl���^:p�L���N�M{��?Y���ٴM��?y���?!���y��;DƸ��Ѣb���������'��<�	ӓ[�`h����
P�(�3��%^ֹ�<��I���D�6}�36K�39��aH�j�	2;���D*�3扶#��bK �m���*C�I�P�|�`ÂZ�+�~!�Pa�Lb@��'+L"=�'��H���Sٻ��p��0O���م �o�Z�����?i���?C��"�$�O���T�J���� ��*�W^����0ID�H0���Q���y���f}���;IF,ѹ%�8h��@AC&<ΰ�� KDV��̀T±��=:���&�ɜcr��F��$XYP1��2H0��C��O���	2u�����<?+�<�E�M�B�	�:D��m�K�\͐'.�%_�H�O�0o~�52x-i�4�?��0�P �$����m��y�v����?)$,���?�����T,�p¾�ڒ�͋L���Z�KHp��,35hW�l���9��]�yNT��஄*i��Fy�j״^�
mA��=I ��9���7R�xĺ�4k|C`cּ@~�@��K
�!��Ey��?T�|� ����NU~��1�*;�y��pQ���T�D�!2Gʉ���'E��|�'K�("ǋ�2@` � ������J>����˛��'��U>5�U��֟�Ke��L��b�f�=M2�H��Nǟ����5�I��D�S�L��Y�/^�� v��n����"?)�jv���~�;T��;E��ٛ����:���K����7��O�d'�"|�����t�1(*/�~���fB�<!��?&s$E�P�^�U�ƅ��I�'f�}�b�%|��r7+NƆ�;�ه�M����?������WCU�?����?)���y'i	@+⡺���"-"@�
�  ���y�%"|�)�� �>���)�����?=<���O����D75����C�~!jm��œ����&B�KL�AWg��>)Y��`�|RaQ m�&�̻!��� �[�`�(���$cn�L	ڴc����'+t(v�'1��ɟ�q�Κ�O��X A�W�VR�9���� F{���҈y�������{R��Bo�k�����OdDmZ�M�O>�f����+O�A! A�CdF(��F'��%pvȒ,&[f�З��O�d�O���[��?Q��K�r���lӮw-H�փ�5J�9�D�2 �H�r����N\�P���.j(����n�u�'�|պ���(�>l1���3gkyFX^�!ɲ��R8D�rgb�Q$R�i��ҋ��lQ��|ҥ�S�����О�|�v'�%F�R(�[����$��O��"��-lyB��"�W�p|ـ&J%���?��$�k�V!ˣC�7?ȪDa]�L�'�T7S�i�'6fI��l�>1�X~� n� x $���	IB�3��?����?������nV��`�ƍ�{.>���!�+��{-ʗjn��f؅5�ం-�-�|�Dy�.J^eb
\r` �kN�ɦ�ҋәi�,+����4�
pkª�9��%Dy2^�?���i10˓A�
�h��Z�m�.�8@� �%���	�@s�e���/frT��o�v����E{�O�����	\͐0�&�6\�!�̐A^�U��{ю��M����?�/��I���O���N֌�x@�r�[�p^ �#���O����%tŪ��O%�b��V,���qF6G0"�'zy�#��N�J4��Y�� I�d�'Ҷ�J����7�p��a�ÄCP�ePIK�"������u��~��E!�hȈ��A�����BL�O�%�"|R��������g|A�M�<��#�u92,�F�R��{"�t�'��	��HOv�	���)k��`�BL�N'�ɨ4��ݦQ�I̟H�����C��B������8�I�ԅ �𭨵�2��=��%��r}�ՒK��hK4(��x��p���3��M�I�=m6���+/�r���J����ڒ�8)<c!
��Or�Y3�1�o�)� ���HC�
UL��!"W�,=��as�'C��/3Yx���O<�D*�ɢ,Ma�\����F텋M�B��j	$b�$�p!�(�/M
t8�і'�<"=ͧ�?�)O�-1�MНE�|H��IDt��Hqd�)5æ ��o�O,�$�Ol��ݺ����?	�O�����'�4AҤ��$o��K�o9@���I�z�� � �� $�џ�Jc��!;�h5��	Ӵ1� ��I�=/ެ� o۪I��jpÉ!)R�F�.�<m��}Q��z��[�+\9<2��?����'�>U��%Y,bu�̊���K����,D�\P�fU�+�<\R��m�H ��%�$馕��MyҌ	�LgJ�'�?9t
Z5$3ç�1�p�!�Ź�?�� Tx��?	�OK���M� �0�
R	ȱ8�D�X� �2�� �ˆ?간���b2��W�';��x M����ԙpF� �|��	��L"�<�$O�4V!2�"� �j�@X�'L�����?q�O���d�:Z��� ��N'*�J�|r�' az�%ƛNY���_
w�dh����?�Q�'�2"%M6|&�mX�L�2mt������jαm����Iu��c�H���u����G�}��L��� �R�'j"�H����"�bc엢e�*=���M�𱢞?e�����=ô aE='Ǹb�)2?�2�D?L"��Ǡ�?7��qh��֎�uW��	P��	����FMr&�>o��44����P����q$H�O\�:ڧ�?)�!��$�5	��=��`S�A+�y�ㅊ8���%�
0�Zm1��
�hO$��O��uG�
5]����P��X(�,��(��M���?���tx�+�?��?����y��W�8��2d��1��ER�dԨA?:%��$�'k9������8H@�c��t�ո!��(Ό��t+"d�Ġctj��tD��N��uقa;��B�Y�Ќҷ��/�^,�/��Kpm-��΁�6~ ihĢLIʾQ��쉉o�b��`�b�O�d�OV�����#@�����
P�c$�<yFMպLT S�E� İB�A]ğ��ɍ�HO�)�On˓%�I�GD<�h�R�C6Y
>�*g�ѶowZ�����?����?�������O$�ӌp����Y��>�Ȕ��&a�Pse�/�N8Kߖv�ȳ�N,P0N���	0.���:��z�T��uE� 0R�
 ����5h�$�i������X�(O�Y`GgC�L)�Ĭ�!b�,9��I(�M�C�\�'ݎ��v�Y�$��@�Ġz|���'��@��$���%K:l}^�l�n򉅓MC�����;#t2��O�2�C�B5d�CJ�N�� ��e�R�'H:���'�b;��8Q ��\�f�:T�W��D�Wc˴T�ArRȂ�	��w"T�U�h�� "�?�(O�MJ����ވ�%$[+g��$#�RS�dSqg	�c.� гb\���Qq"�-�(O,�"2�'��6m|y"��+|D$�s��r0Q;������0>� 3r���U����fA熈S���
�����GZmlUh��W�A��\��Iy"烤]��7��O����|�¬�?#�V!sB(�#"��!d�"�l���?1�*e��� 5���8z+�	�R�ѹ<H�9+ȟ�Pz�oY��s$�V.I�V@�G��0stN��e�5�e+�p��*&�;F��x����S��J �M��o�:��]H������(u}��E�t>��aBEbW-(�XࣅA56��C�"O:���ŷy��e�"��+LJf�P��	<�h��m�VGO:h�%��А)��0�u�����O����"�:�����OZ��O��$~��G	�
yS��yb���f�`�$¹n�b1��'r�0x��_j�b>�	M<	R�Y:@�:�iק�=b�peiS�V��!:�˟E}�}rG/��"I~
�)Z�,i�;3#^q���2�80���^�u����4*���-�&������g�	75���R'�0�@Ѳs-K�Du���ȓRl��P�F`����W�H�X�'��"=�'�?�-Oj�td
9�:��rL�F#�L;c�3m �聪�O&���O ��ں����?��O �i[@T(3��u(-p6'K�A����@ [6����gn@�w/Q�'������>;N�!��#Qܦ�x���L���ʀ#H@��S�D�W<�\a7�v�'�h�q���}����7]�|i�\�RVȦͩ�4����Dx�f�a;�q��G����ר�*�yb!E�I�P	c,ؤ+ϖő��M���T0�6�'.�	"u/(������dU6���M�C$L��+
�&LX�d�O��B��O���y>�Fˑ4] �(��ˑ�WoO� ��̈��(H EM�X�pbX)0&(��������]���#$3&I&��ф8	�����LD�Rx�	il@+,�$�s�#?���D���͉*Olpu�6?��pp����-�r�%�|2�'���`�
ʮRT��Agң`PL=�
��R�\$?	�Q�Hm�Ā�uB�?Y)O���c�����ٟ��OP�}i2�'nPACd�=�V|��C����' B��.����\��j'E4��Ĩ���&���U��	�6kS�>Ul	#1oR����xx8[ee�-�����V�u��m�6���UK:�O�����HѮ<j���g�r��{�O�$xg�'l|7�Tc�O#�� D�I�MWj��"�	�Y��H�"O��BR�M�Jw���W�s��2�����h� `ckȢ[>`�&b�0#Oڕ3Dh�n���O�dձ�F5y���O<�D�Ov������C�\�j(A��G�?KȈᑥĶ��t�V���H>��s��961��$�0��~�MA�&Uۑ��*�q�B.�T$����$p����5(��q����FR-�j����:��&%Q�u��dH�/Y�t�ٴ�剳|q���z�g�I,>�Y�b�ta�B	|����Jzu�R'�E�ubp� �VC�A�'��"=�'�?	-O�����З^�˖��04�����P��@���O��$�O��d�Ǻs���?ɛO5����Ⱥy� �3P�:A�!��/�#^����1��5��"U�/�q��r�'r��"��T�|}~!�則)tV�+�V�g�r���h����K�"��1�5�Zz�'�����*��w�N���N#���dG���?9�iyt#=���dR�§Rd����,ֳO�.,y�"OzM�pb��t�z��3������A�|�Lb�6�$�<��ِa��'pB�� j�hu�B,JW��ɤ� �v���'������' �=�^�	��i�d�h��̛^�rI�L31�,<�����D`P�Y U���bJ�	=Q����'����("C��l�d�jSm�P��D�&�׶�`���9!�2�x��^�Q�����OH$%�x��yi��: @@Ж�zƦ1D�$ `	~��Q`+܌:�.0�sH0�ID������O�]�
�=+�D}80���Y|�{b�|RLCe�6��O`��|"gՒ�?ɕ�_�47V\Q�l�i��3��Ӏ�?I�m��Q%�P44�|1%�=^���V��Sb4}:ȟ� �}�vH�m�5ۨ�♟���/�&Kh��P`�>�&��#hY�z�ri�p�7B��� %l�jv%8Y3
s�j�k~��J"�?iҿi'�#}�Oz��W*��H�j�¦��]���Z�'�L&	D�"�|)�j4R=p�����G[�O!���!��4S׊L���Z�L'JA��i;��'D��Ȏj�hX��'�B�'�b=�.�s���]�6�
w�E
P�Z �'�6SK�����.JQ�h%�H2x1��af��)�~B��%�JM;�&��ap5:�O�5�q�,��dyD���V4( `C��哉k���#2�`ޝ�����r�-؇� z4�t��(m��x4��$3�3��(<��%�$��i� pk��9>�C�	�aR6�����%T��À����'�l/��|H>	@�@����(|9�*�Evؤy��ʟ~5���QYp�c�Mfɾ���=D��rJ�40�����dl����	'pl3��#%�,�ɈP1�������I�Lj�(q�EP��RS@��Ɯ`��ʕ8%��i"<�h��c"�d9��G>���&o�9��Ѳ3e������aR����W�RL`� B"�_� ���Î��'Qa������E(�鈱p��Q��&۩T���:��̸��I_����@�Ĭ�|)�'��h�BI�A�9�O���'6����L���ר6��p,O��R�a\�I������O���	�O�d+/��(�#�V�4(Q���/�B�R�QlD`D��&;0a��ɍ�bF!�a�1�%� 	T/rp�і��#]��$��<O�I�d�Z}�6��WB�	�ȍKc�شB�Q��#�)�uU4ك�V_���vܷ[��S=8��o�^����'�����1x(�i�_�xq��� ���!�č��(͓k� fViq���d�ў|����[�j�]��Aٞ耭A3�F�NQ@���O��ƅ(h ����O�D�ON��D��OTrĠF��*���jS.4����JC��x��k	�*�t� .x.�l%,xV/3}�N�vt)��/��1�<����},4���ڏp�P����)��	q̟Z� ���	�R��(�#�L3%Q��6�$Y[�	�'ʒDA����f�?�O
�	�:���U@�+���
p�{�B�	�� E��%Np�ҽs6ƍ�M���{����'��I�|��A��Š p�w�� 'X������?�BL�Iݟ���ޟ��Yw�R�'G��ٛt��a�.3�
�{�j�.BR=y�☺(i��*ͣ7��0HA�YW]\���ğ�% �	��Lҽ;����J��1
��i=�]�h�
Y���K�8 ,���^�mM8Tx��z��\�M���A��@$/�6m�T�' �4��ܶE��;�3Ect��ԧ$D�t �hM�s̭�`��4ZR�;��<�@�i��_�ȸ�������O��y>��tC�eN��$	̌tL��d�:��d�O �d��NJ�U�����u��'K��A9j�����7B��x�ꔖ_a�b�.�J9��Z��9B��%	��O',��lI�LXL+�m3AT�9@%��K˔ Q ��3l��j��(wy�$K̦IPJ~��"Q<�L �%�E�4.T,�waZey2�'U�,[��>Zb�
t�
�D� 	�}A�ɉ5�P�3�$I���00�˹I`�ʓZ���+3�i]��'D�S09��4���������9����e� ^�&4	�n[ɟ� -?F�і�
�F����FCP��@t�⣍@̧m*u���+�lЦcK(O5�1�s�ɱ̂^:P��E�_u���f���ʰpEEƳ��	��x��?�!�w�8K��d.�҄}Ӟ}���'��� � (F휣26D�r���,~��G"OjX1����Z0�@}����d�OD)Gz�O�0M���E�_�؁��M8N0�p�'R�'�����/�W��'�b���d�'H��փ2*m)AO�<.�#K �.����B���Y�����S1Q:uʁ�>���ܛ����Z"~�de�����MA���2��j��Qҷ��\/r-�O���7��d��t�|�7OM_�CR�Z�"��ʓ6|E�I�M�ϟ�'����d���\������o@f�!��@"]vz��ӣ��U�d�"@A�Y��H(��|�����$��4��,�7��>r�r���ǐ�E0�Ѷ�M�N����O���Ob,���?����4��,d*�Ht�²w��-��ÿ�sȗ>
al4�t.�
1E:m!�JU
�QFy���>���E
�-��A$n>?��t;���,M6�8p�rY9��@xM(�;�q�����Mxx1�A#�"�D-�z� 1�s��DzB�ɸ�����N�j�F����,A5�C�I'�RQ�5��C������Sb�˓=��v�'\�2h<�	ߴ�?������'(`J��Y�&�Z��#
�?��O%�?9��?w#�K\,�bׄ�7˂<a�eYJ��;�͇�40M�S�ěI�dDzPiީd���Dyb��=4�ͩ0�@
s����/��_�~4Y����&rl��p���"�X5_p�@Gyr���?��	T>> �Ū�)	�v���1�DT�M�!�$ۼNS0����߹`���r�\�`k�����	Fy�9N$9��"y��<��������O���Obʓ��*��i
	l���d��G}��HfKIe}�0O��Ħ<q]��>���U:��Ea��8�v����1��Ϧ	&�L1f���խv��	�,�]$rQ6
G�y�X6m�O��h�d���4��O����^��t���e�V48��8A�#���� -�wY�l�ӟ��Bd�ܟ���s�����"���dޥCfi͗wK���`.��R�Y�B;d,b�'�"y�9O0������	�?Q�I�<!�?X�H�@��G3qQ�I@�Y-��şxqdc�ԟ���Yꈴ����d�$�_IL���N��}�`s�R�g�DR��'�,	��~j���?)���?ibӺ��0:�$8�W��\��t!Q�'�( [��?!(
*�?�^��mC��ܴ%"}��*O��삇�v�8T�&ՠ�6c�O�x�r�'L""Üz5"�$mݡ�I|��	���C���`�6ъ��E}w|d�gmA�<iV�ҟ��	9�uG�'F��D��8��i��L8�̃�{!q�7lE���z�#�c�86�d��I�����Hݴf�A�'b�����	�n`��s��aR�@A�/C���o�~Ha͓&δqߴ ٛ�OWL�O�%JU��
��*�&ŞPC�$ ��D�z�(��B�Ӧ�O�����5������O�H}�T�&�<���ߦe`�c�C<D��[�b�����U�H�˳*e�\��<���Y)�S��d�����Ilr�ȡ!��%5bt�(TꋙW��%��O���?).O��D�O����H���*1 	�m��m�Md�r�$�O6���Od��Oʧ�?��{E�q0��+M0�@#�J\9j���ǰi�2�'���y�剶�����]�"��$�OxL�����'�ɡ(FT$Q�/��N����^,L*,��4����O�$]�$V�|�	d?���И&dX��T�q+Z$!Bl��Q�	��0��؟��Iuy�Oy�s��Zb�oJ`|bMCFxu"O�$�ÇZ6A���?#�0�"O�ò�vܵ'L�����"O8@ɖ���\�]B���F�ؐ+D"O�-I�iL�>�:<y��.z
��"Otdb�G' r��p�)ʵ����П��ƟX�Iݟ,0��tEۑN�~a����S��M���?����?���?q��?	��?)�.��g��m�A�[A"P��'u��m����������ݟ��	ӟ�	ԟ���'`�>(�@T	F�xCq �x�j�۴�?Q���?a��?)���?)��?��Q��@�@K'qи��������E�i��'���'���'�r�'G��'phE*e)�?���{�@��F��B�j����O��D�O���O(���O�d�O�q �1�.A ��ߠV�����h�Ӧ���ß��I��t�	ߟ�Ix����`2VF�XQ�� 0�U"2kf���GĪ�M���?���?!��?Y��?A��?1 �V=<\�	-VL8�a�X�QR���'�2�'�2�'���'���'a��1q�\c7e���@�H̤n?�6��O����O ���Oz���O��d�OT�d��K<\yz��Èd��豗�.|�l����������̟���柔������2Ozvy
�恎�t��b9���޴�?����?Y��?����?���?A��8��es4*�S$"��&�G�;l�X�ּi�2�'�"�'���'���'	��'�F�9Y�j�Ї�V�Yd Gț:O����O΢=�����b�N�#f�T��!|R\L��d��}p1��x�I�?ݕO�R�w�P�$(��I5�ce�z���'�"��i��6-a�$�'��O�<��`�iS�$V�R����4I腤�f�ri��)��iS����^I�O�4���	��`$H�\����&�18�R�?9��i���+�OJ�$:� pӶ�2Q�51rL]�%f��B��'�����DY�OT�lZ$�Ms�'i�MI�,hf)�3h\~�炇@1�ʓy��L�F�σ�}��$��;;��S�<yRF�L�u�b"!u�tCFFR�'Iax	��_{"EKp�؃Aրx g@N��?Iĳi�x)Z�'�``����<ͧ�b�i\^���B�+=A�h⦈S��?1��i�Z6��O�Dz��tӮ�"A�U"%�R�E�d�]�~�y�� ����̛�c���`��۟�G{"N�P�Z�+��ٿ:J�v'���ɓ�M;��u~r�'y�$Q>��	'g�=��k�$8g��@��Q=�%�O��m��MS�'_�>�(@��,;�؂�d�`��܊6��M�$��9?�mʪ/�H�Zw�n�D�O8���O��Ė.lI��J���%OJiP�b�.O�d�OX���O��d�O�ʓR]��l'�y2��B5젳�Gz�`��Oɂ�@���?����O��	�Z����ӺC紟��]w�dE�����Rp�^)2���UL½ӛ�9O�7mJ�.D��yv�.g�j8�'R��IH�(%�q� c��`h3�GֵE����E3J0������;I4b����T
�T�0���	7vB��8
3�u�@��4$Zl�ܒ<<=��p�X�F���F���a�I7�X,HWB�[����$�W��@��
˟N�L(S�2y�h b�@�)�2p�S�8���� -|�r$y� �t���j�<�K�)�.yB1�"ђ,.�A��>}(��;rh��"O Z�D�}�Y�� 8N�6���'{�y"��_�D�ӁeQQ�mD'GBYx�a��p"�ى�W
�.��姖�],.Hj栘�R�oA-SjB��d��\zb�Ȃ�Z���	iT!9"�"���0v�Rx���j�.�rr�%�2���P��fpI�kQ+-#r���^/X���y�����`ɠ��P^��u❌,`���	̟ Q�a��ē�?I���Nx�8��$%�r
7����6����?A�g��?1���?����?����?���5��i">���X�
��tIȕ�Z1�'��'��'��'E��(�pa�OT���ڵ���H��'���'I��'���'���5����Y��p�X !�T?%z���W����ܟ�$����ܟ�aP�؟���l��x�4 �A�2�z�x'$֟��	̟\�	ߟd��˟ �jA�ħ����a�L��l]��A�H���?II>����?A��C�?����?��똷=�}h@b�`�a�����M�g�f��r��.1�)
�,U�fo�IBP���%�¹���O�7��a��y 	ĝ��<�`Ǧ���'��'���'�Қ|���7'p�9�ȕdg��� E�^������ҟ'���������31�a���-{�D��'Φ(FV�n�8�M�S�'d2�'��D����'�¡�`�9�N�\|�h4�PO�Ա�5��
���k���O��8W���')���D��q�Āڊz���pVhZ6|!��;)8�r$��^5�$hN�Ll��#�#aL�=����'r���(�\='%�irfݸ��¦jK�XD�� ��{�,��r���{��a��&s �8X�L0���t��{9(<����O��P#𭕢W�[V �,g��u�^�	F�C�E�7(��-��i��XQYJg[*$\�j�}P�r�b��<����	<�uw�i���D���2��� v��	 ���_!F����{)[d
�'b�܀�)��d[�#&q��ط�Q�R�˥]8�3�枋W���&��}7���%���[&cu�}4��$4_�)
4 ڂ4"��(.O�p��'��6��$��N\|�h�1�E�F�x�T.��A!��6qĜ�8'��:3��[�n˟x*�DF�'%�����r�fhp@*�%�Dm��H��5ފ�P�-�	9�|�d�O����OZl�;�?�����4.&o\��U�L�g�f�u��8SH�j��ܱbPʀR�oֶp249`C	�,��Fyo3R$��K���/�8� �nI3)���#0��:l{��{�B�"�o�$8Z.�Fy�ł/�MsV��(.���?����S9g!X7M�Ӧ��ny"�'��O�D�ν:f�`�-�=whX���f�7�p=y�}"�X�O��hd$8@b�����􉇏M�����d�;	�x�O\R�i�
m# ��qbЙ���{��e��O�d���Ov�$�O
!:�E�yO��G��M[�0c��w���b��&Y��p(�J�fb����&8�y�%AO�ws2�1b�<u؎	��0{M`�U��MH����B���=�6�ӟT��4K��6�b>3�cfT2∤OJ��,lOz�*([���
��Z�v+�,��'����i������� ���bE	wղLI,O�B�Ѧ�������O�&YI1�'ߛ�E�� �@�w�nՓ`�R� ���ߐh:y�˒)3��e��%��Q�Ƒ�@�l�&tS�`>������X8Z�d�,OpP��+c��a���ސ3�ʝY�#ö[��BM~Rr,N=\���/�12��Ӷ.�F}�6�?����?1��H�&�u`ȩ� ��Hڙ#��!��>)����=���_R웑R�T� �dUk�'P"1��?Yb%�^� ���s4EϬb�>xR����?!���?�OE�9��m���?q���?�B�qޑ��@�/FA��)B+~���eO@�hk�n���JA+}����T�.�tMf�xA�,Or�i�+ĘEy���鄞,9�a:5ƚ7ܦhX�`D�E�h��aǟ�C�O����#dy�I�@����a��5��I�W��	�&m��� ��埀��4��Y� �	ަ�����x͛��ȀGA��3�<���<�V�@����酨A[�T�,A��b�:�lW���?a��sy���t�? 2-���O=��a�C3 ��s*Z�"r���͟�I��T�Zw;��'��5Y>d�����b\E� d*@�\qGlM�.8:�Re�i2$�V/�2�`	P4�	�P��K�㚂Oc��1Q]�#�8L�p�*~���'� U��	M?;�����x�@$���҄p�>��sdJ�1ẖ:_���b���d*���O��d(���s� ��,�r��c�V?�Ѕx��'9�O��hҦH5[؍��j1~�&�#�>��i��Z�@X&,���M;���?	�4j� ��I�5��땞j�����'즰�D�'��'���Q�h�xb1O�C�jM�#2!�w��R�d�����d���(�c?eHf��`�v �d(�T���!�.�b�����؟L�I�<�;8�T��
6;�V��s`�+H���?������63:�4�B�?ˈ�10"�`;�~�˧�d�$�e8�X��B�?�*(k�aB&��dP3!�XZ���ON�$�|z��α�?��4&ѐ�r�E
�T+~�iÒ`���c�'L�FdZ�v_�	DOS��bu�R>�$>=J1DP�n�������;���i�ͨ>�J�68�@a��E�Z%��!On�ON8  � ��-	��"1���O}`w�'F7͋��(�6��`�P�`��X�+(̘���D�����"O@�����~��A�`X�r�~d��I�h��䢓`<+���Z�ؿZ�"X �: R�'rCuD��C�'���''�~�!l��Q���C$�A�B�Bm��F;��3vIW1m��И��[\L1K ��4?Td�)O�2���| \� S�+4Ʃ��IW9wfi�d��%�J)񢕞m��O&�)kQ�py�OyrX�����k����o�}�4�'���[��5L��2�'~��i�R4E��Ee�	��� ���r
�'�!��{����i�!�0�P�'�"=���?-OR��bF�#��ИS�94U�Q����Q	�OX���OJ��кc���?�����Aڴ\5�b&�ĘN��*�E��@����)܌�"7��t�`���T�a�A:�2Ĭ*�O� �@�i��yU�νN0zq�@�΃��(���Oz�'���	���&���Oʅp��6Zd�Q�nX�AQ�'\��с/��XY	�W�>2��@N�(�ݴ>���\�(�P
%����O~7-��_�T�P�P(%���Z�@<�I��]��I�D��0v�Q��0�^uS�
M$1�j����جuf�Õ��=(�H�Zl߰<;���*P�z�2�0%��
Y��]�K!מ�a]�.{Z�	1e�`�ӎ�D�;8���mӾ%������g�(�0� ʙ`�	[�>�����=�,�*o`r ��gT�2�BQ��O	P����' ��,6'$�ig ��{VI�C		#�	e�P!�ش�?�����I�`�n��IԈKB���;/f�SƊ�ǟ�Ѓb�`���%S��|8��Z&%�p����K��Wj|i�m�>Ŋa�LU.�AX�I�bLh5P��!ρ��^�UE�V*Z��|�x0 X8Sl���
/:��$9�Q��z3��O��mZ�!Q>}�ɦ5�˄:�<�2c'դ~hƉ�u
"D����]޺���.TR��mjqf!ʓ�?i�鉔Y���J��W�`�l�6Fŝ<5�����韈�I�h�tkFw ���I��h���ā�5�%�a�'M���aٶU�B@��!YAw����	ݓ?�i��͏k>�O��ulU@yB�Ȯ�V��4!����ڃ�\h3�mAD7>�+���0p�I|
�d�.0�ʓw�\���1,R$$iE���1��x���<���U�<0ڴ���;+K���g*+I�|�pr��� }��ȓ��C�P,U��V���"���mx��� �4�?�+OnT�����#��۞%v�����ޣ4������O
�$�O��$�Ǻ���?ɘO���'u�4�E��L�������2�ȠZ'���$0�����r�Q5'�J�!�ŠHM���#�	B؞��aӈ���H˂.�b��g�\=��}�V�،�MS��iq�O>`E�� 4H��PG����7IS��yJ�FTr@�O��܍���ŉ��I	���<����X���'a�i9R:�b("��x��@-l�
�#�O�Ñ��O���OR<CT9=�0b�֝-^㤼��ϛ4G@���@̇h_�#?y�#Xn�z��~0�<���G$^0A���%�j�'������?����?�Xw�����f��^3[{H�a�'�r���Ԩ�q"-Rl���E�U�w����x?A�Z8�Pr��S�G���a$�!DB�I�+�B���Iџ���A���K2�i׶@*�/�*a� �K���M{�Bvm�O���5
B7c�شy��V:d���{��3V��P2�)�I�#l�F��E�]�u�
�0����~��I>^�VJ�~s06M�^����Q6A�֓�>}��	�V���OS�=��L3�W�P8�"�O��mZ �M���H�p���?m6 �d�(h��P���>!����D/��?�"F��]�@�`��E�Z�ya%,ʓ�?�ѽi��7m9�Dzݍ���&)t!Э��a����EŘ�?����?�D
�-������?!���?QUe�� vR���,��49���?���4�x�[Ӱ=
ݍ!t,�JTCT�$��`z%�M�I93%"��$G�lj6QUd�CQjX3I�-pN�'��Ԑ��o��x2�J�*u�C�R�#���ct�yr_�P6dEX�*�3p
mA�	�~��=�S�O̺I��AԾZ�2�D�q1���
��z���'�b�'�"`t�	������	�qaָy��_��^��#�J>݄th�!3�xQ��������ǌ-#�!�G�H�L�V%KàϮY�L� ��J0Iϓ[�$mZ�	�$ڐ��_wMxR����P��n�'�'#�'��&"�v�Ss�7���,H`�0B�9D�,"���8�t�ҕ�5<EZYq�O6}��tӚmlyҰi�z7���'����E���s�L4z��h�L���'�R�T?����w�6$�mͰKA�e�&�5O�Q�`h�5�E��:k�ځ�P*J��q:Ѩ[ S���"�S/K��5��gFB�ln�j���ȫw�B�ȓ~Wx���ψKX�$( cp)�ȓ�>A���\�Y���+r��~�e�ȓ)y�!��JR<�����K�F�Єȓ>q���EU���	2b@˸`* �ȓDr�p��ߤHe��Ǎ��kt6��O�����L$W�� ����j��Y��d�Pҡd��6��hW�R�Vt�� P�	@ ��&3"��G���PXxЅȓT�	�A
�A(�PKwe�5t�ȓad��KD$H��Ѻ��7V��E]��81<��}��)=�,ąȓA@��7jK28Od=ˑ�O�pɅ�5 �Yɴ��7��%���Ɉx�ȓS�H𻷈K>��� 玎�tPz��ȓ1ܖ�i��|VB��QC�g2��ȓp���eަl<Y(���,j��ȓDƄ�7�U�7�h��Ed�(6n؅�K|��SB*�?~�e��d[p8)��o|�'�ƪ!��bdX�+6v���.]d@�P����������
�QI bԉ@�ݨ�CE�W��p�j1��N	"d*��6�v���[�� Ҭ��c%�8�'�^����HTԍ:�E"J� ��`�2x�ȓ@L,ca"��n[�~�� �ȓ4=�u��F�*2��@�Ex�z܄ȓ
��}�5)v|��� �1� Їȓl1!t/�o�8�դ�^/
)�ȓo$����<
#��n�DdLh��|  ��7"��Mc�a��_����ȓV�:�:ЉB�_@ɚ�l f���ȓ}	��[C�� 70)1�!Ʒ>����ȓu������Z%#$��@#��3sg$��q�:��WB�̌�AIų� ��ȓ9M����R�/l�0F-5�B��p��B!�M%�5��Z! ��ȓPҬ��FGU�-� yY֢Ȭ<��<��p�������'82�Al �J���v�>���
"�&�T���V؆�.>Fa��� �a�U �`��P��[j$��a�(\Ӡ����C�A0��ȓj��P� J3B�ˣ�F{�ц�(e,9�0iКy�mK�@�!U�!��j�N��&%BLr��Y�J�i�ȓg��Hg�"VB��u(�ą�a�� #�K�0̌��ŏ	x����<<2�)���S1z9�I֣(0���	���7�؊pM���b��
����h�!��gݨz�@P��G�>p���S�? b�VH���&7�Vi��"O�=�e޽�xp�2G�+D���4"O���AO+rԮ%�%��(��q6"OjA��+.���4n�g�6�%"OXP{ 뙡Y�܊�'�*+��U�'���8�!~
α@�G�(`�֑��'zyp�"���
ǩ\H�)��'`")�W@Yj�)r�&�!θ2�'�Vh�gዦ4���x���wr�Q
�'BN�Q�j��3�8r!-�&6��'^�����fx�3,l��'�X%"M�PKμ�򆗯�y�'��L)�-�P����ޥ
��1�
�'H|�&��V�@�3�e^"2�Fh	
�'K���c�+f:e22���b��=�	�'SX z���M��󑪃�YzL��'��٩#�4W��z�NF,H�'����0.N�#�2ѫ�Ąb��A�
�'�>����E�v�y�%�@V����'4P�4�M���:��5I��(�'�%h`�V�K�ZU��M��6eˍ{2�'�D��CHM�$>q	���
��X�'��֤
�[�����b}��`��2�ygD�$J0Yñadg��rj�p<Ɍ�DУ6Ψ���٤����n�9,4!򤋏����,t��=�pc����hO�f�Bvn�L�-��	C@;�Ap"Ohi�"V6=T�ݐ�킘/!d*��d,lO,0��I݄]�LhS�&��<���r�*Ohѣ�>��"���rT��'�{�@��*�
�1��l���'@6��C#0��;��M!>p`�	�'��8�$'c�N�q'H5%�y
�'�z8b��0c��xPBƯ!PԈi�'��<SE�ʄA�6�bf�\�S���'��y�e�U�(�<��`�%=�r�'p捹�,���m�$G��
 <�H�'A���R��t_�T8q�T8.��0�'e��#E3s�0ȡ��t��U+�'-HP��ΑA��P#1�V64D��9�'�ֽ�ݥ|��u�ꍲ^s*`�'J�%b0ʔ X���#��kҰ�	�'�Ҹ�f�:< Xӷ�^�ayP�ȓ�8��G�Q/e�.���
LQbl���t#d:�oB�@l���`[�/�n1o@c�E����{�a��+3yZ]�U��h����UPzA��O��i� �1��hKID�U��8H�"O�q@��E�yƐa�A�f�4Ay�D�2R�����'~�j8�pI���q{1�U�l�,0��N��m���ΪY�r��3���Y��-����gܓHɀ�|�'��k��˼P����W8`���'4��9� Q�:��*A(47r�IB���f9��$fL��O	y�
*�Y�F��(���=@���X����i�LQ�F���c�Wl��ڠ�)D�|�d�{��C�Ƀ)1�B�z1�&��$�X�?%>�"���?�t�ŢL�v�p�i�l D�ta���L��K�A��G�Z �ā?D��Bե͢e2)���}&�ı��>D�(�eP�	y��p�È�Rg��q.+D���p��>K&�������)�F=O.m�$���'� �{4����CLq����'Y�����Z>�f��&�öp�@.O"p�an[��jșK��|n��v|�I`��-i@~��4&Na�<1�(�5��iWBZ�-{�`��"U�"��ʓi���)��V���ا� n�#��H�vu#��ܛd�J2�'�� ��O�.m��j�-%q�Yrj˸'v�E�V��ٖU��I�y��M�2�A�;�"�1!*�
u��>�g�^*
��C����'#���z�L�4�0��!��q]
%�ȓ3�B�y�X�:��Y&���wRdո��B#jҎEʇn������4 _�G��%�c�C&�� �"O�0Q��^���  �ql���
��G���d�03@�@w&*5��3�=N!����0�#7&�%�����	Yg�ə���$Q�pY7ω�0:��а��B�}z�Jv��`��IA����a��{���`"��b^�#>ٓ�Țz\,X)���K�1R-�L,!6��0s�p@m]7Jd`�b"OxS�ɺ'E�LT5'"��3O��S"K6Fh�d1�"-L8|�b�����z婷	D&� ��*�~�<�PoH�z���$��^�$�2�I:	�8X�N(��*ө�r���O�0�@hD�#->%�0��'b��9���'��@��H�G��Ȧ��o�nA��iҮ<=�isH�
h�����'��"�]�I����-�a^5����#_G*�C�I��W;��C�|�q���V����������J�<EX61�v���:8�j��FN�o?��+`��Q��7p�z��iF,d��W�.ܐ�JAi�?�!��R-pQ�`�n���1�Ɂ�!�f�1��O�x�T�8L	J�M?���R苝B�K֑�n�s���i�a"-�<.��p��	̴4P�U��l����R�)��@[�'+�")I.j9��vh�|�+n/��!��躦c� k���n����!5��a�"Z47���C"Ox �vKJ�a�4!E�Q��SC�>�(7���?e��H��}Ȕ)�
��i �?D�l���.aV칳���0��X*�l=D����ܦ3�8�5D�0�Z�0rI9D�I�Y��j�	\8y��0D�,:���<MR R��/_@���(D�z�\�-��@�I�\�AЄ�$D���&�N:\Z��Lޒ
���!")"D�x��FW�ɚ�Ȝ"�jXY�<D��q���O�a��E��u�PX�7�1D���dѦ-F4�a�&Q�J�/D�$(���0ۖ�*�{d�A�W(9D�8�g�3ӯC.����"D������ Im��@bh\�%b8�kǍ D�ܠ�[$1,[������-D�t¥�Wje;ֈG�IS�)/D�`��`����3�X��/D�8`�A�$m	^�k��?H�4�C�#D���� b\�� R�h�.���?D�,� �W��Z����-��U��(0D� C!��9h��^),���Щ"D���#�=����I�8�d���'D�T��)L[�qx���#)�����%D��aAO�%Ҡ�_gPX��O&D�D*�K�#����� �����%D�X���	-�\%��K!u���r� D�<�G��!R��2o�B����#�?D�L���ӳx3ȴjC�^	Yj��;D�X�3���\,^��hھ3�v0���;�s:�U��	�`�$q�㧔�\G�� ���4o��B�#v� 膄	cΘM�wG�)<mlC��I4���=3p�KP�Z�m�DC��=�.͂��Ǌa�L:B�Z@� C�ɒc��{qI��vʸP���ܧ}C�	�&������h��q�����B�c��rG�߲o��a�s��+��C�	\CB��C��L���He��rF�C�I�<5  �J��ЌU־a�hC�I�-������ۨ= D��@���C�)� ܨ*ՠeYq"@�u�:c"O~��w��=u�Ҡ�����+��b"O��Hu��,@�,X�ڭfb좳"O�1��L�#)�D���\޼��*O` KD)�`q�!���""5���	�'p
��cѸ;1���w�̭��<!	�',��0lO�qB⌋��F .8���	�'���2�@�h��X��5/���	�'N0�AiG�=V��Rr���<M�	�'.�U��+ճ;h$�N̡��= 
�'���{��]�buv� ԠȰ?���'�NY�T�ę/;�䳢��,�x���'�\���h֯4jPM��E*l��Y�'� +�.7K���3��)_�Ia�'t� h�GF�`�7&�r�P�'^:I���V):�9p.̃w�R=;�'��=ڱ)^�N��X;taH�Z�̉��$�2�&�t�:���k�h�H�$��.p�s푆i��88UG4D�HYՆ��BT�I�!�<���d�<eNZ�j��"�c�<�P-�X+2�贂_�"��h �^�<ap�I�<�|x2����O�\1�4�HX�<i��~qN	�1���w����#BK�<�A�*�,��rFܧ]H\M@b(OE�<#�  ��f
T�7����̈́g�<��F�,E$�a'�^j�q��j�`�<I�hט�нy�dI�U��^�<a�ϓ�b��H)�lN3mz�=����W�<Y��p��.]�e�}��k[3,x�4��1H��a�2/Wĕ�d��vL=���Y� (�W�8���Q+ ��U��!91#�	6:��tR�H�ȓ.v�`��Z2W�� ��eD6-֠��qW)���.���q�41��q�ȓ'dȠ���ى<+~d0��3S��l�ȓsK,�2#��/K=�x2�A�J���ȓ�P|�P�0
F	�'G� �ȓ"�^@8b��-,5&����HzƸ��ȓ4<�A���6d)PY��cE�-�r��(a<[re��(�p$`F�V5�L��ȓF'����֥fN~-�W�M0�������LH24?�i��j��TL�܄ȓ'�<h��d5yn��WH�]Ғ|�ȓ+1R��7nM�r�L���En��ȓI8dL9�k x0J��/φ��d�ȓLp>�vd�!1 �((Wb��bv<�ȓM>�;'�ۙ=Ҥ�k�� o�b��ȓ�h{ci�[Th[�ė�x�ȓ3Gd|�V�� M���v��;�r!��؅�4^0�����\� ш �I�<���?]P�D@�#^��5!�l�<Q�λqXD ��8	0�))d�a�<�
*����FP0j԰���,�_�<�KȢ�q����g� ��)�Y�<Q�@[��+s,ט��ud�P�Y��F�q��C��9kN�AnB�?��Fx�����@o�>[�֝r�̤����O�X��8v'��y���eS
�����jq�K��O�ư9U߳���Zq�a&K�v��u#U�O�,#�Z��e/�1�Rt�p�|���IgFa3�o��RU���o��x��6��,F��sT��=\��,z���JN������S���@���&#P���X�L��'�P�����D�V�#�@x�&���zQ��� #�tl�8�4O�D�K�\<z��;���B�P5�I�K�%-�Z����Ik�'
,h�'8�8і�5��)FH�L�&h����$�8�s�%�p��W��
��	��<E�dh ��(Z�c�:X�7���H�Of, �۟f�D"���&���O� 5P�}�d��G�3P-.M1�A#AM��G�=$:1��´��S��5Fi\�v��8jW��H �!���@��Lb�g�� .ax�F˥�|��H�&L�0	�N>��@����{�Ow
Yr�oL�Mm6�Z���)� $�u��wx���d�F��� �`g����V7Ya^��E	�<����
Ԝ��Ity�$�S�j3��k.�1	����D㸐0�г2�py�?yR�V\UabU	�p#7h�A��oc����,q����t$߈U�O0�dE%x���3��W0�H��ӱ<����h��X��B�2��! %���"A��p*E$#S+\�PP�� ��ۀE�3X���nΣ+j�h7�
�Iy�Ѽu8��{p�RYmfTc�	;�y�pE��:���EɃ]�B��s '��(Oyc�d4y��{��L�l���H�&�6A�㉦sݲ���*��#t�Go��yG�H�(����I��q?��)~��à|�s���k0�_�BԔPѲ` fj ��H0�	$�(�h��P�(��m� vL��'D�bF�����P�AʕEU�}�B�<!�'��Ez�V0��F��MS�Iڕլ��� K3�J�8�"=H�O������tc����'£�%�e�!��7H`X��B�z�@�!�,S%d�U�i4�PhT�w��܃�4YF~ԃe�	�H�j��!�!V�Pe��g�W�A�P��f?�J�֘��f��㢟�`�4|���-s�b�y�`8��<��%��f(��;*�� �G��.CE2NV���$�����	A�$#ѧrQ��H� {���7��)$V��3o.���L�a
���u�g\�K�H���o.}��$Q�Т�*��z�ҳ͖
/?� 
/N����Ο���������@"�Ntz�ҷŦ>�T��9
?hh����#wɬ�sS������=-<p��w�N㞘	⍍y?��F�RH�p�A�}<�c'�
9��oZ*IN4굧�'>l�T�&���"�"?	�&P>}��&
C!O��tas��@�➐y[b?��'���Ӷ
�P�Py1%'Sjp[�M
-+0@	��'<M��eEw����'f8�!���/OP�`��]�y��]"���x��7��1�O����~�	�.�$��4ɭ
�jŁ���(0H�?�V#I�PH �a���ԈGx��T�?'*`!�Ȩ6����C���_/����j���?��D��:1"��وvA���C��~}"+H�l��F)��Mv��¡L�2�@�,*���@h�j��D���!{6�r%%�L�Ĺ��֭AE�6m߆.����aɢx��Ѹ1�X<MÑ�a�ŕ �U�#[��n�Z@�L�.��dG������;5��w��Гu��3PqV�p�ߙ����ɽWO@�[Eh�ռ;��  ��r�!��&��3�hMM�Ip��d2�S�<��u΋!P� ����%U�Z�k���2R����BN�_~$Bƫه*��B�ǝ��I�(L,�ÁxZx���m���'����Ц�� *S���r$�i�<ѯ;0[�ɸo+��)��х@�PYI���,!ָ����I�R\
 ��Tx*�f�i��8�JOQ�@�7C��{]��$�ӯ��'�y����>�
�4L"%�ށ]\V���	�� �C��Wnڀaӎ���<Jr� �n �s�8�p<�� ٙB4�D��w>�!� �ڵ)��������7ހ	��#� �ϗD�f!�C�S-N�$U;�耧Iu�2�������@d�Z��H�r��!�Z��)p�D'Fs*X��⌽M�0Fz�9r�h���y�,�bu����dDPw��jǫH%&	f9��2�Fuq���6<�U`�h�+� 1�-_^�Q��� iZ4����9}�4o�}j0�$E��PbQ;�ɣ&ھ#?��l�>6��iӎ������+X�iIV������3���	j� ���������?1"�/	��GlE�Ň�,�"1���>���)����s����OQ�B�,���/!; �B�8T����h�&�
x�k��Wep�@�Ꭾp�(c��'�:]C�!�8a�T`�A
�	�Sϓx�Ub�I�I�AcDl���.aG��b�f�7`H��ȓb�FqD��^:\��n�R� �&�\��f�6 �(���=,E��*ķc(�@ʖ�G�]3JC�I27^��#c'k��Z�V%��%q�-X��	�Bʆ���OZ��Q����<e��K!��+��41Ų�JS�L|��{ �HkB�1�NI"����!�TP���
�XhDyr��&qNH ����aJUR��*��
3wP �RÓ/�@���S�=5�2w�k�<��VԍMo0���Q� �Je�5��D�d���
p*�l�I�mx�N�HY�U	^%P"�"?���.~�p�%L >Ǽ�h�"I�	�<B�� C�捩��^2g8$Y�/U�0`gθ�p<�l��xi2�w�����=S&�D�5־V�x���=-��ȱJ� E��!N��p�à��t��$������d���āS�(��r�Iyh�V�4�1�%4���kp-W�KΘ�Fz¤E7�ؚ��::X�4��#����A%P�r�I"�3[X�U��o�U a%�d�8ᵍU�E: �*O�B�?�)� �ݚ!HP�s�N�y��+n^�ۓ�i�hw��	s/t�{���+>������dڹnw@[��[%p3
d��FK5Q���O���S$[�����O��4	����E��s��m��=���]�@���$J;cZАy 5�ݣ��ʚ3r̀V&T�'}��h��m~�T�(z��,h��RD]?��Q�B���r�i��TQՀƖ~�
����#��4b��ȏ�R�����m}�X��'�y�$M�Jj�@�W��!ƀ���U�����$_e�(d����N��?� �(WO�OldcB����Kj�g�L�d�� �J���0�����>f�UK�!�+0*4�Eg~��a�T�X���F�<��*ЃK�A��d7�]�ua�\6��á
� 
�2�$ךp�z	,���T��-[�UK�qh�E�*M�ʘx�nB�,\���&4��6���w���S�4�<��g�)@�J�uOR]r�o˧h���u�p8�<Kq��mV�ϻC^�i� �<_�@c����`:�a����
+�ĸ�#+��'Ĺ��o�m3So��b���b�ㄙ�z5ʃ�)�I��09�b��=E c���)s�n�h����j���ؑ$:��'&^��X��[.o�J �����ɗ�y�HX7�1����S�T�e��Dd�gV���K��';�5[�BZ�@tn�韈x��L�o$Eb
	�a�֘��G���?�'F0,hb2/YESzy��ɐ���n�%��`Z_4�D�C�`#?9�j��#��\��ͅT!p��e���c*�89�n�%J�ܸ@O�=ʈ;�S�)�>;����~��ƞ<;L$s�K�:��/��8��x��:l�lQ�D8�l	A���kY,A0�!�812[�Ŏ $���Z�M�'�%�lC���V��?�q[�P���A� P3�FD8����?	�)B�b�"�> �b$��0ܢ�#b� z|��;eK 傒�Q�)�[�ɇ@��R��>��J�!��B�"9�eqPi�%�����?p�Iѷ�7Y�Y���J�!ș���4=[(p�)��]<���'�hHұ�
9�X��W��+�i�.oh4� R��'�a��͇ͦ�����Z��P� �L3���U�#��
Ic�E�!3@"0
c��]����Ţ`�3 
�`p���G� ?E� D$+���
���ô,�(�@E�V�.O
�pÒ #D�݇Z.&4��'M�si� �%�=.��|��V��c�l�� �8�Yw�&5�OH�h
d���Y�j6�^-S��1��K��E����"n��?-B�nѹS��?Τ��"L��z�ɍ:fF�9G��8e�r/�it���5BO�ST�؈q�@f?����Q�R���V�L���?��'i:����N=��y�G��1���B��	\����Ы�G���'B�N}
V�~-x='��X?/����ƪ���6�cᄔ�>��҃��),jy��V�H�Ke�C?��O.]ZTc��$>LB1 �Z�*%����(���b?eE�X���ȑL�c��� ǣ_�$��J�	,�����y�望y�����h(	�b�4��u�θ�?a���@�D�ih�|}��@����]����!��PB6��>VP����ϑ�2|���+}��LTQ���6)|�#� �(�M{���
�����'�nma���P���!a�� pdr����A-�h)4�2Q��r�Q'�N�Ъ=�ԟ��. :A�Z5;�	@E�[L 8m�%��\�b/�A(�t	��a�Z"?1Ԭ�=?͊4�H�"De�4u�4)H>!@m����ħ�@�0��d��0j���(\6���ĹAS�x ��#p�:�7��sG\�4I��o�+?oҘ9o���'��b?�{�μ?�[ã�.$)*��AXO��bP]��B�L���W��RUh�g��v���O��w�q�����J�as�u��i}� ��|Í����,,y�52IW}��y��a3u�]! |4A���+\P#���T�W34��$��3}b�K�>��0ɍ_|l���M��o��&���ߡM�t` w�'|L�V�˙j���$�
��ů�4��I�M�85������8 �TD���^�s�M?o��F�'bT���K�;V�8e��.Ҙ��'fPQPD��R�Z�{do��&����'5����|,�E��%����'7>M&A�	� ���%"Jf�
�'� x����6����f�>��'��P�#�����с�F����'�|�H�A�=�J�+�	��{�&X��'�d�e�RM�d+�CyB:��'�X����%:i�p���_d�
�'����Q��z����S=4P�
�'�#Bl�1G��p�&�@��lb
�'�^� t&>ljZ�ڇ�ܔ@Q>M�	�'�`��fB��MP�����Z��	�'Y:�cwE�g�di���w����'�Xs����lu|��gI�r�����'1���տ%<����R�h,�#�'�j��O�2�c�ԗ2�����'�dzA���T��L�쪝+������?0�l;��U�l�4��_e�<� �p�@���*����G�[�>z�� B"O����	 ���s�	Y�b֥Y#"O�7E�/N0������9�3"O M!a"��i7�|b6OO���pCU"O>�R��1.)N�S���"@Q@�"O����^�1��	���%E!��R`"ONl; !�=y��yd�&��S�"O6(�A�� �z�Y1��.��@"O6p��K4U\q�!�ze��"ON�Gŉ�R������g+��yu"OL�9r#8t�����l�`�C"OT�k�G+��YD)W�
�f�1a"O�v��5!"���M��bB́�"Ov|e)m(<IU,�� I|��"O$� �O��u��+��~׮��'"O�!ԩ�P��D�+Á(�B-rU"O2�sv���xL�X�UVy[���"OL|[�HǣU$!�pQ�-�"O|%x��3V����`��OD@��"O8�K�I��*ǲ�"#gF�pg�0�"OF���Ō |Y����+��A��"O2�q�F�0oe�E�R��"(%:��B"O���ЦQc���g�J�q;�9�"O�T��0v�>�c�	�.|e2�"O��:-O�n�l�"�-"h�"ON	��Fs��c��/����"OȐ��!οs� A�cH�x��9�"O��� B�u[���Y`2"O�l
EOƵkP�L �jܻi��:3"O�(Q(�"]ҺH��-��� �"O��X'-Ac�+�3���1"O�dP� p� ���P
W.T$�"O���d��^y��ٓ��E��y��;(&��)�Aƞa�j���	��ybA0_�p4`!�,'��xq���Py���	I�R�iA���hx��R�<�d	�3pl0�	!7����N�<y`��1�`�o�	��C!�I�<�2%��l=P�+��+qmx�s��@o�<���H])LbW ��\稡�$�l�<����"#azH3Cɑ$w�:DSB�k�<�p'�'Q���#�'#�`[��8T����j k���KmTS ����+D���Fm߭Sr\`���Q-�PH�
(D�d��Ŕ
�[�]� ��#��
!�zB䉿z��!ѕaS�9���zk=;rB�!j���ȵb�2k�jЄ /lJ�B�	1T�n��cL��&�cv@
v1�C�	9`�,��GWK��1v�;}ǨC���v	h`�\�mL�ݡ�*�.=DtC�ɯp�Bp9��&eV����^�}w�B�	3qQ�a�@`�'N�x�ꆯ�<[�dB䉀_�dԺT 
!�FQIs		�9ELB�	![c|���)�N{i!Dd�9w�C�ɏ�z��!��%S��p��0 ��C�I�Hr��k��$o�tSF��Y}C��=���v��}�X��,P�E�C�I�_UF!cgd�_BZ�x&f �8B�	�Z��l[��w�8E�ҭK�x@�C�	�Ab��b�c�r�r8�D˗x�C��,j�Ϛ
LZR���W�B�	 p��ЂQ�F�s�~�11.;��B�I.O5�XB!i��t�P�h�+0�~B�I�vP�usE�вB5�4��֖}@DB�)� T����A,rQ�$y�A`���؅"O�=I�,�XaN�; Ҿ�^���"Oly��C�DC�]p7��2S���"O:�v�B�)v��Ú�Qt�(u"OV���g�	�B�`A^ :�X A�"O�x�R���f�B���u�"O����!�{G�PF$�� Q"O�0Jӧ.+<@$16�Y�"O�p���]^ծ��d��)v���"Oh���J��0���S蒂w=����"O�����R���93��� ���y��"y���REQ	5d	ڐg_�y�!��r�����CUg��3�A�y�J[0VRd��BX�I�P�q�fϢ�yb�>FN��c.�85,�`����yr�Y�xE�FG *k�=;��ӕ�y2"	��hV�&�D$���:�y�O�3���fd�ܖX��M�y�f�-@� jV����Q���y�#1�*�ɦ�!<y&���͆�yr/�r�Ȫũ��fV�"�BX��y�c�1Q~��H͑�H ���Q&�ybA،q2�0u��1nM����y��N�h~
�C.^���!�y���s-f��BN�Y�.����P��yr��(.$�u/�MG�M�'b��y�e�[��2�g��H6�D��A�y��j����̍����5���y� ;ki긚��{�]X2*Х�y"O�,&<ș#�Ή�D�T�@-��yR�#�^a`�)ƽB��:����yҨU.�����<���w�N��yr�@2q &{�.�Жe�=�ybG�ehӳ�|CN����)�yB�'\�i��(�;tp��lS��y�A@�u��� �G�q=x�+�Bc�<��CM�,[�X1����1����Q��l�<aRM޳�4�G�P(�d�y`��k�<�#�D�8-���&[��`�Q�Ig�<ya��8Lqዕ!4Š(!���`�<���ee��J��8k>�=:�l�t�<9�����$ �qe�,#���p`�Es�<�R�1jQ���	(�"ݸ�aW�<Aţ�
0�����9�0��G�X�<��ϔ�&:*��9�B5��_Q�<	7�K:@����cʐq�@t�<�0�ڑfh	rg�Ș|1�at �q�<Yd�C�s� ��P��l� �.�h�<A�)3B&V�W�Φ?ݜUw��J�<Yb�M�@�L�&- p;ܓ�J�<a��76t�X�E��c��0r���}�<�# ��0�fB �q� ub��b�<i��M�h��3�
�b^P�ɶ`H]�<��P7O4=�B��hx!*Y�<�S��<����M�2uQ��k�<y������{0G�;P�L%1 ��j�<��]��(����XI"t`��
f�<��E�(t&�H�hU-7�P��b�F�<�edE3 c��T-V�k3j��woC�<Y�+�)w
�@�M,:�tak�jJ�<��#�;�(95-��G��E+i�D�<�F���gc��C�#�4P��BI�T�<���Z<���0�聹�JQ� �TV�<A&CQq@��1��B��`CP�P�<� |��ѧڬ>�TՋq	�v�<�7"O�	�/�NlV�إ�}�(���"OH,H��W/q:�Ф�VoaHp[�"OR� BJT/9�2)�$,���P&"O�1�fԫ�� i�l�<qn���"O���m<l���r��z�JP��"OT��O�TCT���Q�[���w"O��g�G�\���*��6��H�"O)CQ��69A^��ꊧ1��d��"O�-@C腃G���F`�>��p`1"O��R��D-����L���
�:E"O�i��j�'d4�IQ>4r�ɛ�"O29�ʄ2H�	@�
�:fU��b�"Od�R�;B<E�6��*7֔�"O`9��%�I�a�M�f% A�"OB�'�L�m޾K�� <Rp���"O^˅� �40N�ʕ�=j��j$"O�1I%�Ĉ:��ؐX�~�Sp�'c�O@������L�僦]�> Z�"O��V��of��4F�j�����"Omѥ�T��xr��[�@�6Y�"O4�X���yz��V�A+��)2"OVii�c�N�Եp���d(�C"O ��C"��|���J 7��(��"O����A3q���I��ZW����"O�Y�Р��H([���>Tڰq�"O@�r�-ן
(��aڨ(U�,�g"O$�Q%dr�X�Um��mT�I"�"O���uMT8��,Q-0\\ f"O��QqaO�2�LX
�J�&��s6"O~a�! �<r��Dx�j��"OM���E3�d=za�չ*�(��1"O��AE�9��)2ɶG��`��"OZ�C��ǓEs��ЂN����2"OVpQ*ܗds�����7��M�A"Ol�H�b6�l����F����"O���w�ĉP|�b�x�pi��"ON)p#D�`�x���]ȀI9�"O,Q���B���}�MПY�i�b"O>�����2x�E���`�^�6"O8��ą��|��H�P:z5�]�"O��"e 'o�Y��Œ䰩�"OX:B�L�6���g�7�~�"O"ǂ>Q0�$�2�2P�5"O���MR	��8�G�$-3���"O����ɷ�(f�-I7l{�"O6L���)�J�(��΂� ��"O<�ʠ����&���̉�j��!"O���,�����^�Q����"O�%����>�9�1��S�=V"O�ň�D6^9t�b����/��)t"O�u������A�c�f�`1�C"O�5���D�h" X��B�8H��yW"O�4A��ԣ�x(A� ڪ}��q��"ODI���G7)��x&B.Wv��q"O���ɏ�5ȉ��O�Ji�`;$"O"	Yg'�c ��&N�21��#a"O�HI��TU�fc.�0C9���G"O D��+R�X �0��'	0��a�"O8[#X�K�4U"����j�À"O�l4�˺΂r�a�4���:�"O�9sŻ2��Z�%Dr�:�2,�V�<YVMë
N$� AO��v��%�ekR�<ׁ�8,�:¡��8H��{"K�O�<� 議6��D�TT�v�6��Q�P"OZ:5����0N̩,}��"O&pѶjF[���h�M�#mb:i�"O�HF閠
��́Q��Pµ*"O���c,����51��O,d���"O9h�
��A/�=�F퇱W>>�"O؄BVf$IҲ���� �2/�!��"OV� O�*y�F�R�T#:����"O����Y�u�p+'��)���P"O&�rR�ȨJ	� g�˫nDxt�"O:s�5u(lt�r��������"O>i�'W-N�.��RN4|�4���"O��B�!QoC@(��cS'T�lݺ&"O�#��
�><v�ӝw �+"OL�c��t%�P����A��"Ot�W�F�;X�I���ѲsW"OB}kq��
U��\���Y�����y'AQ��I��ʺk����)F�y���)�m�ǖ_�N�V
��y2��z��S��;��)�
R��y2��<��@�l�*fgX�E��yϨ>j�%���Y�D �kO�y�+�4S��p���^Ӡ��4ʸ�y��\1�Px)�,e�t50���	�y�V.\�4�Z���U��7�HyR�'� A3.1_��l�eO��1�P���'ڂd���Ʈe��1�n�#^B���'$�-��+�n6�������'��L�''��@�D	�i�R�����"��9�'��Ȳ�A�9��aX�
�����'�l�+�$Q�5�  ����[P�':�QbRnW�PJ��A �λ��͢�'c�K��B�A��!�*�ip.H��'Um0��ݽT�E(���YE�AZ�'���ᱪY"���p�h�?I�����'-*���V�`��DM�C���8
�'��P�.�1T�Nh��H�G�>%�	�'�]���ٕxTi!��m�P�	�'���x��K��Y��`���z�'iY�N��L�Q�jZ�F����
�'}�[����@*􁡂�.<�}�	�')�]�C��wg��0AE@4/	���	�'U* �����nD�a��̱6��X	�'�^��a�ݩM��iv��+2�� 	�'���ç�Ԭ4�V�xUm�
2Ӵu��'f��Ul��^���O�27"����'Y|��ˏ����f�ʬ+���	�'?H�)�΄�o�������	�'��E���/M�z��r�'��m��'�L�Qq�׿���"A@�3 "܀�'Iv@8��Q�W'�hP��u�����'F��¨�	{m�,�4��#Y9xYR
�'���#5ώ5Urt��ʌWMr}	
�'D�u�!��IQ�A<$Zԓ
�'!�kЇ�<,�.��sa��Q@��#	�'Z-H��䬘�ӈM�J��5��'�PQrE#x��mj6�ͽ94�0�'�BxqpCF}F�s�OX>7���	�'| 8@���_5v1�zB��	�'*x!b�"�.��SY��ub�M$D�|s�DCZ��� ��:���%E!D�$t.ηD�e*窑
<ܸhdm)D�p��Z.2r5��@n���'D��� n���l��X�.h��O D�� ��S6�׆:�F��*E%a�xP�"O�  �L 	x^���	�F���w"O�lHD Ǩ(UPXA��)<v��[T"OҔ�猼bd�Jր��#p��$"O�ܓd18�M)"�K2'e�t��"O��� I��Xq�K�l@򠸗"O8�zpKL�.�tT���&J\ Tq��'�ɤCٶ���4w�nKB`J:x�C�ɇx'��#�I*@�����R�nC�	 =?�T�2ꟜKY�V�Հ+/B�I<A���q�ǔ5�:��"�$r��C�IZ�5�@
X�����C��sNhbS6c�ÈR�_;�C��C��1�Q"�Ҽq��� }�C�I�1������n]`�/2��C�	�}��"��OIt���ͦk�V��^��h��i��7�e�2BtT.�r"O̵	TN�93ߐ4�0��\F ��T"Oh�Sָ)��=����� 3
�bF"O�9¨UF��Zc��X�Ց"O�ᒵ�I���=�iG�;�=+�"O�h��U7��ȦG�;Z_��yE�����ɳH�&�[E	C�dìq�Ae�C��B�	�{�����F,s�11�B�8I�4�4�E�*H.�C�k�.��6m&�S��M�!-a��@��A��O�M�<i�J,ׂi��9���cp(�R�<��*U�z��2!�Ɉr����șK�<1"E�^�y�sΓ�:�4�ԏb�<HXY`�Y�%cǾ	��m��]�<��(I9�j�Ç �q5<4J��Z�<A�O�<hd�������l�*�(GV�<����Mg��5�"&��@�v �l�<y�hԟ����c�ɝ`]��!a$�e��<P�}���^u����Ǔ�hp�PD�D�yI �q�,�R�c��4���y�ˋ�_�fibr��d�]�k\$�y�
�yi
�	MF �b�W
�y���)�FĒ�	�?D��������yRލTxd��B ;��0����1�yb��C?T��򠁫(��8QRf�'�y"���6Lñ�(5�ܚ�%�yb�E� �B eҹ9�����yB(S��+��:
}�@�ҍ��y"�1?�x�������򋗙�yʀ�}��%)P	Уz&��+��݈�ybn
0w'"�B�� �puC��¬�yB D!}tv@�T���e�$��E ߊ�y�C�9^�	9��~V8��+���y"� GeV�j����	Պ�y���D�=6�,��%#� YI���r�!�U�S���#D��:#D��5�!��X_d��$c��c��h0V�!�dC6��i�SfX�G�4���#	)�!���&ixBX F �-�i{���
t!��ˡK�X���]t� ��!ʧTP!򤏢NT8�+���x�0�
6!�dJF*��,ՖVm����Oϓ�!�Ĭ8�|qz ψ�W֝������!�O����R=#߸6�J,$�!�$Dn.AkS�	?ђz�O��!�$�l�v$��J���/�'v!�DZ�VݙfIV*Pjj���O�!�ć�:��(��(�*<br�b�-ʝ�!�� ��Ǧ�Y�e��pѩ�"O�ݣS�	�$�)��Ō��`#�"O�X����[D����~�\���'y�äXA�a��I�h�-���p!��Ɨ+�Feۗ��} �A��!'Y!��0n��,x��\#c!��b�e%<�!�ʾ?��TP�D�+[�P��$M�1O���D�y�@!�P�T�^)��b�j!�d�U%Z�����#�>�A���$�!�ď�f2����I�ζ��!7�!�dS5�b��@�O�9�:�
a�W�M�!�$��Q�4�����=�HM�1/��c�!�!!�L������/I�D�EM�X�!�9�4�:�"�5�E��l׮`!�D��Ih��l' ���r�&�'D�!�$�Obu���	�T���`CaY(\*5k��+LOp��3d[r�Rp@� '~L��8s"O���#@o�a�@��=��u"OI#+��M
�nԦ:���AY� ������dF�P���9n7FB�	�?YLŠb�`��9)��Z�L�4B�	1l�8��
ĳl�\����<@$�IQ���d�ą �r���C�@��p�"&�^�BOd��1O��{��\�}B�8إ"O�!b7�G�?�x��vj�Y "O
T!��I������ :n�
��"On���hE�k"���b�Ɛ��"O�\��
�J0,�
Fx�P�"O��w"�{gF�I��D�^`��D"O�Q@��ű#�L��(�\AN5�"O����\n�HmU�P�Rq#�"O4H"B\7GKna���C c��paA�\H<!�.ɀ}��:���*'�� UH�<�Fg�*e|a��ʞ)~�l��g��D�<Q��,cx��֎�)H�ݙ@�j�<Y���3l��ae�Q�Y�p�0�QN�<�&WL�@@�D?���Ek�d�<	�?f:л�/��a��l�V$Rf�<q��ݏF5��*�#x���m�G�<Q�����ՉR&V"5�(E�	l�<� *A�V��5��Ú��كEA��<�q����e��*�` T(��az�<�P�1U�^�:!�r<L��n�s�d!�S�'Y�b�V���V@�A'iZ!?4U��yV�{+ɕW%��dǝBfi�ȓR���É��r��]b��[x�@��{�����ڧ/0�d3!��(8�l��|B�(��28��l�%e��b���ȓ~-��� �r�hCDߔ;�����hO�>�oOL_Ū��PY�e�vl�2,D��T#G�[�^ �nʙ�|{�(D�8z*��V�|(XѮ��Z��%D�\`���1;7�ă�GR2V�B%��� D�<����Yz�9����;Ze*���=D���㨞�~M���@�K>9� =D�|�Ī�"5E�|yȦJ��l���<D��ʤeE�v^���kFIG��F�:D�L#D�ʦ^���1�J�#0G�(�8D��y́���m:�����ЫQN7D�|賫ͩ&�@3a���B�S�/D�j'��&�fԠS��=�,� d'/D�� tBX�&� *���9X��*D�`:4�W�"�3���4�����*D�l��B7���*G �(E� 	�3�=D�� X��� (�z��`&���x`�"O�|H�/ Kخ��d��C6���"Ollc�e���8 @m�|F�-��"O|]+r�:4yda�m����ض"O��)6��BE�7�d�`�a�"O"������������Y�T�"O��[e��O�i!T�ú��D�#"O�$R`�C��ȅj��
��h%"O���PC�F�F����R��I"O>YbV��	W��L���"�R"Oz���ꚹR}L� f�ƱI���r�"O-�G����m���:zh�C"OСCv�Q�+ j좱���h�"O����	K�.�
��<y�J��"O.L�w�ϠqV��T@6�F"O�e�a��]�6l�'�+�(��D"O��HU��y͜�Bo�ro�$��"O@��(�4M��P�.O@Uf�1"OL��g)�&nT
wnY�IPn��g"O�(W�O\�� `��p:��r"O qpe)_`���	�l��	(�ջ"O���� *vNPMʂk�"Ps"Ozkd\�`�����	�#30���"O�Z�%r$���5ƒ�1���&"OP�
0�ȨR�X����LR��"O̔[uN������4" 1��"O�[R>/#Ds�놈M�����"O1�#d�(,���p��=X���#"O��u�O�m�&�*�i^5}��� �"O�[䁔�n�F�3�ǜ |�Ӵ"O�=���?+H�zQ�V�v���"OV��w�K&E�JT��b�0�"O�4�t�T(S�hժV��HEn��"O�)�F�,s ͊Ц�B:�t"O�HpԮ�d���� 3~��	�"O.]y'�17\	J�� u[`R"O����ɼb�f�a����c6�C�"O�x"&�+
Q��/��WN���"O|;��K���O�;dP`�"O�� ��\�V]\�Bv���)o~��"O�E��hޝ%"����(s��"O�#��J�!�d��̙I��iB"O� ��"K t��ԨaK�7�&�Y�"O�LY���*h/�P���%;ݖ�P�"Op����*�fP)Æ����8�"O��� J/>8)�"G/h�J1��"O�[��c��H���s�R�U"Oxe�F�W�`�&=9���YvI��"O��{��<`���g��d?��h�"O��P���NTȧ.�,4^���"O���Ċ�	Y��S-��L�0"O屖��-3�͐A�z��1�'"OQ�@@��
�؄<P�4!t'���y"M֢�| `��E�Y�F�"K�>�yb��� 8����ݜYuH�h�$�y���`�*rR��A��\r��1�yrl�ch�y�ÁNk��YXq�H2�yr��h���$���3����y���>mT�e����.���x��\�y��q����+E�8��B!�#�yrB����H���'Sx��ʔ
�y�h_4yC����:bJ(�e����ybl�DE��c��	�G���1���y"�C�,�8����F�;���x$�ȼ�y
� "�e(W&�K�)9N1r"Oꕊ���k���q��V�k���"O怣��##���+���	���"O�K�c��8i���=_�qIs*O��1Wčj��� �/+�x�K�'���pWgJ.$�h13n�o1ܕ��'7p�[�$�\�	��_7b�#	�'��|�@B3�D�f��*x��'A�\ w�?T�\|�rh	Bj]��'�p#Χ@\��bwB�� ��3�'��PiD눛@��aF"�pO~� �'*!8!���~�6txrG��k�e�'8 ��v�0���\�I	�'�j��B�%�P�� �D-OL*�J�'�\;���,>y\8�W���N���'��Њ��4�d����ÆL~&�;�'Ѭ����G-E�$���]�<QV��'8�@4۾a��ʎ6sB���'L	� g^��^�B��6�h��'�&4h�!�73, a�L�5�t�`�'sl�Z��Ӄ-a0��P?3Yڹ��'����"B⢈S�%ګ'nb�s�'�\���հߦ�;%a�"V��+�'������}� �gF-� ���'���pA��hSNȳ�Lέ�����'�>űC<�P02J�z;��*D�@*e��*-e4ѩ l��6�0� v�.D��#��]�&ߐ��\7���/D���4�A"K��H�EU1<Uj��,D��r��32t(q �M?i ���T�-D�Hi��� V���)4�� �?D�\�KӖ+'zcCX,6��}�h0D� 9!
��=�x�S��S�O�D�[��(D�ZG�.B��UEЅeUdA'D�|V"@F�`���
l�2m�gj*D��z�H��w�pIi����A|)��m*D�ȳb���GEpTʁ
 � �\bC$D�d�"!�-i�(�U��JF"�ZR�=D�$d�1�֡"7�Y--���*8D��hp��uo����Y��a{�	"D�����<x�
���k�4;��q�ь=D�P����6��}rT�Ԗ)׺u�'>D����ӨG�t4�5��0zf�q��&D�L�P�߈E[��W�Z�r���h�`&D��S��-w�|}��#�Z����$D������g��Mx��T�D���rG!D��A5D٥y�8r�ӭV�"Ӳ>D�Z2�ŎB��Sj�X��,�1*=D��9sJ�R0���G�!~���j9D�x@�o��N�gH�=ߊ�8r@7D�`q���5bP��o��.m"��"D���E��<^࠴z�0��!rb D�8��U5Du��	�CV�Q]��>D�У��u)>��U	�m��?D�\����	�j��Ȩ���!��"D��@

 cX��I�DǆJҨq�%D����2';V�#"gE�U'�H��$D�L)��£l%.y� �f�r�)G.$D� ���öH���r`Àq`�5#b?D��P@ǎs�`Ǡž�����;D��A G8"@�@��P�|����-D�����,��h����	mJ��DH*D�4а��:	a���c�4ٚ�{�%D�;C �:���v��f�4Y�'$D�� �$�ƀt���F3�eQ"O{�� 'O�#��D�DB�&�� �ȓ3^��ST�.s�@�$�C�h���ȓ#;&ة`po.0���X�ST��Z���qqn�k�  $Z�L���Xy����-�!i�f�ېDX0M��%�ȓ	��x!ՇV��؀�$W3�༇�H\�� ���'��{3��X�y��	�,:5eA
\�ԭ���)Rb�4���
h��H/l0�������X%�ȓu�=i-ߢkUҔ�fO�oT����J��`�s��2K*�y�i
PFʡ�ȓ#ޞ�8d�N(Cqn�����%�ȓ2iVE�,�;0QN���A�[�z�ȓ]b���@W�3`P�2vG�Z��^�A�D��-.6�48wAA>x����Md`R���6����!B1M�֍�ȓI�R�0n�7Y �x�蟭B��чȓt������Z�LD a����F��� �mS�(��0-US�����P��F�f;�q�fW�!�ҭ�ȓw�ؽ�#��>\ �P@Ѥy�̉�ȓ-�H����_Neѐ�^PB����@yFd�G0bUQe�W�R����*S6�#�P6{ڄ��AY�°�ȓ�(y� �N�<T�U@���W��ȓI������p
 p�9��(�ȓu��p2�ŅN&R��@�+�v��ȓC���㐂���zu{B�� bK\�ȓ�~m"��;"�5��\!�6�����Q�D���k�h�ф� fLI�ȓ^rt07)̍{yj��V�
�Ndh�������M5W�~j�mJ-l(���]d�8�@�'̮��% �8,�L�ȓb���q�]��Б�@эV6���F�:��%#����h�k�I��|��F�F$J�`� 9c'���ȓq��|�K�tx4�c&ԊnO��ȓ���`��_]  IL~��$��$բ�0��^�V�*$8�!�U*:��ȓf��k��
f+D���BP��HH��$���Zv䐤_�<��P�m9���ȓ0E�{��B!J���ERy�ȓQƤ�#c�J-��ЄmI\r^,�ȓ4�
|�����.�lyXF�4�*\��)��2gM ��y���Q����@H��R -يz�R�ȧ"	C�f@�ȓg	X��Tj>Z�@�指j�-�ȓu�b���%(�܉����?��ȓ2Xi�F�Y-X!�E�M�*-����8��H��CRUIb�23V��ȓ�4Z��حGк���$־uJ^مȓgg�����<-����U�*�ȓ�ZY �h�.*w���bHES����a�f���	�ou|([r���.A�ȓPhB�k%'�IVؐR0�{�Z���z��!���C(�U��'A$Pgj���T�l02���������k��`��w7>A��ϔT���rr���,��ه�v���2�A{2�����:�h��ȓ=�Vd�A�BB0�Vϔ��b-��P��T��0���a���;��$�ȓ{F0�F*P�dt鳆�7Qv�����
`�6�x�b���>���S�? 0�K�P<o�<tI�NV�d�N�A�"O�У��UP\(�"o�"��Ph#"OF��f�0G¼G�@�l�:5��"OL٩%䙐S]�����1�"OP�IWB'X�����j^"���"Of))`�Ҭ}�*	а��5����"O^Pǯ�D�,����
*t�"O��0��wg��R'Q�E�x"OX��JU�s�� ����`��S"Oڐ�䬎� %�q�������B"Oʥ���O�W_�a���˄��"O����(�;T�嚁Ȋ�ؐ"Ol� 	�<��	zB�
9tL�r"O���2*E��hIx�*�|�2�"O��#3bF#\`���c@�d�
�!"OD�C�㚻;RL�#ʛb�*Ac�"O��SB�� @pn��A�\�z�
�kA"O�|B1D˭!8\�҆�2 �kR"O왣�bΒn���f�5�B��'"Ol\��,7����0��	IJ���"O�d`���,t��m!Vګ5.ެH�"O�\Ô�%v0Q�l���` �"O�%��H���a;�H�����"Ot4@5���q)��y�I-�b}�"O�=�7�߲)]��1���:^I�l�"O��;U愣4����ӬJ�B�˙ m!���敐A�ն.�����B�!��K�:�╻�n�!D����`:N!�ߋg�4R�)X1_	f4��.K/Y[!�D�Z_esc�<��%��Ԩ1B!�D+y��APP
�*u��q&l�K6!�D ~��q�W�YEkx�RP�2y!�d�9JW���7G½3V�U"���!�D�<�f�I���(5U5 GJ^�!�$��<�y@m�ONƍ�!��
1!�d����d�D�+`���!�D�|�hA&�͠r:��#OP!��u@i�Al�6*��M��2C!�)�>��p�޳O؀0����)a!�DX�HbT���p���ST	��m}!�d�5�X@�C��b�������0r!���>�,E#5���_��X��拸K{!�dQ�F%��&�d���&��-Fk!�$��3����F��� Q��*.N�!�]�q�t�j�/�5������=w�!�$�>/���LD�2���xe�L:%�!�h�n!�u.1�h��`O�x!�D\�d��Ab@�»G�R���@�l�!��RPұ;�L
F�z)�."!�dQ?����K#}�����śG�!�ˈ}g��9T Z"5�$�
�I^7'�!��NMZָ��=4���ڑ���!��7(�|��U�J�0�J��_�d�!�dK�[6�� ��M����yRQ6�!��B $M�d�m�|XA�	�1�!��l�D���O0(���PMѪ/�!�䗣#��J�`߱Mư�
ba@�\�!�dI�rK\�;3���/.5���
�8�!��0D��&H���E�$*I�!�r�x�j�o��DmtU;1����!��S�\(�&�޵e�(	6,Z�1�!�䙖L�.9B�]�v�`�� N�t�!��c�����?�0�Y'��!�$Y�x��E%t��}��Pe�!�� ��,���|�
C$�֠"Oz�{'�^2U���p̋"� ��W"O��#� �$�	�h��`�����"O��G�6EC�8���^*���"O�1�ޫs�"cƊ$ �j���"O�0�q�T�r����'@;��e��"O:��R"ڇx�l��� ��W	^��"O �W���l��"7b/Z�Z�d"Op�q�o�~# �Z�f^�S�d�!"OB`��o�
���T5�`!)�"O~U�j�|����G�T��!�"O��8�`8i��� 3R�%��Dۅ"O������C�t��d T����"O���.��p���5
n�@�"O�-x���y�Af�D�����"O����"\�D<��AW�K��%�R"O\��C�������ۥ>�:%iT"O�S��	�w#� �5LG�p�z�z�"O�ْ�4DfY�R�W�
��"O����W)Fz8�sPĊ!{�`*Q"O�l R�̾]����T5!�"O$$C���"x�$���J�F�Xq�"O�,0�钍J*v-K�ד�и��"O` �'��|dF�
��s�ܑ��"O�D�W)��]�����Y�"O�YŀQ�75�a�t�U>P��"O���/F��lA��O�`Is�"O�9�aI���]1A��Lؘ)��"O^�m� g8��Q�A�����'Z�u;��ʞ���i��K+H q�'pT�4�/<�� u��\[b$�'�������VH,������i��}��'�6Cw��'WH���"`'[��)�'����&���Y�(���ɣ&M�1I
�'��E��AOФ�(�H��	�'\����R�#�F�P1�OQ�u�	�'y���/�{�rU`�F\�,h��':X��$i��F���#F�Q�\�z�a�'*�IBC�/�p�I��
�O8�L��'�
� ���|%ȝ�g���v"OR�bҌ_.���B�0W�ds�"O�H2��ۀ;`��P.S^�� �"O�<���#H�������q�"O
!�1$��Ș������=�"O��ď���J���77����"O:������H�F�3R�9�"Ox�eH�"Od-�BEɽ%d�i!"Ov,�'�K�["�=ʀ�	�SRjU� "ON���#�5-cT����<Lf��"O�� q""Jآ}kQ��$8��%"O��y��V� {��j`���69�Y�"O��@N�4��`���mD��3�"O��#���>�)2��:e�|CT/�<��(R9-҈�j������R�<�CǳH��Ͳ��A�{�LѰ�%�J�<1E
�/uV���ȟ�F�����I�<�5(}\�8Єĕ��i�t
IZ�<�.�P�+�#Õ-;��"��U�<	s�S�V���i�l�6xB�괤�i�<��dZ�U$>��#��p <��q$q�<I��[3���P�Ô184��� EC�<� Ŗ�-��YV�74�s�JU�<�C�J�Y�0�; ��,5���i6��v�<�Q��zBl���ǬI��mP�\�<� ��ckQ�:��ِ�G�w�X�r"O> �T���k^)R�Ei�I��"O��ؑ'�
;��;SjQ�q[�ı�"OE91�ˡ�Hjs)C�~��m�"OB�c���L��������?7��v"O`�h�b��uB�h��A�:D:4�C`"OQ�s� W��ٻ�j��Y��ж"O�0�0f-�"�F�\�əU"O ��l�$>�<��BչO�t�8s"O�`��,�
G�pa���T��}� "O�95���T�[��o`P5��"O���2�$�� ��=Pv�q"Ohă  K%Q�EPQ�o��j�"O^P�s!�[�xMRfL"�XG"O�Ƞ�ӌ�� �oT>"ذ�0�"O�Ae��z�R
6�ѩ3��@�"O8���&Fn��Xe0Z����`"ORp�b��f^���mL8f��Yk�"O�1)�M:n��6f�'Aq�i"O�#v�Ѕ'.��t. �UpiC&"O��sm���0���ʺC�T	�"O����kO�#Ln�A�%٪_9X IF"OMk� ��@�� ��ڸ.� a�g"OLa���F6ֵ�G��Pa$�h�"O�@ѕ���-)�M;iT<�"O�d9���%�3�G{Ch��"Oظ���A)���q�ʞ�',P=��"O��qD*�S,s"�4Q��<A"O�ۅ��~��k�� "��{�"O$4s�",.��d����o�� au"O&�9�c1��B���)��(��"O�$�����.��g T!|�\#�"O^ȋ�b.�Qb@�E���8"O�1Q�	k`�@d�I�e��q"O(���8E��"�n �=� `Rv"O*�0�C@~�h�P1��#1���H�"O\a.�r��|�c�)<���&"OTy���f3���ə�K���`"O��3ѥ�!v�|�	D%�ڞ�Y%"O�D�]2tZ(}�D�0�.���"O�dR"@��t�p�×�E�����"O ��Q�	x��)���	�H�A(�'��i�E"C�-Z ��Wo�L��
�'F6��e���e!I�-ZQ��
�'�6s���G,�U��F�X�hA�
�' ��i��J�N.�q���T^^�
�'�b4B���`Ġ�fT���aY
�'�h,�Z=m�8��^:jN=�	�'�"���]�F.��@"b���y	�'x��Qn�c�b��-C�T��'Ѱ%×��m�x(�U�9=o�c�'��1���]ft�;�&�2%����'l�iw��%i�L����Ժv|����'{\�!� <Z[t0�l�\���'�"Y���Bi���� �1>t�3�'mv�(�@��:d^U(�B.-�Z��'����Co�](qk��"��'���$�>l92���mmD(�'�¼�Dj�T�Ri�q%I2]�pP��'k@=[�͔%9"��&+.ʈ+�'���i"���">��֭�&�@q�'{�A(�*2h�f��^�q�'?H�مdЁ{$�����9[��m��'�t�{Soڀ=*�i��WJ����� �H)w�%'L��:q�e�j%3"O<��(� ~f,��?"�YC�"O��3�%7�P�'M)�i��"O���Ɲ�29�)�PᘋvZ��a"O0 a�;��xV%���2�"O̴B2f�d�¤"O�@z95"O��� ���R�D<K�n�X[NX#�"OP1+V�'p�MIs.�W��Y�"Oh0���ʴSj��7��l���{q"O\$iņ�cHVJAM¾fh�"O�DRD�ΔsO<�Y�,]�(r4�Be"O��ʗ���L�aq�0�&T�C"Of죴&� s�Ѩ�+8� ȓ�"O�hï���ʧ��J,��"O��K���2[$�1�E��m���q3"OF�sF���DI4�"R���T��)�"O��"ĺSI�-㰬Z�XK�1D"O��!��
>;,�E�IX@�1K"OR���j���((4��9=(� �"O�k�L��e�á�>-{�"O�� ��"8萭�b@��I�D"O�A2łƷfF��*$�5����E"O��jR�I�l%Nu�#Ǚ
��"O�a9@/ƼSPb)[UBP�*�*i��"Ox��5�^�f)�[�&R�;V:�)�"O����܋w�r�H0��2 0�"O�R��2z��Q��/�@��"O����+�,B��D(fLM"02���"O��y�2L8���!�͒`oR���"O��:�g�X�GHX'R�m#v"O���\�j�`qGQ$5�n�b"OZ�9����l��cM1͈�!"O��c�cS-X�PAnP�X�\��"O`s�F@'ljh��䉵B��P�"OP��⁐���0S�\���Ź�"O��`���Z��\�3$�>�h	�"O~ţq#�4H Π���$0�D)H;�yR�a6@2wD1Q��Q𓩁'�y����T�:h+�PMD:�۔	�y�g�r��SG����!�?�yB��3-���)�"�>����c�Ӣ�yB٧T�hQ��A�i���C�����y�ّBs8̊���l.��a�&D��y�#��"vT)�NWS혩�KH-�y`ѱtP ��T��Q�ȸ���:�y"VV�<�hé\��8����yRc�$HF Q+�F!f���*�CP;�y���,���J
1�U�G��y2e��"�U�T��vs������y���y���`/ӺXVB��h)�y�nO�,lh�
�8{�B���(�yBmB�'�2��7$whu6I ��y��gL��g�ζ����u�D��y2��l�fq&&��Q�\Җϝ��y2��.Y�a�M*��|�F����y���,���*#�P6j�� B�I�K���#�ҿe���
ԨA�C���Z�(��K�%J��%�&�;D�xX!(�p�j��5���3?D�|�掕#]:P����~ ����*D��
�jP�4X�H�뙿~��H�)D��x�H޹�2�)�'^[~�c&�(D�$�č�&|Ӹy���/?�Ĺ�!'D�d�P`^�b1!��k�=B��@z�(D�� �yC����?,,2��,T� ��5"O�5����`+�iق&��f-���!D���BϱA�\�tƖ#�)	q/?D�pۇ�'ISf�җ̗�,K�3Bl*D�� b�̞,�C2�Vr��Mj��(D�в� 	h+VD��Ȕ�nܝ;0!(D��P��#�F�3��5%н� K%D�0s ��i:i[&��83R��(�%D��R��H�B�0�hQ�R3<ɒ'D� �3� v�>:�.?)�4�w�'D�p�TB�W|DT���U[]�-	b*%D��CMY; ���20ˈ-H3h[��%D��zƤ�4^0n�1&B�I�Ac>D�(�@`�&o���Z!��$^T`؄�:D��{��%Uר����I�~q�8D��z��d�� �c!\5\5 R�e6D��1ej�K�����'*$��
/D��)�(W�D�`�Q/�<g��i!%�1D�� ag�,�����JÆ44�uz��.D���#*�),m���5@��?���H,D���Ǧ��	�JYs�o8I�y�i$D����M?jn�4BAI�5=�\���."D�(h�N�*F,s��W�FbB��1�"D�8IEV0�|�f�՗(�<)[ը4D�kƥ��\i�*�1B�s�%D�<�D�M�a����aM$R2]���5D�0��*~m�q�`�H�]���3D�4Bbm/z0lE��mett(vK1D���eJ��PΞ� ��Ԙ3X\�Vh4D��V���F:�� ޜW�B�'D���+ŁSɎx�X�
�l@��)T� �ϕ.s1�  �fy��"OZ0��@�� �Pf���v͎�2�"O����W4>��+oˉI�T��"O�P
�ʍ%?,H
/\,n�"�Cc"O�}�f��"naf��c��!t�Ss"O��3"�
�8f}j%#�="���"O�p��jŜq]��r�,ΤH��S�"O�q� A�!n��9��L�,h9�P"O�P�
Y�{l,RՃ
c��)�r"OvD�e��<��Q2P#�042� �p"O(�K3��h��q�e��~��"O��i�L�,�QT���R�����"O�dK��Ȋ;ƞ�ap�s\`"Oέa�D��02�q`�?Cָ��"Ou�4��f�j�*B�H�O�{p"O<��B��3ڰ� ���/G���"O����/�3ٚ���?5�T�B�"O��jl�Oժ�SB)���ji�"O��UF��+��U�ڭ*�"Oҍⱅ[�IRR\�B�#�tx@W"O�c�� "zj��	�S�����"OH�A�eH4I�(G�.r���"O�=�7�ؙ,ܬ� �ч&epX�1"O(u!�lG�Aʤ���(K(5,1q"O<��H�-۬�ʄhė	T�;�"O"��d��B�b�@��H�JI欀�"O�x�R�'20�0�x�с�Z��yҭ�\Snh�Sk܉T�� ��HT��y�EЇr�$�E'[��SsW#�yB���sb`�V��K�KM�y��S2#�D��V��B<�����yҪ]|6���!�%�"t0w!V��y�c-b������I��<���Ǐ�y
� ���ŏ�9�����؉q�["O��b.��`���a �A�{���4"O���E��� ��Kց4���c7"O�s6d��`�[�M2S�@x�p"O@�YL�'�ڜR�#D�#�e"O�q9�'� ��+t�M�k򈉡�"O��yp�M��|4Z$a��HQh3"O`����j<$Y8�������"Ozh����!av�+�=ˎ�"O��dB;X	�-��IM� h��"OЈK7�*q�Xy7i�d|��7"Oƕq%�� p6x�ǟ��l<��"O�۠	фgĭ��	�\�4pA"O�[P�n<�Fm�.X�H�#"O��'��]����&�$x�"O�l�P����-I���dW"O�|�1���SX��Q�ΥZF�;"Or�+q��'P�\x��J�aOD  "O��JcA�1[,&�D�Gw��ᐁ"O�V�88�.�#�a��h�P"�c�q�<9���!v�n�Hc"Ɔ!�j�Qw`�q�<�ph!�l���I���9� Zm�<���G�P�bSf�#[��y�V�	S�<ѕ�_��ǋl�ͳ���s<���4<|�:f@�Dh�
��ȓXl
�9�"P��"0A��L~q��ȓ!��� dc�+P��H4HC�#�����m \<b���;�^=��A�k��Ʌ�)r�`{�,�44���I��
>n�����a����${�&U�g��>S�ه�"(��Ί�!U@9ɴnL0�4,�ȓ�`H*����f%�1&e>����9�Լ�K��@}y��M%z�ꡅȓ/��@C��A	�Lx�T�"F����ȓKƄ� d�X�K㊹�u針x����b��3"�A2H,XR"�G�/z�ȓ_(���Λ�lf�Y��Eȋ��%��go���k��S��i���V�`��ȓBe �q1�F�!���z���}�"L��!a"�3�D����	@u���`�j}�� d��02��8�~�{F��Ch.��ȓb�Z'G��\6�{�G
9QJ�ȓW���"��� 	$�s`��(d�ld�ȓb�ְ�F��"W\݋׮�&R'>Y�ȓJ�U@���G^��Sr�ɺIBP�����`�4�$Kw�m�(U�A$6A�ȓ{��I�Vd�{v��X�,ūI�ʰ�ȓ�Di���&Z&,�Dc0V ��r���"-*�L@c�LEC�jm�ȓU^�j䃋�5 ���S�P(�ȓA5�͖<C��t���� v�\U��!}\�qD�wc���"��%$�`��l��D�"OX2(��kT�@k��m���2! �h�L�l��B�	J1SlƫX���R���K�B�I�q ����ʺy������pB�ɛ�(���Mbb�`Wi�%?�jB�	�K��$	1�ӥ18�R� EKfB� 
����o�j	���TG�NB������0|1�"T)
d�n"D� :�d���[��h`��-"D�����_1)�ұ�P��1��Q"�3D�P�n˻���#�|����.0D��s�ǪYyhÒ�P1^1�E�P�,D�� �<{�B��-h:]�&	#5}���"O T����}~z���F�rt�T"O���ҵG�Rh���N�Gq�#�"Ob5Ӣ��%�5���Q&D����"O>��V�̒`��B2��B��Ѩ�"OĥR��i��IS@�0�lt��"O�����H���%ǒq�Z�*"O�#B)�
R��-b�J 
F����F"O�!zT�ل�(�; i���&L"O2�R̉B9~`��Aږg�E(�"O���� 4^"�TZ҆�~I�"O
���h��+�fr}�D�U"O蹀���s � c�/��ev�X�v"O�cAd��n!"GA �h��"OHp �v�,|�R�
J2L�T"Ojp����_<B5r��XB��"O&��D�tҀ��"Ў�L�Re"O$���f�	l�����i�%c4"O.��7I�O�as�G[��v"O���0��)y����HJ���"O���4GQ�)g��Ī�6/3��9�"O������i��ޤM!���"OJQi��0F�X|��İ7��;�"O>��a@:B*�Q�,�=��"O��h��ǎ7���т-�V@b�"O�yB1`�	�#ɁS�` 0"O��h&nT�&ޢ��g���a�"O��zE�UY*4�ȷ�K��!kw"O�M�&g�f A��#�| f�"Od)�A�	�jX\�"a1���A"O�$��$�@���I���[�"O8�;!e�t_�5�����q��"Ondc��#U:H3bl����V"OT)މ��T�Ԡ�7n��Q"O,т�l �z<�qp؊-'l�`c"O��*�GW	�e*�l  l#-q"On��CM�sH� 8K�4)*�P�"O��eՔv{L1���ɾ?��<�"O\{V�E�r�ZdJq�Ӫ|�q��"O�P��خ#FD�����$_���&"O�IB"�!$�\���p��h �"O��D�0S�+�eT�?�U8�"O�QĥL�sIH ��'|k֝Z�"O��yA���!��CVg3\��"O8���s�$���B�H`V"OlU�r��$.x^DP�*Pg��E"ORa� �f�����,�Yj�"O��ТڶJn )��ئ�W"On�� �Hcֹ�4�(w���Ҕ"O|��!��$|1;զU�A��@"O�ջDf�mA8�k�ΨC�ʄ�e"O9 �.���$�`�\܌Ԫ�"O2���w����@�32�"��"OXʣf����`n��-��tJd"Ox,x��ӽn��i�ҍ�X
��"O�4y!t�M����k\Hx�"Oh�����'*�b��� �6'K���3"O܁��KӇt�؁ĎP�|L�b "OX���U:K�^��ƭ[`b�à"O���oE�*��yW6mS�@��"Ob�z��A�x�����L00i�"On�y㠟,+)`M�գ�K�f��"O��{kށ��<�t��pu"ԡ�"O��;6ɚ� x��4�+PK��2�"O� vZ�b*l�����;��"O
|Q�*O�{� ��ӯ� 6�k�"Ov�B� �$l�p��C�
��p�#"OF���F��tdIH\�q&��"Oԫf��	, ��; ���0hD�*�"O�Ր@LX�U
x4!OǬ.<rŸ�"Ov����ܩ3�d�aPd�;%D�9��"OB�+Ŭ�:�@%��b@DBX��"O��P5��"P!�Y`d�V�C#��d"Of�C��0+�V��-Ecu�mK�"O:a���#�3��E�fH
���"OܡJ'�ߍ5��*	0��	�"O��C�����.�z�L?\ �a�"O�A���G 0@R1������"O�:�*J-@���0N�9^�d9r"O�$YӉ-	��q#Ҭ��v�r�Q#"Or%�f�ŉC�
���+"#,��"O��9��YJ��6J[)�Sp"O�q���+?�@��?o�5j"O$)�k�6��WN��u���	�"O��j0�:^l��!d�y�V-�p"O�ɫ�ET�BN�dy��nz�}�"O�l�&�IZ�-�0��Kt|""O�{d�8i�$�:s�M�H�"O a�u�׀<�>�7eͮa�ȩ�w"Oz���m�J�4!I7��#s�j��!"O��.�4w�|8[sl������"O���
i[���0�V?,�:eHg"O���� �/^�b	@�	P>� ��"O`u�c�Rb�p1!f,�@E��"O�@ a���)�d-UMH�J�"Oެ�E� �]n����'6.��SV"OX�0�([��c�g$@��7"O,y�g��m"(�%Z�;1f��f"Of�i��/�����Xj0����"OV�����&p�!�"L.o3����"O�D�ǁ�/!q�Q�ݥ�>D�"O��a0gO�6"ʤHS�TAx�`�"Oܴ�"�@(0� ����?X6^���"O�5�e��>G�� a1 ��i,f�Q"O�s�"S��e�MR�r<�9��"O�+�/[�J���1��
b4(�%"O	䤃�2�v���ʇ�X)v�I�"O�����'�h�0�KL�@,�Q`"Oڑ��]�>�0P9bˑ�,,�m�"O�i��`�<�l-�F��,zF�a�"O0<(�MVv$\ا*�Y])�a"O�!�7�N5������$/[��"O������'���j@�T�Pu�]K'"O��Xn�}�0X�'��s(Su"O`�����j~��O�w}P��"O"���������$�=�\ɥ"O�9�!R^}st��1 ��*�"O"$�ttx�`$��U|-��"O!��_P a!�$7^���"O��̀ �l�#��҈pY�"O|1*����@�#���PL�x�"O���R�ҕt�V�M��ʈ""O5���O��˴-Z��6۠"Ob ��G��q�Ӌ�N��Ip%"O���ì�P�9�^{R@#u"Of�I&gA��u����b���)"Ox`��iJJ�R�J��2y��"O>����͸{���Į�D¸<�w"O� *|sAکq�p2#��M���X"O��"�'p8�m�g/
�)9�mC"O�[��=^����h��I2$9Q�"O���h��|,!�$(�%%4��"O�y� G�~ߌ͋A�_+8��"O ����{�R���`�0��"3"O*aib�xO
��4�UU��� "O�ABc�.vRd=:0�ت5���"O����8A��a@��3��x�"O證�IݪK�ԴX�-M�f���(G"OPXҷ�]�H��������\be"Oڈ�P�"<�P�aBi��t���"O�%��"G�K(괐�G̜Pz����"O�����ߓ����G:{����a"OFm�w�M�Dp����4{6t��"O:�@0A=�-@����zbV��R"ORD+e�	�T�
<� d^�n^b��"O�����K�>��A�'_#M�q��"OJG�B�[ �	��o�/F^Ё�"OLC��Yv*r|
g!�2T7
��2"O����,C��� ���!k�Hp�"O�l뢯�
1���ġ3A����v"O�P�OX=f�;�i5�� �"O���@/t'J��p�@,�p�0"O��SL�*� ]�'JϺ	B
�Y�"OPY��|��a��S�7���"OdCC+�/L�@4�!XȲ̀W"Ö�Q)�d
���U�Qd`�"Ot@S�T�B�~h`º3h0��F"Ox<�6]�"�ȡ� �{1�}(�"O>�Q���w��hQ���t��%i�"OD0`�C�n� "׈CW��"O=Q	F}�>UK�,F�1�JQ""O��xfH4o9��Bl�'����u"O�ɱ�!1"_M㫙�:��@�"O$e;GfN�#�l\��+L�i2�C�"O:��m��싇I���KR"O4I�#o�6*���H��"=�z2`"O|aie
	��"��7�ۻjd���"OF�r@G�+I���s�;ya��r"OT������0�TiF��)�\��"O��"�8>`�"�/^-C�i��"OB\a��W�0���0;R�� "O�u���(u{�xK��݅tF��A�"O�ЪC�7sLU9�˂b)>���"O�8ڣ	�9�tD�A(ʧ]s"O�����TgJ(�d��/]r�"O�qH@�R <-����t�c"O��X�I�3� �pEг{�N(��"O ��`�6�a�vc�{r>I��"O:�S���$�p��#/��,��"O&��D'ا=����q+�Qȹ�`"O���'W)9IDasႏ�`l��"O<Uѳ �����מ%���"O�EA�晿}2&���N�e�:E�D"O(A�j� zd�y�.[�A�e� "O A�j�gB�yC�	p*2"OLL���3���[D $]�6�!e"O�����߿A%�QZDjˊh��X��"O��C�V'bi����@l��"Oz񅢅�m��	K"��iL�)�G"O�Ш�o��hɊȆ�p)pɦ"OP,3'Dą
�zE�'� 9dXr�"O�]�oJ�5K�!y�ģ<�"O� �R��߱zff�alY�3Ѹ�sG"Ol#�,,I���U�6]�v�{"O�ѨWgG#W���$*��iZ
$��"O���A%�!/4��ShЗ2B��2"O.@���(��Ԋ��л&5daR�"O4ԋ��%��Y`G� ���"O��֬�);��u�I�T���"O���ǯ�""d��Zb�Xv� 蚔"Oֹ�T�@����:d�BZ*�:u"O�lZlE�k6�x6+F1nR�"O>��5"@�m5|�Q0�7
��*�"OR)�rM�f���RgOތ=�4I��"O�}���ߧq3�d�C�:ҒѠf"O�)��CW�A����T�V6��C�"OΡs,,L0R )'b\�i�ԉR�"O�q�3��0n��i�@��4疅�#"O��5eY��eC#��{��kw"O6y�c�4�i��B~�́b�3�y��
p74�!�L�y)P�:`�.�yB�@�YV@��a��|'^<��!�)�yB�l���u�فw��!�Q�(�y���'URD�&�, q�$p����yr&�)20Q� BH�І�y�W!F��Ť
���ɋ��y"�@ *M�Q͗6�� ��L���y��tWf��##�4t1AĚ�yB�(9���"�aO�y0�P5�]8�y�NT�Xd�Q����y���yĎU"�y")<3��%��%�E�F��+�y�]$��)33'YF������y2cs������dbG'�	��%��'�lh��H�!�h�t�(za����':ЭӶn{����k��"� B�	� ��]�L�1QU��uLǈ4�B�	/M���ǩ7{��T�����:�C��+L��iZ��P^�`C΁y�C�ɚ
>�cw�G�XU(�#q�E"�C��Zd 
�(J�^'��ڱ�ʺzzC�ɴZ�V�z���?����升5��C�I=Drx9
��֮�j0� Y<mYrB� IT���e��s�!cᘝ<6B��6m��i��V�]X$� �XQ��C䉏V0򄉧(#K�P���U!~�C�2!C���"69���!I5�jC�I,��������Z�a��pr��-ʓ�4�xU���a�L��b���\��~l5��яN�x����(�B���F�֬A"J�:Z����A-���ȓ#�q�f��a��yZ��ʕ{�*�ȓ5q&�:��̉a~�+�G�
Z�Ѕ�|��)BB"�p�z��#X2��ȓ~�̀�GQ�p�]bǣ�"Fmj��ȓBc$�y��	0�T�*�A�,��Q�ȓ���I�㋤|V�
`� ^�8P�ȓq�F��ъ��`H�#�=1�A��!m �J�ꖁ���/Q�n���ȓ 5v�j1$�
k��!���D,`=�ȓ`Z��( �.p��1t��3��T�ȓ	�� h��)�E��\1��
����R�/)R�@�,{�]����)bW��[	�t��A�X�p�ȓuc\d�%ܓ48t=@��!"��$��nNH�J ^i���UK	�J���ȓ|T�53S�äu�6��G͞0�����S�? �=S�FY?���#���R�y��"O���d���X����a��q��q�"OV�ʄˏ�/�&8����,Ǌ���"O�QCƘ�\�=�'�W�V��)��"O:���49�:!�y4آa"O(��B�-ZͮWֿNr$�KQ�BD�<�T�xV���u�_�D=x��C�<	�D�+	�y��@�8����⢛@�<�7c�8��M�2PdYB�c�s�<���C�(XAA��G�4����m�<E�e�@!ĈK@�d�ϔ}�<�O��}�=��e��e��! �U_�<�qI�!�B��W#b���	���U�<�A�7��U��E�%h��	T�<���*��+�l	� :�P��
�z�<�G�Y,[FJ�3X@)�g�|�<����D-*�j�����`�!�C�<���ӂ<����	۫k�`h�@�T�<q�BU�j֠ȣfl�� ���!�K�<�I::�����l^�)
�4�E�<�f�s4p��n�}x^�õ#C�<�F#��<$:���F ��	p�
C�<�W%�j��̀'�Ё���)ӂ@�'G�y�`Heɜ�{bė�+> dH�M���y�ߑ&�,	�%/˥���Jb`�1�>	J���C�1D�����C
��1����0�.�	I�'��)h!��Q���X0/�#p`1;��ٵ5L  A�#z8B#�?s�qOL�=%?1�3 �')��I:�� Z�V�J�L>ꓽȟPI�c͐� �r�@q�&��93 @=�S��yү�1��P�]�e��\�%��(�I��$��M�����4�4�I"]'��x�JZQa~2k�>�fO����a��0ZVDk���E���'�Q>��7lضm-0T���&:�@p�<��ē��\I<�R���V� y�UEL.};.U'��-[v�b?`ԃب6�0RS,�7o4eӒ�y�E{��i��x|�4)s�� �p����T� !�d�'�Dm)��+w�=+tN�	Va{2��ҟJ;Ɯ�`��4O[�B͆�W�(�ē@l�f�޿���1v	���r���:�瘍0r��Q@A�Q^|�ȓUR}e�M�G="���e\�IH���h����E� ��i�*��.Դ��=Qߴ?��c���J?zD�-URd��P�K+���pe�>D�H1��*Sj0��a�$o)x��B�0D��a��ٔ'�v��+��lTt�q�,D�������t��&��cz�SD'�	j��ħ7� ��mM�0<X��J$��ȓUh��j�fX)����1��>�
%��U�f��H��Y���j1��`����sfX*Q�4?ъ��S�*�����Y��L�b�C�$CL6� ���p<A�!yI(�@�5D\�R�*�I�	�?A��d��H)�U�A��QseH1<�.y`0$���p?Y�'�.��g��8f*�ʑ-�%Iq�|���'��=��/ȠJ���!�qG�@2���'��m�U�O�R=y��6�+�O��kU�����x*0iX�
k�|��`��|���n=�ڦ�DxJ~��kS�[n90H_/�QJ�H���e�PǍde���4N!2bfMM����&��6���D{����i�����^�b�J�I������WX���d=}R�Y�24�2�ց#�x�/Z�֘'��	k�O�Le���+�,�k������:��*�S�d�As�
����.��1A���yr��;a|@ʓ��||�Q�nў"~�S�? fqI$�yS�X���!`��Ӧ"O~ě�Cךi�80QS���(�%=O0���nRt㧧�\�9*����!�d[��Z��!hM37�=Ґ.��	t�',�I\�)�S00�p�s)V��0�c�&|�hC�	��T SBN�T�dI%i��/�JC�I)��35 � @@~�J�a9�8��D5�DQ��H0Z�R�~#�HP̛�H�!���71�m9A,ƈC<-��PR�"O�Ġщ�\��hz3��i�T��"Oh-3�i�)x�"�hf�F$�6�"�S��y҅�6��b)ً}$t5�Ĭ��y��߯0BH����Χ?��WŅ,�yB�RF��`�	<F���Ӄ�+�yr$R#q����:3*����"�y�JD`)�H�%�P ��ڻ��'֎#=%>����d̚��d�ÿ!�x�D+D�x�$I�X���u/�����5�HO?�ɏcṉ�d�U����hI�v��C�2:&@ s��G
f?��)ȗc;�B�I
�pT�F��/r�Ȥ���� ���}�u���y�x�*b�h���Xd�Ի~�C䉐BX1J@o�@�@�1����-}b=O�4�}&��B"O(�ݺ#�[�qZ��&D��6Ik����Z'�$r��)}��d3�'�2��ӆ���J�G�#�� R	b�+U�C܊�j7B�o�	��u��XU���O�����	�4Ɇ�	R�'�����ؓBl���gdOO7�'3.��'I�wA`�s� �Ac|�;��$:�QYz@X%�7|p�3j�6|E&p��I��R�\�)�zP�U��VMx��ȓv�z9�HB��E���z譄ȓ`�d�p�_0?�!!4L�Iw��$��F{����Dp<H�'�
pr*�Ѵ"���'xR���O��#*Kt�@G,}Ů�"M��q��xbH>LO �3�M
�"���HҮ|�r�Ð�L��	z}e�,�.����̄���*WO� :*��d�<1ņ����6�M�ɞ�1S,��<Y�'��O�c�a�n�x�A�"'�6��e��GD̩G|�$?���!#�0���!=�1���@i� ����O��+�d���D��H�������'�n�Ex@�	M@ d�Z�E� t $m���D.�Od`�3�N-�
��� �Pd��i疟D~��'��	�^�vIP0 �<>hQ{��F�`C�I7>�*��Ӷ��X�Fk�c��oH���j�""/�&%c&��*+%vH"c�3D�C$���|~}r��H�p�05r�/�1e��Iϟ���'��O����ލzJ�r@�X,yr8u
ԑ��F{���V�(9�YYWC�Y޶L���Q�����'㰹i���pP!�7LϑvsB�:���(}��Ɂ�X�; �#6d �B��v�~B㉋9��fR�?��ia�fY�*R�9�O�������O��Èyr��9=y{%�W#����7o��yB��:U�TQ�	�	;���	��~"�'3�%�t"��0�Xᅇ�n4)�}��3?!��IȮ;����"�)H/H ;G�G _!�$Z��T�H�dƹ) ��M�vS�	D}2_���|�'2����N�̸8�@� �ᱴ44��ڇ�A&A�6���%�D��٘�� p~R�i�qOV��~̓GF���$�p�=ʐÓ)�J���	�<��� 'SfF��V�;���ISi�<yA���Y�^,q�g�)���2��Y�	D���O���L (1J*}�
��|8�]�'a�~
� �Aѕ
Y�,�>][���1Q'��7ғ�?y���M�R�9^�nQX6�ݎl�$(�`�M�<iV'Mg����Gv�9�D.�E��'�`��I��Y���X�,�����j�)>D�\�N��Lƴ�sÂw���X7c�>y��铹X�1�!喦32�K�mȂ[�LC䉸�a�Qn� �nM�0�G'%*:C��uU�0�1d�__4U24+*l�(C�=�Z��G�P�$��s�"��B�	:z��Ͱ%��1~�*R�ԕS�B䉵3*��p��?$�&�E�k��C�	 x�Ɲ!��U/ZP� ��OŴ*\C�	k=��4m��5�y��G�:KHC�ɸF�&Y��ꂇ_=�;fGR�@C�ɢWr�u���L���B �9\�.C�-Rr��C/�`֔$Y��/B^�B��$j�ِ�_.|J�7)�(F8�B�I%儹�c'�k5�'�-{.�B�I1@��c-�Nx�XX���?wXB�I�L�81��,R��P���r�B�	(S��A�CZ*/v�J�,�$F�|B�I�-�\a�@�N�wj����bРP{pB�	�X���Br�.넅+D�#S�C�I�P��ِ�ӄ&\|���IL�B�IP��p�
l����&A�.�C�I{m�8�� ��0���9fÙ	+_�C��90]��2�
�S�ic��5{�C�I�3klT+B�?u���#����t"O�u���=�]j�e=	�4��"O�P֨4�2`28���b2"O��u��lh���udد�h8�"O� �sO7����a�گj�ZY9b"Ol�&��#?Bj���)I6H	��S�"Ov,�h��eG<i��	�Tx�"ON���@���YhJ%Bʼ@�"O��㄂���X��ӱ�0�b�"O��S��0�j�9F�L.m	=�"O����}vL�ԤՉG�L!r"OL�k�%ӑ ���FȦZ�HU�C"O�|��әN�����A䖨Ч"O�P�t ��T���$�Ē6�tU"O�����g�h S�M���@$"O��Z���R"�|�eI� T L��T"O>Mp��[[
�E�4�^	K��t{�"O0\���HP��`���ȭ+��X�"O�$bӃT���j���q@�"O�=�6�E%|�RQA�m���X�"O�@2�j�%z"���c)��}�����"O�L5BJ�cfH@��GmD���"O�T�,�/7t:3bAH�0�J�"O���ȽF�P�9��F�X�b�"ON\�S	�9��Y�H���� �"O^�*�c��3r|���A_��ty0"O�4�C��(/ú��d	h`TX��"O�8�A�ōb�h\���X�x�"O*��V�Ȣ\;�qE���"NH�(c"O���`Z=;0I����D�T�1"O�]!�S��$T�&((2�|���"OfdqR��@�Ry�B��"����"O�l�4A2H4�Ӱ�\�CA4���"O���䃟�l|�P#�C��m�r�"O��Yw+��B�ӠS%V�l�C�"O�tۓ`��%̖���߅�0e�"O`ՠ��ݝK�"�������ZD"O� ��(�O��o;؀:TAЛF�bi��"OT�¦��8%lll��fߖ;�h0��"O�E����C)�%���%Q.�HR�"OX���c�d���Ɠ\,
܁�"Oܜ3p Ru�5�wf�@;�	B�"Or8kӅB$҄\�WL�P4V��t"O����@��8 ��ӥ�պd~�!�%"Od�z�&L]��hQ�J L��i��"Ot��l�|=�"/ђ~���!!"O�k�I��+�y���9��[p"O��eT\@8��fM��W�Z��"O0�H�l�ϒ��Vb^�~dR�:�"O� H�1-�<��b�ʬL:(���"O�QzA��I7�)��E� !6�H�"O�A�D-ڣ$�����]!Fm�"O���A�؇" �e�B�38J��'"O�L#Tb�$��b�<8> Q "O��B�a 1]�6�Qf��|=�t�3"O����Y�'Ep�YP���n fTȢ"O�*r��s��I4k�:"O��J�AY9�jD ��Ҟ|�����"Ox 2�D�9g��̉.�-;����"O��P7��@�4��e����1�"O��sg&�fX 6(\��q�g"OF�@�e0�$�Q���7W��Pj�"Or�P�O;8�S�	
8J��E��"O
=@�ʂ%B�D���#j~ܐ�"O�M�U+�7'@���F芭d����"O��à�Q��Y���3�F�R�"OR��l��f�$)C�.��2Q"O����NA2��p��f�F�P� �"O�0�&�X0f���v��(�.�
�"O<��c�ђ}�(s�4fׄ�: "Of�:F��&tB��q"�΄[.��'"O�;sc5z���w'F�.�Ȱ9"O��"S��	[I ��u'�9k�"O���d�Â��c@�\��!�"O<=3�j��L�ॎ��he��"O��cq�O8$q�L��N��d#�2d"O��ʣ�ǩA,D��k��7���t"O��qefU���0�I�-�|��"O�L�A�|&���A��m��ԑW"O��i�^�7(�H;���,�ꬳ'"O��#�*��\&J���-�J��!"Oji�A ���`��B���J�"O��Q��"��9�i�o��!�"O0!Pg�d�h���G[2U0�i�"O��AEV3j�!��e�:t���"�"O��0]7(��1j倀4F�| v�'=��L��f��A���H��ZB�>,`��aQ��?UH(H��e9IS>7-,����G R�p1'� �i��q8gG%D�h� ��8B~l�ъ�?���sr�7D�l�I��d鉊7�b���H8D�H���ƫ<Ў�1D�F�~s��q !D��z�N��W>��zj�X�]q&�=D�`Sd,�+��؝Ɗ�"2�<D�,z7M�.ϲ<(`�<Kl��.D��Xu"9�h�##AA�c��hI��.D���,3Oo�̳$�_)(P{��.D�4���m�� 3�a�`��e)D��*b��<[t��c��A<k$'*D�����AX.�R��f-H�Ԡ)D�(!"���eَp���?0v�m��*D�� �4{ �ԄW�J�y��1�R�E"ON��Dc�(�\�#�ɋ�IO���P"O��⣁��)��h2%��$yKءcu"O��`��ե|��y�i�`\ZY�"OF�DM�#:�=�H��dF����"O )��.�7d.9CS_�U�XI�"O��r�gZ-zư�q1�E�o�ʖ"O�+3)P�j�@`*DfE�-d>)��"O��:�ë4[P���n�(�is"O|���X5bc�ݢ�oB�z�*d"Od<Q���O�F�ԭ[H�9�"O�}�	�m�9�#c����bC"O��A�K]���Բ�@�НY�"Op�f㈁�hh9	R���u"Oj鬲n�n����6�yV��A�<!�M��EH�e{�e?M-x0�(�w�<��/�U�� H�D����s�<I�$�:�0� 6����`��o�<��Ϧ+2�a�
�g��ID�Rf�<1��;.ā�LS4��8{�ORL�<��.U"z_h%�B�A2���Є@m�<��̑d�.Qu���d���`f�<Y�+F�8�
�G�-��aQ�i�d�<y�HG(M�|���
�b��f��_�<ɶO�}{:����Ab(�!u,^�<���R>>�����c�n%r�/�d�<��h����V��?�>d����z�<q�釉8�0La h@%%��NKs�<�fE	�%(�pQ�욐ں�4�t�<�EG��(�J��Ro��U�b6�Ā�yr��)m����eCU	M���A�%�y��*VmVE8FG�.�4�+�b�y"�XW(�A!Q#�r�Jj�o��y�a^�~���"@��6 r7!U���'�az��,2�L�Z��{?�z�-&�yr�K%��4�q͏!!;��COF��ybn�v�8��B>jB��R/��y�`W"K)���Nx��
q��-�y�M��|E�a��w�>l�qeJ��yR�R8L�����4oD��X!M\2�y2BL�.+��A��
a��U�����y��	<%���1�̩A��(ڂ#2�y��2`d�����	�}��n6�y��Ms�^�1�mZ�|��=�����yB-�0&0H�ie�]^侕R�mV�yr�8��+G]�X�E�����y⮅�cN���Ϝ4]ӄd¬��y��O;�|�V��\�^09�H���y�%�g��#�-� ���c0@5�y���?L\,�!Fd�1i���c�dԔ�y2$/��Y�/�^�֨�d��6�yb-�3/�dqdR[�n�#aO�	�y���h"0t���W?�HS� Y�yB�c<\d����HHHDە�V��y2�
�>'�)��)B2H&J��QiT���'Oaz�����K���=k�ϧ�yS�p}��I��P	�hO-�yE/v5����I��*l�-�y�%G�����cƺ�@ዴIΪ�yR�5D?F�b!i���LJ�)�.�y��
�(e�V��{�J	(��#�y'�P�1�%�׻w��;U��y⊛y�����q�c��0�yB/�[�$Ejf��aM�4�nǉ�y
� � 3�� .'A
AJ^&3>��Xq"OxKK�mQ<�a�^-V�~���"O�Y[BX!?�$�wd�E�A �"Ot�6I�	m���4Q�NH�R"O�x��U�{X�s�c��1��"O��X3�֝O�Q�!D˪ud:<��"O�@�7� 9,��2�V�T5� "O�9��P�Q�v��eݠfL�)�"O��~N�Q�Ė�p�r��"O֙cP�Z�w��'%�ƈ�v"O��إcŧ]6>�Ǵ3��c"ON1 ��ٛ(QƤ�(�"���"O�yk�L�U��}�r��77bm��"O���Өa!�� �L��"O� "���rM�"N�.˴:6"OMCG�R*�頢	_]�M1"OV1Y�� ~p̡�2�#y��t"O�H�6��1�0�J���h�=pG"O���[�]�A�͚xZJ���"O D𕡖�!T-�#'�wB0� �"O��@C�W) 8x�B �ӘH'̱c"OD�N�WZb �������"O ���n�/ӌd,A�65��h�9�y���#�� Qc��S0F��F��yrq#�c, �t�x�f՝[�!���)xgvd�ҏN�(������tY!��ɅN��ٲ�
^7/�ḇ��rF!�$�-ZJ@
�%֔Ulr��P�c�!�d�= ���tDީ�X� ��!!�dB!:u�Ȓ&�&.|l}SC,�Ll!�d#Xv��L9JAj̙�@ɇv]!��М���酀[�*;�b0�=�!���\dB��$�DO��s��T�[�!�Qh��P�oO�?6����m�J�!� G7���N
�-26p�D̒+!�$>����ٳ$�z�:���!��$v�С$�gK��E,�<87!��.֬��P�>I�����w!�Vd!f��"cפ=��BI�6Y!򄐓P�\��n �`$�a5��^�!�DԹ_hE��h�;.>=s���!�X����a�*UN��!�@�:�!��_+8p���p�A�B$42��M7	D!���(^>� ��2�r|�`$T�0!�ċ��u��P�<�hf"�>	!��ɏCoZ�9�&�
Wf{B�"�!��HY��̕w0����
�!�d=*WH�k��ء-ܗ |{~���'�4���.��|��ѷB��)�f�:�'�|)3�L�$^��FI>!���
�'T��t�8>60������H��	�'(9��I\2����"���8	�'��H��)��f�%
�L�'� ��#لQ�f�ٱ*d��ZpL�44��2�ƑrS(�q�o�� �H���/D��
��-B����W@�v�j7�(D��c �"�,PK�WR�pBC&D�ܲW��f��(� ��1Q�)s7G'D���#�8%����ƚ�w�^T�@�8D�Aç��)=�dJ�j�c����4D�������+ $!�ʖ�U�`�$D��I���P�K%ָOC���f%D�����.$4p=`�U�5�R���"-D�d���� xŉN0&�(5iQ�<D�X[��@��T����)�ܘJ�G:D�� 60�a��B��8u�[�d@���6"O��!b��.���I�=3�a{r"Ob%��C:UwrкS��=:� SF"O�Yf눲�<)�'%v����0"O�Tr�F�8���	Ӈw�
p3"O�}�I�'N���j#(A�_� �v"O�q���'�n�A�n/(׎�(�"O����J�]B�ضo�k�N=��"OH�󡇖:!���
'O[� ��!�"O������� ��$Q�ly�"O�������Y�N�p@��,�d2�"O��J�k��7-,h!�ˌ�@��|A�"O�dbqN��l�� ՍBqx� D"O���l)L��ѲS��ef�*3"O���S'[�]���z4H�h�H��"O8!���<C���Ƃ��SC~	�"OB�҃�B%7�
a�UgӞ-v�"�"OKM)c�	�q	�1�	���<�y�㛂	
"`��lD=��Ԋ�����y�	��
�dRe�W,��Mk�	X(�y"�ގh�"�a4홋&�P饬��y�L��M{�4P�L�a޾Բ$d���y2$U:jx(�vk�M :�� ��y��k՚xQN�jκ�z六�yr*��t	�m��E9v���snM#�y�R�V�Zw�ڶa��Qӂ��yBM���z�k�	]|�H��؍�yr	�
t�4`�FD�z1��Y��ؽ�y�c��9FH� �~���֦�y"�T=�&͌e���aE]��y2&��GV5z�bS�B�T��O� �yR��)`�t��%���V�4��C�9�y������S�j���b��
�y�l��{�� :�ND����+��9�yB�׫%p"Ò{z���ϸ�y����6s
0ca Ј`tƅi&�D:�y"`�;q�z@��KZL�q`u&�0�y�k̵U��<�Њ�b����)D0�y�� '8.9�RD�x�TX1f���y�*��H�3��1c ��%��yraE0r�V��v �h֏O�ybH�3r�2�:Sǝ�{p��"����y�oO����0R!�e�^��e���y�����p�ˍn@��@�kR��y��D5(C�}+��o2�H�s�ɘ�y�A�H�8)�,�?Y/<hRbk^�yB���h��40D�IT(hJ���y�
�t����"�w~�H�DI��yR  ^����		*�Ԓ�	�y�.��WL�E�$�Oz�l<SoΕ�yro�W���k��~����C�yB-��[�\�{b�J�l�t`�e��y��@0��b�
R�[%ZIB�o��y2e��ؙ����@���9!�'�ye�#/c�	1`�v�4��g�� �y"Ł94����`�b��6�K>�yb�XQ��ÇįY�&y�u��y��<�6�R�V�0�$�-�y�nȅ%�lRd���O~�s����y��[�(x(�$�F��9���yR��v�Q*$Y$3�V�1����'�a{�ǚq"m"A�����@g��8�Pxr�iؼA����5�
ظGB_�q�@�S�'�uȔ+X�����t�	+h��̂��HO� ��y��T����9���h�Iq�"OP�c�k�^���cсg̵�`�>)���	��.�[���y,v�H��DH!�܌����P�	 m2RH�79qO4��DƙB���w�ˎA��hѪ.!�ē9^<9���ē�R`#p�5�!��$\B�����1��<� �_l���ٴ�}�b�U�8�*�#C���ybkU�o��*Vǡ>�]˶�
��y2F��1��	����#AR���<�yb(W�J�-$�X�Z
L�Z�fͰ�y2�K�,�\���G���Q�4�y���U���@�+��1D�U6�yB��'Tb0�0�JU|E��)�yMF�:>����GD�h�B̉��y�l��kz�����6o�3��1�y" �C�9H�A��/� a�����y�FMۦ����C�!�^�tZ�y'\ϴ�xD��u;:y����!�y�˚Hu�)x�G;c�l����'�y҇ނi<�̛�5bt�{5����MK Ǚ�p?#n}$^�[P��L��W�CJ����*�rI3�O�y
c�ϟ:���!�]8�+�"O��bZ�bP�6���H<�	�����%���çN��$��;�d�wA�,j�A�ȓ��i8WbKO���V�H�^��9A1,�G�P���|�'B�pz�NJ
��T�#(���"�
�'��Ñ�N?%
(�	�F\X���8!�?B��K
�/E�|2���!�*)�f�F�x���"H��qc�� ��*ۻ%�B�ꀏ�</Z� ���?D�T d��+5J��a���Q@�|�WH/��"���?%>e�p��."u64 �ϝ$B�RHyb�*D�X#Sm�S�
A���T9d��!-D�(��,y�a@�N%8f�XM,D��;$�!v_�1ܾ-��q'D��!6'����}���\O��0`�%O�։��'��!��A��0U���.�	HV��'��S!�å!� lI�.�~>N`�,O���E�:m���0I��|��	(,z"B� ]�ę��QJ�<��fZ Z��{5��>7@��1e�^)i������gԀy����'@5�0�ӡ^��dP�!G?%��
��o�Dy�ËM��$%T 8p��ak،"�J����L�@P@��Ĝb����Ȉ�1�3glֿR�Q��9������YC���r��ӫC�"��P�L'q� E�"C�I�Duz����T1��M�b���	(~ED� �cd��F�d�O�Je wV'��4K �U;��!
�':ĵK�"�0\K,x����|�Z�s"�:5.����P�Ẅ́����I�Z3ĵڄ��?<��u�d"��>WP����)����ϖ�8�G���!�(.L/��Xa!�|w���W�>�tQa�C_*\� T�׎˯c��R���,/ `�#E�	��y�O�n�*�A���Q��瞢���x�'��Yå�����L���Q��H Y�'��AA�·Kr���iD$��?E⢃^�"��\��J�<��� !D��	� )�&��4�+�V��Ti�cv����O&&�R��ĚJ�2�g�'+~���5W����+F�Q``�(
:�a#�,oM�5r�A��E��)ߘT$>(�f!#��a�E��y)�o@=	����B�Q�F|�h��-b�)�����'�X8C0Z>]�Ӥ��A<�X�΍%�$	J/D�H���D �������h�B��,A��"@���7cǑ+Ja���w��yba�!M@�yȡM �y��rO��i.���aCDtȖP(�'tM`5�Ԏ%.����O��E#ʈp�QH�[�u0#�'ŦI�G*ƃe@!E�C���d��p��)� ��"AQ�~�%B0!K��ɔs���ra��,��Or ѴL�'P���O|� 6���(!
�H[�<f|�2V"O�qn�?�D �w�@(Eш4���>I���Q����?aY��F�V�(e���t��a'6D�kG�+N\Z����:�@�X��:D�УuB�@x�Ps�v�&x�5�9D� ��D�6q��B�$\��"��9D��Y`��@`�䋦�_[�y��1D�0xBHG�@�Er҃`9D���.D���Ud˩.Zp�#r@��f���Չ)D�@;dę�\�`��c�'Wp�kB2D�p�u��4���SF�I7n���Ј%D�{�`/X{R�y$��<2a8p+-D��h�c9���H@��'V��q1E*D���$�J�Na���1�����n-D��s��ǧd]���.(II�8��!D��jsN@,� q��4`򔨵�3D�BT�V�{�p�p`g�W1�j/D������)lW�`�R�_��%��,D��qd��7dl��#ڑ\`�QUn-D��Ȅ�ޜ�V�Q�l��y�t5���-D�L�|p{�����;.��@�'Ѣ��!��C!t���g_%
ҹ �'4�h#�#��%��aa�͠k��j�'�V[)ѡ
QA�`M�_��H�
�'Ԏ�YAg�%�d��IP�[�'��]�C#ψj*�X�ꃓ@$�9��'�����ʌ-<x,zw�N6 ���yb��KK���6�Ǵg��	ׂԈ�y҂Q���z���)����I/�y�o�=��Sg"'C��á�ޒʸ'H��XR�'��t��<��M{�_"����'**�AC�	�j�ѲA�POr�1�'s���b�H�t�Ģ�MDb��'��9x�&J\$x���ؤ	�:�I�'`�٢�к
��@���@���'&P�Ke�Y�~���g��E��0q	�'��4h���+e.l����	�9ٚ��'��aڣǟ�9kAGS�;�hб�'ւy��֐!5]{&� f8��'jb�W�V�$(�a��䔗E��C�'�Nm���#xc��b��ֶ>�n��	�'�`�ABQNߦ�u�1�ȴ�'@쵳tD?�z��"]�1%���'�\mb�!Ed$����	R�)��5"	�'^ű���r��+7g�#d��'۰�J�&q�@�ND�1��'��=#w ���`B�BV�t��Z�'�(��剓'v-�BgU�-����'� ��-_v`H��J�s�d�C�'R�("��EĎ���cή�>Y�'- �XӀ¯I��8!HM�#�8���'��Y�7c�D��!��Ǒ�&ڤq�'��������AQ�a�8+��`j
�'X��A��թ+_f�x&&̃Uബ[�'�zE���!m��)��ȐTT�
�'p�����;&��ݢ�KE�N�l�8	�'�,x�nC,G��l��W�LF�	�'����r�2������R�<26t��' dk��M7z���X�hO�b%��'�stb)Ne|��l֡~�<�y�'����K.e?�	����v"���'�zmq�		T� �HSF���'k�XТA=|&D#C霘C����'���h�9�ر%cɫ1����	��� �ȑ-W5_VN�(/A�Q6�d�R"O�ٱf�O�)��P��Q�b����"O��u@Ͱ$����W&E}H��"O����T%���YC�٦z��1"OzXq4n��J�\�*�	D(H�"r�"O�D��.�D�&4RP��c�2�R "Op�)�MJ�K��)g@�]�x�
�"Of��&E�)�r��4��1��T�a"O��ؒ�2N�@I	��֣Y ���'j��f��$&�8Q�R�
��A9
�'��|�6�I(� ���L�&>�D���')��.Z7�����J�/v�'t����T�#$4	�ףU�`�9�'o�<��Bn�x=��$z8�ɰ�'J&t2é�b��=fh��&-t��'���̕�Q������Q��'Z&��$ �iP2�j��F9����'Ж��'é[�`I�*�(��'���`�m�G $YIҎ��d�I)�'�(��"�&.�R�!A�;����'�<I(�D5V�$���^y��'�xy!C	y�<��E��#�'*�%�&�E"U��Y����t6H[�'r(\q�Gٛjd~�;�b�qI`���'�v�x���l�ȴS�F�4m�,���']�����-m�I���@Z���:�'�vh�[��6�3`�,^3����'z�����a�m�R.N�J���*�';��·FN�gޜZ�(R��|Q�'��M9��ĈOxR���@8NZ�9"�'{�ii0cà{R��pǅ<�����'� �8���򝰒�3@�EZ�'uv|���V���1��N�<|R9b�'G&��CF�D�(�3��Ѹ7��:	�'�¨AJ�T�ȼ� D)o��2�'���A�(.ǈ���aǻY��
�'JL��C��F0��'��k��:
�':�ዅN�5�>�C'�a �X�'S,��ӥ�L�:�"�1���'t(��υo@ܼ:slQ4�(a��'#b�#��j���cZ�&��I�'d=i��H�a�dUYb�K����'x�	��D��H%0��Q�Ͳq����'t�Yi�� ���1�G?GH<��';��u`�3&:a��O�$.�2��
�'�f��EB��XYB'�9쨋	�'���*A�֓08�
9��`�	�'�5˃
J2u� c"Hē���!�'i��:���
<AӁ��4V�J���'V��J��]�iH�ŉ�E�n�C�'e��0i��[�<S�+
a�Q�
�'*���V�Q�a�L�C���6fd�1
�'yƩƦ�96��P4�G�4�Q+
�'���a��j�+�[){,�	�'����#�&X�N���>�R���'���㔥ʳ.�z]��V$ -�x��'p��p��ՃI$a��.�~��'9�Q� -Z�M�J��X��'�tss�O{����8u�>!K�'P���F$A�T� 
o}vX��'>�p��B!RZ�U
a�m�'?"`�$�>Vy�r��Yc�\a�'d��"�J�yN-��"J�R�x��',( ����P��e"'YJ��]��� �FX�VՆ쨆��l�*��e"O��j#�$M3.��dK�?H�""O:XA�lBE9A�MR"�"O8�h���Ȥ��vb�2�`��"O�1�5/Z�;T�l��-��"O�!��÷f��4��iz�Q"O.�Ѕ�\%,��9��͔kRy"O��񈔓\�6�`���A���"O`�q,Xe"|!�ۉK�V��"OD���͚�����wl��k�4�Rr"O����J�4kЎ�@`+_	U�y�"O���T8[�@���}x$Pr"O�Y�4�O�U��T�G�x��³"OQю
�$Q��E?K0�]��"O�Q��V8*�0@j�$<A����u"O�U��,rs&���E!:Ӣpb"O�{��!'�bE�S�üxw4�+w"Od�(�G� L��9q�*\
8w�a"O��4L^�w���(H��	3G"Or�����v�B �:@���"O��s�)
,B�5Pd��5Y�\�"O� ����%)�TѰmE-MD��!"O�1�DÌ@���B�>Ȇ"w"O�x��
Cl���,�E��"OЍc�L���(�7� �e'��ڒ"Ot�1�C�3|n�H�7f�
S�&"O����R�T���	T	�hyR"O��%��.c� \H�gS����"O��KM(Q#f"q��9vP�]�"O��F���A�P����.	HzI�"O�����A�+!� ���L�U&�e�S"O�x��l�`�T��#�$?4�f"O���-�1��)�gcA.]��"O��8w⇌�QS�?4^�;*O�� �<z� �u)�-�p�'z��S��
7�tHōW}�6�
�'���0��67x�-�t��<nU2�
�'�x��N�8�$��5�LAp�'��Y���V����&`�Q�X��	�'�����%�2x�񤓏H��0[�'[�����t�A��=��A��'nr����D�@l�Ni��+�'���G*V�?��Y��DP�޹��'l������	N�(���:EX$��'O"-p��@i�p���ƵZxN���'�����B�K���q8(Y3���t�<��Ғv��d�t�"��PQM�u�<��M.u�ڌ2r��M�0�#�s�<��@ݠ|%ʙ���R�>�x8���U�<)2?�,Y�M
i�����TW�<A���K $t���LqJ��V�E�<���Z<zP�1�H!P�|���|�<���K�8�&��@n�tf^t�<��/�#�R�1u�Εkw�,�j�<4�q��h�q�?����SC�k�<1��E�N�4�e�޿8y����!g�<�A��(_�y�qg�;vz~H���Bu�<����]���.�T2eX�Iq�<A� p�������F�So�<0�A:v�0�Bm͛8�:Ͱ��Xp�<�3cޅbt�5Ӧ.������
J�<Y���|,p	B�hD�i1��HQK�<q���Ҥ����V�v�
`@���G�<���,H�&���`�BlȐ��B�E�<� ��)B��P�A!Yt�J�"O�)�P
.��P�q/��luB�"O���\|�(}kG����X�"OԨс�=���S@��^�X���"O��q�'-���s�P	S��P�',6��F���t3�A��Jk��'|,��3B(h�.�!���!^�zI��'۞� O�!ʅ ��MC,M��'s��Z� K�J���ޗq�@Mc	�' RUX����`�HR� n�(P��'�����"��zf��wP��'�bq���_=3U�)J�GN	�D�0
�'`�4"5ӷ{�A��+�!���
�'��B�B�IX�`b`��b��'�Ɛ�5��08O,�xҊ�As�=j
�'��](� ȠMx���k�*Lк)��'U|�J�\Z�Ļe�@Ҍ	��'Y����~?��
%�%C[H�p�'ۚ��v.ܶP�hY�b1��!c�'��-YQ1X�lyA1��H��'��0���$*�T�Q��G�T	"�'�&I�d�~}�mH��C�4��;�'{����0G� }�#��,��9I�'N$m12S�] �x�ċ/N��h�'�HY��*�Y�E!��&o���'w^0ye�Z�SO0�!���Eӈ�R�'~\1�i`����hԮ"b�H��'�D�4O�N>�(����++���'Y��K`!��H9���̐pش!��'��5�擖^�z�Z��?4<�	�'E���#��"���*�fD�:�$Lb	�'T6�b�'��\
4��$DD�an���'1v� C�=3���d��[����'s\u���݅r_���(��B�k�'�>�R��ʖ!��(ZG�¾2o9��'�|���cB`�|��Aa݋g��e	�'<�L��B,K�%��'*3�<P�'� ��"��~F����"z�vI3�'�`أr�;n���y�kSrJ�9
�'o앉#aL�*�òNM�PM��	�'�:�'�Yh�:EވJ�H�:�'����v��[�ܡ�q��t��x�'@���#g��#�r�XfA-u�K
�'�ֵõ�ͨ
��� 	�n��	�'��3D	 s�
e ��_��0ͣ�'9����&U#$�h�zDM�:j;�'�Vx���_ �$ˆ��|V�h��'�����ǝ1�l��*�h�y�	�'�F����Z4��ۄ$�:���J	�'�D{R��x�t�HT�&P.���'\X��0m��+)�m{�/Ȭ�-�	�'��� �*D��H#� G�qD�3	�'�F��	L�.=2,xߠ���'��`��̘`�pb�	zt�}��'
V�0c����b�l ?q+@�I	�'�(��#Q�)p������/sQ���'�1�ᏖyZ�U��קm���'��i�v��f���p��)b",��'�������]���pV�R+X��5P�'�{�	�<��ub�P��b�'�����!�>�\�� Sw����E�p��aLR�Y&�R�>2��[��ppc�=z��ԳAN�ieC�ɆHH}�G
Ȋt�:�6�؟G�&��=G�i�$c�֝_��#��.N�ș1e� �2��c%����A3<a2���� 
�	#��9��TBu� @�TArV��	�Rj�Ӻ���g^!7Sj$��6J�1�� �,�M#�F
���ȟ�0؀I����Ec"	 fMAԢM��'�X��iW(Q�Ƞ��&̋~���B�=\$�O��a/7�)��G4E?(	��ϊZfA�4*"�'�Ȋ&���ɤ4��p�\4�R! �B�?�I[�]�?E��ك`w��[�Č�i�!��o��Ms �γ���ȟ<X+ǇI�cx��ap�ͯV{xx����5��'Zڣ�� ��CC��J4�`ӌ�*��'%�0+�j�>o�v@�S$L�A�(Ք�y� �	kV E��î?��|d(Bj
ҝ�v%�2��S��W�S��im�:B-<=� �Y�SN�|`�'`��9��Sl4q�t(���aT�(��7�ͦN���"z�%�0|kQkۘ�^��9�l⟘(��2�|ZCi�3>-�D#5hœ����F��r�xp��J|j���Y0,L�� 9$�^\����V��I�rI$�ԧ��D)&N5|u<`�w�^�MH$�)�X���!C}�S�ON~H	B��qrF̀
0B����P v��?E��^?��Mi�$YK����Ҭ�"-����?Y��=����;Qʓ?G�N1
�-G�/,P|�>��K�����'0�΁���4Mr�3c��L�"�&�� �41�O�&q�F��e.ārEx  $�c+�͡rA�=�B��,%h�%HdC߸@Ztq�b�"!�C��!^/�u)��R
���i�%k[�C�!7���+�&�p��7��6^B�I1	`T�$C�-F�<�b�J��T9B��"?��sLL`�rM���k[B��DJ�d�%��KfPA�(ӂ��C��$'�`�ڧ#�27�.��F��8cd�C�	�)��<�Ed< 8�X����@`C�	+`K�ђ	۸����7� 6�C�ɝA�d=	�M�QT�� %"�< C�:Io\�0�/��i?Z�q�K�n�C�/�nYza��
WP2�@HF�!�\B�I4�܀�e^���J���9ObC䉃oI ��S�~%�-�Q�G#s]:C�	*Ԇ	i6�䄭xf�2��B�I*t����=�0U�/�6?�C�;��P0�@-gn�鲆@�{�B�	�P�5�F�@���A��G��-�B䉔3��B1�=NzU�T.O�B�Ɍ+�6P P�B,V�B9#ʊ�dxB�	��t[EM�r���W�*%C䉣f0a3(ݭ%��D3���
�B�I+�Hh��F'uaU��yB�I�� ȹDD��w�QK4�
�]"C䉭+�
u��
� Y֢Ձ+��B��h�ȴ�m�#6C��  B��@��#eW�[�9�񅟣g�B�I�'���@�;~�H�0�)��C����Tт�^�0H��FF�ԂB��:��T�tf�l D�#�8_�:C�I�gQ�kB$r�p�/9��!؀�1D��s�@۴u�m�$.He�%T)0D�@��)��j9�9��m���|�J,D�xr hJV�\��Q9HѢd�(D��;@HK7\D�0�2�J> ̬��'D�8�cЯ9��u��.D���S�&D�tSWGM5삉� JX�^\��Ї!D��kUMV�i�ұ���א dέ�Q-:D���D�o�.���*�lƤa�a;D��ђF��dQ�dT�E��Ģ3D��9fD�<�, Y���*qR����0D���R%�UN�H�sC��*� �A2D����@�:?!8Qm�A��n.D��  t�Ӄ��q� ⢉�LpJ�"C"O�y�!G�w���@5!+�ڠP�"O�xG�NG~yS�� 2��t��"Oh�X�F+}�$3�!ܥ-���f"O�4�«ɠpF���*�Kr�]�C"O�)��N�*ra�H���ڰ(�Fh�$"O�@�̈́�D��p벧�* �Z܀�"O���'E<Sy:�����a���!"O�Q���V����':�"�x�"O���ÈiD0�y�;b����V"OT�z�Ƅ1X�Aa�^04�
""O�`vJYN\�آE��`�E�1"O>|[��ܰ;�r\�E��:� 0$"O�q��P -�EҔ��t�q�B"O�
BA�
���f���J�\iS"O��S􁝜?Xdh�*	�J�k�"O�U�C� �RPPQ�#Kт`�5PB"O��#$�	s�&I[dI��$�Fy*�"O:�p�ŃHG^, V˗45���3"O�q��F��)Xh�Ѣ�[-")�u"O&|�!)�����Fv��+�N�<�@ �+���j�*'1|�}s�%Bb�<I!�l
�<8&
6ԅ�VC�a�<Bi6�*���E�+7���1�Nr�<��삁y�"A�Vn� W�1X���n�<��#ءq��\(���n�t�C��n�<I%��#~J@�G�	����`�i�<iQ��&�M�š��Ԝ���BFe�<�IH+(�����+Y&�a���{�<q�f�7n�xC����{t�v�<ɗIʸ,ք�IЈWGЄE��*Gk�<ad�Z�����"kZn�@�NC}�<�'G�rv�ç��gv�p�Nv�<����:?ZpCAk��R�xA@d�z�<�"Пk�2��cD&���k�z�<qE銏����L80��]3&�Gk�<�Q�� ʒHB����B%#��d�<�!է9�x�"��k���Fi�a�<�c�+j��d���QJ�Z5�s�<9f	�P�`��0�6,�L�!S��T�<ieo�$E.�sf�=�zmA��P�<Y��QD��K���6]���X�<��
�87��b K��U�Ơ���o�<��L�&�[&C�6*<���df l�<��'Lt����V�zخp�!��h�<)�۪>��;��4 .��$*Gf�<��ں v��o�2]�~��C�b�<�t��M��	@L�ת���H�<�A,9�)rTQ�=� A�$FNE�<)p�Щ��:�������$�Y�<I���"UN��
��W� �"%�ėk�<�6Mȓk"��F��,Q)fT�t�[�<�e� -*W���BD(( z8i�bW�<���[�	�6�����9�hup[�\�ȓ
��(�FS��	�6��'��h��l��%r ��=Z�Z��٣'�੅ȓh3�9�&.��'w��҇��!]j@%��[+X�#�k�C-�9Z�ᓧ"�v؄� j�H�+
��
��#0辸��QVEqqȗ��9��ʤU�><��
c�(k��Ԥ?9�¡�M�[���ȓi-uh�oA56F�)��噈F��ȓ\�c"�̡:Y|�K�D���>˪�r5�яGL��`��&=��S�? @1C�F/Q�rD���җ��{%"O��s�UZ[6���C8I�>}�"O~U�!�O>f�s5�-}�6�9�"Opx�U�N�tJ���񀟋`�^�4"O�!��n��V�ە�l�LY@"O�6 ��u��ĳ@�Tш�{"Ozs�CWe,t<�2�U�M�:L�d"O.0c�g\68u�-�a�U&g����"O�ݡp��r�j<§bN�鋤"O��{�	�1i�zu��bإe�4���"O�Us����~���)��7��"Oԋ���5 ����ەi�vkC"O�m`�N�,vw� ��F�@�֕��"O�\����Fљ�뀙u�<���"O�=b����a�*�6��|��"O�=R��ؽ
�"�0d���_�.5@u"OZ�S�NJJ�f|�W@Z�`v��BQ"O��ćO|��(�蕌d�ir5"OiB1�)#Nq���P�d�2��"O2���:2�c�	�$��]	�"O�U���	�f��
���Qe� ��"O��9���F]ZQJF���9o|���"O�d3�$R�S��p�gF�jE��"O�Kda�h�����e�<�>���"O(Dc$-�g��%��O5;��u9�"Oj{5N?0!��W�G"^��|q�"O�L�ǘw\\�Q��F�*-"Ot�ʑh��X28��Ŏ�Gkt���"O��I��ŷ �h�b��ibP*O��
C_$&�uʱH�+4Vf) �'b�X8&��<?���������Y�'�8��&@et�	M�fT���'�B}�S�̌��Ij�iQ�A�\��'ͻ5e�	X�f\�r���J��9R�'$Rd�6��UF�3L2/� �
�'�n�ku#K�%%��:p'I�(�����'0@5�ÅX+yW.�A@uc���
�'�lP�e�� ���e��i	�'^1a���/�r(�L�a36%��'ȼ�!%��5��=b�@P5`�x�h�'?�pc�ȥj���B�ǰx^���'0d@H���Cg�`�EΦ-�
!y�'f
c3�@$e���&ƃ�}��]�
�'m��a0'F!�N�T��_@�Y{�'�����H2�T�l[,�Z��'G)��*Y�Q<��/�($��'2DzB�ӞYm�aRM�"�i�'8��B�Ëg�re�Qo�MS쉳
�'�|��G��Z)h\⡁B�G+N��
�'�p���A�V�h8��E�*?���P�'��K��D�'�5�Ed�&���	�'9並��3���9d�ȃo6��Z	�'��rA�PU}N��b�6��D��'2e �a�$�r�a��+z��'�"HB���&�	ŭ�x�̍ �'nYxv.��OK�%��#��[�2)`�'���Cp�U�&L�VD�+\'TC�'T��&��>H,�AՇ��#��=�
�'�`�a��7:��q)a�  �
�'��l�rn�7g2����K�H����	�'2~x��7{Xd� c+i�6�)�'MHF�2\z�:���'\��!�'��e�k�47H�u@�n��A��Г�'���:-!)���kV�+A$~(��� .�I2+R4j�Lϴom�,�P"O�w +��{P&��U�t
&"O�Q�E��pY��W<t�k�"O�H��@1w$���m�ر�"Oh��)��u�"��VCU9����U"O������$\u@J#�A�����"O�3�j��9�ȹ��f�M�^=�v"O�L�GK��Y`���1&�6n��bR"O,݉!�C�.�>�Q���}��F$D����I�c^i�HŖ$y�z��#D��Ksb�?jz�&�ei<|��@,D�T�f�л#��lX��@�P�����)D��i&i�
��ԑuߊv�Yҁ&D�p�����Y�f�-V�0��bi%D��e�7�Fe�G�"�6��!D�h����`���z�jA�c��h�� D�T�Fd2"9��e�/Vގ�b�?D�4R��ԫO�h�yWf���>(A(D��c�Θ(��1�w@>�; j;D��q*�'z�Fȉ�DK��Ţ��>D�d��G�l�hn�m���L�{�<TA>X*P��@"ǁ =D����O|�<6� Z1�mrt%޷@�J���Gx�<!��ӳK�� @�G�4	�Ѓ�y�<цC�>e6���FB4%t��Țq�<�*�,�nhQ��/s�Ƙbu`�n����ɰd��˰�i��v�*fV����ô��\�͌X�����O�$������O���%9��8Sτ�h�4��� Y������0��ɷGQ�DXX���+�8Zt����I�\�F�]�~0�Ʌ�1'�ves������ƫ�Jv�r�j�dj^`���&/�*������H��D#_gd��  �uo4�q.ݩ2���?������'�>�� �j��]��	*b��uG}B�6!ƶ�!��]L��U�l��+ɴak7�iܔ6�<Q�o�Q뛖�'�2]>%ū�5�|��s�M(��hva�,l��Iߟ �	Ex�i�u(%&��D�p�ɤ<�<�A�G��X�^�;y�j(���&rܐR����%��=�>1aƅ�O�,A2#�&Hx��0��1 
T$*��H��T�J�"��P����p�� ���ܷ1�msӌ�$>9�O�h|X�H���@�-c�p�!	!�D�O��<���T�QbH�E�>4��5d?!��4�dal���MîO�e��-yA�Y)W|4j��p�-	D���M#��?��|%`W��?���?I�4ת�@�*�tߜ1�a�$M?:ш��S#�ȑK�(
Jy�sw�T�x]1�Z>u���dC�N
f����[�i'ĩ���6^�z�A#�o�ri��Q�_�v�kT/�R~r�>���w#�x8�%�4r��Q� �ߔJ���6"�OBU�	���IBݑ>��2����A�湩��ܧ>< [��'ea�͌�bk�M)�9Y�4Z��]=��	�����4'�������O��Աi�@�P��đ1��yu'EB��ի�N�O<��r&�izJ��O����O���O��i��=�o��<9>	WE���Ciҙ0��Uˢ]+I1T�(#��4��!x�4�(O�pj�f�q0@��4/�U��oN�N��xI�c��(���^�	���u�'��z��_y�p�����2nx�C�!�*wh��pl����IWyB�d��&��p��`	���ߑ@ɘ|�&L9D��Z����c?Pi���3gt�%���u��v�|by���i�<�$���!��6�ib��	E.����!���$'�%f�O��$�OpLK�@�O����O��hD��<2h�5E�f�xInSf��d�eaP�`���ʍ�A����m�oxQ����]&Wʸ�C�̉ui��a��^��]�R��H����f �1Lw�`굮�/kQ����O��lZ�I��90�n�-�� �!S�Ju����>����?ъJ~���Q�I��qr��A��]�b�
x�#=Ɉ��w�~yY�A�r{.5�'皌2���-KЦ1�4��$��Ӽ$mZП��Is��ᇵvez�$�Q9�|kA!b��Xr��'F��'D �O�<5:��s!#�hy��f��b֝ƺ{��	1Z�<U˕AL4v�Fر��I�1�9{r P�7����JY��}�b%߱@�
�ٸ�$��$G
�*�cWLd�|㞼;F�O��l� ��'���_%b��P�E
Z�V1���Q4J����?a�S�O���9I \�fK��>	�p2ʒ��\�]�޴����J��@�O�Meؽp��[j����O��D"��"ғ^�x@� @�?   6   Ĵ���	���1tH�>+���dC}"�ײK*<ac�ʄ��iZ�Fm��x�\c�7�	�V� 9bF�	�|���$���k	�K율g�5n��M���[ ���b�9��(F
Ht����4А$�<6�ԹYX�y��M�Qb�syIQ@0&T�@$)}b��t�L$��H)U�A ��"��
b��
���'�܀I����)�'hl��kl�ؖ't�����L4��HNK?� �p��	p�Tv�xRcA�@<��$��p���*J�a]ةJ��Y"����c$_2���N�\ɷ� m�t,M���чO�r�@��2��(���*���vMJ3UlXhW�'xT�V�	�$Ԣ�'��(K-�sI��$Q�<� ���t�q���)�#˝\Ѹ��O�=��	f��3�5���!U����1"����-zuh���ֶ`��'Gpa�-W����<AA+6�b�f�uI��Z�����@:,���z��'&Fp�O�{}�-��,���7wN��)�2�T�dؚ$p�k_�|�TPa�:CӜ �4�%l��-O(��PoS��dH�<��S�$���DQ�z�.�"�&VX���F��o��-� �#�9��7q,K��>����bE�C��>~Z|+d@P�`�#��O�����`D�9v��6�6r����=.��ʡ V�g��'�V�p�����\�:Q[D]�<�T =F��cU	�p]:���L}r�f����J>)���b��%�ءS�����-��h�W.,��Uΐ�P��3�4�yb��O�œ��Y�B3�d��<I��ϙޖ��U	G�7Q�R2-�q�S�X���id�N/)�B���fݿ0� 0)Y�A������~�&@�}�%�H�34�@Ӂ��vd��Z$��<��$�^��$��� ��	VXO��BBCV�� �(�ə�ԅG*��k^���':�q�lֵ��'*����M01�.e���R 6(�9R I7!���p� �  �y����qIf�,g���р���yBؒH(��KT�c	�}�ǭ�y2��/�N���*�&EY⍈W(Ċ�yRiW�$_B͘7EZ?� }�v�R�yB� 5��#�HI6,ؽx�Mӂ�ybG�D�<Ҩ+�8�`A䂶�y��sY�L�c,6xD�I���y2��e*����̪~�j�����y
� Z���B��s*hU/֊3���"Oj�Ȕǔ�%��y�+0c�"O8���̊=.�~����� OV�j�"Od<�Dh�94��+��"0P��#"Ob�ޯ4V�sq�R�b%�1"Oh|�r�ּN�Xi���#DtB�pR"Oj�`�W<ڢ̫CTA�m�`"O���s	1�c�ȹ"�\M2"O�͙��ҋ*�����!�����"Oe���2	�~�pѫ˚f���s"O���`Ϟ.Q��1�%��8���;1"O��`��S�F�Trc۽��� "O����F5��h#!P9w"���"O�����k��D�@��.5��0�"O:k���[ `z�$�y�41d"O0!���`V�t)��yl�3�"Od}`JչE3�8�rK4�T��t"O��2WCߊj:DU f#�9&� ��"O�E� �U[$�u�B�&?�����"O�Y�*�%}�TPQHՠ;P�bS"Or���Kӝ5pZ���f
q::��f"O��ش�@E���a�F0
;̜@�"O��m��+!�L**�$"OX�Э�(Aܭ;��P�=���h�"O!R��s�z d�6UJ
�"O�U�5JU	E�h��K�'�:���"O$`�!��T�fy�3&U ���P3"Ot�"d�Q�K������tF׍�yR�ޥd��q#A4`�V���DQ�y���71P�jTLȚU>V�ႁ���yb�^3��yD-�? �B'���yb��e0�D14�ŋ	p8���l��yR���S�@=X4�E�Ple{��T��yR)��9��Z�V� =RlЧF�y�	8$� �,I	j����t�<A���0��a�
�Kz�y��DLD�<�3��?��SGD�>��cu��A�<��t��uDA8�b�2$C^z�<�q�^�1��,Y�(�3w �,�t,�s�<�v�k+��bF�0@��	jAr�<��C��!�Υ TiB0	�|�Y�X�<����}$ہ�_���ȹ�JW�<��(�$*m�Y��Q��D��Q�<a��sD,I��O����y��q�"���~�)m���To;��ɀQ7����O7mQ�cz�D"3dݎPHɨ�  (A��<cF}�Ӄԑ|d@��$��	Qf�k���N��OQkl�@�P��I��-��9(��Z	�6$�R���ڳg*1h�A���5u\ umi���A��y�ҙS��*KҮ`�3���@ ��O �oZ���O�>7M	�`���ö��Z�;���!9���O�㟰Gzҭ�o	|���N���dg�ڸ'[� }ӼXm�N�I�?Q��)�n[��3$6䈓h�.f��홂�'r ѥ3{�v�'���'rit��I��voF�J���*�ԡpwiE�X���(��Ȫvp��;�	ՑL����'T�ʔAQd�0���W�� �f��'AL1b�^p	��ӉI�M��JǼA{
���
�~�ߴ0êt&��N�Z8��ǁ0n�)� I��?���S��?���i��$����OR�R*��7��^�L�����wDT|*�)�矴3C�\7^~ zG�J���KFBG�L��fKj�ГO�������ʓM�ވ���\�zO�D�pn5h�l����>��b���?���?I�P��?9���?��j�p�Ub5B�%�x)��@	n�슰Q�Y��p!�Y��@�� ��2�=Fy"d��cذ,A"�ԝ(��Թ�A�m<�4I�NJ�x��|���yoD����
=�z<Gy��ǳ�?�SB��|��!�J�T�o���U�x��'!��T>aP('x��X�vꔇql���'�����GH��X� �󢢞�@���¢��x��4(�\� �5��M��?ɨ�6���͘5/n@iS�턆�R���jӱl�������I�9�޽��M\%��r�� 
(���L�,X���z5U�c=V��+Ĺr�\����"�)'�|�f�Y JU�\x�-�F�����6cL�����ŖCh��駃�;/�
��&D3�o@4��ɩ�M;����� ƨ�v��|��-���֙�4X�1e����'���)�矔�6厭~%�uxan�n���CeI*}��i>i�ڴU��&�i���#�_XI����f�ް��'�*!NkӲ�D�O��'J�A���?��4>(6��*i�E���[q�|���y�r���\�qZ�-(Fa�Q���^���?ᬱK1T�ю�4Þ-1�m�*-nLlZ>AL>�Zq�Ի�VMFc�>�" ��P�2q�k�U�nk~�H4,Q7BV8�OG%,��M�/�?���'^���'-?7��(��x���rJYZ���3����Oh��dM+'�
��5!�� 0��`�3|qOD��˦5ڴ��'�b]w�.��N�:t �Th�	������Od��W!Ғ4�S��O����O^��Ӻ���MK� �&l`��"� :&"m�'���$[�ku!	�}�(���&[� (I��OaX(S� D���cr�p���
�C�i���Д
���J�A,���{�E�6���#�Cu��!���j�%��B�/��¤�Ȣ�jl�F'�>�G��ş��޴W �'r�'��	 �z8�4��?u�x Z"$�")��>���#�L^)Z��YJ�-�);��hf#K5b5�7�@��Q'�L��?�'��oږPO� �  ���D2�H��I%i�����`?�$Bt�nhT�����?��9���@
X��=�W�H��O�oZ��MM~��'���4Fby#�E(�t!g,'ZH��c��'�^9;�`^p�"�'o��'�d������æ%D&I�)A������Iׂ}�gzS�����j�0����%d�af8�?ɖ]�A��T�w˛�3� �kөCĢ�ɢP�Ļ�J��t�4	�סoݕB�����OT	��#�����*B�;n�0�տivpd`����j$��O$�D3񄊨:�|�Pn_:|���C��D�E�Q�T3��d�~"�+j�hV"�q@4�c��
7-,���e�U������2� �  �o9�r�-8j:���\c)�H���*f�:tY�&H$� �ڴ6�I�M��P���=���'�1%Ƣ%����)'^⼻î�����yX��+�d�7�mK���<���(��Ɵ�AݴL���|\?� �f �pu0��eIG�'� ������?)�� ���)茊�?����?���(���O�7��~��bحx�L8���<wC�L�C��6l ���@G�7�}R4�K�?�����79��OB�Ar�Uq�8��T�3o�)�"*�.�5��!�^�X%�q�ի����P�'�|��ˈ��`y@a3x�����4��$K
)B(���&���	�,�'��4�Q#t� �y7j�tپ���'��}R�io
9"���$��dZ@�!��U��fPܦ��ܴ����<��d��M����I�/\����cү	��t'��?���?�<8��S����Y��U�#� |V~�� c��G���2Uk�%wvΈ����4_Byxd���d�F�;�!!�jn�@��^$=(���c۫Fʨ�
X+\j�8�t�^Qj!kTJ�1�f�F`'ʓiv��I�Q��� S��j
d*Mb��v�i����'��I� �?�O<pҕNݷy��� ��&O��'�2�㔧�<�X�Gi��ma���O�-oZ9�M[*O���������Oh�@Q��J&�:��"�׳\G,�ˆ&X�V�����O����)XL� ��E=��E�!呪i2�@���a�2�'�U�N8�l��צX�V����I��ꝫD�Q�z]�ܛ kڦn��9�����J� � �M,P��I2L��%c割0�4�$�Ʀ�N|��4���Ò$\&j]r�)��[)(���'{�O?�O �"`�L�<�<Mh�g��zu�:���	;�M���i��AL&#{���t��0B?���2���͟��e�IA�l� q� @�?�Z4;6��;y\��cŔ�7O8�)�iLg����8��0s�̍�V�����ŋ��U����o��)n��a��_NP9٤���=�d�'_�r!r����ԙ�mٍ��(%��#%L�OP�mښ�ħ��'"�$M)'��	����$IR��?��Xq e
��ő5�z���Jƃ=���u�i>�X�4S��ƚx��ފQ���*a��);�pHa-F�t�lZ�����ğt�,5����	Ɵ��I󟐮1#������Q�p�r��J�i_3s�X$$�$����p16�2���?m�Xan�;e�'��Y��9e��T܆2������Q��!�R�ہ{��H�L͖�q��$h�Aܼ�2��!{��!th�#P�
�(.6��yyR��?�}�I���nZU��u�E��9y/�JCEN4:f��L>�7�"���M\;!��H�����oK��?鶸i|\6(�d�|:�O��р�"h�`���E�UU���]\j� �N���I���I����O���1G���C��5�B�J��R�{sL���&=<]x M2#��e�t�1g(��1�*AruJ&H�5\�֔����y����e�C����&C�g�@�M�\.��K���>t,�ڷ*T`ݪ����M:q�Ģ�OR��IĦ��5�'���d��_�z ��C�Glhz0jߨ3�!�D�-�X)��'�,=u 1��7�4ܔ'�"�`��lPy�Ͼc-6��O6�i�23�÷N<^���B�Q� ��I�e�ݟp��՟���k~�x��G�g�`(2�˦>��QS�&�����!�W�[�V�ð��!n�<q ƛ�
�4�f�[�m���p�]�a�^� -��P�ْ,�}�E�H+nN���u剞_��d	Ҧ�[�'j�P(J������M��}��'E��'��O�vM˶��z>U
�	�8I~X��R�I��HO������ ֥��ѻ~� ݁I�'z�̑7o]��M�N>���?!O>Q�O����	  �,J�IKN	8��'<�'��'�'T��@ �������с]����/Ͷ�(Ot�"���/]%lZ'��n0��Y��27C$\�5�9�\�uE�F���bO��(O��ֲi�X��C��Y]D%"N�^��0�%��蟠n�Ꞔ�'o���O�PC� ����*�V+~$
�'��ĹQ���RvΚ�'�Pa.?U ���dyߴ8��F\��he����M����?Aش9��q;�\b�}�5,�!q�J��S�'+Jy ��'���'��J¤ДPrH}�g��:a�i20�,R,�)��ɐ��( [#JC���E+��V	�(O���T�#���r �?��bu[	�X[n����X FD�/6�Ĺ�A��(O�*��'7�6��G�Ƀ�o�n���0F@xd,K7m\<�	П��?E����Z#4K���1}�$���	и'��"=��Yg�L-l�$3�`Q<
Fb��4hZ p��]¦�|��'�B�|��x��
�/ D  ���3 ��{�q�+ �yita��C�=Mʧ%0���L�<ب˦(�s��%��Y���O(�Iڦ�	K�'T��x7�A�N���_�*�"��=!��°<�q�A*�
 �lϪ8
l(��J�'p�g���m�A�S,q�y��M�JȐH[6́���9��iB�'�r
��`H���'���'����M�n FA�4ʕ� ֐Xc(ݮk�D ע�7nS��q����I�O���K�C�,C��Z!TM����+v�(�T/�X@�W� �vPS��JL�Ӥ�L.,�Vm�}"Q�n���( P�B�dޕNi�D�"�Pk����4n��(�v���'��i�r���E�?P$�:c��!l����o!<O$��=���X�V�"���_2�EO�R?-�Mk��i�h6�?�d�4�I�>Ip�:�v �fD����
WˀM?Y�S�Z� `  @�?˔��/���_�=��˧�u��7C�l��KP�Yn���թ����dI�n��M
�I@�z��;�i�_���/7��'U��%y�]t~�JfJ�+��˓uC�)����Ms������q�C� ƴb�V�"���jU��?	
��
]�.ҹ?\ȁv̑ 6bXDy�'v@7���$�d�;�j�K�J����@'߈Ct&uba�'���'���Y�M�>�B�'���'j6ם�����.�,g~�C�d0�XA1�ܖ���S ���kd4�C	�=���?%q���~O����a�DK�5�>0zAe#�Ɛ����"��יY9�����w0���SrA:����;)��u�J[ξ���χ(q��)On1���'��%>��O��dzӎӀ#M1/���Y5,�C2v�)�>��RV�����g��� �ɏ&�u"�'�`6M��&���O�� c[T��*�e�$y�����=9�D��kS�X�x���՟�I��t𯟎���O ZFf�W�W���3,]94����Dϙ�g�8u[6��
��K���~�t-��	�k���ZW!��5�)bmN�0�{�OU�pN�J ���h��W w���x��Gz�7�S�j��8[���ȓ �'�>����Mc�����O
��)�J�p��&.��a���v{!�$�Z�R��T+S)%?���ϵm����O6�mڈ�M-Opx���ަ��I��Lm�2��i�1�X9Rt[s�E�!i�-���B�i	���?���~�'I؎dURlr�lH�8|��Rל3�8��̛8An��� �B��I��iNF�'�$��.(5�x��͹u�Z��3o���1���P�0*�ܒ��܌|8D��,�x�'�&���r)�6�3��̮g�ޭ[��5�TU;AI)K�����O�⟢}*�IC������^�&٘܃���`ܓ/A��d��5�M�r��-c,��i�fU�� в��`rK>���?�J>9H<��(�; "  �� P�|ځ�'	47-ZMy�����;�q�'�5"c�:D���=j�i���'C�'ay"��5N�T[ı~�UBu�����ɟ,S۴&!�f�|�Y>�mZ�7Wp=�cBcL ��B��9t�${�����@]�?����?��lD��ڟ�mږ\��@p2`qjE�J3{����f��(��Qr�/#t��Tl�\�vA)�)�@��[�����hj��L�w����M��S�˖��P�-�ʺ����E�|�DR���I�޴�W臫.�y��B$}L,��|���iX�^���	^≊q�����%�d��` ��C~$B��V5�!HT	 P�^�x�$�R���`��i��	ޟlxߴ��/O�%y3�����nڟԖ�
r�^�(p蔸��i��?���Xƀ�c���?9��r��t�f��!"p��@���AP��:�gA�#
�샢b�
Ԯ��V�C�(ʠ�1�De�'.��㡀�~9���N+H⅋���z,��ZF�@6�	�g�"6�� T� v�'F
`��5��HJ'r��xgD�7H�����T�v��A�O��$�ON㟒�����s�\�.�1T�x@0��HO�}��%�$�Fm�s�RŹ��^��0hŰi�7m:���O&��=��v����`@�?a�LX��t��B�-)�T��#ۦ*?x��G�c8ܱ�2K$�S�,����w �|馄��g�|Ѳ��K�oت��	֟�l��8�Z���)�<i�4>%��I!�g�@�J�E[Z����OF��k�0�\�G��F��Ec��On�Mަ)ܴ��4���i��T� 0�՛th� � �QSē�)��1 Rk�b-d��!�'ob�'��i~���ߟ��	�@R�#u�K�l�P�`%iQ>�LA��ɔ�vu�����`�Vm�`l�
�	"��'ʓd{��{�Z&>���GV�HX2�lL9sq�U�a�Y���a��I>�Dz�A6�F6u��z�ɢFڮ8OH��l�ԟ0@ش
�'G��''�O���ӏZ�J�B�����J4��t�d[f�']�O6�Q@mԘdT�b�#T����se2��ʦ��޴���?����!��i   �*O~�����O��-J*����ͫ|k�9���8/*��$<O��Of���
�0VP��E�-ufA��>Q��zE�V�s�f�O&�)�6-T�\@xǉ�r�J�d�9����>��� 
  �Ӭ�P ,d1_>���Vi�`E	ά �Z���2񤒜Y��k�<&>=$>Uҗ!�;r���s���mL����/}R�'��|��D��C�"1�W�h��-�Cl$E{�O��7�C릡$�`���EH򠺧��Ͳ3�\�ӛ��'���'$0�ô������'iB�''k�P��A��_�C�ꔺ4��c���R��k�8�-@3V��D2WHH�D�O��S�:�?��m5.J�x�fRʒ�{礈�.�����Ɲ\����ϿyT������� !��]�.�X�8 �V?�Y�#�#B��e���'4���'�p@r�������b�P؊LJUc��Z�i�fP�3EH<�� E�j����
��22�0�b�t?���(Y�&�k�X��|z���ڪO�2%��~�(x35��A�d�[&,_�Q|�I��	���I������uw�'���'$�U ��B������+�P�B�矨%I�,yA
<h+։�ӬY�41S����(O���AAJ.,��`"�]Ũ�2�K��^�t��@�8
)���J�W��8�vG��(OR�!�� �����(I9+��X��'BD�m��u$�@��؟<�>Ë�6��չv���#x�zf�N�|���%>�;s�A ! ��&���r�F�:'B�=����6�aӲ�OP�D�O')5 l  ��m8���#݄�q�G�L?�a�zG�F�'?S>yq���T�	ŦQâ	I�f���6.90��t���$�B,�b�[�∪��C?q;T����� (L�.�`�	i�	�¥�2{���q -�f$�jbHe�"��	��.H��rC��j#Y�CF�U���(��\co��ʀMC|��	�`S��H�شP�����MS�W���1�禵 ���)|5���J�pΰ�A¥��(��Tx� ��'�̤��oɕ��,RS�V!0�أ�{"�'��7mѦ%����ٺ[U��@��@��Ɣ�+�riAGbX�U�'�a{bip;   ��&?���ߺ�g�Wؾh[�D*�t��.Jyw��'�J�P�����'���'�
֝��4m-r���WFB'O'`i��A Ys�P��.]"ER*Hj�FR5K;�A���wcϼ|��&���fJŇoNj��M9]�:�2c��3Z��؁Ն�
R�d��t�6#���Ԗ@��M0�R|�qk!Lجu�`��1N��s���`�z��]Φ��M<I��?�O0mN�^�D�Bvl�9�pQc��ɐ�HO���6�.�v��(]�l!�!�N�:���i7-6����0��kӒS�  �u5�j`L�~��E��^:��lZg�q��5n�uPu�i7B�'���̙l�d4�0K�I­x��� (�<<Y0A���?Ǭ���t���EC\�j�i�0D�����M���IAy��uۑAԹ=2��ψ�r��'(�D
vZ
>����	 ];�;�aJ�m*<��OF��4�\�2�:�:!�]�i�K<)eB�� ����M{����OW���)M�L��q��M�%Z4컊{��'Qay�O��-�� FA�� T���<��O*��U�i
�4�ħYS��aT��:X<lYcࢎ��m#ǀi����O���O�*�LЀ��O����O��Db��H�  !`	�4C�,������e̒pb �U�F�}�F}!��T��A,�R�IF�UO��k��'2p����n��u`�kM�8�s'�*+*q��*�?jn(��U��;q���"�EƼ���D�'z2Iׁ^'Q�3% C�h�J6mAsyR��)�?�}�	��l��z��YQ��0?zM)W��^��8�wqO� &��*"H��y HB�)w�] �OZ�dĦQ��4�䓲������Tm���pL\�w�P0��ûJ��1�O� ��	�  ���>���O�6�F�?�
��E��r>�{�f��n����'���&%�20��2���8]2�Y�'��(v��9o�d���?���i}"JX����5�Z�
phQ�I��~��'�ƹY�  ��Y��m?-'��r�nF@���.����F�i"fO����O ��i�
�,�{���41@��+B��j>��H�~��mG)T�<Z�G"W����[n��ȦM�ڴ�䓉?�����DE/;� �  �R���>˓�Ms�(k�|�7[}����e�='7!�� ܭ;�
��8l��b��Ē-�Vyr��O��Kզ���4��4���I���a��%��%£��H�M�WS` F�ޡS���1�'�r�'$2$c�I����X�I�R�[���?]C���_@N�I�-]�]�T�6�H&YU��(G��N�U��"ʓO|*���Ap�p!dF3sq��6ʖ'6�
}��atO��2�!@�W���+pn=���c %ϴE���CdۨF��)2i
ޟ\AٴM%�'lR�'��O6��Q��,���pG �<F��C��dN`�'��Ow4�@,c�H�c��	�H0s'2��]ܦ�q�4���?	���5+��   �����*��ҎK�c�(�"˙�|�?E���q���س��`�P����
Cϔ���I��rش7ś6�i��`8r�Fc�Ρ�F��)M��;�'�h I�d�|���OV�'	ipA1���?y�4{�!�t�W�sڐ͘5��<w8̲�!T(z�>�3$�Ԍz��|r$O�Ah,��7͚�D����?y�1� �iG'�NM��0#�պQ��	oZ�0�{��� *$.̺UsŐ�8� ��A��;g��+E�����Y�7�&y[uC��7�����k�4n��韢"|nڪ�8��*�]����+X;v�	ß$��	�~���"��YH���k�� A�e�9��'J��ڽo�z��?��;i��� U�wǂ!��ȥ�����|��'7�L� � ���Fx����@�Iϟ��[wOr�'�¢Ѓ�@9
F��O򌝊�'�Y"�+�W�s!r,�tHղX(5(�$"���J���гP � �� �-Od��b��&_�P��EB��F�L`�1�[�:�ٛ�I�hPV�����z�? "|{A�.F�zI�����E{����&쟨hܴ$މ'�b�'u�Ot�x� \�V�
Us3M�e���D�B���O��'jy�R���xW)��&t � 6�DF���4��D
� �<�n�̟�n�j(=5�ɯyPP۴ �>O������?��AZ2�?q���?�'D4<?
�ʷB�|�N 8B�^��*�� ��	�2���g��5	�HS�h��Ey���.�8�EM�^�<��o�Z^p0���$� Y�%˭�e���i�­��d��~s�z�v�n���q!4'�&Y^hs�+�/ɠ�Q�%��D�O��b>in�-$�mc%Ŗfܢ0u�9VC�I��t\pR+Az�Q�,6��!O�%�M�-O��h	�P:<���O�ʧp���8�4B��Q�"��m4��� %+���!4�'NR"C�68`���� xf�tPҁWRv �C���,le��C�W/0�Lx(�iF�]�On)���i����֫�C-����P�=v2q�.��|� �$`�I8��x><��xBN/�?1»iG����)��ȣis̰c�gޜd�D�)'���O>���V����j�7�衹��8�*E{�Oݺ7Wۦ�%��I��Q@H�[Q���R7\)@ �E�ca�6�'T�'�������.&��'�Z�M�^c��!*C&P�9r�d��f���c�Lє-��a��::( cF)N<���'�SJT�����I ����*�(���0'�J���,�+#��8 ��)\�6K���[�'l�N� 4��`j�kZ�d��Y8�(k�������M��Z�\��@�Oq���'��F�۹dT �0U�X8��������ēO,��ē�@؝0�τ	rf
E�0��ev�$�O@ll�4�M�O>�+�p�4�t��S�!.��() ̀�$�$�I�,ԙ w���r�'���'����~J���?AV"!}ց��EȚ�a��@�t~������#z����K�KȄ A׹759Fyb�_�z�@Q��NY��Iac��'��9q�	'e:�p�'6��+P��'TEy�a�h�T�C�ȣ--Re#@��3(����5���i�S���	D�$XV��%�(>� �j��A���ȓzLp���O���3��_.��aW�|�I��M{t�i�&b>Ji�4�?�4H�:�dM�8�*����3B�Y��'Q��� �"�'�$�#��S/��'6�5ߛ<��S6oS�S�H��W��y܌�cpF�U��	H����P��T#��K�T@�@<�P�qH�'}mb`�ڴ��p��8 �ă���<H�"�z�h��Ot�����&A�T�T!��
�*���?i������O�(�Z$k�����nюW��l���D�E�'���բl� �����K
��ǔ�^3����eӼ�O0���O��OT�(F� ` @�?�E�JH:�,J<ql�$�O���7$�lD��6:��+ea�p��K���Fo*�7��M鐈2�����ԗ8�Q�L�PM�	ZLR<��	�13]�Q(bO�
��Ա�$4� �+��@4)��R6F�Q�lk��O �d�OB�d�|���ܽn�$��F/z�r(�3 ��?���9O���W��]}ܹ�c��ɺ���'�O={�f�{f�P��"]����O"��#�R��"�'��8T: �	ԟ����9x.�k%�ޞDr���Jː7�yQ���`�l	�J>�Oz1��B/Pj���/��d����Jc�@��#۳x��O?��X�,�x��˙:�ܩ0��J��MÂ��O���OX��9������FʈRl��5.j���w���nx�XA�*C9 :�U;�Ǖ� �b֍1�&3���'c�͠r&'}�虲j� "�A���?Q��V$���y��?���?a���d�O��P�Hs����flͲ%\�r��`D`(�I�N�&�Z"f�7z��̢w<��;�y\�c�K��B��dC��nU�5���~Hx Xa�]�vS�T��i]j!%̗g��c�`X�O�4a����	�,�8�sL�Ɵ�Y�Iğ��	֟��<!����1V&��i�%	�Gr�D2��^��!�d�O2e�f�Z�%gh J�d����UǌI���T�'I�I�1W~��4T2��!'͘b�>�!��Z�^��)��?���?y"��?)������= L�@9F��M1�j�l�T���H�h0H��݈D�^=p�`���Ey"k�����0�������d�թʠ��0cV�l�X|ZBM�yT��
��2Z�]Ey����?���i���BG��1�V|�1�F�/��u��l���� ��9O
��ET�]��@�O<E"��P�'�ў��5T1��b�;c�$��� p����4�?),ONHi��z���'���hz��N�<��kG B n�@x�&����I�Dx��ğa2%����,�P�T��Ys��1f��R&,�� ׹g&z�y�KL�A�\�<���ۑdJl=(���"WU�7Z��h���,	>`$z�S����Ej�NA�<tFy�C��?��i�*c?U[�J�T��[fA�+3�8���)s�(�I{x��4KP�)΂M��BK�HcJ5�O�'���LE�Hܺ4
D��
hti��5}B�i*���� (u���+g�<9�Dʌ\�� s�"Oj]B��h�ZK%���t��;3"O�Qrʚ92n�@�7�v��S"O
U��-�1F}T=�q!yr�Y�"O�f��b��c� `u���"O��!��%?�-�w
�5Oz�d1�"O(H���o�!K�"�	*v@��2"O�=i�͆�|I�-���E*vm���%"O�aHw P���8W3��t�"O�i@DQ67j�s%ܗD��"O�`r#��8���T @�,q�f"O~}1F!C�lۜ(i�o�\f�m�"O>3�I�^:� GO��|��W"O<�E�X:� ��3��
PszyҤ"O��iJќH�t��ƣ��*rs"O�x3�#��Jy>4x@c�# ���6"O"ai�{~N��.0��P"O�D�࢘�H�ܪe�W='[�"�"O����<F�dp���M�I�"O�h8��77�=�u"54���"O̘���ɼn�����7ep�G"O��`$�&E�J�J�$Z)��m��"O(�t�P�d�b���A/]����"Op4�� ʹP��`J��&(̍K�"O�� �E��$���� ��F){�"OV��Ʃ��H^4�{���&(L>]��'��$�	�!E��7Ƌ�46Ѐ�
�'O��Q�ɇ<m;',B�:�b"�'���*�e\�/R�mv��7a:�!R�'�hU�B/"+��x�Î_��U��'�ę� �
�6��Y�����H��':Jx	�m�5^~�C��Ԩv �����@^�˓#��S�O! �X��	�,�+k�ּ�@�ޔR��I�$)\X���$2w�-F~"6eOx�ǥCn~`���E�I[P(O�L���O���'u�u
�'9\��(O�U�c�	)C�0L{1�d��$85\|�Q��0ӔWCPlCB@\������:Bߐ��tϓ�q��{��˹eCޓO�y��ۙ%��"~ZC��8%F0I�ȋsʐZ�/۷Y���'g�#� O�/�����(f) {M>��o&���Ӯ�>�h����[��b
[k�3H��Χ~m��w��.�'��xumƅ}��D	��� �Z�`�Wf]ڃB[��������&I���f=ڊ��"�/�nl�`����AG��b��J��;�Ӽ3�)���Ѷ)֬� P}�dCn����?���)��CF1"�K�$8r	G.~���6��p�"�"���+���Ԓv����D�^�NA�ʁ9 qO��y��,�I��	 �v�{л1�������?�ju�S�I���De�|������f�Hg'�_�qO��� �\YX%Ǔ(�^ͱ4�Ƭi�\�X�pk�Ժ�,�K+�y������\�:O�L%&	g)�v��8�U��Sp��Pj"�?c��P�%�1}zZ�)C�-{�����*U�rѣ��r��Ҷo�(<�Q�杁,|0��g��<x~��FA�ow2�'�������I�1q<���ތ%ʦ��2l%���ē�]��Љ��H�,zh-�R�w�����C��[:`�oǦ:���[p�'}vm���L�E����+��K1�P��aҶel��
G�ϾZ�Ʉ-K���O��K�)��	�~{jΓ}ty�B�Pkc���c��s
|x��7ktt�'��(���T?�~be6�L�O�����ԪOm����ܹ-gRQ��˚h�L����ʾ^�a|�@B J���+�띕Q��B� Φ�$� �r>�X�I
d��mD~�;�U��DR�Z	��� �$�f�"O��
r�ѴL�:3AJ8\�j�8�!O���O.5�r����&I�CCT'4����={-Z�c^�J@Eĺ>
��$F"j���S��� e���5.f��*T����e_�p�4k�<!�dr �; 2H�G�*ғ(���c2@\�C�ִR�%7H쾑Ey���hp��a6HL�,ֵP�-��d�/B<\����S�[�Ƶ����pHV� ��ը({<4���	 8����!��$�عÆ�oz� �K_�J�")I�ɞ�{�l�����i���]�pU��:uG��i�Ȩ�`�2*T��'St�S����3&��yFD�(��H�;FY��9g
9��?�{BL&EH)��@���$��u��7>q���qO���b�3��?����2�� ����H4`��Ȁ��I!^��R��7$T&��I��ܐT���B`,>��,��#��r԰�ad�����ÂO�S0t��?Q��������LC0!�]��	@KFQ���� A�<h�H��H[�@4d��ΟJ��O���\�ذ��&��a�B���E��Sq���i�"	�"�(ޔ):�i�aCDQ���A!��x�dT�Q->}�J��sp�O��D����<��JC�S�$��xI��\$ݨO���Kۏt�8�If$��4�׏	�(W�9�6Ċ?}~v�6-��qO���2���K3Ѯ}��1�T�'�|�pƅ�D�I�<���(7�\)H@�S/�������O^���&��YdL�BNT;Q�~}��+�?>��;9|֥s�)��i�ȈhK�̺� qt��PWMh�X�2�݌k� ��HW�Mup��3�	7*��]��dѸ��A-C	`�Z��2m��is�h�a����D�~�E}�w�~P�s"��lA���
F: �H�|ۆ��y�S�''m>1!3Cؽ�b�����5y�Eq��#�r���9�!F)n8|]A�oL4'e.3Pjً@���ZV�X$58T��� ��'�T����$�z��Q�%�V���gJ>x�� P��$�$X���xC�f&�2H"�NӪ2�M����5���?�Yi�U)�g
�L���'�����` �%��>*��<}2Nӓa+Vp����Sjܠ�lS	Xc4<�j�IQډy!�,��ʩ9���.�3W^��!V��������9mR8q��Y<"u�H��H[@G}�wxraiem�>'����7~6ܤN>��5z>�� �<9�C�ǌc��%6���QTO͔8�>YtĘ!q�JX`W�8u�M;e�B�K�bH�3a�o��`"u/��qQ�����D<�	w��_bI�+�2"�9���{�8��N�G~r ->w�ph�+��O�p$SB����'�v�c��4�(u�@�}C����d�`��"F�X�FP�P�|z�G�P�3�ݒ^">�����U��x� U3��,�!�Sh���O�T�4f�)r�����NQ���!l[%��� �M�,n�+�/Y?��O�N��|F��;�∅*���(g'��S�'6ў�>	�V�%J��%�����=>&H�Ɔ��.�Q�X�@�J�Z*z���k��+����A�6� ���Sv����f�'<��c�#���J���J�v_ �`�<,>�: g�%��c5?�qH�(0�J�I�H������#�i>%�BB"&��`"ߕk	�Eq!�]o�1O�Ds%�-��T�kW�'��M���>#[�*�M�8`n�`)�'����hFy}��,��b����rv�L�fؒ2��1p�#A�[��)�6`�9�,+�b�>�G�A{0�>�;t����͝p�Y�DeȦ1�MA�?�O��o��x�.w�vDЖ�WT�x����7mBQs�O����;D@0�fS<5�V *��G38=���AT!c��P�j�+�5�׋�>��8�T����$��bN$t#� J�1v��'
�����&��=	�'�i(�LRҘ��tAM1�!���P<%�&�=q��5�HdT��s,i4h��Oȩ��Hb���h&X�S� �J���3K/L?��b��E�@�j����~�c�"~��4A��`-8����~	����#6�B�Ўӡy��m�h[0-��=`W��	@m8�S���.<��2��G�;�n4��?���� ��˕
D�4p���|1�L�[G���	��$���ҹs��������O�ș��\�_,(�9��P��G��2z������A�A���p�i!�c����	C�8������\�����&r�8aa�F�Z����bH�G�#e���3�̀ _�B�l�ډ�P�,�I�-�j�p Cڳ1N���oa�����'p$=����f!R�d�mj�rOQ����dc&}"��e�I���Фa�t �:2�R�鏄m�x�����>I���"�������S�H�� �%8�(�����^`�)4m�4_�P\�7�B�O��� GEبd�t��ꃃ^|�R���9�'�|�A�ΰ�PA�+F���O~Ҡ�5`2�� a�?+�8�OMZ�>"�.P&��c���E���&� �Q$�8J��I'��)f��9�e2l��"�C�PJ|�a�Q�ʧti��'�@����<c�@��,S�p2|U��CX���$I�zad��×� ��x�c �#1qO�A\�zs&x� iN�	��(#����h3�l�&�M�|qH]��u�M�T	ʬl۠kO������v�`	���X:d*��G����j���i|���>�VT�4KF�`���3G�	��"_d�H��0��;w����8#�M֮>!D��Qj�Ł2�V�~����2kXE���OP$�m�>�S��u�. Z̧%��|�4�3.`��`BlϠ�0 Z�d?��^1�NJ.fD����}�1�ָ�j�JQ�S-Q�j�9ŦQ�<)"�ϻ0��S'�����|�!ҟ��5�ƘZ�ֹ)��L7]t4rSl�^��'��jྸ���܁hָ+��\x��?�g��= `��C��E��k���?,��S�̙�ug��}�`�����!b�X�R�r�����q�Hna(h� E�i���JU�|�S�'T4�	��H��ڴ��(��x��C 	B,���U�]��s� y��Q"��iޝ Ѵ �zRٶn�8��6}��-]�O���Gj� ,d�b���\s�E8�����OH,��\��� �c�H�\����Z�$(���ަ����R�˦E��|+�m�B쓒�a��L$a�	��~3��{'
O`�D�ū>������� JЖh�0� �K_��?� ����hG!F�fmKFȜ6�^x��'I������
0�1cKf�C�Z�T�5�W�-�R��s���t#���K�#x��f$����h�2����S�t�Xu'��pj� h�$S<-�<4K�'Q��b��n�&�2�<��� \�6
J�H�6	��#X�E1g�>1����O���b�Κ:�d-�� G���S�h�fj��<��C.d,�� 8��Q�0��ip�ǡ��C �'S~�S�'֜M��G�>��D��M2�< ��	
/w��)['*D}�	���x�A F�Q �
�.���HO���W��ю�1cC�91z�[�剟u����S��UQ��3gK�;y�z���%��>���O��	D���h�!Ҏ`�a!�O����6+����1%oO��xц[HJi��`�<^�b����H�W���]"{Lԑ�HF7Xq�DR�2P�C�&���	�C_/����t�m��i���ɿ ������
�h����������+�`����V�f�^����+|Oh�jR��
���T�]��q)I =�<(P�睈O=z�@��xR�����a(JQ�˓7�>��'[�����+up�d���C�f\%s�?���P+O�<r����/��^�l0x�L�����).,<H���^=Q���g�?����ʓ$*:����Ȇ��c��Ķ{�|��!�T�mJ�&��Nm��� �"�C���w�B�ie/��M�v@��A^-2���M��`�\�S��R�����S3?�}�0�øP�t*%M(�>"����ˤa�Ƅ�����ʈ L^;m.6(�l�L�Jd"�)#�I��2�=كߟ4d'H�rd�yj��?0�D�	ʄBZ�\�'�j�H �)y�m�@�mV��{�'ER�ٰ���P=�vBJR�R ���#i�^�[6V1���'UNI�OXA�+�-'���9�B-Ev��ʑ5d;��p�"�S.*c��3�	FT��C��w��qˤ�4RMjc@H���dhzce�:�H!��4��"�̓.ZFݒ��YY���ř>�!�M�����O��T����RV��j��P/x����$&_u�'�0h(aX�=�c�������$L���4�'}��w����'@� s��k���	�������] w�a�+>�tt�1?!C��9�����e�ڼ	��~�?e�媄�w��\hF�\��z�B�l@�.J�Oz�@�dp>�ycݥ&��T%�>!f�J<D�� ��m.B c0��1B�>b�J|�@:���3��@���ün�~a1e�K�_bB�;�C�k�<���6����!�i�ёU�X.<RY��D��=>��qf�<Ia�r?���̟��������+�<!�� B�$��D
s���
R&�E���?�PD�6R�̸�#X�����u��H(��Wv˝=�%�GҚ�$	�K�<i��~?�3?�����P�X;|28�f�'j���@.8D��I�+�� OR��$%��E%�}�`�7D�`:2%��w�$@����ŤaH���'� �)�JS��6iه [�P���'5�0Y�OɿR�������6m�X�'�^	�$�]"X|���!̧-S\�r�'V�xS@���w�"Ȅ��U|�ى�'��������%b�Q=�u�
�'��	P`6)n4=�W�Q&46���	�'���#GܶVJ��gC����B	�'��@�
E�?(�cnUy-�i��'�.Xz�i)�px��X��4 z�'rsfȥO�x ���<X��'14��pŝ\W�M��Όt��=	�'����P�J�_�F̐U �;�N8�
�'|�B-�m�,� �˦^	�4��'�j��wL�n�� �m׻'6`��'$ZMq�Ga�ny�tE�$H$�9�'Ӧl٠��2t)� �bӦd�=��'ڄ�P�
Q+�j � V�
jI��'�>}zW@���%�Z��8��'yPZ1��$aF~U��mͥ����'�Vl02٘�^i�Sɘ;}�2d�
�'�d���IB.�����D�x)��'	P� �n��d�� !ឝ>E��'��X��D��fP3��!;�|,{�'��4��̰�U�El�$ii���':�y���!|]"��+ cBd2�'�v��v��;�*� ��Y����
�'����̯t��]���ŝc�t�r��� �L �H�u�8��ͅ���<�c"O�t�ѥ�WZ�e��N��n!	"O��HC�ڀ�(�Vc_�K�H���"O����H �,o�����'�xI��"O��xB�U?���� ���:���b"O:�֭\�"s2�S¦˭K���kg"OZ��t�	��y3Fѥ��m)p"O�U"$��s�
m:Q�
6�5�t"O��"H�4'��۷j�:m�����"O`5ʰc�z�bQ�ܓtoZ@Y5"O<�E�-/:J!�"0����"O����À�c�X�wK�� �E��"ORxb�m�2r�i+�γZFx�"Ox��'� Dy�h��[{�� 7"O�Dp���+qa��RIɃ�\�"OҤ�F)�Ȓ�b���4pÚ=X�"Ob�)�#P�q߾�;ġ�N�l}�`"Olj���7�a#�@�s�����"ON-�`�	��*q !G3�<��"OT�Iˍ7]��N�^'VD�E"O��+v��[T4�1%cY?f�ʹ�"O�`pg-� ��9�̤\���*e"O,��3ȓ_ȼ�PP��v��Kf"O �B�!-��i"/�%I�nQR4"O�9"d�R�R7R��E�aVzTb�"OB\0�e���`9�d/��,&=�"O~0օ� ~C��a���+�,��V"On�kN�Pg���aBPJ�(|�@"O6�%�x�E��<A͔�1�"O��s�J�6�L�#�I,?�����"O���S��h)(��*B�#��Y��"OVy!��*/&�֣ٚ�;d�\i�"O%���=y}�u�0eS-A�q�"Ot�r �'[6�P�Fj�cO��"O.��G�-d���a��@+D��7"Ov@����Z�����Y�OAhtQ�"O�i��HT3	I�yy��E 4��`d"OpMV+̥U�1�#ѻa�][�"O���gǂ'1<�p�,ϥ]�����"O����Bԣ\�$M�,^��qS�"O:D��c޶$]���'Ć�?x�\�%"O�I� '&%�@�Y�X@�*O��@.U4�����,R�*1��-�S���XX�6d!]d���t���y���3GZmr,R�����؁�y��EN�i���R�F�ѣ�Q�yB��/!�R�Bb�$D*`5�����y�J׬ޔ�(T�HI_P"�	�y�B�-&T1{!.E܊Ex�iƾ�y��3���	ըޢ6x�T���η,D�=E��)���xSo�T_�h���
�G�q�ȓ
dDu �#�k`�4��A�d�fy�ȓ	���*U�e�bḢ_�.�̆ȓ �(q��~�2}0@�u!7fAt�<���,KS:)
'!�,mJ�7�K�<�G�1@��W�FTqq���q�<9�#�B0����C�$qӍ+T��[#��DAa�8,�2IK�/D��:��#����M�@=�Y�Я+}���&�'=�E�e���r�Lǲ�>�ȓ|�����; �����F-dΎ�ȓ
��80��8dq�ٲ� ��4n�x�ȓntH1mЭZaBURr�b��]��oȮ"�*G-��y���c����S�? 
�o�;\eL��W�#G�ܹ�"O�L�T��!=�>����5P�T��"O>��!ˇ�9;^�� M�(c
P�YP"O�rB�٤
J)�!�^��q���f���	�?Y�0��af�b�D���s!򤁉�����Ò*�b��ՈD
l!��MT�ic��̛>��(J$��/k铉hO������(]����Hи1��Z�"O�i'.C�i��sʋ�hp�"O\`J@�	n��A�@��n30�1"O��)�� �-�i�)Q��V"Op�vi�?A1-26�G16��"OB�t/�d�Xp�@CL�U� P�"O��C4��j��LX7��b�XH9""O0|"SC�"v���Ѩ�cG����"O�)Y%គ|\�� ա��8��""OH򃠌9Ot�}#�!��T`��"O*,7B��D� �c�U_{Z@�E"O4��^���r@�Ҷ]0ѩw"O�$Y��r���Q�K�O*:�3�"O칪����W#V��W��#XI�G"O�q1��2{�	:#m��H)���"O�͙�L1s�6=���c����"O�c�Ȥ�(�̲y���kE"O�)��ä<�����X
W��$B2"O�X҂+$s@:ݨ0��&|6��c"OX�;ae�T�@,XS)��3z�� �"O������%#9������.xde��"O��q�
ΗW��I�
��+ô��"O�y����!J��{`)\�_�\�"O��,��.��C��Ը�P��"O��j'���W�6ЛG]+m��p3"OTL��ְb��ȕƐ�'���"O��Q�,��{��J��F-8U"O���E�n���B{Hu��"Ot�'a\(���ĈǆRt�i��"OL᫗������H�S>M�i�"O��+�([�����ǄF�~6:�y�"O�KU�:Z[�u �eZ�m˪1 "O��k����Ly����>Lb���"O"����<YxXS��M�a;�"O�TF8U��x:�
37�΍�a"O����-*>�	�#�y���r�"OFd�@��D�� d��z�v�a5"O�� WB�`�Zh����#�x�"O�lQ.îX[��	"�UvX&MS�"O�5b%B�*D>X8s,� {=�`+"O�ճ�ÁL��x�4��m~Q��"O�\��!��&�uE��q�A҅"O�1���,�.̠�e��|�Z��"O
�k�!VtX����Ѷ+6�pv�>��Ob�=�O6N�àD%����sJY=#ǎ �	�'�l�Q�,�mXqh�o˓����'&D��W�)/❻�,!JQ���'̠�Rk�wF\P�B����Yk�'1��,9W`M1�O�@ 4$`���y�<i҈�-E �y`�G�D',�Y�Dp���0=�Î�*���Y4;�ڹ�E+�C�<)c�5 ��m�f��,ea8!S��C~�<Aw�99v!㥈ީ$H�3CV|�<Q �ƧQ���ٱr�J�b��t�<	Ɖ&H$Ty���C�.�T��c�f�<a��K��E[�-"�#^p1�ȓ}~��c�_��V���+�9��S�? ��YƉ�n��Y�4�~(��"O�=�2�
�>n8
MGpbmi�"OBL�u�в>�� �=����"OB1�s��&�z�X�"O6<�CM�*L| ��Bs�$m"O��fFa�(,1�ǁl�v�j��'��I�F����9���"�Q<��C�I=2<X3-ΨYBݘ��&Zt�C�ɀa� ��:�U��*��z�XC�	�9; fMH�vװ�KC�Ҵ-�HنƓxJ��
V)�]�  �gɋ,Fq��!�2P� B="\�bF ��@�� /6A1����.|Z�r�C��D����ȓ~��݁T���<Ľ�
H�c0����~��Y�ȋ�	��Ptg_$U�}�ȓ*J�3� ��-�p9&�G�`4�ȓW�P��+�Eb��$���;�a�ȓE�k�*�)Dڱ���
:�H��ȓp��,Y�e��qb�*�S�4��KF,Y�KY�0ú(��F5y�,����4�"��R1��赋�^"t��S���0��:8t����. ���ȓ.V���G�;= �(y���U�h��&�l	$��
J�*���<=�,9��9(bH ��ֆ�l� �$
7��<�ȓ[�*C4� �K9���pG4O���ȓb`Bp#eJ�=�R5�%'F37�
Y�?����~A-�|p(�:�n�\�DD�@�B�<��RA� ZA�����FT�<��N�lSD/Z�N�͊�lOM�<A�n�)Y��P�R--88BBJ�0�Of `6C[*Q!�50��Q�A�`T"U"O��� ���F)∡mP�2of�R�"O���A��;�f�2��F�RZf�S""O@m��Cڻ��iiÊɏ4t�B�"O�\��!�:5/m�Rj�Y�)b�"O�,q��˽-88�	�2O����"OH`��o�T0�ڡ׊M*X��"O��J/�5d�y;��o��`�"O����
��Q�Ѭ�1r�$h7"O0ey���xZ�ł#\Ӛ���"O�|�a��c V�)s�" ��q�$"O�<�IW�w�m2���]�$�3!"Oa�4.]1	V,���L==��0F"Ob�Fj��gA !iE��$Cg̼��"O%Á�ìZ,�H�
1G^��5"O,ؑ@�)���JJ�MHљ�"O���㫏
�F$��h�9u�:���"O�LP��
���zPIS����)�"Ov ���ʬv�T0Dh�"4X@=�%"O:m �*W	n,Z�ta��$>�<�2"O�8��[-������%2-y�"O>P�Ǜ0��+�G |d}�7"O�`�dkH$nl�E��(QD,̙;�"OH���dُ]��d
��]�'r~x�"O��)^i��d�$�">������[}�<�e�N9.e1��ۚt�Hi�`�d�<���[�P��l�Ab^�$� AE�<���V98 �u) ���66�cP��@�<A���EAt��@FRSz���X�<��W'!��ٹ��ӋA���!�FZh�<��!R�K��PxhYGu�PQ ��\�<	��R�h�&5��e
�b�2�(�@�<Q���p��0HԠ}�\=���e�<� Nuy�#4���8�4T�.�c"O��0c�.�9�H�'v��t�V"O�)�cj���WJ�Fq<�� "O@�Z�KM�:��0!F�{h�{�"OȘ�'*}��y��HV���"O��Z	X�cfα�c݉���K�"O���O»O���#� �S�40��"O0����6�0�Є��R��\��"OR��"����)Րu�t!�P"O0�V����u�U(�.xahh�"OH���,[�<}�GCbM
�"O��7�6 f��A�H۰[3�hae"O�Yt�q�̥R�&]�+!�asQ"Ot����pT�a`��� j2I�Q"O�����O+ˆ�R���D�
d�U"O�0Q�C����Y��$?FV�J�"O^(7��1>��1���N��)8�"O�}q���;�HJ���i��a"Ofi��a�Ⴕ�t��]gH�d"Oh��'E�r[��"#�6W>Ւ�"O��p�V�\�XA$�\�{GT9��"O�(eۜ���A䗭=V����"O�	�)=8<�5�M9em��ڣ"O~ P5fL;�Ʉ�ݏC��ӧ"OԵ:�I�Zpأ��ɸ�N�R�"O�q��L$D�6`c�ߤ5���xd*O$��کf��0����h �
�'�0��ɁV�ၳ曑\G��+
�'>���"%�6�ͨ��!x4%��'�n��2��e����)�7tʘ���'M���M�v��Qr��L�a�&���'�t� f�9�:x���_%.���:�'UZa¤�X5L`��"�!;����'T���f�X�9
��#_$���'��0��,73��6bB>$i��h�'�J��&�t�>D���
��ԉC�'K"d�ӹbd��C�� ���'�x�+��V�3��H��P}TZ���'��X�K��6��0�
�p0fTS�'�!��nO��'V��fQc�'�E���=[��;TM�vxI�'=l%ۆ�[�=p3�ő>Ԩ
�'4t�6(@�l�Œ7�ȳ)Ǭ�	�'Y��3�G�G.�x��a�(�R�Z	�'W*@�qGQHf0H&*Q�^P=�	�'��tqE(�O�V�2R@�(:��'��)rt�����4G(Uδ��'8��2�ϔz+  �ŀ(��y��'�$��O�n���j�d���*�'�(i��O����˟�B]x
�'K,�S���P\<ps��pP�	�'� ���.סzd�Ҫ�����'�%�'J؀7[>U�RbF��D�:�'�֕��l�$Q;bl͵yu�`��'�,MC��V3FQK�MC9lTl��'�r3� et���!Ye���	�'�.sR�Ω�v�㢫X02��	�'u��% �>1�2��	"~�ɣ	�'�v�kҧ�"2��rhIBE`��	�'9Pű�A˂d��)	��ٕpF�x�'�2	��ޝV�@�8C�$o�$ �'8"5��Ϗ�/ ʒb&n�i�'Z��㒋q�F %��	j�� �'���:�DQ�~��D�B�h<�D���� �Š��T�e�����i�9Ħ ��"Oڱ(Hw�rM��&b٤��"O��P�oAh؛R�03 ���"O8*!Mۍ^� @b�5RP�(�"Oܸp燝�@6-i�nͪZ��U"O�M��T�W(A�.�t�V���"O�P��R�?����mP~q��S"O4�BQ�󀁋��ћ6�\e5"O���̓�yk����(��&�Y�v"O&|ӕ(cjL�`�Ӕn�R�Y�"O6�6O�"����T�RB���p"O�9�&a 	�:�Y�(0f1�a�B"O�`��Ř���-��EZ<{,��5"O�Ize�@��h�D�/jvm�D"O:���n0\K�qx-�����y.-&[���1~S����y�i��)n6���W5q���"�;�yr�H���d�!Id��x��_�y���O����cb��+�`$��8�y"�HX�8�e��Ol�(e���yУ�(9y�/�*A�<z�hI��yM�GR8�TfN�4��bI��y���X�� y���.:�|��'���ybl��~An�0W���]y��>�y� �=0f.�@�P�s�����Ø�y�Ұ��a�J~�$�xFe�ȓ��$B�II�U����p�5z���ȓ4$t�Zf��?����j��qV�����*�x�C�'?+L��Ӯ�q�|��5겵��!�I��|(���C@��ȓ� �ʗ�<�E�׈�x[ d�ȓ�śFk�:^�6�C"n�k�����+j��
�&O:��	ʔJ>\r����-?4e�t��!G�<AXpa�b�Y��c���ӭ;	�ٻ��]2m)�Ȇȓ (�E��7>9(D��fפE�,Ȇ�I��c)�biZwm�=�P��k���'�zY����+�2��ȓ ���v$҂���1+S�tl���ȓi�~�J4b^qD�Y'ğT�`X��]��,����>8��A�cn�"��h�$ �Ԩ�5�ա�NA�[��ȓ1�H�����ٺ��@	o)d9��[���b�E,g�:l2�r}�C�"O>��lЧ1Ύ��J"[`�y�"O�+��]_�2���c�>	�ʣ"O���� �n�Zt��b؈�,��'"O���5�,{$�K�5���"OZ�z�lW�W<<�Bf	�C�����"O,�Vㅶ=�R��C-����"O�DBR� B�����@�R��"O�=a��D	I��1���B�f��"O@��`
� 	�4�L��q�"OBha���DD�U�8��cl¶6�!�č3�e�Ѧ�*��	���۶?B!�1`�whY v-�c���!��K�\4\�#@��D�
E�u	��0!��
Oќ�8�,���phfj��!�$�T�0��&�L�+�l1'�G�!�$L�Jڰ�z Bƙ��8qrE��a�!�dة[�n5 aֿ]^�1k�4�!�DL<�
�Q�Sj00+���<�!�dӥ:�.�صe�+1l�(ڗ��=+c!�d�z�N���_�h]�����A\!�� ��	W��M3�!��!C� � �"Oƽ�Hޘ=4=U��J`�Q"O�}�#��>�& GO�0p�݁w"OH|��b�H^��"���=Q��R"O^i���R�{̈�f�=dN�옓"OpDp���1hd+�E$E��"O�9{�NW��P�&Ϻ�N��C"O�9��`���S��$�X$)�"O�T��M÷x�
		�Μ7V�mz0"O}�&�WD�~���%}I����"O� 9%#�䔔;��wK��T"Oލzgo��dR-�ЇǺzתEˠ"O���+�%Q|���E?<r�$+G"O�H�zɊ�(du����"Otl�R��v�B�y�)�7e,tz�"OVA2.�>_�HL	'+Bi���B"O��Zu��T�̥�ŭI~�{"O,6�Z9Z8�T�Vě����e"O&��VG"�b�s�y����"O�tZ ���$`r��ȥi7"OPi�͒O��;G��&(��"O�u6��s�*�x���&I��D"O�
C�ѐ-��hQ!��)ҬA�"O��s� ?cb�P���7���(G"O���W��:#ڙ
�?�.��"Or9;s�H�`�DCC΍�aqR<S�'u�]�b%M�iF�����$3n^p	�'3 �I�A2(m�ywN��x!���	�'<2h��Ē�D�E+��i4<	�'7
������i�u��N�Q���x�'�f-�&BȞH�tY{�k�J8bi[�'fLE�bH(��P�!��IMR�@	�'ݖ�ȀM�,^��rD�
�L=��' `Y�E�,=�(ڢh���f��'�֭إ���L�����4v�t ��'��ͣ2��H34�j�$ۤA� ��'�TȊ�Nԇ4aB��hª4U0��'u���
\|H�$��=�$1
�'��	�� ˲0���
�X�D���	�'��i��	-���B.͊A+���'8Px�df���a���;�)0�'���i��I%�(YĈD?f����'�� $Ŧ'�n��o�&b���'^���Wj�+V�B 9�*[�$�R��'�d��F�%��l��k�-��b�'Ozy��N�6[�ġ���d����'T���b�v5#2��4�
Q)�',�0%��dhHL�/B�+�X�ʓ`�2�e�=w�l�8�eÓgbZ���3�dM��L�)�p���C ��m�ȓ5��G4"U����e؎VT(܆�},q�$A�.�d��C9����ȓJ��Ug� `*��(�`��$a�ȓ�}(2�LP�Jm8�h�?o`���ȓ[�^M�0
���^�BD�[;l�b��ȓr�(�0^=\�z(�!]s�25�ȓ��1�@�06�U[�6S�b�ȓ�bQ��k��8T~��a���s�<Y�ȓu�����1tV�*�,�0i�M�ȓb���̌�0��ibDI��}>܇�#����l�6N>H��%d�!n��ɇȓ)O��	��BN��&*�y�Iw�<�$O��Y��X�}KH(��� s�<Y�F�^���A��@rpx��Tk�<� �@D�( �T� ��U�)�|��"OTuiC9]j.����D�(��"O����'L?W��e��Ţcƨ�Q�"O���fj�k�d`J�txڇ"O"A�E�����Cbm(@jt"Oz�[C
N�i&�12�/���A+3"OF�DIفS�&��POW��)�"O0��%L ��\�g�EP�0]�q"O�eY�p,��,�$]��i���yR�Џ.,b�y7��Q��-�%��yb�K�j��I���U�7F �Z�AJ�y"cd��O'(�T+b-H��y��ƥ?�lи���o��;���yB��tޱʅ�ٲ3F1���܂�y�hE?�2<CU� -G�){�hS �y".��2�y�aG�)R` p�&ʝ�y�A�#"y�h��'I"�����ƛ"�y�cS=�n���#K)�ѳ�F��yB�R$B��M� -��!�*�p)F��y�	)?�E��W25��@�yb '�V}Q�׵\��-4%�y�*�1=\T�r��4Wqz4�Cފ�y���E���)FI�x���!�y��\�0��P�b��G0Te�$(�y����R�D��I�$E�b�#D�Ӑ�y"dQ�:6��H:AO��Ԍ�:�y����|���Hό9��I*�L�yՃs�� � I�8�8LZ�@C��ybe�5O����p��&3VD+�@R��Py���~�D�CB��S)|�:$��[�<ٱ�C�.��My���Y��C�KV�<)�l٥$YtH:�����s��U�<Y��Д/Π�&	�1tZaH�`�G�<�wJȡ�0��0��98�`E���B�<q��m�H�8�F7��8�׋NE�<�1��?=�^���a_�
~^ &�J@�<!�o_c*��ˆE\�ib�U��a�<���

�(��<��Qr�O�]�<	�@������Y?�4T�w��\�<qW�O�r��!��g0t��#�N�<�F�,)\a� 刷
�tPkǭLU�<!BL� )��#�[1<�5���k�<�!њ�B��(�`M�� }�<�W�T>B��2��4+��u[���UTar���ef��v(ؚZ���ȓM����B!�y�3���W�(�ȓP����@�.�b@@1&��A��`�:���͎�! ��E͚,� a��a0l͓��|��1�Oȳb	�ȓ|�^~�d! �B�3?����X����Rk�X1�aM�}_����wo�e���0��i��lh��d�ȓx����a��j�-��٭���2�"!6fF�~�t�3n�=
J�Ņ�S�X �%�+��=�.��15��ȓD�̝x�)�;@�hk��F�h��<�ȓ/7f�� _�|�Z	���K{����p�a���W�~x��̔���d�ȓ	i��%�
�P�L�H#^%	�V��ȓ~var���2k��1�V�ybH4��J�@ȳġF�6��]׀	,�Q����G�� f����L���84���*D�ة����,H
�� �8�,p��!)D�옇�ɝm4`�.Q8��%Q�9D�� vD a(Q�`��@;��Ȓsެ:B"Ob!2)bY��f�6]qJdr�"O��u�F"=��}!�/͕Nz0#"O�d���^Q��̔g��"O4P�&H�,�$��D .��"O4\�%��c�D��h�:^�`�C"O�����˦u����>K�~�H�"O��
t�� 6a>�b�R:�x\0�"OxIZ��f툣�� ��a�"O�Iq�Es� =�EQ��%�"O�uS�ϟ�2�!4 ڗh��e۰"O��E���Q5����o^��3"O�p�C�0T����N<3P:t��"O�iF��S�rY�#P�A:��@"O|�p$'�* ��"��J�"O�iӣH�8f�ܸ�뎌U��H�"O�0�s�- �H���ɏ.8?��a"O��a _:*�61#�uG�J%"On-��T?H��k��Q8$֨�ф"OָP�Ĉƀc�Ԕ,��Y�e"O<��(4���"��F����D"O2Mr��U's����V�V�9��+r"O�TҧM�61\���ա*-p���"O��t(\�� ࢮ�A�Z��"O�y{@���Q؀�)�m�3T�����"O�+��F;P@D�!l�xt~��"OR\@�A�#$a�pJ#/HB���"O�٣���,*�٪��Q(����"O�2� [�2�0���C��TPQ	"O<x�P���t����nMXL�r"ON:s�ͫ��H�F/L���"OT�п!F������2�\��V"Ojx�pO��$�yӂ��dq �"O���I�9=J�u��͖)EE9�"O
t��	�/ˤ��U�9<vCe"O@�����v[�Y��� t	�"O2(��Ŝ1|�=�'^� �*��"O�����&|Ej-`B��
E�"O�Єc� ����e׉ꀌ�"O|����o�\��C�)�����"O�aB��~�����B̾	���"OP�"�cۆX��Tk��S$,��͂�"O��#��;k���8��:;�B�Yr"O�l�D)�%�� ����Br<�Ɇ"O�S�ɛk2��e�K�kp�k�"O��W�>h1��X�B�H
~���"Of i�>�6��&o�,-奈J�"Oʘ+�n��G0A��K'M�*H��"O8<b5��"WB��umZ�`���"O�}C�:zUJ��6��; ��0"On�`�'>e1���X9K���)"Oh����5D��Hi���A}�d��"O��� ]���P���wF>�a�"O@ŀ֮L5�l��tf�G2�`K�"O쳅⚞c�] B�ֶW�� "O���#�'gQ0�+�3{�ԝR�"Ol]���FS�	7eW�^<4pA"Oa�I�)c �D#�ʸ5�R"O�PQ2��]8��H�����01v"O���D�>o�p��e��1�"OT��`m�j"DԳ�mφ
� ���"O�j#H��G�:IɁ͓�sB��4"O��g�Y	xCZ���ar|�J�"O�9��MZ�J�]°{a$8!�"O� �D�$�<L�A�G�U_�k%"O�!�6#~hܢ`.�3\[�"O�L��׶:fԣ�MK���� 2"O6��d�Y�H��$̓!d�Ԉ�"O��PC
�i8V��!l_:E8�@��"O21�"�_@�sk
{Q��ye"O$ec��2�.��D N�Ȁз"O�	�LSq29��E�j�
��&"O��šY'��p�v�_(D���:S"O`=��V�g�·��P,u �"O:Y�bf��~�Ԁ����%�б��"O	�u�9�6�1��F�+{^��"O�up"�'mnHbw�3�n�[�"O$uZ`G3�J@F��y{���"O"ypn���@@�<vG���R"O䔐r��)'G<5[V%�>9
�-�"O.����f�L��d�2@	��"OvH�Ï܂,�����Q�@�K"O��+t���,� 4��C��S%"O���4s�mif��yu�qp"O8	:��X:>6
qV�E4fD�`�'"OF$)�§c�Nd�5Ȳn4]:c"O�8�P�R��]��B��	T�@U��Jd���N�&w"�A�Y9pg���ȓ_bHs6�Pr�9З埞�ȓn'��`�'4|f�}#�N	wT�ԄȓI80}�w�U;$D�S��ӚB�j�ȓ%����ቂG��,���ʕ�~��ȓ�P%Hu�Q�Fib��ُ{o\���M��PR2J�"BJ��D���!����	�AT�� GM��#�z ���4t0�1��3j���K�I�=xt�$�ȓg����PG%d+�7 A�!���<y�
��Hl�%A���y��ȓF|X��(�
�؜�!�M�4����<�>i�O�G��� ����P��x���E|rhs3����(��u/�0�4g2�,�چ
�*�Ԇ�Ha�Ѩ���_3�Ȃ���.I�l�ȓ=�&q����p���IT��=	i�ȓBݢ�⮄w�j�qD�ī+�a�ȓ���±��{������(mb칇� ��Tz$B�>tG�<k��ݦ
bL��*n��r��Q�
��k��"D&��YvR�"��Q5zj���qM�7g���ȓ�qI�'�U��S�B?+ �9��m�� .\.�0���Z�4�0��@���{gM,2U���� ���0��	@�TC�!�0�?P���ȓK�0�S�ԧ^��E����:Xr�مȓ'�����CYF����f�!.���ȓn�pѡ��3|@S���;�Q��k �DR��]4PJ!3�_,�ņȓn������D�rf���^�0���ȓ[MzX�C�0�ba!�I��G/�5����C����K�@O�dq�ȓ`)F�{2(	-Ŋe#q#�|;|�ȓxQRbh�7�t���L%~:�م�S���H�aqRFQpQBȣRV�ȓ �6��CC���&AB�&S2Ȇ�*j 8�����hS�	�2~K���>�q��S[H|��
�,jA�ȓ{]����ۛXRl��>Tژ�ȓ"ؾ����4��]( bI�B}v���S�? V�Q���04�9�@�Ʉ(��xc�"O�8�tiAn�I�!������"O=� �T G�2��4�w��R"O�y��żR��#�M���Xڧ"Op ���T9���;��iJ�"O���3�F!�V��rP�>�R<c`"O~q0�ȫ_�L-0�c�2�̉�7"O�$���[)�1ң	��9AД��"O`���ȏ6l-���ǞJ6&)!A"O����%z�`hU�^9,�I@"OT��m�� \᫥$V�	A�`�"O4�C�����, S"S:|P��"O�5������B%�A��"O.ś��3�bi�q��4l���"O���(Q�=:� )�@N^���x�"Of��0kشE���Oè	�8�"O.����I'��æN��ma�"O	��e���d�H9�l���"OfT gd
E���� ��-��(�$"O������̨�J�h���Zr"O
�{�a��d\�c��$qҭ�F"O������3(�M!�ݜ8	���"O<��ӎБa�BQn͒r��Z"O^]�W�P�ـ�U{�� �"O8,��e?;u��s#̈e0�z"O��صT �Z��<)p9P6"O��ѵ,�5\
r58�Ü�&�r��"O�Y�X�[u��@Dż� �"O�u�ũ§/�����6}  "OL|
�M�hALY��ڀ#!t܋&"O����J� )���� 4E�xy�"O�Mb���'h��%�DA�夵K�"O\��W&�����g  +ܘ11t"O:8H%��09��i$��V�px�w"O�T)R��1^��M��N�3�lAr�"O��s�K�L~(���%�S"O�,xa�K�&��t���S��d�x6"O������,C��]&֘/��͹%"O$u�f��,����EP��vm*�"OX�q�lS�D�إ�҆D���8�"O*�Q��H�d����r�ٺ1�Α�D"O�i8�!F�%숙�v�A�����"O��WD�{��d� R}`h*�"Od�:C.F�H?4q�2�@�'Flcs"O���QHE=;�=0T.��)9ڑ�"O*0���
1�Va`��L��-b�"O6��U�58b�)�԰{b����"O�=���Cjtp�6p5�M�"On����*Y��q�`�ӵd4P��0"O��p��ޭB���.SF�"O��"��
���g�� 3Y� "O0]�D	�*N��ӷ�X�4+ڤ��"O�q�V,F5TH��w�.��7"OzA�fZeKn@ӕk��V�zhKs"O�-Á-C�aqJ�
sax�=p"O��R���t����% �a3w"OP!��!�h:�oZ	�Zx�"Od����'9~,@$���ֲ��3"O]�Q��>C����\5O�V�2�"Ot��'�Ѣ �X�����-�t<9�"O�Eʐ��7|A
"�9����p"O�Y)��V�|����Y[}��qT"O@)��^76	��+�*|��"O|�b��*.I���*��g�<�"�"O� |ܹ�J�2� \!a�m�	�"O��� ˳A�؜�b�I�)�܉!%"O�Q��D� ���P�P81�$D"OL��S&RoB� �B��|Ic�"O��򖄈<�P��5K�Gv��8�"O�ad��E̐����;.l Ii�"O����O�-eꤰ��
B���!�"O���$L�"cԈca��� ���"ON-(���9^n�E���>�(L��"OXmyP�4�t�3��8�=c�"O]a���V�(�i��a�)��"O)Y����O���KB�
s����"O��CFܤ�n�XU� P��&"O:uK�lT�I��8�bHH�$(D"Op�DhL�Y:d��H�t�F�R�"O��B�+_�9��T�s��[��ܰ3"O��	 $�rLdm>�()�"O,%X��[9� �00˒'���)�"O�tg� 6�	G�3?`в@"O�|��b��s~�� �
�w,�q"O�<�5���:BΤ�T�Q#*���"Oڄç=�X6���A��W�<!��W���D����P�)gH�h�<�͘bx�I��o�=�(���_h�<aӨX%^�*UI��V3o�P;�Fz�<Id��	���ӡ�	 ��E+J]�<QjѹbufTYa��T�C��	�<A�G�C��� k'��U�c�<qG�������j��R��Vb�<�dΛ�0��$��C^r�99���i�<�F�0��Y�pCJn�bM1#��M�<	GS7���3#Z�P���m�G�<�vDK�m�FE�ƭ�;�>x�j�G�<Rl	�9��J��ɸbz}h�	n�<qe�1S��؀G���R�ʱ"DoCk�<�ι<¦��`Z�
����5�O�<A�dܢ6�PU	�j�d���r�J�<Q$�|u��qL�I�|�S+S~�<)��G&����Q(j̽{��Rb�<ǌU�uGz�ghc�DdS�Du�<�.	=:���	� N��C��Up�<��@�)�0`@�'V#S����[e�<�]7lGF��Ī�t�[ �Ye�<Q�L	�:���8hM6qj�@a�<IU"�(.tH����%����FX�<��޹}Jz���ň����#�T�<�(�$Z]l�q�l��z����,�e�<񣤛;nւ�Cd��"<���EI�<!�A�s4��r�&�6�%x&  F�<ѵ�73��"F�P�<��S�J@�<�2���J� �k�ʦb+�,t+c�<qv�0^���%��B�(h2 KF�<y�&�X�`���a�-Fqb 
V(KK�<YяX�`��-�(A���b K�<�1��E�����/$צy��/B�<�v(�3La��+�+)�P���@�<�%�J7x�8p��=C��8)Jz�<yA�_$d�9����tS�]�C��u�<���"X�h�H�5}�8�pr�UH�<���:KO���+T�i�x� b]�<���mLҢJ�,IzZ�@���Z�<�2�n���a�V���QS�<����C�2K*f-(7E�K�<Ip�ܼg,��r�I�� �x��B�)� b�aӎ\xTR9�0��=�m�"O���a	�9@Ё��j�)Ӽt"OD��#M�4֚��樜�V��"Od�u�w��:�g��.��U1a"O ��W�B^!��!�����"O�P�W��65�p�X�o�="��=�U"Of�9r�P�z7l;�k�%*�x p�"O��a��D<uhT��I�l22`T"Od �o0m��0�!K�T��2"OD��p�n�y' � V�����"O���&��^l��,ZhIK�"O��$�ۊ:g��aC��Mz&"O�1k�X9����B]�[��yD"Op���F�C������Fg�n���"O��@U�V�b▩Jv��,�ƍa"O�D��N��� "���*��i[f"O@3�O6�N���C8l�,��"Oj�UOU�Y�Ĵ0�펏d�P"O8��3��P�(K���z��q"OT�c�>at��b@� ֨�R�"O�8�!E~���N<��Q��"O�MS�l$�<�
@'V��Qˣ"OP���MV�w����V&4���s"O�U��b��8;�ظ!��1�"O����'�W~��H�$Qpr�8�"O�%����wt���!��b a��"O�U�(V�� \��ҏ/��b"OPU�@"Ջ*^�a1r�8tn8a�"Ox�AK��U��A�,Ra ԉ�"O�X�E�ŋ+N.a+R�D5D��"OJT�6�X�;�Z�sKO�R0Tx�%"O�����	y��P���,.j��c"O���޵D�~�ą��wʠ�F"O�l��/t^���DNY���"O�ВE�Ќ#wFx�2bԾ%3j�g�<�R�!x��� F��W���<�1LB�R@h��)]�ua���a�y�<A�m�?�h�j��8X���j�<q5����䩤�O�:ʑ��Hj�<��f�PP�S4H�R�93f�5T��B ߸^kVX��$�#0>J�Q�*/D��R�m��/�r�:H̑n�*�V#/D���q`7B�`�l(�I'I8D�xa��Z%H���b�.2]�T���2D���s�!*�:�3��N�9�i� 0D���a@̺*�z%�6fI!&l�5Cqk0D��:'A#.����A/w�ZQ1�O+D�Hb�lN* 7(�����L�J�)D��+�I��m�qB�j>6��c�&D��锋@�*w����&s�4-9q�*D�<�$9�  GD�Bl��Qt�,D�؈�	P�V�����N֎
��y�6�?D���F��4qpU�5��ۘ�#0�#D��q�)��<�����N1��{b=D�H��c�in����΢�\���L:D��afgyx^� ��G9X�9��%D�a���"Sqz9�BȘ3#0I�P�.D�� C�[9
6\8#g�&�M�e�!D������?<t!k���L �$���3D�h�%H�'�]#1��f0Ĥ��0D�#�+��&l��P�KZ'ؕ�C��y� �k���n�^&�k�d��y�גq��Q��M2F޼�����8�y�$��yoĠ1P���K�h�!�� ��:"aK�hU|��$�@h��Ř�"OD�G6sD��B�;a�~ !�"O�Ha�D�=�bI�3"Æ �D�"Ox���dY$@B�!�@ţ��͈3"OP2"�r��وХF*ͼ(�T"O�4�f��ir�S7H!D�:�A�"Oȱ0�c�����o�������y2�D�R������X�:����yB���#���-A�b��yD:Rf�'�|���H+�y�KE��ܴ�L�9m`������y"DM�Nd�̀�Z-6T\[*���y�����)�M�*oY�P��y��Ң��E�q�%�1B	��y�C�"�ѡ�/�<EʑEJ%�yb�8:q*����$iM�Q�٭�y���,Y �;�J%P3��a��(�y��/i��Y��<Cf>�a	���yb\�0mH���cU�4�22 �δ�y�䆝J��aAe�6.�
�`�F�'�y�c��f��s���)ʽ��K�y�c��s�hv/Z�X���v�I$�yM�n�܅Q�F�\��Ժ6�&�yBlX4P���� ؚiA�A�y2b�4)���P(��	��,�c��y���#+�8؂͆� ��A�B���y��3m� 	ۃ��|�a�	��y�HG�bBES�!M�r�ĘaA׆�y�U�5[��i@}� BQ��yrE�Xh�92�J[�c�\� j��y���)��L���4E�4!{%V6�yr�ô/v��`cG�j傉�Q�B��yR�դ}���Ǐ.�����a��y�+�3�=�R��8(�6�� �y'�"{A�p�O8(Ҟ�h�㝞�ybD��f�����D�H�~��e~8��-N�ۄP����5cY�S��ȓ�(����I�d@�3���>���"����bI�M%ҭ��~��ȓ.P3Á��~�h�#fK�P\2}��(ָ�DH���ċb�̀�xP�ȓm}0����\<�܁#�:C ��ȓ/�|-���>}��y��<[�I��4V�q���7-�*�����R�Z<�ȓ]��(�3�ȧ:2�T9�$-e�h�ȓ]�`�I^��e�'�J'���Z�,�FĈ2r��@�.LV@��ȓ"� qPhQ;�-	�AG������<i�s�G�!�@�,�$>�,�� Vx�3�y�$8F��/�x�ȓ!���PG	g�h�艘hTd0��$Zn3e�U~�޵����V�z@�ʓ!�n0y'C]4��K�o�%�B䉺qV�D�Ç-��X��[ <�.C�I�uv( p��t:J�X��ڇJ�$C�	>s�F@�s�]�RIB��UN�glVB���8��e-Y� �\&�C�.~��� �ۑ$� b26%<�B䉶��Ac|.��T�UL7C�	),� X��0_p�-���#+�C�ɓO�2�(� b�Ѓ��#m�C�	�=�� (e��-($A��@�Vf�B�	�`b�q���Q{���0k�C�B�I��b�¡	�	q�%��;AdB�)� �ը�G��F�P��a�p(���v"O*���X�PG�E`�S.ol$�؀"O��S6�?@'�H3cꆲ?W����"O�+ǃ�'�x´��.OV�Y��"O�y{`��;��#Ɵ?h�¥I`"O
��n�-�1j$$/�����"Ot����P.O��iKd���Z�Z�"OȈ�'쑽 ��M���9�nu��"Ȏ* ��+hJ���&=�zv"O���u�T��eB��\��Q��"O��AŊ�4@������.��"O�m����r�u�@� �`�dR"O�x��a[�+�:{WnL�#@��"�"Ol��֛rFL��s-
�G,���"O�q�i��>+�K9	 b�"O4��������w��gV�u"O�q{`��MA��a"��h��=��"O�U�t��9РL���G�X�Jk�"Op��1�/Jŉ#�W�8�ڌs"O�Es�	T'3tZ%����4A�,�� "O��A��+o�^x@ԫ���z!�"O,�Q�EZ�N��ɪr(�Lu����"O�5�A�Ԛg_����[U�)E"O��1,�,H�N1H��G�hAm[e"Of9�g��4/�;��=�!�E"O��Q�B{��hbk�{)�d9�"OV��H�I����A�)��1�"OV1���E jaȵ�˘x-�X�t"O��P�"A���m=|�f�kB"O��"�(��~,�i���vTE��"O8�	EEޙsdR�J��F�|���"Ot��WD�V{������n���S!"O���o4~7�	���pMI�"O����"ST:TQ�$��ȩ�"Ox�;f�ߕz����͈�`,t"Of4Yj�?-�����FFR<��"O|��E��C^�Y{��->@�e"O�i!e#X	�f��g-( p��"OP5�W!ӽvՂq��ƍ
bAZ�"O�\	�@3X���R�^�J��"OJ����U	+ΠJӄ	�>G�!�4"O�ܒG؎C��1Qv��-�6���"O�<�mӀ��%R�&b��`Z"O�ku�<%����'r�~ig"O2�ȡ#R��)#ٻ5�z1h�"Ol��K	8��A�"���J�"Oh�s%)�r*N�)eh��Q���"O�!�H��sќ�p�n�� ce"O:�Qn

I$VM%���"O�����K$��+AΑ�U֚+u"O�i����%A�X� �텤O^�q�"O �1㛥6�,8�/���*"OV8��Ê�<�n����i��A"O��Z�O�H����E�Z�,sq"O4Ā!�\�M�����&�����q"O�,q��c���kĒk���ɒ"O��r��=z}z@H`�S7f.���"O��sۦ#8���d�`�LM��"O<,*`k�u(A�Ƥ���Ӗ"O�)q���>L����G�m�Ȩ�g"O`raCQ��GNZ��RD"O��K�"=�diXd��+i�0�)�"O0hQGɘ�1c�	��op�8#2"O+&�ѹt�Xm���=�8��"O� 2��=_8`�s��y �}aA"O2e��l���A�G��'=����"O 	iu(�r�lZ$�&$����"O�|����: N1���R �م"O�\j��U:I3RU�˔V`<p�"O29{k"��Lh`�ϖx ���"O��Qg|���
R�M�+Q����"O*͉!��5;(�U���%hLV��$"O���U��6tuL�УE��{�2�"O�)�+PE
L�x���M���U"O4i�E+H���#D�JkV��G"O��ɔ7^���r$�&r�pr�"O��� 쟓Ut�@�RF	R�LY �"O0�R��\+ P<)�.�/�>���"O@٘�	�yzJ�xd��R���s�"O
�@F(P��� �!�F�Aа�"O`|��q�r8AR�D�t���'"On�(��4y6�9e�
-��ڇ"O��ZS��(���c����y�"O�\��R=/���M�yjd@��"O@$�tN#O��Pp*���ȅ�G"O�]��
��l5����XEF�:�"O��)����>C��`
�xD�ɪ�'8}���5|ؠSm �����'u��Q��D
5�4Y�#��dD�'�0İgO�}�&<YZ(�l�0
�'Q�|paA�({�~PR�Ɋ8�"�	�'_Ԡб��l��a!���?T1����']lh資C�|5@����#da^]A
�'z�gI8oB�����%0o20:�'�Zͻ �P
�������6ya
�'��m��.�@�2��ԉ̺�Љ�	�'$v���W�x�҅���j�PUA	�'������B1��ՆHn2�	�'U�y�a*�R�q���'Zx�	�'PP�be`Y�j����4 6r]`�'v�X���
$�R���˯���s�'����������$-���̊	�'�����؇i��]���M>��k	�'pt��΃?Y�HqU�W�3�4���'
^���k�?B�B�I���'-K@�8�'C�qB��/m̫�R�*�Vi��'v�P%aK tPs����X��'󪍉e$ؐ����ߡ�j��'4�=s�ۺPk��B"��0v\�h��'W4���ׇWN�H���g� ���'�z�ɤ�ĳ~�Bܢ��J
7�,�"�'�6��B�Ku�z�ڃDҪ.�:��'; ]�Aa��d�0҃C��*�zh��'5N1a1H��3Z�BS�I%l|}��'����ɹ$�%B���N~��s�'3��ceL�o�l��b._A��B�'��hF)S)�؈����	(��99�'+ h�4#�����L
���'K��b��Ѵ4g.��!� :��x��'l��S�� ��=Q�[�̂�x�'F���!�Â<F�4�%=���{�'��TBg�G2*"h�{"k�3 ��
�'���a
Diy6��bK��)�M�
�'���рD)����N6N�q�
�'Er�A��2o��$(�lO'PhB�'��Q�%���Y�.�1O���
�'B(�a�
V<lN�#�g+:�>�!
�'X�[ �B]%z(�v)+�T�	��� ��#!��^��Hb&8Ơ�0"O:�
Q�Y k1�����,|0t��"O��О~��`QK�7i!�1�"O���SKa����I֥q��S5"O�:���6�^����Ū|�4�c"O`�b�)�5��1 ���H�"Of@у*Bd �(��%Q@"O2���,�A�j,q����s� �
R"O2�Ȃ,����W6'���� "O���#R&@)p][r�^�Z��(9g"OZ�" �S~j`�S�����"Or�ء�@O�$*1L�< �.�[�"O��胮Ҝ<)���U+������"Of-ju ~՘lyC�ڧ}�XA�"Of�j��F*DB�=Ȗψ�H���"O��Zf%.O��i�&�F2d�X�3�"O�Q'�ę(J���� ��Ȱ5"O�x���V�X|�eGCd`d"Of��l1Ks\��B*Kf��@"OF��+T8KH򙚧���AO*��"Oz���ޭP��Pƅ�9�P豷"OF9��F
�>� A@������"Ofؚ��"b����������As"O���6�BD�I����+#.�"OxxE֕c`��K&�B�G4���"O�d���ѩi�MP����z�PK�"Oz)TJΊ{���B%ftP�1"OTH�1F�UM�E+b-wa~�a�"O؈��S�5l�hFꂋpM1��"O�xRT�K�oc�0(#$�6f$��"OD��s ��$G��͍'*^&�A"O��rC3W�)r��'K>Vl�"O�H!�L���{�Mz3D���"O���B�g\���`�Ƌ)).9Cq"Ox�F�O�|�����_!@-��"O�Lᓅ��~X�k�5|A�#"OZ{1C�Ғ1�
)K�~0c"OB<: �D�N=�/،��"O�0+��͢z� �-:n��(q"O��h��C
~�^�I���r� ��C"O���CD̯�D{go��L��$bf"O�В�φ30�H3� ��e�V���"O�i#S:m[&�[�����"O�є�_K��R!LW��p�h "OV6K@�t��Ɩ�E7�H�l<D��;�n�}�R�ڲoR�DM�H#��/D�Di0B�온�nd☰r�/D�P� '
��W=g���&�O��y� �	{7���5�%8<ZY��KΥ�y �>5In��A.��c��I��͋�y��Ư
&䠢�H�c ��H���y�E�E��ئ�S1,:�����y���juJ�� Y0#���t�(�y�,D�U�4�q���j�,����2�yR	�p)H�Ԡ9\��CM��y҈K�Z��ea5>����B7�y�"�=lN�苷'�>LvqgBP���'!v��뉏k
ݙ@��38��X2�יX��C�	�X�4�a�J(Ё٣�!^��C��<>�1�&��4������{X7--�S��M�ՉL� �:ԅ�|�pY#BJ�d�<��@�cO���Bl�)�T����x�<Ѳl7V���OH-E��"��EK�<	&g
��Q�G��a��#�K�<� fl별��t�! (B"�ڼ� "O���$�/���%�T��O`��@�Q2��V�N�vMнB�kʨ6�!�Ċ�`�"�&R�0��Z��ǫ9K!��i����$rȘ��+i?!�d�64��]H��K38���n�Q)a|b�|b&C�3�ĒTn��wj2XS�[��y��IIJ�(�̘EƲt�l	ٰ<�򤐃_�H#��^Rv�PO>�!�H�}�`u[W�/�>��`�}!��H�WQ��b��u�p��ϑ�Q�!��Lq��J_8U�V�)��V�!�D����pYpDP�v���-Y��!���X �A���l 	��m���O^��D�cʾ���M0���J�~G�x��I���=�!lÇ&�v�����G��B�	�i��Y#�Z�}���R��q3�b�T�'ў�Ӽ0�e��aD�~I�e�3�����B�ɡ_{|��]&<�Yj#�M�fB�	#��apt�[';)�)
`J� �N��hOQ>���(L}�!y��!"j6�Hn/D��1C��W�H�{��A�n}D*S(+D�X���XJ���&�=z�"��E�.D��Qv�6T]��rI	]8��	��G{��邟I&ڸ�C��:ih�:#`ƶD]!��+<�M�FDۈXTZ)�5��zI�'�ўb?�+t���N3�d��oI&k\�cP�;D���.G�qC@�� ������c8D�����]�7E4(ؐ�_��|����6D�����[D��|���\�g{T���*8D�Lp �O%.&�/�YT$"`�w�l���S��M�'�P �� q���MjP@t��o�<�Eb��~Y����4^����'T��+�n
l���b�#����2D���A��Ѣ E�)B��`��H�3���
O�8GΔ��zLh��6k�aCV"O�9!P`��3(�<��"ٽPN�=�B"O���S�G/⺜���r���@"O���
1�8���|��1@�'J�dO�Ò���>~n:�B�^*���&�O� 4k�+s�$u��]�u����ژ'�A
A�����c$ǘ�ICʹ��'���Jf��M,���$�
��p�'��II�	Z�O��+���v�:Q���.81�=��'c>p"�k�4�D�Y����y��'�lH�L>�i>˓;��i�>2}�Tc_�ELІ�H��Y�˂�7������^�o��Fxb�'�V��e�=i�<�isO���њ��d�>�-O�b>��p��%{p�Lz�̊9\�6c���xb-RG��Ǧ�(p�Y0`e�"��DRG�'�6���,�G�Uab�	Q���q�,D�lp�d��m�~�R������)�ɕ?Q���(���Сh�fD� ,͢|l(\zs"O<���4�Lez��C����"O�����	\tѱ�
" ��E@"OVi�
A~� ���*!� "O|!�v�	%����oL2[7�Ic�"O�@jb"�1gvXh��/s}�tb�H�<y­��̍��)�3p�< C�����4�S�Os:����u ���� CUT�`	�'k��y�4C���'� 1z��[	�'r�QyoZA����B1vcb��(O~�=E�#40���Q�M=S�>�[�
��yR+P�;���A!]$� k�(��y
� ��jD-y���d(yR~���O��$Ml�L�Pt�ʹ?Ld$
4ID� M��xF�Ģ�P�D�x�aK*jjIkA,��y2�'6����9,�$����y�hF)4 �%�H,Jl��⒃A��yR ��aİr��B�o����r	��y��R'lp� 	�A�<}�bT)�%�1�y���T�3�*�))��(�1�=�y¬��g��L1en�1'�8��V��hO���/L,�HT�tH2�F�!#�!�Úe_TU��@�/8<Ւw-Y>c�!�d�p�h��ӣS�5Z�&���!��W�n8�i�b)����R��*^�!򄉣+(`��N'5�e��G�2��$1}�H����av��	��G@l5�E(�/J��xb�	�!V��1Q��?p�r�h�MX���	P��h�亴�S �s��_�\dq�"OJ� 2�K�S���2�%N�r+�^��G{��i�&�f�"Ѳj䐩�GF'x!�'JT����Ƙ�1��P�!���x��9�.E�r�H��af�~�X�$�7!<|hnA�I��K}n|� �+D�k�eO0T^*� шW�ZtAc(D�<b�G֒3�< ��֥.���Ц�1LO��,[b*�OXi�"��:J0D.��(�SܧZ�%�
ѷ]Fxۂ�eS|I�K<��O�ϸ'���@�d�=ID4p��������2�<<OX��=fh�0W
�5H���"O��D��d�8ȢQ�8204��"O�]��H d��UP�ǝQv^���>���1§2�mZD�"  �c�ۗ#ތ4�ȓx���y��,��-� �{��}��dF��k��ϥZ�$y�	��?J��F{��>��|���Y�=�`�rS
	OʈqT,
p�<�IE�2ֈ�D*@�1a0l������T?�Gy�*��}�v��U	,G�i��#ԏ�y�&X�r�4�����z��Ac���'��{��Epoڭ6�U*m�li��з���hO���=���	myh��@�]ąS�"O�Z	N*{���!-mO�x�D"O6��"��I�}�`�#lH�h�:4�����b\v0zGf���P��:D�8��S`TYґC]�u���8�&-D��J&,�&��8����	PK��P g)�'�O��`R���|w䙫��ގt�H:�"O�a(���HP�x!n��og�ݹ"O��Q�+Z��pLӪ.8�^�zW"O�ѷ��n#���!�xþy"�6D��W���E�G�:y�I�B$5O��=�'��T����1�	�.���z�l�P�<��ƒN��;T+�� 0�dS̓�y"���٦ �V��p$��L������G��'�ў�>��@�ԭ;0�UJ �j����e8��|���On
��s�7=6�����A����yR�)�eC�Qjv팕^��ɹ#r��y�ȓzֲēb/� âU�PN��@�ȓ*@`��/5'[Ґ�v,�1	�X��R
�C��=Hr6�r�H$�H��\�%����c���AQ,Twx8<��*��C���X?X����X@�但ȓ@n��� B�$�Jr��V�>z����v��(���՗D;LE�āe$j���St�io� *��ra�/+��'�F�Ge�'\?�a#G�t�x���� �@�� x���$��j�d�0�"O I(1���Q�a�	��L�r"Ob��d�=D�:ģGaL�7����G"O���!��C�-Ebh�P"O~%�!�@2����FFe�Ҩr"O6hQ��M�'=Lđ"&�4p��EY�"O��G۾\b��ˁ����Z�"Ove�T/��
.Z)h Hα"�vP��"O����%fݬȩDm'	ج]pe"O�0�`����$����d"O|Y�wA\"�Ա��@�X\� "OzA�a+G6Q��Mr�ڞb�nIr"O��`�H5��f�C�|!�"OF���F�f�J�G��'aG\��"O���O�6��Y	�,N�Zh��"O�|�$�Ɂ6[��d
O�Y��hpg"O��ac��"������c.���"ONL��.�;#r����Q�P> �e"O�aZ�/F�.��G�;Z�7"OPiB��'!�<�Gg�|p�}�"OUq�JP����G�PV`��5"O�S��Ln���F�4H
i�D"O�$�6��wP�q$��7aȼa"O��#b_��Y"E�@��@+!"O���J] M����-�5*��0H'"O�����>�0�to�j�`��"O����C݈f�,�s̓?]��%)&"OT�� �)�a'JH#u��{a>O0 �� �5v��*L?�Jɐ��	�4�V8Bb�;l���B��^LB�� ���2�<d,D�e/�
nhC��&���;
E�,����(
�-�C��%���R�ͦ�f9S�	�Y}bC䉀[�"8{�Ɗ�$h�csқ\Z(B�	3<�R-�#��3h6y���D	:B�ɍGd);�ź�%�
�)ੳT"OK����,H�(���+�(�A"O85�T�Ǔ6�4�aBJ����"OB5���p0nd�j��`p"OE����B�i`�,F]J��'"O���`��x��k��)
ji�A"O ��#'��4n��P	E�q��2g"O�0��aسkM2SAHW�[�,��"O�[��ȱb�D�	Q遚9�X�v"O 	j��|}�T���Yv�|"O4�
�T�@��cBCR�i�"O�	�pF����!x�/мH�H|�V"OZ)؁j�_���˳��}ӂ�
�"O@��U*��<X��߈��T7"O��yS �M `Z�EK�N�Ĺx�"O~���ȀE�h�aV�J�npM�"Op�@	��x�՛��Nc�J�X�"OFq#��5���8�&7��"O�ѹ����I�9�@є?�0PB�"OL z�m�4��%�ɺW:	�R"O�%�iN�6��cd!>`R��q"O>�qD��i<�Qd�ѱH��Uh"O�����>}�0Mšp��E��"O�D�5%�"?�5s��	5����6"O䭺�B�r���3�ȧ�H�I3"O�%"tJ�����)�?�� H�"O���N�4=�j��g�5ۢ5Q"Ob1��iF&7�>��#���6lb�"O�D�*��o�0Հ��3��V"O8��BOC��[��3G����"O� ���үɜ(�V�zw�0+��(j�"OL1�"�>m`5��1q�����"O�L�u%�2|e��hK!k���"OL03w��&@#`���TIf�D��"OZ��r抠�ą��X�dkИ��"O��D#I4$n��`v��k.�Ä"O�ٛ,O�y*�� ��y�)�"O���D��(,sC�[�
$���'*<k"�� (�>tɶ�A5L��F�u<!�$�aj&��a�L0&6 !ԥN6~+�'N*px2�]�S�o�LL�F+G����'�%�ꭄ�+C�]{F��((X4���L�z��(��{bF�?Dgb?OV,�K�v��)ف���GZ(�9�OJ� ����fI��;�/پ��U�7���'��H�f�6�ƣ.�,��J�>X��IDW�q��|BB��R�`��#�E/l�	 -���y���JEP��BCB�_<��Ќ�ē]�(@p&?�)��	����J_=*}~���.@(B�H���s�ļ>C:��ťO5�D����Fh�)�.�X�X�!ʑ@��P��5D�(�CΓ�L+R�UN�+���I6D��"t&;'(������Vt�m�"6D��z� ��P���1�ݮ��y#�+D��9�ʫIA�����&T����,D���bیo��ҡ�Y�w���*O|��b�>=�e;��36�^Ւ"O����瀌5�갓S�(.�P�"�"Ol���#�4h� T ݅cZl�7"OBH�b�U,Ov�{_�$�bg�y�d߅l�9"�E��r<� ���yB��$q	N�:���T��\�P�VB䉆E�n�7∅J��,0�a��~-hB�ɉ>��e�p�85Ƅp��b��XB�	S1P[����N't�)Q��V��C䉎yut����T� -KO?Q�C�	�i�<�@�\�xM�p���H�B�I�a#�5+� Nh�|ތ���ȓ=n����J�|>-��%W
�Z�ȓ4�ٚ��j4���O��F��ȓ+��]3�e�?'�����s]H)Ey��|� �=#y�}J�%�e�b᫒�u�<��#��|��c�v�)�h�?�V�Dy���';0U�w��|*l\���C��p��'|����S��P���8�Z4 ��ě�c>�(����W���
��e��1T�لē{�R�0R)�\�� J�ӄ4�Tܚ0�� ��@��	�f��e!��#Q>؍:FB�8^'t���L�h�P�0G�8�$�L )�� ����8A���iz!�.�R��ꌂ�1��+����5�P�I�C� %/0�ӛ�����C��b�R,k�lC�n/|=p���y���jD4��Lk��8�Gٴ`�6�È���:S����ö<��0��/Uo����FX�s��3�I3|O��+� �=A�<!��o�77�ޘ�GU3U�@u������P#͘��?�w��
"P�w�'y��	2*�L�,`���r#ވ4� ��+���J?!rǔ/Vl,+�ʎ�nz���Q�&D�D��1D��m#%�0F�$)"��4,�kt�\7Q�
,;�Ί B|�|"�g����E=�@�i6]�r�r�RSC%D�8s�Me)�#˫f�AQJ��=���l?��Zv�\�,�Q��n)��=1�I9A����"�F����s@
Px���b�D�����ʑD���q�N;���3�g�j����D��X��="~a}�N�k5�B�F�m��zF���m��Zm��&뤬��c�+P�n�֩�)f�H�=�]�g
�h?B}CR	�3��ȓB�#��Əprd,k�
 C��L����<v�|�@�g���<.ЦT��$�)� B��X�;'|�Ȓ���i��%3�ػ[�4�ē?�� �}�h�lɸ+�%�-�>�9Do�+����Z�WRv�"���G�m�R�ϐ�(Oz��E��	w#�hP��}�v�xC�'�B��@`
��łA拍R��9@t1HZV�RC�?&Aju)�@_����Ձ*4�|��0;�Q��.#���Z����]E I��*C�;�{�g;V���dX�4��O?<1z����">�Q�$��D�2��'G$m�`5ZT ��:f$�D���i��"G4��cFlC"e$?��Ɠ�y"@�� ���`e�����ܐx2B),p85���kl������i�\��Ǔ��|���Y�&Fbu����.v6)�q�ɛey�A2F�E6�(ɥ���<��Ě�i�uik�K1�AS�ζ�t����6
��M�#m��K���Ai>��y��o<�O��H�C�Y�A(�$��6:^�{��xr�I�;kz�Bg@��jP�kV#,�����Ǫq��Ȱx�(�sE]��*=��å�!�D�B��ꄝ2ej��� �#�z�h�J���T�I���nd1bP����jj)R =�R��!y�p�uިn^���O�H@�d�%|i�I{�cQ4t�"�ذ���UIVU�'��B1u#G���a)c��U�a��<�t���){>5�%�Q�K�`-1���mX�xz��
�U����Jڭ^�X��q�ܶ8W2P0��>p�UQ�げY-�M��C1YTm��	20���Y�KÃMp���`ꜘ#�NO��!Ua�82@̽
�f��;�bA00	ϝPF�S�?�"�e��K����r��&~z��L9D����+�^��#��L	�Qؕ�T�]�"�#����>9py���^�@��ś��@�\�F��#Oڐx�R+�C�	�W�;�8C�I7t��C�D���i`m_/{�$J�A=cFhr�π���Պg�R!6|��#�	S50��������x�dX�7^^�����P���4YP	%�%SlTHp��>fʹ�O��}� D���(�k��nxCB"� 
���c���<�6Na��;*F�'#>�� Mh�49.�vd�0,�W2�%�PF�U�A)P"O��.M��xQХ �?�~	*e-�{���pI�^j<�s�W�R�Q>:E=Od�v�RRg �a�U�){p�be"O�L����8�PԠe�*o��)�N4:��[��E�8T�����3��.�T��$�Z�P-�5�I~)���	�^���^ V��CӃƽHI(�B�a�4c�� @MB�5>lԛ��'=����/D)t���p��e�N%r�����E�~D�!)�Q�D���(���+gt���<�N�P��6i!򄎍S.,A�MY&�|H�0�� z�f��%)��!ۤ�ݏ)�)�禹yPI��T��bD������1D��3䄗�[�|:ˣR�t(�#D�,�e�Y���b�žK`赳�!D���dGo� 
��ǋV��t���>D���mO�*&�	�i�#F]j�*�+;D�p�Tg�k��Is3(�.?�0e��,D�����Q(�i�S��D�%{��!D���BI�$@�(I���̃{�����"D�x��mJ��i4E�f�r�� D������Af�pI6E�&�h��7�-D��˥�<o��lq�a95 $D���(D���dK�
y�l�0`b�i�rH�FD&D���5�%7xH��`m�$�:Y���;D�0z1�S�y>�qJœ9d:��qa7D����':�<mx�#@�xY��8D�D�T�R�ҌaELL ?����:D����ͩ~\�t�"m����=D�`A���V5$�Z􏆇v[�,8�;D�|{��D59$X�@�%ѣ0�Jq�bG=D��r�HF�j��uS�/ϝth��x�8D�܈�I#uJ���N/�&xQ��$D��C�[�=���##K�%:0�x��9D�� !�����$
�t~�ۀ�7D�8`E�M�q,|$`Dj
���#)D�$@�.3B.t��U��s���K�%D����e�jT�AMX#��i9� D��p���9���ס�	S����v*D�p9w���J�xd"� �Xh���/D���o��Us����&�!���k��+D��k������D�ugT�S�ڬ�EA'D�� �1���� ~ވ�y��*uAx��"O���`\?z ��B���hMh��"O�}*�����L�0�� 1�axG"O�L����A)����Y%D�Q""O�\0,�f?�hQ@e �`�,�"O��! F�=>�S%�ԇ��p�""O4��MJ�&�x�EH2"�Dh�v"O"�d#ԗ0Ov�R�Ń츥RF"Ovrr�V� �H���ȇ�qк=z0"O,���+و){�� �(]�&ҺHX"O��k��C�9�I$Ƈ`�|�3"Od<s5�)vՐ�R�dNo:AY"O<dȗ�L�Dy��;�B��8���R"OV�C�D8.|#�G���-B�"O�mhPl��O3R�Cւ02��P"O&��BԄOG����"��$�]��"On���B��u}�}�'�!<X]{�"O�9���A�v���Je���D�5"OZ�� �Đz��ؓ��	�,p"O> +D��)��*S�Ҡ���s�"O���J��k��dpk�1'{��c�"O�0�B!��R�2A+G
�^l��"O�-s
�&N�-
��-l��܊�"O�T��B
=a �#v)�F�����"O�頒��~��h�En�lS"O��M-v���s���-d�D0��"ObÑ!	.l��P���a�:ժR"O�X��
���K˽�VH6"O�1*u�,{{�\�GW�����"O2j���"1r��KV(�hs�"O^(8qH�:��!J�q#�)µ"O.�SfHN ;� 걊A�iz�|(&"O~}���~؁�)~W|��"O~��D�]5�v@#��U�>_�j0"Oph;RI� $^Pe�b�*2>�d��"OH�����E>V��2���C!B!p%"OȠ:փC�$��Q�� T�*��Q"O,e��l��[��P��l��<rС��"O��z��� o�����?Zo 仇"O�X&�O"N��t+tǉ�2mݫD"O��(�N�C�Á�^�^�%�W"O�I[% �	���U���{�r���"OzQ�nL  ;�щ3UU��qf"O���6��C�L���A�D~Ũ"O-q(�2{"��iZ�)�(W"O�i"@�U>9I ��w��K&��"O��G�/`��(��˰l/�T�p"O\da���'?ĉZ�� ~�"O�H�r,ڮrT4��S.	#S�(z�"O�X����0s���G���2�"O"l;�.��FVJ}u�ӯv��a5"O��2�?�	t�ی|�����"O4H1�JƆ�X��c�Œ(��A"O�]��d�d:�̈ ɏ0�B�'�p�k�*P�}�Zm�tȄ�WF$��'+�x��iC#ZB	hԇ�?U��+	�'BE��!Ug�P��3�\�X�K
�'��9�L��Uo�#c�V�$�f|�'���b����s�Mآ��8�{�'��%Q5@�>8����O@�!
f� �']
tJ��y���1EŃf��'��	"3�V��.�B���
�f�
�'I�=����VǬ4��/L�y$�b�'��D�J��sU��Xe囑o����� @eEa����JƶU���b"O�D	ǫ�0��(IVR)� �.D�|��_.n�e�F%2�Ф�A�*D�[f�M&"lP�*5!�tSt+D�ઔ� h6H�v���pX���Gl)D��!s�R>MÖ�c�H#!�h�	��&D� �m��X$FKd(	�e�L�Je�%D�ܢŤ��ꘁ�l9n8���'D������hW�n}� !򄃡W���b�H�BwT�+�D�X!��Y�k�x�[�bD' i�X!l��MS!�O�N�����7dYv�`.B�s�!�$I
h`q���Q5��1H�Ff!���(?�}ړG�<=��("�̠G�!��d��=ҳ��*�		b
q�p�� :t�d��#P�0�ӄC�]ML8��oo�L�� ���\�`@��jx�y��@$���.�e�5S��$3�ȇȓ"|K���&��
$�D<QN�هȓ<��P�%se���b��m��ȓm�|i�̈́�/�Ĩ�6N>me�Ѕ�����*�12'ތP4�H�gi���C9N�+	
s�,<b@K�����r�i��L�q%�ĩ���DS���ȓd�L j^�^GEarNel�ȓNT�3�S8=�N�JƂW�J�<��������	�Y� 2���(�C�ɖ��	�Y*;v�'�R�ZA�B�ɺSp\I�u.Q�A~���� �rB�	&8��M�2�R�_�X�Ҕ'�|~B�ɲ-e4�hU��7��#�A %nrB�%�(T�AO�%��a�����"D�����T$G�����/q��!�� D��b�M,*�H�اV%Ts����2D���$.�7l�1����>*�H���>D��2a"Y"W��@!i��kJ�����?D��ǫT�qȼ1Į�5]�D�;D����ڮFi^ukF�O 0���4D�P��	�{�R!�O�X��t0�5D��3���v���k���<��#'D�h���V$*���_-C�hY%�)D�4�@"�1OK���1�@0w<aQ!#D���H2&�h��p�ݛ��lA�
!D�D�1���Hiv#X�����F?D�8  cEE>$��l֛��*c!<D�(���U����s�ڱu7���K0D�4�'�ӛ1(���a��P�D듧1D����`��8+W�ɪ���+�
@��ufZLE��O��;�+��\��"w"܈�JX�cO��BI�.o����+�2b���F�6�
��v�'9�m�|�r� v��
��\�
Ǔ_������oS��X!)H�H�8�*ރA�ȓ[�$X���@xh�2��I�6]�O����.�ʓO� �A#��8]kD��'� I�A"O�*.�;M j�.H�c�H���i�I6`�V�B���|��H�W�dy٧���>Zs��H��PxBDO)I�D�P��u�Cd�	z��a@tmN�L%D<�
�Q�v%���+M�F�Z2��X�����&q�*�CA�	P≖X����s��?6(i�!*�(B��9/���T)܅ z6��t�W~!t�'�Dju	�-'�ɧ�O�H����tj�����FJ�� 
�'6 Y�e�9���C+՜kN"t�c2�d�hI6X��L>��Vkm�`�e��=�0��
 mH<�%�ރ��e���2��2�H7A��!� j�v؟� j�� ��!���Ԍ�漸��'	�@rf�|N�x��0��F>e0�|� ���y%[�9@|�Rӯ�B�M�d��y"�T�1Ͳ��<� y��!��y�L6�P ��-CM�X�v�Ĩ�y�a-DQj`�����T�����k\��y�1p��t3��*E��E�� ��y�̐>�P(߅<V�D1�"!�yr#�kv�� �����R5'���yr�� �4z��M$.��D����y�� )����e����q�D���y�o �\��ߴ�Ȑ�f�	�y�k0�2P�(U<X�H���NU�y�����j�V�̠�)]�y��_�:0�clX� �`�8��Q�y�P	/j�`q6m!��A^��y��
6 ;��8�)M.	��!�@�4�yb��=\���g��/(s���`�C��yRC�<0�!SR��%]l�`�%��y���B�QJU蚝A����Լ�yBH޸��]��K�,�a�����y�A��_���S�/I_iL����'�y��W0c-j�5N�ִi@닠�y��de�p�����;��H�IF��yO�&蝈nB%*Y���%�y�kR���{���4�d� ���y��N�vA��q�U�]�	Q�
_��y�Z�R9j���� L�t�f ڰ�yr�̧>�X@�i�2���Ą�y�Q��,�nG/�b���	C��y2	w���q��W	ʤ)��9�y��# gjk����&Q@�	�yҊ��5*ze;�FÞ}`�$�S�:�y¸����S1�0�����Ĝ�� *�	�q�N.1*��Xg�)	�*ɆȓEP���C��{nh��Tjˠ����ȓe9��Q�e�#a����
O7['�P�ȓ�e�Ck$����K�7����ȓ O�%��O�D��C��,���N�TLZ��ؾ6��p1RnF$�ĆȓmڌZp�I�%4.� ��>�d���+[ �+���!>^t!�Kܴ\B=��l�t��A��I�6=y�,E;ۘ���%t8���ŬF"��Цg�+����C��Em �|�!�#�2E$1�ȓa�@0� �{RR�[��	 5���l���W�ʄ\��a�� s�.)��29}�V/
`�pAU��>T8�ȓ�D5ˑꇶ#V<Ɇ�H;����ȓK��A4��8ov�`F�ߵj��{"��Xց��8�֑`�郲AUt1�ȓ	w����!><�|@qeJ�;�����@�P��!�HKL9ȳ&���
!�ȓQѲP�0�؀@[: ��P%���3N��a��jq����e	�@�ȓS�x��㕩>!�D�Qeʖ=
����\�h�)F��-#n&葡K7khP�ȓ+��P'��+�|ٛ��M�ꍆȓ&�4���\�i'�<��c3&��9��[�rq���([
����oܦ'����QA� � �t�7آU��ȓC�Ѓ$�V)���#0o]��r�ȓ9��#��ɘi�|�P�N�;�ޤ�ȓ>�n�&nG�✱��M��5��S�? ؁
dj��QF�#8���"O�3���EJ%R�dD91�@��e"O��(�۟3��
��W�Q��)�"O��*�X9Rznp�K�8��i+!"OjAS�(��D^����
&_��"O��	p�3WxP����E�sa�]s�"OJh$�O��DCwj$@��0"OU)�%Ė�A�
�u�2�:Q�4D�7��K��\����j�Hӆ0D�x�R�-:֥��F�6��p��� D�t
S�:2�U�S��(��s*O4�
���W��bU��~��x�"O�R!�-vb��S2�O/�riZg"O��9FM�A��x�,߲�VX�s"O(��͑9[R�����'����"O �"��֊q|e��B���Qa"OD��iJ�]��f�N!`t��#�"O���BG-d����́A�\�f"OR����3)M"�"��B9�˓"O$� oU�M:�ˆcT�_�xR"O��� B�B�L����I���"O�Aq�̟#9�B�'ȯ�^�8�"Ol����]-:A�=�D'�&L�.�x�"O�H�申(3L�9T$�	��Y��"O e�
�*K���8d���G,��R"O����,�Dt��jA? Mj"O�8��(A�HIpA�ގì�p"O* BiJ�?����ă "�<UY2"O�05o��.�J��煅�eS.� "O��#��7�0bp��v3�iD"O���#�2 _:�k&LZ8ջC"O�)	3*��q������8-�|0s"O��!�l]�`0���hO($8R"O�l�c�C�w�2a3T'ɷ8:8��"O�$�v�]l���RJ� ��"O�e��D�k��1��v7��2OR�Ȇ�DoT��c@?.�Y���O�$r��͸�ICz`�&�G�9O���v��9s_BB�	ϟ���ρ��� ��I9"W@@S�4���Q��Q� ��>p��(G�!��{W�xb�N�'�c>=��\t�P3g�&d�B�yT��>�å:�ӺGxH�dfhiuf�m���1�ҙ�M��)�'0�`��A�:U��]"7BڔY��<��	j��S��˃t_�40�K�4%���wE3�hO�����`N;&���ɅH�O�q9���	�bQbv*��I�0���"2��I3S�Q�"}2T��,	4)�+��B�0б��ڦ��5�)�'���1b.$ney�Y>�|�8���GN> ���<�8����.�U
V���'������)4�s��my�P�.dҠ8R�V�2��}�G�xb��m���O�����U�]����Fw���O@)�����G?J@�ČM�y@���G�A�7���(O�?��1)V4�	�!bX�Q,4l���@X�'�
��IӼLT5krǙ3�İ0�.G)GI�OΣ=%>A8�'�t�L ���3<I����&|OLc���K��,b^�(�T	<̘ـ��<q���M��fPmJ`c(�\�r)��f�R���&�HO�>�gH!#�����QB�@Щ� S�JpQ� ����r>u9Q�_1mn8���!��%-�� j�Q�� �rU	�#U8��$���r��#�x"�'Ҥ�&a%xq����%�D��X5m*�I*E��PM|�ţ�<ͧ=�����Ņ"���C�`��vQ�u"O�����,�����R��E"O�i{�.W�@\
��	wpR�"O�أ�m͌R�0��V�B2<u��j�"O� �Ó+ǧ>����T�V���r�"O��b��@�R�i�% %1���r�"O�$�+"��E�5n
�0�"OH�"�mӗ"�	w��'v9|+D"OF��D�����>8ҥ�R"O0 *3����0C�%[$H��"OpSQ���oCV c栉��0�g"O�����+����Y���a�"Ot-���g[8K�%郂
��y�%^̺!#J��-�YHcC�y�HE,i��p��_?8�����yr��&n����'@&P�Y���_�yjU9���㉀"���@��H��y2ݳ8������ ��|!��R��y�OS�^��,��)R�,8
�E��yR��>����Ʈ	�T)HfF"�yb�
�a��<P�F�;���*�����y"E����a���frd�1�� �ym�� "ą��S���9Q@.�y���d�q�녅R,�c@���y����-](�X@��Y���Dۢ�y2�ʛ�\ڒ����Y[d�Ċ�y��u0��ܳrDҡɓ&��ybJ�v�*�&��<d�왩Â�yb�+$����.V��Qz���*�yBJ�X�콙3䁥Q8*�����*�y�_jX��u�
2R�"���T��y�/��B犩x$��� ��}�`����y�m
�L�,�g�"�E@���yR*Ӛ��]R�����2Fև�y�,�j���`ro\7>�Piæ�D��y��J��lD7)X�ͫ6l���yڒ43~n0�6B��ʕ)�$�y�+_!��(���^�Z�SaԤ�y��'B,r|�s�P�j�"��)�y2��$�:0�L�P�F����!�y2��k$K��V�Ge�9�$����y��\�L"�EyKڏ9d� ���y��P?8���Wk��>�BhY�f��y��%ZAz�ɑ�����3��y"c� 
s Z�%]6[9��#fˡ�y�l�����9	�4
v�\_�!��Zp�	��͗�>���ȳW	�!�DS ((�􉏧D���P��;bv!���*Fx90`(�$��=cG�-3�!��֗���s�( }�:�fS��!�0h0۴�_�3�(PaP'�<�!���>�d�կS O�ѸF�!�!�D�Nx�홙/�t٢e\�:}!�d�'~��C^�h�T�)��@mT!�$��1q\���Z?H2�Ւ�
�C!�DK-����ԮX�l'V92���5@!����%T����%v�aa�.C(I!�d�;8����ĠJ��R����9!� XYd�����<[}�	k$� 9!�䀫��	S�).ji�As �TZ�!���!Z�0=��a'.,�u���=-�!�dr(x�Я��p:^u��ݫ9�!��$8$�A�DH��)ӊ�2ǉ�uU!�$�#w�t�1��H�[b�<1΋�ve!�K�E� �v�/G����lG�1S!��=F}��{Ed�c8 ��EC!�D=z�I:��'54�Lb���Mb!�DT	'b����Ǉ8>t(�u�źN!�� i3�}�d9��ڡ�n}y�"O0\*���+C�dUx�S;"i�C"O�ÅOߨ6��ݣ6AP>r1��R�"O�EC�H�i�,¶
I�)Fȣg"OpX �MХ.�n݈G�� 	��H"Oصᠦ�wXF=JtG�H(��"O�$��L�"C�^�h�d�>lꀴ8@"O�\R��ב6�>�1�����9��"OVL3���@�F�`���,LLQ��"Oؤ�7kJf i� 	#6���"O̵���@�5��I��]��cU"O�Y���$�d���B�3�I�"O,,����.j��Q2ũ�]š�"O�aPQOúqı�P�u�����"O(�P�U�Eg�4���_�L�Ɯ�q"O2�A4�ݜ5����Axj���"O�
��	�����z�L�R�"O�舱E�U�|�	&%͖
��� "O�`a��n*\2C�тau����"O8��5iG�y����v!�l�SA"Oz�XWE�����"��X�l2�"O�љ�L��6Kt�)�AY�p��4	�"O�5+ũ��[���Q�ۦb�4�#�"O�$I�G�8f�%�0��#w��q2�"O�$��*�(� xCl�6Q���H"O��@��zWx�3��춵{"O\4@e��C�R`�����Cur�R�'f�H��. �d�DJ��U�h�0��'�(�� ��^i��!G��wo P�'��z A���Mj��L �Z=Q�'VZ�2���S�6��W&C`��Y��'&����0z��kV�$��'{Е�s͊���9�!�#h�'#`rKX0?j>�kぁ�%����'Y����b��_͞, ӊ %�iz�'�����X�9�.1��a�l *h�	�'&~�y��ϕCe�9��'��|5@	�'�pT�uE˞�)g�к�	�'�,\GfK�-ՌE�$1}�P+�'׎����?s�bE�f�I5�����'�j�����Q���{��*=4
�'����@�X/V{x}��HVIb�=z�'
r�͌��Y���O�&����-W�y�ʄO�4�aPi?%Y�pP3f�y2D2>����V  r���2j�.�y,�M��@�D�b��(B@G�y��K�B�b���.n� ��B���y�2R5���iJ�ބ;s����y���#OB�I�E�À���e1�yr@ y�u�d�ߤ����g�V�y�b�`��@[���O�Q'�ݕ�y@�z��@�|�ik5.݈�y�c� �F#�P h�$�$���y��4#~\�wˏ)�b�(���"�yR��~�qC�N�!�4Ȼ�@��y"F�B=�I���M��ϟ�y�M��g�VL����1D��� gX��y���m�Z��Wd�)I��a��@&�yRF�>��\�IP�N��`�9�y���6X�@0��\�}�[��y������!���i��M�1*B�	2��A"'噍I��U���s
�C�9bw8�:D�M�x!���a&��,3�C�I$Cx\ �Cj��~�æ�!�XC�)� �-�5��k��k�*L��c@"O�$*��U�TBL��Q�)�F܃%"O&<[�@׭p����d�
Xib"O�ș*Z�9�@��`��4����"OZ"rh@D X!�`�9^�l�3"O��#��ù���:Q��!0"O�|)��=(��dH���%�"Ox�J%�9G*�J��Ĺd}R�.�y��V��*P3V)9{��C�m�<�yb^�G�R��62%�R���y� E�u�@�g,�Zl@"I��yB�G�^E���&[��J�ߩ�y2LZ�r_ ��G"�1�z��� ��yr�$�X�H%�L*Y�(�Q��Ż�y2�ف����C�KJ�릥U��y�3*}��fD������y+��w5q���4� ��$���y�2 [��X5Mɴw>n�r����y"�ٕ*>8D�Q
ۤz���"���y�)�-$���k��j��4�C�y��@�>m���E�\� 9�A\>�y� �:���� i̶E�>��`	�'�yb��0�	�P��/=�>r7њ�y�ㄇr�v���Օ d���v�ر�yb	�tܞɳ� �h��Z��y�+�7uh�1���rh�5�[�yr���;����ɸ��lB��y�jKr/��jqm�~5,�˛��y��ҬB�1��,�!z�}�Ӈ	�y�Z�[k�	����e�$H���ݟ�yr�֜9R2�(Sk��dM��A��yri�&	B|B���k���S�f �y�gZ��`):B�Kd��J�y�g.Y�q�`�Ӂ_K��k��y�I�J�"��-I��� ���&��C�	�'7n�:�̩n5Z�Uj��0kxC���2@�e�S�a3��/dVC�I$z[����Y0���:a��*��B�1�N%���i���afO�/gB�	�"d=KI�?fQ��V�ȒY˺B�I1�C$ʆ��,�qN$;�@C�ɚOt�yC�T�)����6	�dJB䉽h���Aac�W�����9�8B�ɨ���1g�ޛu08��/B�I�d��@:���>a'�J���)B䉑o��}�1'I�-�)0 '��El�B�I�����ħ��/��0Xc�{kdB�	"��eÆ%�"+�<rǭ�"8B�I<�P��N�
$��;����C�ɛ	wh	 ����!i����L�NP�C�I�Og��b�N��L�3筑�[��B�	P�*��'OM�cY��I>%�C䉻r5r`XS�G�x����͈؅0D�8{�%�I��,�&+��e��=D��Xp����x�@L��Шb�	<D���R�	�X���mS�(-D�TIuŝ�
�h�5D�N��A� D�� �Їq����G�N,C�4D�\q��B-�Av�m:��U�0D�t����Rh:8���^xK&�1eL3D�$��G9�0 ��>[� S�o1D�	��{�")�eE$#�|2�%.D��.		6�~����׍\{�a��>D��cq� �1�
%B�#R=1�>2�;D�� �����Q5L���,t!��e"O�a0f   �      Ĵ���	��Z��vID:F���dC}"�ײK*<ac�ʄ��iZ�Fm��x��_���6�-?>�g��{��Y�*�:H�t��0q��l�!�Mc.�5��0t���I�:�2���柼Pe��J@�䑗�7��E�s�Zx��I�W����K�1d�P�K��k�jţhR@��cG�J3���B��8g_�H
@
��)��I-��Ha��8Io��(a��aҤw��	�B� �H��\ͼ�CR�FD˂e�,H�j_@t'�@87�A�D�@�d����>̶l��iX�Q�d����3i$� �+}�FU�,�E�9}��&j�����'�ƄI�iE�U�*9Y@n�G� ]3�'�t���j
$?���'�X�~F�ď�<���D�!����!}:L��C��9�r�q≦Zw(���P��m�lB�eJ
'|T�#���6:H�	 �3�zOT� ��3x~|O�TT�*+h��x_R����63lH�k�dձ+��0�ɶE�4�C�'�䆓?�Zp���Orh͓'�jYh�.��[�ܳu�]���� HD	�h��P ��� �TY(O�	��/��Y�2�i���8�e��f�x�A��05D�B�d]��C�m�ŢI>al؄i�<��O�z���)$k�AfgܔM(VH�QI���|	;�G3��#��5���|"��-�򭙁�T2D�${��[�F��Ҭ�O�	�9;H�h�-7�Ǧb����8Ot I��˨L��X�DS�,�����X��y&΁�M�`�OT�`�@!G��'�z@�7�E8f�[�=N�~Aa]�b��6�l��;�2���R���K?!�O�h2��2bP*r2Ȉ�L$�k�  �d��F���!!�i�؅0���R��q�̟���u�~Q�I�#� ���T#���͚z&�51���or��A$�db�j2�Dû����!n�J��+�"7n���L��|�S!�� ��y�F17�0��E�Ֆ^�z �Cn�劊�B�}�<Q��C5 2  ��g�<�#�6 2  ��N�C�	�R�-zG![�clP�`ԫ(ݚC�I�ht�P�6��E�blX��YR�C�I&gyN��k^xY��Oغ�B�ɋu���B5�X�Z�8ͳ��Y�:^B䉆�*���Җ-�6��REԘc�B�	�>N�l��CWU=�6	�b�B�I]UF�/�8�h�P99�,H��+D�bw�*��dr�/�9*9Iӣ,D�p�֯�%Q!n�A2&ڂ��0   �  o  @"  �,  3  E9  �?  �E  WL  �R  �S   Ĵ���	����Zv����P��a+zX�B̒!r�V�C �{�`�@-7��!:7�Ɨ 2d01G]G(�B�N�S�����Ɲ?L%���9/�T�y��О���G֬U.�-cs�q�`=9�,����*TQQ[�u@�3�E��!/�ia ÖŒ§��?)B�(��C��h�I��,fVis3���H8�8����A�������؏+B���Ë��≓�%���@���H( �]�ߊ�#('��c�O�-b�o�)H(����(jް8#��[S�8c��ϟP�	؟ ��$�u'�'��1�Ҁ�R�l��4�P09Rb�$:�D��OG�'�d�3l� C&ې]>a�À*"l�'����3���G�|��_�F�h�MF�P���w"՝�P�I.��@�q ���( �đ ��	
r�� �؍^���'!.����?9����'2�IX�Li����H*!<�ͅ'|�!�U�o1x����ɖZ���tϭ@%��9��|����$���)�+_������Z ڢ�"��G Q�����O��$�O�;�?9����o�q/Vm��%�7x2i5��t�B�a�tA�ejC��yּ����,	FYEy����@.� g��HM��p®�� �ͱwG*PdD��N�Y�LH��z7cr!�'��r�^#���3�J
�t �AC��<м�C��i3�#=��$���}�� �8ua�B��7�ay�剑JXP���j����i�~�^�Gg�V�'��I�!dy:��N���?i�d�ǳ���O�:v���+e��AUB�O���OV�'nc8����CTx� �z��XXt�D�B	,ęsLL=ז��D��rYQ�<YԂ��u)�\��B�2a�L�E8�`�c`B
�����	�~���h&t�C)�H�I�hd�$Ȧ�+�����6�����
=J`������/�O����WAt�<+U�?� Zt�x2�i>%K�O`��b��b,��+5�٩��۵S�4�Rn\��MS���?�(�"�@5J�O�����&&(����+���y�"�6iR��l�m�ԸÀ���P�u���#,��)�ߟ�b>)2w�Z�;�$k�(ޙ}<B5�k��4��i��A�<��ةJ˼�:4�H���S��;��U���W/�(����O��#�'������&�'�V]�����7_\��.�0qZ@$�'���(V��Hh�cǣlT�}Î��I�Ob�:4(^�iԜ|H�JR� �p�R�w�����O<�P�M�d�"�D�Oh���O��;�?��ԎX��+B��=PN�=�'�C .ܤ5���"��Jb�;N�|L�a[>Ì2�Z���8���;
��`�o�6V̔��\.R��ʊe�RX1(���?��)�2T���2�gG3D�0IsVy��?��hO���%(l�У���A<p�	�؉ Q�B�� x���N��X�9���|��6-�b����'��7�y���'D���Q�C�J�������1��ן���ٟ�kZw���'�Iـ!�D:5�ݐYfID�#~m�`�Wn\6 ������ˊTf4�K�A��J��r��D[6�5�6 G.U4�I�=	��xд�@01S�e���Zp:��}oڸb��DM+r���'+��	CD�\��l��.Q>yf7�Z�'sQ��1C@�XBxxġP3Y2�`�*3D��0&���7B�$���j��9�vƼ>镻ih�X���#�J���i�OF��.�8+q�;V�`��,�!%�7I�P!����O^���!<(B�z ��!0fd����67���Ӄ->�Pl��؜\4��aJS�M.b� ��%>���c�U��0�b�x[���3��<J- u��?g9�A� 	�95P��7��-|Cb����Qً�D��3���ZG�-��͈4����6�O�,��łwr�V[TBpZ�ݤ��>C��h2�]�{ �=PΔ�S��� "��>9���<Y���?i,����1j�O@��:n�0�(5d�D�1b�4�ll"9�n�[snY/u�2�C 91�l�;�LĻ6�
I�|a�A�`:3��U��:#:U�I�i�0��Q.�R!�fzƀq�G�Neq�
��6@����b��J�IǮy�B�O�[P�' �6�SuyJ~�Ο�Q���$�X-�v���,��"D���Wd�1 Ht����7��d;ғt'�?��o�6.��ʃ��-QU�]:� ��M���?qGOL�������?	��?�d�����NݴiIQA�z.�3#,�=q=T ��я!`�����º3�|@��k��H��1��'� �ot9l��i �K�&�j���*�,8��d!�
��6���F�'s���c��6�đ1?~d���`F$�U�,��	:^
.�d�ݦW@�' ���	��mA�j85���7'M��!���{��x�2-�pA��S��?��� $��|�����ׄ �Zy�	�V��p��O���Q�H�R���$�O����O�ѯ;�?����?9��	�I�f�{얗5���`ֱ褀3E��T.q #$�e��*2G:�`Dy�G��;��pB��r ɣҹ23�кed*$6l��a�
� 	�Pµa/C"0(�'-
k���.�"<�*�yD�R,17H�ײiު7m�O˓�?�����HR,\�uP�D��=WD�p�iWџ�Gy��Na&���(<��Akf���$ed}m�Uyb)ƻY(��쟄��XJp�s�
A*4L�pn J�+�I�(�h��՟dcgf�9�B�W�ЫZ�(7�٫lg��#�V.Y�<����,. n|��.ŷaM��<�$��n�|E*� �1L.4�g�K*S#r5�� >�C D۠B������ 	hG�$6h�[w�|2a���?�U�iN�b>!q �">8�ˤ�
y�4�(�,�>i	��cx(l��m6��ٰe
���E'��G{�O��]���塊�z<@%	&E^)"�A�'Y.��
i�����O�'
LY���?��
�`r� a�A�>WVMx6 �'f���-M҉�6!Ƣ*���c�a �r��\q�ݘO|1�dа�T<$`���j��u)�[��{��4!c��z:T$�('s���i17��>�b*Ɓ	5X831)�O�X�! ƚş �P��OR�l=�����?XU@�o��%�O�N�έi��\�<ɱ)٪	� �� �l�4��a�t��?a��i>![�+��}���h`J�m�H9�R�Mc��?�v��.>~Q����?i��?����Ҿ3�踫0,/a�����	�DL�=K �D�3��
�휯N�BI�n��.ԮI��'�������}�-x6c)4D|i�$&�0JhT1��n(��2���Scb˧Uhzqy��
l��5��'����`� !+Rx� B�%8��.O�D�e�'^��'��OV�?K�����A��6���!)^v�^C�	�,��A`��O7X��X�Ĥ�)q�zucݴw3�����4�'` d[����t����� �Λ)K��i���'���'��tݍ�	�,ΧF�ȅJ%C����B�b�g��-��� T�)RME�B�  UN�9�^�@�#1ʓ=X��3�K��Lx�j1a��mƭ����hOZ��a$Ш}��C�ᒢy:~]�bȍ'(�5�J>�5b�͟Т�- ���d��F3�xi���MK����'|�>7MI�8H()�
&E�$]�A�ע:ayB�	�)�h��AgOA���!1��� 6�E���'���R$(��p���?M4(φ�FmBƫ˘Y�ֹRb�|Ӿ�s#�Ob�$�O�Ղ֚���ɛ��b��㔢i�V�	Uf�eтI��)��	��"�)gQ��k���S�\�H�T4H������s�;��1#FȀ�g�������1!hr%rs-U)U��'ot%z��?9��$��#/.�A�.��D�`Q�C(�����O"���G!fX��Js�<h讽2RfS�uN�'�ў�S.���C"C����KQE�`���D K��?�82�4�?a���ɇ�+A���Ỏ�6�>�����H�)�����,����1��G���3�T *xq�4놱v�Jta@P�'6?��8�	^��\5.mDm*�����/�c�&������^9A�j�N�>���قBJ�y`�'J�<�$&00�$�O���#?%?٥OZ��NŋW�����HQo. l&"O� ����T?|�"`)�;& �́���#�ȟn��P��ӮYq�jҚ}�ҸW�����	��,��k��h��D������֟�{]w���TV`��D�dO8�X��C�	��A @���a 4��F%�B��d82j�|�cj8S�On�����?V*p�!:��m�!$0���	%�(�0,�#m�$�Ԭ�A�x�X+E��X��3t���C�%�򄁜2%��'K��ī?�aGCM�vaR��W�.��->D�(�Q���v)�;�/�4:$m�{�4�Fz�O(b^����g�*�.AZ���\V,7�B,>�6m`�i����	ʟ��ɫ�u�'0�4�X�{gLX�[��%)��ȇ�9XgT�csPŋ�EO�AlP�y��O@��0u ���(O"�[B�Q��Q�X8�lęlݕm#���

F
X5n�#���u�*�(Od���'R\���[�vi���3@8Ra!1�g��Dz��=T��šÍK ��k�#+<��D#ʓd�Z��`�#�j�1� e)t��',P7��O:�E����Z?=��`*Ӫ[��m3���N1��1�$J�������p�IȟA��Y�J�u�e�S\�� 1������&z�|i���\����B&�'�hO�Ԩ4�S�0� ��Y9�Jt�O�r` ��'����c�>%������Ľ\r�a���|���"��=�X�J�q�È7pq��q����q��@�d!#)>=Y��0�O���'Y��3�ĘK5�A��VA�>��O�d+7�����O�ࡁ�'��@O&>�BIʢ�B���Tː�5[in7m90$��W�zJ�9�����x|J��5O�c>�J�*ۓA��H�*�@mn�QքC�(x���.	��  �cH�W#���ꕊv��z ��I('����#�D�@Z�I&����Y�LhӰy���'��I��{�Xh*$T�>dp��!Ƈ�ru�B䉏]Ј��hK�!&:�wK�`L�b���ɬ�HO�))�X�jMu4��q6Ǔ�2�\�lZ��T�ɳ�T�r7`�����|�	��ug�'=,��5�?���P��gT@@��h�P*"�˧�kV�J�L|<֝�?��OO�O�FO~\4�	c��1JׅB�A���Gf�P��5QՊ�{}Zh`ď~b�S�N� �!҇L7$̓g�����>X��e����@g且'�dU��H���`=�D�O�����Xڲ��2F680��_�Q��Q� �>���SG���Y2}�|AB��
*؀�ش$J�FIdӴ�O6���2ʓ*D�`B�ޙq|l1�#���ME���2��=wM"�����?���?�������O�����!t���?�}�6��>�`Yq�Vd�D��B�ԺX�Q"@��`��9��I�e�LiA	Y#焜
a��r,����\� ri�k�40}i��B��[&Qr��ɤ6kL�dp�? � ��e/����r�(F��U�ƽiZ�"=���dP3d��	�e\�6�^y����M�ay��I1?�!�'��a=��5"�F��.���'u�#J�PM��4�?�����T �nfd�ce(U#c�>Y+��P(�MÖj���?9��?�uJ^��Xh��9s�Z���!l�ր`l�����¿d�X�[�L&FϘ8Fy�h��,�X`u��,Tۊ-Z��A�r�D8JRn� d��aa)�#�j}�#N\X�H�Ey�T�?!U�#d����P�zh�eB��15��B��l�	 w��#�9�R���_X~� �_������j�8)R������@'7)�Pn�� �	C���*L�2�'$~��R��2V1�X������ch��Q��gu��Ju��҂�F���S\�'bE x#v���oC|�i%��Ѿ��Jx,���eҘH�C*ŧ&$��Z��1k2N�S�J�|^��R`��?g ����$�����O
�S��{��S�����L�n��}��I�*!���6qE�I)��� ��AڐN�p ��|���i\��(��!�T�o=��bwM	%х˦��	���+ΐ�JŴQ�I���I��h�^w�R�W�sĀ�*�Y��Lp`%Ѣ?M��c�A �<�9��D9ޭj��|����A3Av�d�c�κ	\Z�cƈ�r���:�!A�
��|�3c�	 � �_>�b�P�$Z�Г��]y2�����=��e��'�ў<���JQ��L��eH�-z�ȓ9� |2�nM4**�	�F���J�n�;�HO�I�O^˓f�`��6=���Y�J�'.��Cr��Vp����?a��?������D�O��2y>��B v��]Ф'=�\ڐ��X-�h`fIzZ�]@PG�~�'�}`��v��ఊc�LtЄ����,��^�9�����J�}�џ"���Ovq[PB�����q�f��o+z�ɰ����=��T��h���M��v���I��/�x!�� V��yr)��3�2�K%�ΏZ�*�끊���$�զ���zy��$@���'�?��O�F�bc�.aa��G;.��rܴr�1����?i�UݨES�l�^L��N�n3��Y&>����a��{4��#IFVN�4�	4__�h�	�� �6��R�_}q��'_�v(Gn�!A��$R a۵\�¥E{��.�?Y�ܸO�9#��r}�=�s�H0h�4��O~�!�O�����k���h�kծt�h0��'~�UTڽ�O��VҰnK�.@n�')���U"`Ӣ���OJ˧K������?i��C
Z[��p�M����|��H�R��F�C�*J��i�)]�-�T�X��h�ʡ�V7J�1����A�"w^�d �oQ	/����Oڔ���ڲ֮@'�PXЄ蛨:EȹS�ÎC�'�J,��샾?+�u�c@:i�ƭ
��>��I��S�OX좄+�c�j�ڡ�,U�����"O��,@�Ri��j%gX8jG��`&�Ɍ�ȟ@$Su؇'L�[3E��1.R,������I��x�7�Ϧ?
p�����㟜XXwZc����W�+3��a̕G<��d&�<&�~Q�#c��L Z�H�!���	�1�J<	#	�q9��0>K����N��Q�Ý3`D�P��8A(�O��| ��Z�	~�zyPÎ�;�KnE�|��˓Y�^��I�0=�%) $�%�ַ(�F���"߸5+�C��1��tQ6�_�OJ:��S� 97�x7�c���$�|���@��Ֆ�,�(�	tƨ|�%�Y6/��'�b�'�v�ɟ�I�|� ���]r�(A�(Q�s��DjDǛ��>]Aq+��V��� d�A�|�����ӈ ��<1pk��V��=1�ًz]N�#lP���H��%EP� 9�D������bi�)3��<�q��ǟ��N� ��Ro�0&���ÖEQ�yBE\�d2�i S�:��Y�&�yB�	6�y���f9��w��>��d���%�h��N'�M���?��O����M�M�^&B6ogh�4-�t�#���?��jv����3%�b�SEjќ\���"D� ��E���]�l#^�KK78>�H&��o�'e�M���S)[E�Bqm�7L� �d�/!r���El�Rt���X7g�Ҁ���a�'8���(�>R֨9d�t���T�*�m��2D�,���F�S� ����;ְ�#��#�OR��'���K��T�KDAϦi;�@s�O�L��j^¦E������OA����'�bEH#�d �d�H�b'�%�����6MQ���9U.ɣt� iK�gӋr"�uqI�]�Lb>�А��Ո�Z NϴbT�P!�	�ϟ���į<�*�*��v��,���ː,�`X#�����X�>�B�i��*M����eH�D@��.T�R�.���'<����}:���p&M�rV`̄�zÞ����ħo$v,aC�Y�I��9Dzb#>�''n�1X��� �(��iOX3\���i��'V�h�#����'ab�'�f�]��֘�S9�T���Ǯ;���V�Y���#�#B�K2(��`	щFTE�ê�|�Cm��pH�O�10`֝>��!D�H2�ZeY��b�ݡ0b�JM�#�e>�������xRʙ	Hu�\�%���@��[���N�X�Bj+LO� ��af/��m�P�҆^>BK|I3 "O�h:tLO�R�������3��ixp"=�'��L T|�d̗	LN��X�J�w���G#@
KѰ����?9��?�E��&���OL�d�0[4]Rv��17ƼC���Zp �� �S�&D���bR�2f�}X�	���c��ŲNPu�g��+PX���WD�0X��|;���{G�%Ճ�6J&����KϪt1��$�����On�����UP���p蛊�lAh��	{ش�?y.O��3�i>Uo�&Lc��pK�RoN)�4�͖q�'��O$�<)�l�5'e�%(Q�E�����'�E}��~��mxyb��2��7��O��d�?�As
�4\�X�V�ɲb2�aR�`�6���k�O�D�OJ�@��K�6q)�H�	_q�܃��ٚh�4�`m�3`e��.L�1s���$�<;�Q���@�3SE݉GHsd�cB�<�^��h�	cj<�P�HΎ0>zй�LZ5&��I�?��\��X����݊��0�+TÚ�s#G��i!�ĕ	RW`�8R��+Jf�p&W+Oa}�3?���EX�TDpaL	?�8�
�&IR}�d��UxH6��O����|�e���?��']�hZ��u�z�A(!� A�7�i�|<��H�#B!�H0w�?�L$x׈��N�V9R��)O/L:,�����^@h��s)M�V�$��[��1��BJ��:��E�ɵvL�<е�W�Ot�ۑJ
�!�j �c(q����'��`*�#ɧ��R�`�¤[�X��sŃ �H(��!D�h3��\��y�E&Η]��Ƞ��:ғB+�?%�DO^^7�|��˪6r������M#��?	�%ӅOϴaH���?����?�������X�JE�,h��+��_���|�-�(̀�x���Z��Iai��2���������x�� Cn�� F�؟G��B圼'�����sU��1��Q'n9I�)��P��%��=n���H�陥%�<p�H���<��gן8�	�}�rу�-B�e�8�t$���>U�ē_���/�,@a���O�0���i"=ͧ���p�ї�D�Lf~�	�g�����tˑfF������?���?�#��&�d�O���+*�H�IV.���
!�Q�00�C�"��p�=H���2$s ���;CH
Lr$�	�pT=0�S�Y��1��a��%N:�c4�THO:�3f,*yJ)p!"�9q�����ɝ}!6�$î?�(2�aŃ�������r�>D��*\+iiC	�|є�(��(D���!�[��U.�(�t(	�>��i��'��up��c���$�O���%}z��Ԣ6|]��e&"�7�U
�L���O�d��|��%ѣ� |�D�X��
?1
�·II�p����V.��F��5`�g�	!I������7�⩢E��  ���t��"lqV�A뗜1Rrؒ�?���	�YZ��FX�O&<��E��7&�0@I����,�y���P��ڜ8J~'�Ɗ��>�瑟t Ab����dM̧9Ͱ!�a+�>yB�,l�v�'��V>�������	�}���`厡N�j,����2~��@�4Frl׉R��AP1�����)��y�mQ����D�刦�Ar�$�c�D�� BI\�ZJ�X�I�f*�D`�ܒp���(5b�Sܧk�Y��C'3�Lh�L�� �\z:l��#��S�O������v^����I�|"�"O�rBS�����*Lx�Xr�	-�ȟ��p�葏K�t826�3G�ѩ�ETͦ��	ޟ��C�H� P���I�h��̟��[w�Zc�.�5��9I�^������ tP.O�5V�';RԊ���0�� j��|��M-ON|ҁ�'���� �{Ђ�gD��w�l�-O�Q2�'�����C�O��)��,>�xԺ�
�57!�t�Zik�QN]܄�e[�7�v�"��|bM>���z�e��y�>X�P��pBu�'T��?9���?��'��O���j>�pC�O*��7m0?1u
���	9Dl�B��Bx��;wh���3S�ʺT;��",^�$kr)A��#�O|9A��'툤x�"�t�5q�jؾ�p�ƃ D��C����pyk�+
�mbT��� #D�8�0'���d�W��oS]��ͮ>12�i��'n$"�Ep�<���O:��4x��૲�'$ d�@�n7m	�NQ����O@��^�^ �ǃ%v��L�;#�<I��G�\���xᎦ)NNʷȆ d�
�F�ɠ\�N��9��ô��9Q���U��
�p(�
�V'��tc��W~����I/?�|��C�OW�Y���S�!nΑ��σ;IQ�U2�'x����$A�(u T��<�<;L<و�4���'2N|��IG�計F�A�&�8��O�D�������Οx�O�J�R`�'�K�=0Al���l_>E �� D��9�6-J�P�$$�|�>���_(
�b| U�N�'^8z�m�����3�*�S�O�����%����K��?j� P��'Y��[�� �ɧ���į�i覼bTEM�T"�1x���y
�  �rM��<ٖ���gΠ],����	��ȟ�\�c��%B��V��6?���
�O	�\#f$�M�a}bU�$�l�V�#5��l������y"fB6,� 0z��N6�Xm�d*���y��8`^ ��G�!C�!� .�#�y�.R�Af��p���BFr�Xw����yr�F�WȂE ��	7t+�5p�-���y�
>&2i@��d`@���K��y�j�3$LB��.GV�T��/��y�"��r����u"ϵM��EQ@�5�y�*����,C�������y¢K	O\lIġ�sn24ґc	6�y�I��Tt���� ,�����Z��yI�&KTPRK]8)B�[s���y� ��U7��Så�\������y��ʪ2]�� U�9Yh53����y�#V:��cT���:?�4C����yR�݊;~\HbJ�.��a�0�C�yrd3>�9�f"�(Y�X�S@'���ybJ�o�@|b�+P)X&ؠ��N��yr�W)|j�Xpd��U�L��H&�y��%x�6M���Q�0ٓ�� ��yb*C�N�h�2��Y(��\��`ē�y���#e0pRf�ˤ��b�?�y�NҌ[����0�ϰ?nJ1BP���y���g"(&�2��@��]7�y�לlFp�3��.'����c�/�yr+��O_j� *$"�)3�6�y���4AR 
"��8p*Բe�F��y�̉� �2E(R=���5��	�y�/̰\z��h�NC�`���Y�%���y�[� WD�z���Ju�N+�y�E�7G91�@�)E��a�6�y�o���|K��	92���	�y2�$"0�ċ� ��P ����y�L�5�h0E�W�ׂ=�����y�S]��P�*V�����@@,�yB��4ؐY�T�T��!#s���yf��mN ��	�. 
�(�%���y�)AtE��8���4gf�Q2�ˌ�yR�=G��B!O�&�����ײ�y�,��z�R�� �^�v�%�å�yr���[-�1�W@Z���3�H�y�m� ɔ!lغ>��*��۞�y��ۑ1�F��ʉ�-c.zcjP��yb���5���)o�3�����K���y�)�6t놩�O�2�8�:�m��y�凵w��@��	܃V��\�l���'���ˁ�;ld�'���0,��'�Q��ɕ�;���R.K"�yR�R<.|����m�va�Y��cя�ybG�^�D=K�Q�:e\t��fK�y�k�\��ձ� |�J��DJ��y���E����bL�1{J�s�m�*�yB�ѐ;Q�����l�XI�'�K��y�G�5
b�۱H_�p��]Ag�D�yB�c�rLP��,g�^���A�:�yd�7~��]��J�=`i:��'ꎎ�y¯�3Z4}�a�g���癙�y2�q���L6sz��P����t��~Π-�2���/��J����.(�A�ȓ:��qI�"�yF<�����+)G�9�ȓe�Y@f�mo�����)��܇�A¸d	�� $�r����B�7b�y��S�? ����~
Pq�[76W���3"OX�#��1U��A4��9K�4��"O���r�J)[��$��)I!R���q�"On�q'�Ƌn��w� �(ye"OL�ه!���x��kI8:�$�2�"O���$bH�b V8FE�u��!("O����a)	d����-����#"O�8S��4��Xt�@��Mz�"O�	'��=/zX��eݨ�U"OX�+�M�'O�LE��(*�r�"O�=IDC:$L3Z��
&D��ڗ��(z�h���H�0B��'D�H���HSG&�h���>|��a��F0D���sd/w�8��p�бd\����>D��ru�Ƴ_�-�`B�Q�s�M/D�<�G�/4�=����?M��W�*D���� �CW��?�q�%#D��c�g82E�������Z*4�p�"D���c"�
H���K���K���r�d.D���V�IS����ɸFe�Aq�*D����B�Z
�
҆H�e��$C"
.D��FN1,���P�F�TL섚A6D�P���;�Z-�/A&���6D�<*���::�������o\�1�2D���5��K��	F+���yj��0D�\���S�Jg
Ղw
U�Uw�q�,:D����U��� 
��Z���P7�9D��KgԚd�2��TER�f�0�a'D�ĩ���<E�dL��+�lh���W�#D��2ʆ�/E�큵G� ;^x��$7D�8:��� [�T���W�.���m9D���TJV�����7��:ke���m9D�hd˞�n.�*!���w��EyS�<D��˶g �.���S���P�	��9D�@⎞/jEӅ,X�]d��EL,D�೵����<��(�2[�1[`�5D����
�<2G�A�i�a���o1D��b )��va@��m<T��1�<D�hc�%Y�	�]�`��.�b�8D���g�) ��IS���1G�|�+�1D���v�֕�y#ы��Zb\���4D� �C�ݺD�"���㗖INV�HS)0D� �O�0�Vmp��T�5]���l2D���_Y��bv@w)�ݢ�F>D� aׄ���!R�c�]Ҕ�V")D��*�O��������#p<{SM7D�x�6��6kJa�fiW�f,��y0D���#�Ź�(�b���N�Aqc�8D����,�#"�Y�a�	�/tع��8D�d���6]�y�f�B�>��M���1D�Ģde�9�dlY�M��"�V<9 +2D��zd!�<�:�ѡ� �[�>L	e?D���gڙ<=�s����.�N݉3D�����Ұdᐑ�Y�@�,��O#D���@aY�8��(��G�)��T� /=D�,*Db�y�t{'(�*MK$q�%D�P�"¾o�6�㱉�-� X�%D�(�Do-)[��A�)A�����B%D��Q�U��¶ę�b�Nm0�(!D�x�@�W�mQ�j��	�.���)D�0�L�1]���֛�
يd�4D�d3�����2����Z��1�2D�t�+@�a�p�&��g!µ36�>D����)�4���Ҟb���ӆ*D�� FA������0�OZ����@A"O���aD` �̹���9���33"O��q��f�i "�-}�e�$"O�(*vC��r8�댡L�����"O��q���i�ò�9C���g"O�u;�E�1[(�e��閩���"O�Y�֥YⰭ��/��OF�`�"O�a���#J��,:�9>�I��"O~b�D�!��"�m�A��"Oĉx�O�?S���E4=�R`"O�0��ʔ�Br�	�ĕ�<�6��"O��4�F��֝��J�K��%�T"O|�92Dޗ#=�!1D�Q�W���j�"O���S`P7+`NY��敨E���#�"O���iP*U�*}`�D�B����"O0שǆl���Q���%ڢ}��"O�xU���=���'��_��m�"O���� ��U�N���6;y��av"O��A��I�JLd�B��ڨ@�\�z�"O"Px�鑑CZqpӢ�8Nxa"O�س2�7��:�"�0B�<s�"OZ��@��X���񵡟����5"O|1�A> ���͘�= �I�"O����H)!�:(Ӂ��5f�*BC"O�ɸ4�	X>(��b�:�XKw"OR�:Dƌ@ǘ���[�P��i�"O�0%��'��1�P`�?�vmx"O���Tn�	5ge9��:y:9C�"OҀR���(S�4�kɶj$vq(�"OމK��6�*���	:`,$��"OȨ���7D ��(^�2�`�[�"O$C'F�~�#q� �K=�H`"Ol��0��-C����'#��=��"O�Q�TJ��oc�e���G?#�	H�"O.��B�ߎn��%H�L(1A#�"Ofxh�"/�l�C��/�L )�"OD�����@���ӵ
&�"O*໵-�x>��3q�J
��I�"O����v���!*ŧX����"O�RNC�~�.��4i��Ah�eBc"Of�B4#��q��d�t��%�@�A7"O�4��e�5Z��� ��"O���g�ht<��e�><��a�V"O>���E�X���*��% ���"O|!�b�E)ךa�7��x�$0"Oz�7��F0�h�W�б g��8"O\���Y-|�hH����|�yS"O�;���@�%���M-i�yS�"O,{QA !�ڍ҃	�/P:�"O����2��ɥ �#�j!��"O��:��[�	���@ ���2�0��F"OX�äJ˅$m|a�r�ڬHʁ��"OT��b�E�S]n�b@�fo$l��"OBq�Cݒ:�p�N�*v_��9Q"O�1Aw.�Cupr�B��W=�V"OԔBaǞa!��1v䐋�}@�"O~��*XT_*�2��2D6�z0"O��xS��$u~ta���>A���"O≊�i	��L8��ʗ>�܅8D"O��󗭓�\�$;�@ęm�����"ON麐I�}��l��'G iBp�BW"O�P[B��"'rZ	(fP*���K"O@-Q�L��\��Z��y���pg"O���7ͪM�fa��jN;2�|���"O� �e�� ڋm��Z�I�]���7"O���	�$}���J��G8~7���A"OF0�\�ȥȤ���6��"O$��Q&˪@���3�#G2�*"O$�1¥T2(O�(��K�ꔛp"O
���6q��H0π_Ԁd�A�H��aEIXXX��y���9>��p8¬ֻNaвA:D��(�&��/��*�f�"�9�6D�05�ǩ0��i�kP�G{�)Xp�5D�`ʷ�\8dj�+�3�ry F�&D��CH�=6򺬻���>+.�چ�(D�pZv��>|Xu�v�ٝ7�V8{��;D�4�g�еk�ԥ�W(�\o"|�#G5D�d��Ą�&wQ@��K���D�$�4D��!��p��PgÓZd��?D�����#X��ȋ�D��AJ��;D� u�5q�Fas��T�x��@,D�� �)S 4�<ɠ�-Ǉ0~8��,6D��/թ)8���/��@��U��2D����C]h<0v@�4�ɂ�0D�P�d48�B� hKB�0c�/D��(�Gݷj>1���L/#�,:E+D�DH�jީ�Q)D�I�Q
زR.D��y��)^-���D��x����J>D��4��v��C��T�y��B D�L`�R
jCf� �nȢk�t25M:D�` ��
f�j%+�JBv�J�N6D� X!��-^��F�%d��f�4D�h���V&����kC o@��rC4D���#o�^U�u�AIm>�aRe0D��!e̩:ְ��%�f�j��d�#D����NAJ�F `��X�N)��	S#?D���G&��[�i BN��Rk\��@(D� �5c@�<�lɀ'�� �@�&D��s�����&�C+K6� t:I)D�Њ4JO�&��Uٷn�~��DX�C*D���R�ʗ1L\���мp`�$a� <D��)`���[���.�q�jԹ"�>D�89@$�o�|y�@�ʉ�N,�U�>D���uL�:Q-��q2�ӆ9�T���	*D��q7/��c�\������}�d+D��s��/E���A����i�*D��cW�XX����d��ܱ���)D�$ٔ�W'_��A��"J �5C1�'D�L0��T"�.@�C
S�8H��&$D�4����jA�*��ՖH~8 P)%D��v�O�*g��A $(l+M$D��F�	K�,�恖2f}��)6�.D��QCYL���ëR<�a�'�+D����@M
�aГ��'a���p�*D���`�O�`��R�85����'D��ԋ*��e���Ӽy�T�Ф�'D��C磗�gs�HQ�������XT�7D����Q�S�ീ��@L����6D��Sd$�]Rx sW_oh��f�&D�к���t��'A:me��[6#(D�`Z�C���B�X<�Jt��*"D�x(Į*/�킧�Z�lڼ�W/<D�xI� �
���[�Jٜ(��D��
%D�,0A��4O�|�����3��@�u�6D�`�Rc��H:x@�!<p��8'�?D��!4��G\��4�����a�1D�t���f��ؓ�d^�v��xˁ1D����H�H�<���۳9�^�* .#D�� �Ah���l�B���&��P"O�y��6�NaXG"[�u���"O��9��w>��e�ڜO($5"Ob�{4�K�2Ԙ y��]�yR-x�"O`9�gG��� �{b�G ��""O܈Ҵ.��tS�T©z�qh�"O8��֫ O�*���+I�\Az3"O:���!Eot���E����"O��ȕʤ"�0��h[q
�"O(��*�X�&�#B�2-@��G"O�ĺc��A��)#�Ф4&,H�"O��K���Ȥ��oI-`\�4"O���*N�S��K4���q(���1"O�(�b���0���9<qшp"O aA%A�"H;vX�R+Ƚ[s�DY$"O�҇),5��8���B^,-Ze"O���O�I�\Eh�(2f[�Â"O��Q��K Nx`�ڥ��O<r��"O.i��疚�x���J�@���"�"O��B�G��,������-3�
��6O����%.��ۃ��X�g�E-e"�|B�1}r�C1��-���J 1�tI��F���y򬒗H��) /ƚ1*L8���]��HO�=�Om�"됇"�Ȭ;�a�XL0,��')��{W,�/�l:���%>�<���b��~b�W�Su�$�E]�b��&#��y�g#4K�Ȃč�MD�H�R��?��'_����o�$�M�l�,���'��{��������*vƒ���'XQ���Øf�t��h>��'�yi֠��5�, �
�[J<���'4�Q±i��s$ 8T�ҬL���
�'�� Sw��`ON�����)*
�'g� s�ϑlU�����#W,���'�����O�9'MʨrTaV�R�F�a�'�`�rcK�6{��Qs��=Hf\�Y	�'"Vy��L�)��5���D���A
�'��� �!
Z�j���=�q�	�'WDi�&�H����%#��U�'((�'NIu&��q��F�h�$��'���tĚ8n.0A[��Ě,�P�
�'<���@G>��$ٓ@z(���h@ډ�(�:c�`U�m�G�\���~����>v��!F,^���%��s��"�	1z�Z��Bݫ<±���tE��G�2��"�͔& �ڕ�ȓg�0�UK8�Āے��4A����R�p�KC[?L)+��1�l)�ȓh�\���P 3X�U�A%U�`����ȓ&� 9�T�9c��e�	��q�ȓGy�`3�� G��X%�@�U�>Q�����J�J���S钎$�uiT���y�	� tw�*��M�*�rFn_�y��9Mr0�[���L�>1#I�'�y�m��"a{ ��52ъ�s����y�/KG�@Ỵ�ք �LI�'A�p>I�"o�䀝��|�6�@����B�:�!�d��x��*��T<\�81 P,��OxqO�����+�V#����+xD� a��_���dj�X�<����,B����M ���M�wD
�U�b�|��z���dw ��3Õ�] \��&�:^(!� JH`�@�֦o�T2���[�
p7#6�OH��6-˾0Uڰ�C5i�Np0��'��d��Cy|h�@ǌ���	t�A2'~!�� 6��i�S>TH�a�}ƴc��B?�c8�'wV�t��@=g�04��Q��*P���h ��) %Y�>�۲���^�L���$8�g?�f�K�R�~��F�δfb~���-o�<�u��O*0V��0��Ͱ)�t"%�i��}�%�E��fE�	]�D�������=a�J9��>K ���fe�j،���-׼�y�ύ{(�0׉�"x��1�������'�~hDyJ?)��]&[�.p�ؠZ����<D��Bw_-Z�pY�W�6���@���+�hO?��F{ R�c�͑<��BF��t!��[%)�W�ƫ#���P�8!���Nл1�{*��'o|�!���FsFm�6�W�i�&��'ť�!�$˶����W7�2�3(	!(�!��3C��1����n�F�ͩ�!�DD6"�(�U�J&�ņ^�]�!��<Hx��DZ�v���+2>�!�D��!Qά33	[�Z��҄��.{!�DN�K}HK�̏�o\�z ��U@!���i[������"1�mA�(6!�DO�B2�C��U�H3�bڋ0!!��D<K�y &��-����1��!!��b�-Z"M��6 ���V�!���71���F�9U����[�F�!��5�����à,��k1N�j�!�DΨf�d$����#7F�h�䞸'!��5F���3$)^/,�
P�`!��RTJ$��G�y�1s�H�Oe!�>�b�5�H�c���F\�7!�$�qk��p��
F�J� �ȇ�!�['|�h�i��O�<�Z&g͂f!�D�A&��v�N�H�$l#�]<1u!��ܝQ�"���?f�@� 
�R�!�_�jx�Q�K�gd����&:`�!�dN1:�f4�A�^:C[���ԃ	�!�d�7e J%e��o�bɣ�#��!��5]�Y���3�$lH��!�!�O-?���9$��>Ǯ�Kr�1�!�䝘.CZ��A�/�� �#N�#!��[��b�J��u�p@� �^"!�D�76L�S�M'%y�,�EB�!�DYx�ЄC��Au^zb@+!�X�X�|��ENoK������$_8!�dO�E|&��"�G72%4����z�!�[Q�� )�-u �YA��"�!�D0F/��AjKJR ��$.�5�!�=j�-pk�.v`p��6�?W�!�Y#{��6�!A���ǎO%>�!�dE��ॢ��כ�ΐY�D�!�ē�w�Ţ�!F�?�d`qf�. �!�DОt�@R4	�ik��ФXj�!�d\"�x�f�;C`J w�H��!��ڞ�4����ۇ#5lh�On�!�$�9�v`j� �u6N����ԏ'�!�OeVЧ!�%-�l�'�)�!�D��K�L�'�Ɯt�8��d]�TY!��+�pT���H��B��`dҡq!�d\t�U�s�ɣ�
|B�L֧>T!��V�P�����	?�ܵ� n�/=�!�$�7_�f�9e��TԜ�i�'�M�!�dY�F^��IZ�5'�5��&��o�!�T?T�<��k�#~T��P�M/i!�$�1s��xs�:QfR��3�@!�� ����B�Fv&Zs�=C�#"O��9%a�:*����#]�s��0�&"O��p��Ҝ�˴!M�;��x��"O  xu��~��Y�e�]�x���"O�|P$D�7;bl�Z+P�yQ"O���S@ӟ>~ hX��_�r�D"O&�GeS!]�P3��p����"O���Eԕ�!:�^( ����"OD�+��<�F� ��T=-����"O,�yu��;>��
��?����u"O���  �   &   Ĵ���	��Z �wH>Y���dC}"�ײK*<ac�ʄ��iZ�Fm��x򄋮:�6MN9DX1s�"+kd����KQ>Cq�y�#�ɹ6,��nڞ�M{4�Qu^��I�3&�����Q����	֟�i�%ڔ/%�\���I�]An%��+T�Y�Q�<X�N��m��]�N�����?PA�0���0DU����j��{��b�BîC��ɤ1@� A"�EQ��I�͜��<��*O�H�2鉤mE���ш������C:4jRd��P��'�h!�v��'�cdBA��\�Ȅ�ċ�x���Ɯ�3-�A3�>!�dK�	th͙V�>1�j��>����Ma�ր�N� ��ES��AȜ�W3�����݈EC���A�"̳����T�'�z1@C�0d�^����{$IUf�?EhR�SV�PPyB�=
����B�PAy�l|{���ʡ�0{�1�G/�i�E��(�E~�!�8���Vk�J��
X7$�����+� F�h)l�rR& �g�laŬ�ӟ����Ҹ('2I�g�����B�.~P�d����z��^�1:0�߇Q�}S���肔��4��| �~���ՈXk<(O�Ɋ/l�Lx��iDU82j�]"I�u��6BQRP�d�b,	%�d<�N>ف��<!�Nh�Of�@�ME(/"0S��R����n 0@Ԅ���(�䃮 X�Q�|�('�3�鈞"��S�a�9m�����d�I�F�R���*%�䇖?�r�?O���ᇶtb��4@�4$��s�]�4��E5&��O������,��'�bA�$�`�Ydh� �Zș3%�>~�z��ش�y���O�xJ�sK�d��<9��;/X�A#�EK�a�RTc�k9[7���֫ 45]H�z�$Y�X6�K%l���,�ŕ(B��QE�9�~�N�ئّ ���t��[��#�R|�q�!�I.^��`�5�>�:l3DU�D��bR�#qId}ҥ�P�'̺�Dx��H�+���b�֎$9H}��m4�yb��)_ d  ���� �
�  �j�,L�w�(?�)&i��y�l^�?1�Y��e0x*�A�]/�~b�'�~"=�'�?ɭO��%*�	-�.(xr��'&8zI��O�>T�tPr5n���	͟��	
�u�'�B5��R���$N�*�b�рZW�P���(S�l9��lΡ �ީ�v%/�13��[8�(O09��̈�am�9�ȃD˪)k�a�)n�^Lk$�]�D�Q�,��fs8`   �  [  #  .  9  vD  �O  �Z  �e  �n  �t  {  [�  ��  ��  &�  g�  ��  �  5�  Գ  �  ��   `� u�	����Zv)C�'ll\�0Kz+��D������b��G��y����yb�҅w+��ZGo��$*<1��	C5N����]�P
�D�x�|u	 dS==�]"l?���ӪE����R-�ЫAED�58�0)�DȅeV�E�Qn�1a�R� BtK,�`�$6hr,%��t8�����?��F��Kv���Lm�r��2 �n�RA��9w��ȅQ���I�z��6�&C%���O���Od��izQڐ,�*�B���K]�n�����O��oچ!!�|�'�*�V���'a��-U�(5SU�
z�/J=���'��g� ��<Q���-�;u]X�z�I%Z��]��#�&9��D���VX�ș�HI����2?aHH%�(OZ-��:����� @E�M�1N� ��듔yH*�Ľ� *"�ǒE��� v:�"qK]�5��t�G @m�8b��'���'��rӖ���O�ʧ�y�+�/�0x�Q�E2l q� ��?�F�i�6M̦�9ٴ�?	��i�dk�d�  ���F"���2q��5���!�<91%"_j�'�P���aM�t��t�è�B��6"����_n �@��,�Pp� ���@aθ�����u��$E�z87-U٦ٓ�4���O��:�G��M��;��ǯ%Th$���,tV����4/�`�x�d�`�H@З��+?@st�ȏ?J>����i�7͉Ϧi���6u̅:׌����k!�$)�H`s�=s���Kش8,��j�T���9m�f!8�/�wL1�DP�h�^���,&<
a!A?t]�q����?z���*£E֦��ߴ	��͟�G`mё����u��C+~�m���-;|��ҊjlF@c�q�����e�/hf�A���](5�G��O����$�)?�B��w�1�"颇)r���?���?���e���'I��R̦�Wh�:��l
D)�i��'aʑ�`�'�"�'�
%KԠ�2:�N�#ǯ�y1D����טX$~5Y�Т&Ϋ�U��� k"
�<t�R�V����B�c�\U�u���xe
�R�ŏ�J�J����&����\�5 �<9p�Gyb�<a�̍B-D��S'[O����L�ʟ���Ο�&�P�	�'$�EG�~~�� ��F4Yژae�+��'Ŕ����R�)��';������Od�K��%��!�M��\��|1��'@�IJ�"%�۴�?����?���qP�� ��!��U��k 8)� 0`3#ӥKR.h{��?�(��3���G�']�H�h�-M%������^>����l���	G�T��\�{j�7�R� �f/��H{p��xY�a b않�M��Nh �و=㖸�b��X>TšB��8i#E�O��nZ��H�Z��k%���$��8W���FG�3%莓O����O��d�O�"|v')u}���B���$s���׎�h�'��7�Ԧ5ϓ�MC�OO���0�ɪ.x�ժ[4�&9�ibV�� `)@�?E��ٟX��My�2u3$�(��dɴ�ևUW. #�^7S�(qK�K�}uW>�S�0��� s��ǤJ$@����t�r��k����c�{��Y.�?Wr�c>!(���`�$K3�$�[��P��u
7c΢1"�6��vyb�S��?Q�'���|r�EA�����'H�Qq���cCAR���)�'KR��h�-C2�qis��$�B�P���?�S�i�j6m(�4���ɻ<%@3%��`��l��%��dZ��9(��t�SmF��?���?�*���O���O���
�/���*�L-;KԐ2宒6x.�� ��B��x�ひc�����F��Q�00B��)�H�#m��-���Q�֍'�����+����1E�.���r��0>$Q��C7�p3GaO�k4��EXn�H����E"��d1�SC��b%E��e�G�/(�*�'a~�F�,P���Q�~�N$⅊T�����q�V�UL:�鰾i���'���r
��l��iK���9�*h�5�'��#(B���'r�K�[\B�+g�N�.�)ģh��}��>}��;��٧� YYwf��=@XL���7z��P�Ć]7*�`�ht��4(��0����5V����Z${�
���v�9�g�(�r�'�0���O��o��M���jY$�hu��0Ou��`g�p�j/OD7���P$���%��h� e)p�gИsc3} �8'����X��ht���P��
�q�@�	f�
*�����JΦ)�	�M/\�j�f�T����*O��iJ٦i��5��{�X�t��1��OI�L�rI���p��U
S�2ԁ��5i�hS�C�q�$�Q! �>�*y5nՄXh4�$�$?���;��YM�
F���Q8Ɔq��́�%�z$��'a���D�/-0�b�%�+���')^`��;T�V7�i4��	x�J!-�?NAX݈2�/C���O<�� ���Ov�d�<�u㊾f���	7��K`JՙGԽ\?����M���v���'�"ҥ	�(�-�h���:8s�r������O\�$�1��q��⟀�d�O��x��:��(�r���H;\1-���~��'�|��rGV O��3�Ld���J�C���g�GMP�s�C۳=��H��A{$(Y��a̧v�'?Ly�C+�y��z��$�Nth�i)��a���IE�矼��ן�T*��Mn̨�n�98i��ɐ@x�����NQ�$c0�:��ɍ}`P `��/v��	�M���i��'����O��� 5�.� F��:+Z�Õ�ܚg(I�Q���_3&��	�����^w��']�錉M�U��LcT���Dfϸ�}�!k�%7�xCĂs:h�Aj\�-�僌�$�&qX��{7��/A8� �OG�m��O�P�x�S�͛)e��T=}�&|z���gb�A#�oČ,+��Z���`�'UR�'��O@#|��:C)��;�g8o�`�Q�KR�<q!�G9,�
���p��Ѷ[O�	��M���$�XvRylZ۟t���s<D8�O)+"�q��o�+1����ǟ�S��6�iC� �	��\�'�/,�@���%a� �x��#�A]���&�MJ��yM h���
�@9F���ɑj�H��"��KmT�H��͊���9d`ƐhI�H�U�C��y"ȁwh��O�y��'��6-�Ry"�	7�����,鰅��䓃�d!�S"0���D��)6#���.`��N�C��hO�i���做�G�8�2�¶[sʸ�p�Ӧ)�'�^��"�}�����O�ʧ����h�V�V�E�(Ƙ�geS�8((@��?�� �L:�u�����\���K6;D���$��)P�`�)��!����@�	�Q1��"Γ!-Y^�;�E��@� &���/��-�L��A��"�JX�8p����'B�����?ɏ���OT���c�uMl���%t@6�)D��) �:�2h1Ѐ��N��4�)�[�>���aєwR�ˤÜ1u\���J���lyR쑵L�t�'�b�'�剢r�衃^�(R�i@�W4}X}ԡ.�������`	��GL��Oi�4�f�F�~"FŹ�i#��¼t�樋�#�"8� J���>��L�d���QS0Sb���#��$��Mi�Jd�I���ڲ+w4�{�/� kE��ʇ�I��*OT+"�'��Ԝ?�O����'@4�(p��1m�=Y)�O���<a����O���\�h�[�#s���*���+�h�D�O]n�$�Ms�ja��[>��m��"~��tU�dXh��:�x�wӌ���O����<Y.�Z�� !���b�
Uj���2&ġQV��s+-D}y��S!B�K6�W��J�2��-�)��gȀ��A�ό9k@�⓺M}T�A�#-�"@��ƙ�s(𩓧aL�Fv�'������,A��Jщ�;CG�IP�b�b��$�թ��-	<^����H�BQv$9�ڭ^\���IJx�<�<A�0`�D E@�K^X�q�@���M{�i���E�H4�4�?i�t�}�eh��2�C�$�y�Q��?�r�_<�?����?�EM����j�M�0�wB�R�p�2,θ%P�S��~$3e���H��R�P35��!R��7hp��AdX84�Hs�%F���F|Rm6�?i4�i�(�|w�A�?|�D�W.W,�%� ��	/|>�y!w�E!�*8 ࠀ�rN����=3�igƹ9��V+}P�`�`��w$�xC�t�����x��i�R�'g���X1��<�dm鄃�<E���CF|�����Ο�k��E;
$��(G3%�$��'%@�w�B����KA�T+�5!ਂ���
�s��Х����>&���C��h�u���o���h�:���8Q�D��EDݲ~Զ 3���3��f��u��9��S�O<�0RV/��)!>�"#E^�u�)�'q>�A�a�`LL�����|���^x�O)J� �n�=ۢYq�"fo͚��i(R�'"n�H����'=��'��:�0�� ��kꄤ2
ًR�|�� ��'_�Q����6	��	�Vm����?�JL>Qt�9'_J)�rg�%���u�H3U�fE�#��ƍ��+�<^����|��A���$���I�@W��A�i��7��vyh��?��'���|�\�F���>p�H��MZ�OL��hO�=*uc�=�)���3��}8Y�8��4����'P�7��|������ޣA�:Y�Q��`beSv��d��8J�,�U}�'��V���O���!]���w��I��MP�׾q��qbP�LW�����ӄw�E�$Ζ�6a�]���䔞A;p a��΀j���"҃߄{@P�@��1� �e�$X:���b
1P��`��d��ZA���k�� ����J4�4	 �'X67-�s�';�O�,Jp�P�*`JGE�+��PW��OL�d�OL�=�y�#�Qp�,z�jyj��$�����c�hʓ������?)�.�Z(��0���!�A�{��"��?�ш��?	����g��*��l1�G�2 mSůE-��}�U�<8�B�I7h�U#����nrў�� ��9�ΝcS�L�I��a��,^a&�����|X�ↈ�5Uㅠ�R�'MzE���?q�O4){�!�qd�51���Z��LiӖ|�'�hU� ];��h�W��Xg��
��Q"B'wPr�[v팖}���seT�?�/O�)�
��%?�OB�Ņ&jeȠ��,$x(s6��T;B�'�l3Q�G)T#A`�%ȅ67��a��v��͟��[�Z�{xݠ�h\����p�7?)�-�*��ѡ�ĢA �v��2)��]�):���ސ.���&��j����w����F?z���h���E��9�\�SdlԕO��YS�T�b��MT�|��'���'�?Y!�kF3B�Z�!1)۫�:X���7��?af�iͰ6�:�d�h � ���� ]�vK�K�9)h�lПl���ԁV��=$�4���l�Iٟ��;��\_��:s��"����I�`湸�W3��]�ү\�h�1�]������~R���sG�E��c�Z ,�2E-�u#z-Hb�@T�u�֡^�S�t!��4���d��������؂�V�*�0Ԓ#�t=V4�ٴ4Y�I%т����H��$�Ii`6��g̅�B�2�s4�A0R���ȓ5�d��`�0ei�	��`
�>1u�'=j"=ֽi�2_��`��\�a�}Ղɗ&�-B�ϻ4[ܵ�%��ԟ��I����I�?y�	ݟDΧ44a�ա�2VJ����t����]s��R���10j�y⯛���������� �����E��j�j˔:u�U#�NJ/y��]0"�xL�PgP�&�j�=����mp���f [�Ra�C�d�� �IퟤE{��	�I�\M�č�V��ۆe�~ߠC��<*:�2 B���cpվ�^�OnlZ�ܔ'K<��t��~"�IQZi{�I�h{� ���w�H����?iT���?!����Ԭ
rj���w��0�c�U�GƮ����µ	���(��'��-+1�
 M]ў4�3JO*K�e�`-�4Q���rN(�N8��,c�f`��M�<�t��(IJ�'.�5����?��O�e�Bް.��q!$]�ja��2�|�'�~���-8N��s�	�;�x�+�=}�3$���&J;�H����?�+O�;���O����O��'0����5D`���rᄀ�aK�,g��aQ��?��/��H���7����Ϭ�K�,���9�p�Սnt�)9�/��D��� B~r�R�tp��EOۓ6y�ˢ�N %�Ap����U?7[�L�9-w"� ����rzb�'&�>]� �\�r)҃5Zx��6f� +Q�Ї�Q�����ҟx���Ϟ$V�4D 0ڧNqj���\�^�����<�� �	ܟ��I�����qb��	��\��؟`ͻ!�����~���Zp	X�(Q��8��q�Ԍ,��1aKP̧-��$*O���Ã1I�h����N�����U(X��Zs���~�TP	�+K�11��PA7ͧ<�'G��D_n|30ת�>d:�+QƟ0�'"�}����?��ğ�'l4��ѩT�(1;����qRB�	'CG��`L
#-�1#� B�ʓVs�����`�'�x��AؖTɬ���Q,�p���P�Rx�hE�'���'���O���'��隻Eg �(���p�q�Z�4)v�	Q�9�#*˻*�^���V�Т=����=��)Pt�C/e��{�Z<zO�8�C�Yv��`[�$t�fŋ�D�hO&�kV�-c��)'FֲY�jE�u�Sa��'Sў@Ex�$�X���2F��l@�Xz���yB-�#	4�9���?�q+"�G���k��F�'��	&	Q��8��ˁ�bm�s�[�w���W�F���$�O =K�@�O4�Ds>-�0(�s/8 ���Op��)�-$9"�Dz��Ϙ|�����k�8f�ԓ�Ă}�'�������&��sӮ��䰰�)	I����Z�&�f�jw�]�3��d���I
2x`���O���pY�AW8tA
�0�נFP��%����	*�,!�%�h>�h±EO�]\�����蟨��$��H?$�	�G �=�~h����O"�t��{��?���i9h�����]�\HX,	"Ѡ"���U*����O���c�����Z$&�=4��bN5	K�M����	�*l������Eby��L^�o��I>�,x�!C�r�E9��:V� �0.�u�ӎG�,��-�g7���c�&`����n8�I�xG��>O� H�Ӏ��H�a%�2CL�@I�*Oh�Ճ%x�;��-2�:�!����p�O���e�F�ot���Gѡ!Bx���?a���?A��Q��J�z��?���?I�w�Rt�6@�8F���˴�Ժ�r�( +A5YbL-�m��L��ك����O��}��[�ܫ3D�"�D9��Ɲ�n�F�0{�"UY�&F
H��\@�z$ H�f�I�,NJ�ʓ/V�ՙ�����um� 7�@���Q~�ڼ�?���hO���"J�6|z<�G�/<1��/D�p��O�7���Y��Lf�ap�F�<��i>���fyb�^)
��C�La���AE\�d[�e�_=r�'k��'��'J�0�V�����?-�ieH),<݉��+f"Dr!���B4D$[#$�K ��*�$,ړ����W���,����W��<r�j��zk��΋�mLj�H�ģe�$`����.���`�!R�v��"����M��'9B��q�'V��$��8G�����. �200	�'��sr	�#�^�9cON�$���.�S¦!��[y��ع,��'�?�r�G��r�D��C=�@ہB�2�?���dJ�xZ��?q�O���U��r[�`��ĕ(�z�I��&IM��sNP&Gx�)�0fϮ/n���]�< b�+��dB�� -�[���3��=�Z ��ςI���@�W##8�4D{� O��?i�����+vvL��#h}��Oq�yM>Y�D=����À\�����^�D����?�N"=j�YD�QH?$�#A!��D�'�R����'�"�'g�(-r���	��h��@6C��a�n�����ޟ$��o�q�����Y1"vTP���L�q��X_w���:�F����;�d���
�{�*�-�mF��?S����A]3g��xc����W9����$E����Q�c���' 5���?Q��io���"៳�2�@���Z|Ԝ�� D��	�J�,��dra��6] ��F?��Wb�>YP����gƌ��C��~���o�Ŧ�I����{4�%m��?���?Q���y'���B�v �FD:T4��V ��'s2l ӓ ��� �����22�˃�~t�<	��Z��� ��P��V$8=���%g^>F9�!���8��^?F=2����k;�X��D��K�(a�Ã�Q�!��0ˀ�2s%�3)�@9k#�Ph2�	*�HO�)>�D�C�ޝ����+S�Ԍˑ̈́��l�S�
,��d�O����O�����?����T�#L�D�@�q楫!�L�D����W�Nf��0t��#�$�I�
M�Z��mGyr���rA�ղ���"=m��#�a]�3>����ھ<�x8�P�!Kp>�:��V�P(vUFy�W�.H8�,�X�	C�ld�S��	�?��i/"=���	6 U�T{���x$q��f��>o!�d�#]h2%�N�V�1�&F�Lk�'f�7��O|�{��mJCY?��I�p��Y���>RmaK��	Y�i��ޟ�S��ҟ����|r%���P�Ĕ5-&!A����BT�Ioǎb��y+F-�]�n��b�`���<)4��V���E�K�aפ��EƇ+6�8���BG930�ˠ�䑁���t�<ypK�Ɵ�ش�IH$�h�t�R�e�pR��!+���O������Z��5��@ۅ:�u�aZ0^���D�O<9G�D�j�J�X�"B�a�%�^��Z�锖�M����?�,�rq���OH�3��ЇvQLi�H��D��p��O��Ć�P&p�j∙�$ �����L(l��.(�F�'�
t������@��֦-�nq�'^(�:Ν%z=��ˁ��W^e`���%��a��JMk�N6�.ԉଙ�l��E�@��@�A�Oxo7�H����P�4���!V�~c��Y%m I�8B���h�Q��k�ѡ�g�= �أ?T�Ӂ;�I����\	`yz�@,%g�m���	��2��$8 ���ҟ@���Lϻ/�N�XrO��
��H��� �1iܓ��Q�� JR���.�{̧}vRD�+O�(q�݅gn�*��͈Zeʀjb��U(�Q��\4~Ȏ��FGL�6�1�P<�ց�t}҇°K�m��I��G�Υ�Ѥ�(n����<�E.�ğ`��f�L>�d�K���c�Jܫ> b�8'��y�%ۄ�p3�O�/2L��f,���$�@�����'��ɥ~�J��e�
r��X�kڐf���3��݄~���ϟ������[w*��'c�i��B���(��?u89�fB�%�����m[�E�Ƒ����L����ʗ�{�di)���F�xX��"0#h���fL�8��!+Q��"-@p!a��@�Ȗ)"������D�9d�xh��E5<F@�J�9~nΐ�f�'�z6L�'���s�Q<]ꈪ�L�V�9k�%:D�p$m�~�[֧ރ(%:!�F8�D��q�Ieyr�K4(`��?YEMI�����p�n���oK��?	��NV i���?y�OX�4)�C��O�.�jV���|�� ��~۶�z��¾B'�@�3���/���A$�t�'�����6uA�P�����li@��30�6�æO�!B�6�s"��'�P0����c�'��=����f,�<�r@C�_ �@�GP�9�"��%�_L�IZ��*�+���L�4��3$f� �#�O���=*�8JT뎹80tD���C%t�r��<�2 �.՛��'trU>��v
���bK� <Y<u��Vj� ',�ꟈ�I�����C�=!�
�-�51 �Z�(  �On¹�L�TF~� ��,J��K�OL;�� 	7XxK��B�EP9x�jD�'��}�ť|��%������ٟWX���S~Ri��?�e�i��"}�OX�T�� -o�,1�F�%����
�'3��ö�_*��"/!C0�����u�O����W W�\�!��$��:�i4b�'�N�"T�Y@�'��'��>�H��',��� C(��9�ʌEAX Z�����!��p�A�@{1�h('� �S��:b�̂�B�:pv��a�	(�j$� 5h\���̫�<�$?�b�A�#)���]!7�}�R"�8��i�g�ۥa�Xn���=K��O��3�DY�`-fH��>���+i�nM���վ$��QQʔ�&�~�  � /;�剖�HO�i�O��'���F�Y$T"�@���d}����'�U����?I��?�F��R�$�O�瓎*-X)�S.A$(�b5:���)����C��5��܃�Z�Y�4;�K��k\�"P�94�<��q��&�Cm!o���儕����@��^/�R�SE�@%l/�r�	��U*���ՙ������藋�?�T�i�"=ُ�ĝ�F*�ly��ܩ;���k�&�!��&�ȳ����FE��[Č��q��'�T7��Ob�6�)��^?���f�>�����g�vEeB�-TD����� D�П��I�|��玗t�>�(�
�>Y�+�Ɍ8}Fr�HQ�Y0&E<L��ŕK-���� �B�<)`Y�7|�%��wY^|��%�R��i��@��W�(�*ZLQ�戒�|eh�<�g����ٴ`��I�d����W�{�|�
��K�C�Od��DαF�
dx�=]�j������b��OR��I��b���f�C�s��K��'��	�+Z~i�ش�?I���)�Z����(�h��dԍ�="n�*W�����O`���퟉�j1sDh���L;� �.��`�H;�T#62G��rCɜ�(�0��GDQ~��#8 �扌��Q�`� ]��s���]�IL�D҈yaT�7p�M�����>2�ɨo��d��銋��g>� $�`��
�E<� �ʜ:8�<�"O`T/�.�FI1�_/-�������h�M��*,@6��K��(챹7�x�^�D�O ��7A��-� ��O���O���eީ��G��
	�)"��B�p�ArGZ:�h�f�88!,47l�y*b>�i$�^>ND����^'�q���J�u��i�Bc�h�'$�B:�8b� ۧ)��D[��W<�4�*�')���(����MSG�S<|�����i^6˓!��q�I�?i���kWVě�*��O���b�+�_�v�X�'h4`2�-Z}nD�2��X�\�N�/O
DFz�O��^���B�R��
L��_N��T�QBį+x�A�)���`�I�������u'�'HR;���fX"w�� R�)	�Hd	��\="ڀ1Q��R�(A�c�I,�m*�*��(O�=i �M�]r �З	�t�XTb6냑@p�����_��8iĨH�Z��� G����(O@ؔ#������S$t ͘A� �=���i�^=Fz2�ɾr1*����#������9K�C䉏��T�@D^�F�t�����"޼�O�tlZ�,�'�Ԃ��c�>�D�Oj�	q/NJh}�bNJ$|.a���O���*����O�擔}z�6M؍{����U��@a��Q.mI���Bŉ�*��i7�5�e�7�zI��B'�:i&!�
���%e�dQ�2�,�%�"e$ۆg<v@�#ʓS:0�I��ID�X`v#�)~�0�	�,\'�y�ȓt����%[�oL�s��' ���?Ɍ�4�*X�	.�8S��3D�b�5�."3�ON�2�N�����џt�O��-���'N֩a�VC�JYB�	j��J��'����`�bx0A`��&y(B�[�ޖ�C�.� 4k��b�Ru�v�O���,򧢐�&y��&wTE�H�:hmz��K�6:���9�gX q����OuMzE��(	E���q�W&3̥
�O� ���'�6-�Y�O����/W�������>
�Dr�%�x�!��7n6�!��1W(��A��6�џD"���n@D�;�GبTb� aU�\���6M�O&�D�O���#�ؖ�$�O�$�OZ�]C�|� �*gh1���_�� �`�?:��\�"Aؘs����A7擁D����O�̱��]	G"�qꗖ1�%�3��oN%9�Ǝ>)�<Aa�m"�:t�W�|�W��*E�0λ=B*���	�	QɾT�jЮ�eOZ�	9U�z�D:�3�ɕ7]�����Y�.%҅��4m�<C�
E��a�p��]������O6qGz�O��'Ӥx)G�ݡ �Xx#
	�^�9�EGʕs��M��is^%	Wc
�`��`�b��En���SM��z�nT,7�J�CE��e��� �7
��$�g0<���O���M� ��m��7�	8���~xXw��y�3�C"D/��ģ��)������D�%u��Iu.�2*�� !ec،(�:Y�;Uv��X��Āhs�4z�i�M��]F|Ҫ�?�����O�;WN\=�<9��>��<k,O0��$�y�X�*$/�<N|�8baI�0��}�<at��좸��y�Y��G�tyrfd7��Op�D�|6ý�?��-�2}
4LW�\?�5rC"��
.9���H��5��W+ B���Cd����Ǌ�?��|R"A�7�D(�BI%��0@�L�<�A�ʸ�D�a��FQ%"@ 1�Q ��>H�o��Ud:���K�j�B�)m�CE�ON�$+?%?��'"�Af�3T�jQ[���
�'��0S5I����*�J�*��z���T�O��D��M��#^d��`��{�d���'���''vlB��i���'>r�'
��]�8��C%W2i��f�����Ǯ�ON����<n������N̞��OI ��d�x�D̍%V�J��5z0h ���ݱ���X�0�T�BF�<���ß?��(�7��&�8�Bl��1�fQ'
|�5�'�ޘ����?9���~�lzU+�8g�Bр��G�Lit\�U�:T�$�G��#9�pHO,�0(�'�2"=�'�?�.O�'��A�ۥ�H?���˃b3!-d�*��O��$�Of�������?I�O�Zd9����� �-S,�E���� �*���K� �ؽ��h\)(���pQ�I-}"Pc��ʹZߜx��эO�h���Ϊ1Vzժ�h=��e�׭ە
P60G{���?����-��I0˳yv���C2�?���D$�90{�G�y?N�k�B�V���ȓR�
͂����a��A+ĆD�65�'�x6-�Oʓv�q
�W?����|ek�@��@�f�5Y��A��@�w,ǟh��ȟ ���_>H����eG�/l���R/Z8f��;��G���
p�6<L��ڔ$Y�hO�QK��˿}��\�KB���E�Y�+D�+�����uCU�S��<mX�(�!����	�4�|j��Cm�4���?�6��DNSy��'=��B��)i�D;g�\i��3�u�ɡ.����R%>:~8{�Ly�(˓B�8�y�i���'���Xi���	��B��j�"�E�-.�:De_ȟ )D��h*P�Q"
�u8�����X��Ͱ��\J�'q�Нx��Rjo+H�PhJUr�	}��2�Į Z�\U����u�S�(ʆ����Uܧ"=\�hC�$�H��q�T�_��5�\$�I�MP���T�g�? ΀kɠ^�l�e���KCz���"O�q�\��X@�u�������I9�ȟmhU+�1b��ܩ�g\�p��@��O0��OL�4�ރ<p6���O$���OP���Of�YE��$��3��CN��Y�BۀCq�}Bᩅ׊�#��P�y͟`T�ӡ$�����Áj_(Ǌ��ba���xyX1��$*���r�	!<yj�؂�?�r�ĕJ�	�u��F�'(����	�Bt �MS��	��PF{b9O��[��I&I<����S�
#��2"O.�	��݆;��w+�u�*�!�'p""=ͧ�?Q-O4���S1>�,�(C�u5q���ۆV��Ҁi�OH��O����.�$�O0��a�~���+O�z�Ȥ�Nq��x*E��0�	�z�0���7ɮmD{��ܘL\����m�5Y�q��Z�<Sf��`���s��L?��cc��hў���Ox�����8o�,W9-\�щ1h�#�?���;�x�0t���״^�@	�d�J	�m�ȓ]��$H��ɕ�Uɡ�M��L�'��7��O�ʓS0^!�%_?q�I�|B�%
�?�zYI��X�
`�ɟp	�-�֟,�	����'�D7�2�x���h��X*�l��f]p�@� �qy�t�5�ۊ~���4E��hO~�aՏх0r�ͺ��:B���{REуX����!�!fZ�
3�
&)�ƔR�'ړ����	՟D�|�T샋*t	�� L�~�񑂝xy��'h+M;M*�`QI��%�Ȥ�� 9�O6Y�'�d�ص%Pye�8��	%�L�-O���O��$�<�/���w����#��G���0&͜�*֜�`³>��'�BT��)�Oq��8��K	��ĳ�m��d�~ĹW��{�OY�N|�f�PeƽR�Nޠ j̄�r߳����'E��P4O|�{��'���OJ5O�b!�����,�f@����I�6M�O�����OR����W"@�s��nR��y25���0G�GZ��$A`�T�����	�?I����a�'��n�O��D�F��r�l�"!�!B�pH��I���J2���(����O^H8��O���I!A��s���	��yb�'�:u�$,�+�&�pg��r��IS��?Q��p(��X?q��˟p����(�dƑOb�
w���d"�H����?��fߟ<�Ɏ4q�$����?!��PMn�.o�<���J�n�n)ba�ɉ2f,�z��.�M+��'&�8����?�eĜ�!�Ҳ���D�O��	7.��k�%�� z����U� /r�©�O��$^ź���s2h�
��ܴIlΘ�!B�.6��I���dAD�#�m͹ ��6O�����n�rn��:�͓�u��O|�� �%	=��	4��|hɂ�49�6MF�1r��Ɍ&Z�l�+�M{�'�?�#�'1��Q'�OivyJ�)S�.A� ذ+��դ!��it>YR�h�>��	��m#���M��O����?%���g�9ʐf�'B)�����y��O6�X#�`���M�"Q(7M�O�˓�?IBY?M��ɟ ��ӟT�T̓�S������"��BA՛����<A������O����O��	�#0�%���R�	�C&�#^m>6-�O���O0���OP�d�|J��?�O�-[��U{3��2�h-�ZHYói�b�'.��Xy��EPL ²�/������w�����'!�I4�A�N�"&���Х��P=Fݴ����O����h��[�`�O����!�)��I�ʈp"8L
p�i��'���'�^��u�)�7랠�RGb� �5
ڄ�!�DZ4U��Q����,���\:*�!��ŉ���pԇ�.s�5R�KC�m�!�D®<R�`ЄOR��B�Z����!�d3�����[8��U���M�=,!�4���Z�ڦD2@<�s"Y�XI�O����Lƕ4Ʃ��,�(u��` ��'>�
dY#9=����M(�L$�3�[�kTRq�����b����<�F���#۪#IqS(�(�|p 0M�+q�E�s ��^�d�aB�8Kd�̛X{Vc����f�W�t��Q�!�2���L�e|N����Խ��Hr�&�9���fƒ5MM�F�;H/����X�=[4��)m������6��6C�>D9��uOK>q�t]8f�
+���%CB1U� Ւ�^�}�
)��(ΕV&T�`�,�A��p4��6�L���%O�c�f�*��q�JM�#�p6p(�.� g��a���ן���������H���% GD��ȽS����O��5����=o9�Pw!ܙR��1%�T�тd�������;<db�$qv*9P[>�(�'"'���W��A7.�X�M6�DH;6�2�'��>�m0��TP�bX+����g�/��'-f$k��7�	���A&�aǓ0#Q�h{]V-��M�]�Мj�ܣV�~�nZ�4��ʟ�ӕD�P����	ٟ �	���NW�b;�����Z�1 �럴74m�aC��3��O�J��=�g�M�'x�킔E�O~�sS�ׯ �(�Q�I�!R�@&�&�)kC�V�7kpl��	gS��Ӱ�Z4��i�nPN��;o���q%Ȟ/��.��G��y�fNz��'�<���|"ʟ�''h	[��	�	6��Hv�7[a�m��'Ӭ��Gӧ/D=����V��!�'��6��|����$�$�p�r��STH�hG�
:�}�e�w� -��ßh��ß�r]wZ��'z�)�S1~=Bt(��t2�� +�PЙ�"�#c�n����4 a��iX��C���c�? �d��"+�d���9j{�HR)�Z��#d��X"<؊��g� ��6
�9/��N>�
֥�zMZ�b�\�\�j�n�`��ɲ�M#���E�a�)�@G��4)�P�ͦN�F���	O�I9L���T��:!���b����/�����ry�$�q�(�'�M�b�N�t� L�E	�/i_�}��.�2�' �`���',R;���+�Ć-{ n��D[�2P����(,�PS��4;X���Md�5G~�c���8 ��� ���
��h��Tbr�ŭDB"<p�F��h|��N'�`-n���͟��'ô�� �!?���#�$��3�4�"�{��'��|�0f�	}H
0�g#��)Ҡ���'��L@p�P�`�ɒ5�	ӏ]&5�6-@`�'��	�<�<ڶП��d�|Z����M��3q���P��}I�(E�O���'!�}{" �A*��`��.J� !�$�w*���|0��D{H1�d*��%q���מx�,Y�$>�9��=h,��tN�R�c>��%�N��E#����ċ�9��=49��'��>�n��~N�0�,=_�i���7#�nC��/y)
�[�Έ&V���[3U�t��D�'�ʅ	U�T8v^�� �@�mۦe�`�^Ȧ���џ�	+8��Ea,ퟸ�Iٟ������_.F����G��Z|3��ܢKIt���f�{d��` 
�0 iT��|J�,��4���0 :P}�%E�䦙a6MU�lvZ�2����m>�)���|�~Q�vg<�'^�@�w�W�#:��J�ΜOH���怚��us,O�pB����d�?O�5�5 �!ݪ�"�(ıw��P�"Ol���k��0��ph9��(�O�Gz�O}�Y���d`��e�:�A53�N�X�!��4zt�Efͯ�?q���?���%���O���i>��bס9�`�õCD�4\r�K�U��J�s�K&L}�$(�gM����"+��Q����j�a��;ǪP�M��tR3a�<�|h�ǩc�����)> f�\�MɬV�Q��r�$B,����dd�uk*!�'�J�4M`�Bꦁ���d&�I�y�������c���@�'¹1��B�	a5���T��3~y��&y�����4�?�,O ���7O�~�R�yB�M�c�X�Z��_	8V&�:&UП��U����	쟄̧K���)f
�v�[� �.����8�L-��_;.5�2g��.FJ�p	9ʓ$�x��V��l���a,H�{d疓_L�顥NM�\)DŢe'� u��6�2ʓh (m�I��MKg�O��CT��wDP*rHO�o<�ȨV��&lO(�����_�h�3�`��W4� $
O��j#n�G]��ڿ
�5���@+h�4��<ٴe@$ ���S�L�O���2��i#�-�ch�%v@.�pa]�����6"�O���Л b�8RJ7|eh��`*�<C5�ir�
#��'��L�3��k�8�����͚�$�0�B�:*<D�����_bA"*_�!9>��"W>�;1;^-;�#D�2���)"�*�d��*D�r���E�D����ҋ{�(� ���2t`Ks"O�$�-J� Vp��O��'!1�'��<�t�G'���@�Gj��Z���]�x6��O����O�|
%iJ4�d�O�D�O7,مB��Ő0����wo�"�x�)���	s�уlDq�����
�|2��*0iZ����@f*��p^���Bf�� �"ly�\Æ�#�!
�̚kÓmV�A&�˺G9�5?,^�ؘw�T�G�4���0��C#\ͱѬ���ݴ�?��(À�?�}�' ���M*t&̠F���졠�D����"�S�ODRkGCL��T�H1��v4E�'dR�g�^�md�ɬF���E}b� ����Վ�#Y��s��A�n�st�Yn��d�O����O�Э��?Y�����+ܺ[�0x�Ǉ�t�� s��i��SU+$Hx�d+:�	!�G�'o���Gy�(Ù6f��QF���$%J�u�xɁFK�'w�5�p Ay�P|��N�	j|{2@	9`�'l�1ů�~)�Q ���7&{<�N��?!��iO�#=�}R  �B����㑘<�q�R(��p>)O<y���'J��PB�2EeP!c�	B�MW�v�'�	�0�Q����6��Uߖ(0@I�j�6��6�߰A���ƟȪ�ٟL���|����6}�~!�5��wx�psV��'|���XB�ّa��Z1��h����$�F�<�C�V���k2aQ�^����ѐֲс]rz<Qو�l�Y���\� dۇ�7|88�RȦ���'`z��E�M�I��L� �"(j�{"�'���0dĦ@ň|ZE��}$U���0��|"4�¢`dx5�U�\�*Fh��rL<mtZ-����d�6a��i�O��W>R������B�7o�a���d���z��?y�^H��8(ѤP? Aȴ,O�/ ��v��	^�us��J�[a 
��H�hW�F!Hʒ�R��x�ˌu�L�S�"W<G\��D��/�
T���ԩR>�1{�� �f8���2'�%�Up�HMzO.O&8���'<R���A�`c;)3�t��/mt�⣈���xbjU�C����e�B!sw���q�Z�=�'�Q�@���CRx@�V�^��*x)'�̇dʛf�'���'X<��ЩV`�R�'g����K�Fʀt�n����9�1��Dh���
6^���1'I�Z�
M:��Dj���K���L�{��8rf
�3�-��.,��	H�}�4"fC�'	�����H�+�26�|�tb�=��� ؈�`d�%�$,�,�d������'Ƞ��|����'Т���r�x-J���lk@hK�'���ܦxl���gcK�]$.a��'���+��|�����T�,��+�w7a��*I�6�HY8��}/8���럠����!\wm2�'�󉖜a=��Y%�ڻ_iH���A"5S�H�f�ڞr�`=[g`ʇ>j��� c��XR|QX��ݝ%����E�.'���`�&�����L]�c� ��3�gӰU��	��&�H�fGb�����b�b"E�5ahvf���O��2��d�'E�r4��"4o��e�$�(�F@��	A��a�f�Q��3iZ�x+u�R�B�Dަ�Ivy2 �|F�6m�O�7��+��A�gT+�ah�h�T�1�	��R�D�ğ��	�|�e�Y��H$�p0��<�����7{�ћL;,Op�h��dK�P�~�B��?F<��oʡ:�ayRZ�?)�>����v�.��+�-�,���Aq�<V��;^ߢ�s���1�rjAj(<Q��]`0}��铥)�|���0�B�N>1Tɀ<����'"2Q>�D����G�L
K���dM_>g0�Y����?���@�*U�r���2�Lٳ�% @��R>#�PP���[g]k�(��AO����맔x�g�)7ڑk�I�?C,8�#��);4)�3Ǟj��J#��PvCj�X�4�]��ē7�$����S�-�89T��a*�Za�H)x��ȓo�4���\�R¢e"u�R\��M��	��(O����H��HߦTB�>u[�ũ���M{���?���G8x`1�i���?)��?���߹PU L K�ucF%�4-�h��U��bc���\?O1V�b��R�� Y��DkK�h�&��������بb�~�f�#J�LHb��P��J�U�E�MW�'3�`�(10� !����)�!#�իi�yY^��n��򄚄CG�O��3��^�JE������oR �!�HTྍ�7*K�F�����=����O��Ez�O�bZ� 
��¤N�����_09� C^N��e���?y��?���I�N�O~�Dt>mX���/W��)0&�n������9�JX�s�5���e��2��<��'b���- 3�5@�뗹>r9��5H�&u�!e.�aybB(q����茗+����sD
Jw���?��&6ғ��'�B�8p+�xPP�+���"��(�'�V��$�
���7� �Ls��h�{��{Ӻ���<5�z���ڦI��#�'J��kV��<V2}�˕�?!��t��C���?��O���i90r1�6l�/Ir�2�f�-�I3���3n�5�a*X�L�C�o�'�U�ʔ��yH�ƃ�kx:���d��Zv�̊e���q��8�s'��+z-�ACw�'2t���5��F����jᣈ!�0ʵ�$���f�&�P؞��n��.�2h���V;�@�p�"ʓ�hO��[�q=�,�$�T;6��R7i��Q_�\`���O�˓J}�Hb�iF��'���MJrm�Q�����&-elq�n�< R�@p��?Y2b<g�f|a��q�p��DJ; ���6�A���IN�.g�������~���N�y�'k�u�B)BQ8ȩ�c�D�޽��#X%�`\h�[:Μf�J���M�DS�S�t���+�D	�20s�~M$>e&>�`C�2�ڌ��$���#�&4�ԟx&��>��"Έ4VRSf� B��a)�A/ў��MKW�i��'�L�@w����1P �8+�İ�E)NΦ5�	柜�ɥ]b�Ax�hR����I���	���`�j��W�=wh����)f�Q���Gl�5���|�8���)^�L�΄���c�x(B�]�w�����K;�B|8�	4�*��A���.��ԸO|���m�QD(a� i�/Y�`~�1e�	R��I�<�ÌQ��SG�L<9��+�,#��1�Bq!�(�F�<	�Ϡ`��M෤��e�#z�$����Ҏ�4���D�>�֣�S�D	��+\7�p�p����l2֤���ʩ
�r�'\"�'�D���4�	�|baDP�-���FZ0�D���61/ܵ�a	�1RD:Q9GP0�j�]�-���<�`��3j�F-�%���(49���64U�y뵬�k򠌰�&��RC��:��*j��<����.	���$`M�	�#^:.)������p?9�c�����Z�i�7�h��o�D�<��)��!
:p��l����X���y�#9���|b�U#4\p6�OB7��`���F�I!D铦p�@�?q��r6Ę���?1�O�6�d���O�T`�(L�� ��r��Bv%ɇ2g&�;�l\/aTE��ZQ��ԋՕ?�q��)A� ��H�utpz7��0\�@:�āq���(T�N=@�Q��#�*�O��O���[�O�̼�҄ԑ\�y�"O��z�ߋ����+2>\�����m���$��=��2w��b!1��!�Lp7�=�D�?^��n�� �	X���?�ꁟj� d��XnY|���n�!�
��O�I�UC�O4b��gyS�N�4(�&0^7��t̚4�ēCӶ@Fx��$�C6<L0I#�.K6Q��@8�"Z��o��I��S�g�? �H�Ůr}8�I5Ȝ;	F��"OҌ��aӍ}J�c藳l�8p�u�'Ȁ�<a��j�4����͜e�x�$_G��7��O��d�OJ3��M� ����Of���O7&�U^���D�-\����Tn�YC��X����8l�dS�)�~��q�62�i��޹2���h�!��/����F�?)��!��-p2��� TpE�q��8}���0�GiMQ�vP ���6e��d9?�p�Q��ş��>��%��[YN��Q�?C)vĠ�Bk�<�ց�̅@��>x����!	�@��v���$�'��	9ZA��A#���dP�P`�?�֑{�jG�\mt( ��?����?)7���d�O��S?, ��"Q��}p.0���,0"\��&E5$���FϾk|�u�`��Q�'�VP���:N�JHa����ke�tTE��-����!k�Y;��@*p9џ�z���-x�.����U�[�����'d���O��!��Y�'&��������f��Nd��H7D�,�ɱt���*�4{YX��4i5�I�M����d�?K��l��o�%OK��lԤ�5	��:���q��؟h�Ic��������'O|�1F�۠	3\]���ր��UZ��V�@�L��5�|�v�?2�l5�B'ʓ@���
.,��q*�?�Qx�D�,Hj��m��he#��P0!�|�qb;�#���ɩ��I�_>h���5��Fԁ)��B�	�bhh�Ę_��\�S �;�*B቎w0Ի�ϼ~z�$J�Β1Q�lҕ}�@;
T��4�?Q����3N�7�ָov���A��K��؇2�j���П�)���DX��p"\�YU]�vl�yW�G�D/��f�p2��|�"����ē�����'e�r��a�@t����`�Ues��' V�$R�,�vt{��<M���&����J�O��%�b?5Yă�/B�^1Q���0C�9@"�3D�8��$�=�|���Sp�Ԃ3O��Ey�C�c����<G6tsQ됻hu"�n����Iן(.��&`���������֟���!T�bd� 蛊Sm@xbBD�9*�s֋.8�x��V �=2E�-�P`�a̧+������7m�<]=��`��b(ʐgI��q����3/���@��xN��7�'2%��w�%���Q:#�r5�}rʜH �V�ɞr����x��\]*<��&O�V'� �@O��y���\)p"��� R���U��:��	�HO�i<���(0���E<�^��F�`y@��S�?CnV��Iӟ��	��_w�r�'��	�&9�2)k�ޚ_H��a a*.�u�޵q&-���G�7��rd��2�j����5��H��	cW�Y2���Ж�AL��V Yd�ѿ�����$�ƀ����r�!L�, �^�p	��ّ�'J���ĊZ�*D0��M=F��Ԃ� /P�!�ā��ip�	-ΎС�`Y7u�qO-ow�1i	�Z�4�?��4BX�ؐ�#O<.�$0��A�p�@�#�'*b�Lm��'�ɇ'"�l�W,M7V���
�����h�9	WM�b,�Hw��0|�+��H�'�1)TUJ�1A�(|��ʑ�Ň�8��!�!RJP٤N�.(��|�o�c�'��8��Y�A�X��a��%y��AF)7�fŇ�y�
uc�წm��@�rI��TW�I�
z���q+�����ׯ��_�fu������+K�Q��i?��'��S*���lZ(�&����v��
���4A����?�BױB���cg��!��!���	
uv��M����G�(8Q��^�m-����N/Pމ'����v���i����`#ʺ#�b�FkH�d�1�OM(|�u$�V��hH�i>~� �O<��Sß,�L>�~b�\H���!-��'��{���D�<91͈�&
��Sn[�h� �jC8�dӋ�dחu*�ѯP"",����\���{�������˟ �	� v���$��p�	ȟ ��ﮩ�1i��#�p��._�m�t����V�-�"�AX�	I�,�a�r��O�D��)dV��u��}+��BU@���X-od� "4��*���)7��x�'�Z�M��)P��c�d8�w�ֽ���VZL9K��@Dd���6��B�4�?��#��?ͧ��Y��o� hd��f�]�c�E�7����}XJ>Ɏ����ɉ('�Z�r!HP�5_�e�"�N*�~��'�6���%�p���?��'����-��+��@	&���*��H�H�6��M��	�O����O����ٺ[���?)�O���j0�<e3x�aU�"�TY�C���t[5��-\�����GaQ�YK3��l�'�4i@��f�R\��Q�)τ�[�lW��>�%��6Q�5�*!Lͪ�HCΕQ��Of���}��!�7oK&	�0Hee2>G��;�OTm+�РN��5
�N�#="����"O�,�?�0H�8�+$ϋ���=i�i�'�|��Wt�
�f�Z(+�._(z��F�U�񣖤E�����6Z�TI����ΧB���M#(v�U��4 ����ǔF��m���� X���i䢟�i��� �M3ʓQ�����;k�r1'�[��xR�
Q�2����
�!��<CC"�G���ҥ&ʓ/Yj��Ƀ��ɪ5 �z6��j&Y��h]�/�C�)� |u�F���x�0/�(��s
OĈ���+'d��C�Ͱ �@� 'D��ҒO���%����I����O�RAy$�iɄ�u�D�G0v1B� ��2a���O��dղ## b���Z��u��rE��3�"N0&�0�'hw���-�	?Y0 T�%�.�%�<�. �;-Ѝ;P�ʟ*�^�8��E1�"$�SR>=�ֆ�+�����$0�^D���>��� Ifr�-��)C�Z��Q�������a�o�!�$I3)v���4aD�QҲ/�>5�,G{�O�̢<Ģ҇e=��2c�@ ]$�1�(K�C6(7��O����O��Z R8=�l���O��$�O����)��ah�$�'+AvĪЬӿ_�Xd1a�2-.}���=
�Y�u�!�==������'�n���ƍ:|@Ar������*U��V88j��kP4r�MεR�q��e���Sp�G3Q����p��x�p`Jt�./Z�O~pJ����ē*u�M�FE =��Ͱt	��0oh@�ȓZږ�R�.�+
j��p�
Ř0��O*�Dz�O��'����ʄ43�Y�l�+3 �
 ��e��Jr�O��D�O0�����[��?Q�O�H�ڳ�N�&�b���b��B_4e�i��5��1/Rb@�i��c��=��jCZ�'��4Pq�^�q��4� ؓ����g ��`��˒QmX�Yb�]�C��qr	SS�'�85{3��F���iӾHZH�J��?9U�'����+OT��k�bW_�
Փ�'���*@��u�(<9���"!<�x�{�n�>�O���%���U��������:H�"�BA�K,j$��sd�߈�?�J�p����?��O���MI�XB��*��+l�}!6H�e����A�?����ۗV츼�h�q�'��"��Oi������V�h�:�S�0�\	Ar��"X��Ѣ��(w���p)K�'���p����*9������Z��/���$���Y���B]'$J �6���;s�����Rs����O'En���@<�����ꃰi���'��ӷ>���o#WX���L�?vv�1UOZV\1��?y� �?��y*��0V���%L� ��c4�_�QtOάr��)��1s�=��A(rˠl�3*���O�Q��'�*�O���l�5��I9R��5aB0}��y�"O�%�C�΄;/���ӎ`�͙U�'��<�& @lC����W \~dݫ��1L��	��I�7�y�ƅ�ӟ���ǟ4������$R�l.��V�t��x	����Jo���!\1Z��Q!���	6@��O���c�q~#�'e�AH�A�rk��I�d�u4� !��V���)����6\���$�G0��$�CCڽ%U��%	Jb�AF�iN7M�Ov͋�b�O�N3�Y���1:q�LAS�/co<H���ٝ*�`t�S�'y"�'�
Ҫ8RD�����sԓK�x�ٴj���'67��O�������'M��@j�.�e��1���=��-�D�i,�7m9�����O�@�d�X1Rm�4-��ߧ�j�
�'��1`�@Q48M*�`�L�prX`	�'�0m�L��so4�P��=tVN�@�'�XIc�Q�!���f1x���'���܁%O�U���S�ˮUj�'$�����ɎP��0M���Ĝ`�'� �	Q�ɤ�����f���'R��v�Þy��%��NEj[H`��'�MaA�-؈Xxf,
��x���'P�EH�i���h�z�LԶ%Ԙ��'�,e	���.����'σ32gր+�'���x�
;$u���?VPde��'��ჵLI��pw��7t���'ς�yp�P�Y�l	Q��ғ W ��
�'Y���rn�+~�%	�iAs
�'D�g��3l��#T�P��{�'UpZ0hج@CGx�|��'A���M�9�L�`2��{?���'8(xلHP�V�ʙY�鋬o)�!�'�4����9R�H�TD$j!��!�'� �2��͹n�m(5�Y�b	�'p<�{�m�9>��9��H�jv�R	�'j��P9m���E�	[&Iq�'���Bٵ&�M$Ɠ� v�H	
�'����(-M°Z��@8-����'��'F�,G)����92��	�'Ql�g(ǧhR ���.�+	��� b�� �	�$�!�Bπ-��0"O�	�u���؂'��*U�"O0�()�h��4��=6��a1"O�%b7a�.�ډc�_�Rrl�Q�"O�D��+RmN&L�eF�4����"O�`��] 8�����Z��z�"Ob��FE��E��<J1d�4F�,��"O*�#g%S$S�
�`c��~	�"O�Z�%�� ��8���ݩl^��B6"OZM��BN�v�r{��F�@9 ĳ�"O��@�בb�8-�B��h{����"O�%Z�gӒ\e����;({�|`!�$�-"���5�T,��ӱgU��!�ē�^�b\�gl��a,xL����$YB!�$�5�p	��L�@���F10!�$���YW'�;�.djg�X�!�d����Iߐq��X�s��9M`!�ۭrZ����j�t|F}چb��8H!�ę	e�Hj%�_�8eș�7���E�!�͵K�h��*W�q5�!�EF�!��Y��a�E�M
�5��_<e�!��[�l�&���� 
�����R0d�!򄙡I#���4�^pR��_�7�!��	�4� a��$�����G�o�!�Ć�-)�
L4kŴ�m��E�!��+@=�͡�/�	'���բ�1t?!�@v�6�aB�P�=�������f�!�$Dm-�5h���5��)���Ʉ[m!�[�Vm� ˑ�`0�,��Eӌ-�!�$׬r����m��!���*E+�!��Ρe���P&�X���WHػ;�!�d�:H�>Ѳ��M��b����9&!��L��-0!J�/X�1P��T�'�!�DNS@�I�DD�,;�5JևE�f�!�$�.�(QiG�Rv��1�'�Ȉ�ӭ��ok2����K�~58%
�'$< �5ז{���ŀ'B楲�'CȘ��%Ʋ�`m�.����'e�͹��N�q�@��k0���'g�����+z�U�%�%J�y
�'��m�����e�S�U?�I@
�'�D�'ȝ������p�M*�'�1�Vb Kޘ��&��r�0�'�*���h8�����?B�*�'m�c*�)T�ѨU$,�Ѱ�'�Z���9MJ��U���Ghx
�'l�0���U&6�6}ҤGЗ(�V`1�'6�z�<l���B4�]�"�)
�'OU`����2���
4����}r�'p�!Ԩ�p��6��0��'	|�$jן9|yqfMNy���'s�uQ@	!)�Z1��w"B4�'m|�a���,l�9B��ߔg�E��'��@�̝�	��5�"��&��
�'4X�!G��x��W�|�D�9
�'}^�;G�px��zFˆxޞ�+
�'%R��;E�`TB��@%mO�A�	�'�0d�� �e��y �EiE(���'v�,9��!W,�`d�&]U�)�'��№�Bp*���5
(p�R�'��	"���J)PĻ4#��ze�p�	�'VR]���1j	3d�˒y���	�'�p8���B@��`d�I!"yrXx
�'<@t�'R�<Ėx���)Tu)
��� �<��LP�N�z�RP��z.�g"O0샡�ؕf�$@��	�>qֹ�G"OR�a�Ѕ~��`i3��.6.��"O  "ŘMS�|HԪHA
�YYd"Oqqfd�tJ���v�I�c��
�"O�mѥ@/����U$�? �$+P"O�Ce�9~x���-Y�m=t%�D"OX���+�<Y]�P8"ΐV(�0[B"O�]�P�"c^0(��ψ9� ��"O�=a�!��r�T��E�j�&��U"O�(� i����ta��/q�HkW"O���L�![��q����V�9C"Ov<:����tMH�/H�~}py�"O�A� A��r��$c���s�PpAg"Ofx�m�j��<q�� �
���"O<trãW��P�Pa\0	�8��"O�Hb27yv��e@ҁ�̜��"O�X ���	rj�[�ʗb�h�k0"O��"s놓4�B�����hT,T!�$�d6�<}�:5��X�P���'�`|8wC[7l�Axk�5�|`��'#u�āI�aT4<b��]�3����'� �7?���HD)^�}�>���'*�-p��wަ� $��F3�$ �' H�+ EԌ����n�iiQb�'�]�����4p��c��8��'�镯]�<����adͶbh�8�'VT��1��$���Ój��\h�'�6$�%�N
]���p�\5b#�̰�'���L"���x'�ݴ��h�'���k�����!׈H�|�N�x�']�Hq�J *�4��'Y�mz��'R�Q�(��J.L��qϚ�cJ��y�'A0$������SD��0*u y"
�'ݺ� n�xl��k��,@l!
�'B� )�� ��t�3KΛ0�| ��'%(�`2j�!�T�ÊZ9��,q�'I����.�;7��ɓ�M�Yb�'�-
W��3�L�v}"�C�'X����&��,����0D��9����'�ҌYS�Z�y�U����5���'4���$��$�ZH�w�\�3�i�'xM�� Q��!x��r	��(NQ�<��7v�4��gĀ>�bȳ�eGP�<�TgQ�T�s��?1 �CeGO�<�"ND#tQ�䉐��8ߜiS0� r�<�у�}��,{W��2z��q��n�<��%��Y�c���7��r� l�<9�O�^p�YrL�/|H�Ej#�FQ�<I�P�x�`C!$����p��b�<�Q �F�}���W�fX	uCH�<av�&[�uIһA�1��Z�<1Pn��}�T|i�n91n4SF��~�<qA��=RP�#��
X�Q���WO�<y���+Da��������N�<�'gt���"�L�}�*����PL�<I��[�p��Ĩ������!T�<�#�8���[`&Fב�Y>�P�'w������A
����_b%05*�'�6=��� 6����gж p
�'��|���(aA:��1��\Ix�	�'& ؊�fվ}�.]�Q芈kdC�'a|��v��b��|�@@�Y�P�Y
�'����#�h�"�ޮ ��p{�"O� ��0M�?��*�˛�^V�w"O4h�����]Xh�p�ˎoZ~���"O6�Z�N�@�>��π�X(��$"Ov�B�*C/XH�m��m��+U2p�w*OV-��-�7G.f�nԻ�ȹA�'�|y`'!�
A�&/^0_�6��'�$ԫ�KW�Y�~1���ҩd�0t�'�r�{eC+w��@k`�Ũm��'MP��U#Q,Dj��ONv�(�'n\k��A[d-���HN�z��'���`*�0i2�F.���`�'gB����c��d[����,�
�'v�I� k˓o�$���"d��
�'�0}*�A±h�s�L�ZYH���'��MSH-���'�٘Jd�'~=�VD;, �A�G8J�`
�'}��EȎ�"'$�W䔘I֎ b
�'�x�9gc����1���(D�L11�'�D�sbW�%5�DB�D�#/���K
�')�i3&�@�*����W�+6����'kz�r��<!�� aۘ#>�1�'6e��K�4�Ze"�M�J����'���>~���W�R�#��R�'��0)��L��4�R(v}Y�'�m[����H����L�.���'���!R��-$X0�
���'(�0��	���Da0��-F�
�'o�9����+LZLQ�ː~_�L	�'���QW�N(3ј�9��T�HW2p��'L��3�$x�f�ʦ!��@�i��'�H ���[��vᖣ>*H�
�'�R=a�o�p)�%ɥM^�5����'����0*$qh� t�$/_�H��'BF�RrAK" �R�+C�+�2 ��'����͹g��8��-��B�'�u塑��H
�N�+d<
Mx�'��l��䟉MvF$��	^,T,|�y�'&,�	&�|���F�ǅX�y������t����^Y�	c�.��yrA22'XH���-NF �� �y�Џ/h��ࣜ�8�2�	����yH%}}f���J�0���3�D� �y�O�<I�x�@����C�чp���d��6�r`�_�%K,�2a���!��.��`��׋jZ�eA�đ�J:!�d^�\Nd�5���I,�Y�+��!�dJ9�����?)>&�YEkX$!��rzI���3{��Q�֛:!��[54�Q�*��4�D�`!�D�(+[:�����4jp������nf!�X�9��Hs�*R�p�i��D~!�d�F��q #��%��(���~ !�G6.N���b.9z��$��!�D�6wp�ʣ(��4aFaC�Đz!�_5t�&��7�D�$A��j"�ю !�Q�Xf�1�U9Q>Qg���C}!���Q�긚�	!���@�E�0r!�dD�D����#��d�-�T*�+!�
;5L��%�_�V�\XA�T�#(!��!\"�ɠ��$y�t)���[�v!�d�,E�.�&E;V�pX[�i>n!�R��y��H'LÃȈ!�$�7T\t�U\1]i�11�ź/!�U&��}Ҥ��\f�I���F�k�!�� X(���^4 �4=8vcZ-�~��%"O�y��Lf-�P�����<�0"O��d�A\��-1�]"h��x��"O
�`c�To�0�0�aV<z�|`"O`��.��g.�0Z��әΤa�"O�]#jO�b��غ$@T2
5Ȑ��"O��Y�-@�Q'ԑ3�B��npk�"OЈ�C��GDTHJ���(��T �"O&! bcT%����m$��Q"O�]� ��XLD *��y~�Bq"O��u�#��3�D�/b|�@�"O�q����E[pܡ�kK.��t��"O��3W���7�J�Z���8Y�f�"O����%�X9� ZB�0*��$�d"O��3��!`��`��II�¬��"O�����R�\h|�˶:#��C�"Of@��H�\�P��$�
3"O&��J�<@�uɇb�5�pba"O�I��I N�2��EB�8!8�(ZC"OԸ�	ٞ;���AY�
rQ	�"O�a�-ا��ҤO�;ܚP��"O�@V��h�!4��
	��\�Q"O�"UL2y�T��狣oϬ���"Ot�s�&B;~Y�g�ĢR�Fu�$"OVAi�	�����O�=k�()�"OD�k�mMQr�)��4�"O���t��\�|:���FΉ"6"O.�3D)��$�d�����[��rg"O��f`��/�&�¤@O�vV9@u"O�Hr�n^,HT�s��C���,a�"O��l�;?��Bwd���0;F"O�-��L�][��
$�|#BTa�"O��Q l��U� �k68Q��"Oz���fY�`6�m��mˆ h���"O,��D�[�i�:�XC�2%�yA�"O���� �Zx��Q��=s٘2"OD��H�Rt-
�FRi��"O\PӐ�q.�ЩǪ%t@�y*�"O�#�ĺ~W�T���M�_�0���"O 	�BDL�^��k�"ԋ<T��"O �:�n�/�F}���L6V=��"Ol��' \/@�)ҩ��ZZQ�r"Oƴ�6�0x��d�'H��Ol���"O~�c�<E�pa(�:f9x�I�"O6љ�Y_z��L��	X8�w"O�0�JS6 u�	Rtʐ"N�&�#"O|T�S�G"H�ӎư_9��3�"Ol�bCE-5@,mx���,�T�"O�����;9��y�c�M%8�A�"O�e@�K��L8�� 2�M�l�p�"O�})����a�ސYr���o�@�<��T�y�8(�  I�:U93��r�<Q&Ɩ�>�:ẖ�˂=�֭����L�<Q�(ѽ`���M����$�N�<�dË�j�h�㗫Ւ5^]D�WN�<D��g�"���-V0(�3�Od�<a*��#�~1H"'�h�E�~�<����^��9�!�>&Z��
Bi�^�<��
�V���&X��3��DZ�<)wA� �0 2��8)T)p��Jo�<yd�K/���t��3f#��Y���f�<)V#�#T(��`� �3PS��A�K`�<9CM��[TސA�a��a�$Fw�<9`�C�@?�.T��F k|L ��S�?  ���i�=lP��XË�*�L�s"O���lI�g	�Ų��?\2�� �"O�@y!-��C(j���m�-z*K�"O���&#W�p�?yԅi"O��j��eT��j�Wz���B"O� ��8�V�Pv�I��*e"O*̛g���'�~�I���7h�ЋD"O���%n[�ȸA��5�ưiv"O
�"Q�̚:����Nװo��PF"Od�F�E�T ��mZ6j�@���"ORIb�-Q���M@{;�lG"O��%+�28w^ [�P�a.Ȱ��"Or
"�ۉ��P�(8d!f��""O�l�`F�3h�Y@�鍲$�!c�"OrIzt�E�G�I�H׮h��i6"OL��E��Er*Ճ`���;��
�"Oj�����2c,0 !e�i18�Х"O��b�b>�D(�C"�3v.L%"ON|{Ei�$ .E�7#�t(Ia"O�H��,�N^1C�ˉm!n)QB"O�ys�źy��tk�23ApU�a"O�̱"AE5UB�[C�*�*Q"O� t+E�3Ҙ���k"4����'<Z�0a�ËP�L�
e��<DFԥZ�'���e�X�13^��7x)�+�'��(g&Ҧ6T2$�=^ϊ��'8
����8��=�g�4J�>�q�'�Pa#g�b����K
9w�}K�'���	�����Lk���)���'w�Q�Df�#}d�J双G�6�K�'�~тWǩMnp��t�'C)2�;�'� �Ⱘ7hl����V�sj8�r	�'��u�҈K��A bg�i�j��	�'p�A� ꊤ4���i��dlY�	�'O2 zg+צT�LH�g��!о�(	�'T0�GĥMP����nM0u��'��E���P�o��i��٤Y��0�'exa�v�N�����T��|�'�0$�яú�^�a�#��yK~�!
�'�lL���5n�A~Tf0!
�'�ڬ�o�J%@��Em�'u�����'������C���E��m��x��'n� ����A�pP�e$ɢ5Թ�
�'�tU(���m����D��&����'%�	�C\D�oX�]��8
�'{�\` K�*X`}���ݣ=/��y�'!P �
�\2�y����/�>)��'�^)D��iB2$H��."�����'�,G*�=gDx9��"V�����'����%`�*)�`xulŰO(иa
�'���H�*V�����߯}�h��';0��GW-q�����	n?��'F�I��-�
�A,��De�'�*���䄳h���z�I�	�v͹�'�R`j�k�u�T� @�F�?� 
�'�̝ �'� ���Qc/�#�����'Db��ȃ�h���BS�Klp�k�'}�� jwL��z�E�=;ލ�	�'G��C�k �ha��b��2]��0
�' @}BF�ʊ?*��w���v,Dr�'�nP�F�j�6�b@l�7e���'ۜ(bl��k���S��_4h[@u�	�'�Hi��EB'}�i�ӅӋVl̉Q
�'�R�!���8�Aq�aڿv�$1
��� ��ڢj-L=Z8��J�|و��"Oȁ�ȑ3'��Šπ�=��ŨB"O����şc���+�Le&p��%"O�9���\�I2:���F	v(�ʵ"O�$��NY�
�X!��9Z�f��u"OD�!�@Հ~��u��,��� ��"Ol5ँ�4H{�e?�e��"O�D"�#+�����#�A,EK�"O$�(�|�� �B,8d;�"OR�d�N��)B��`B���"O003b��6c�p�Ig�X�i��ɹ"O�T���^<�4ygʮV��E"O���UC�:#X�H�#��̈ZG"O�]�JD�CAp�;!ҫY|�S "O$����*��MK%�/xc�-P4"O,��Qʐ$oZ��ǡ�"JK��"O r�k-E��Z�#E?O��h"OF$�60[��A��
���b"O�]y0�F�V- �Cр[6v��4�S"O-�Ԡ��c��Ձ�G����A��"O��prm�I�BDB�'JZ=�(6"O���Ā�d��)e(E�.��a�"O���Y�7��i�O΁s֖�"O��!d��L*�}x@@�^/�C�"O"a*&�۷= ��k�\;
�<�a�"O�]�M1-�^l����Y��9D"O���˅�m~(h�5�N�B :�"O4�!߃,y�C#T�k\J��"O��w�D8� agZZfY�1"O<HX�f�dR���&01��=� "OB��e �w*�-2��@�e�|�Cw"Oty��cE�\�L5�+���ƴa�"O^9x��By�H��GغXѢ5��"O�=�6�]+�52 i!���"O�ͳ��$	 ���&I.K��U"O>�ۑ��1Z� "�5Ę� d"O`��B�@!{v�!�Ò\��"O<�8�ꊩ0j��_�]Kx�� "OP�I��Ĕ�Α�aџ~���#"OfE1���p��DAׂ����"O�-��e��kg D�A
�:9�p7"Or{���+ŀAk�	�*sLz`�V"O��Dg�$|�*Yd*�v���z"Opٓ� ��j�B슭�p���"O����m�	?�αб 
�P�D���"O��!�i���.t��Ę.9e�e"O�l�c�j��)��S�.Z�r!4��AbΟq�Ș��^lLxL�h8D���EB{�.$���9Zb|9C�#D�؋���q��h�ǧ5j�@<8Q�%D�(���؝r��8`�N��,vE0D����aշ1��dj���
3+�5�WD!D���q��l`$�[DfD�;���Cbl D��JDlG�R|�2�)l��b3%1D���э�&�5���g�I��#D�l�*(< F��`���=>f��h!D�|(�m٨P��Q�ҤD�oW�\;F�>D��`eH!t�
���m��
��p�?D�P��bN�C�2d�2g�>�D�9D�T��gAz���-�����I9D��R,O 9C���ȯ4��(�<D�(8��P#����1|T��ӄ&D�h��&��.:�"W�J�h��L%D�lA�ß��ԕ���_���S�o#D�� 4\�tfJIj)������B"O�|Xw�T�
:��UϾ�9D"Od%9f�	c��`D�f�Tp�g"O�=�El��<���cf]�.��-aQ"O��Oܙ+�C#��T�:�ن"O�Xu��r*�ɺ��""o�	�"Ob�ѐj�>�<8 �f��cl�g"O�L�`��GCX�H%,V*|I�B�"Ot1с�m1�uXX1Bޥ�.�j�<��	܍Ͱ`��I�K�V�@ q�<�ɈHP�T�wׇ"z�.�A�<�c�N�[Ө����9D����q�YD�<	�Bg���W�2L7� ��@�<Q�λ0IzHé.�z��BS�<ypCV�y���Ck�-_t��`$�LV�<�� I�Z��-���e -�]�<�,)RF��#,ƶr��U��ȓZ�<a��z�Ej �w_�k�Fb�<y�h�8[�{eܣL3� 4G�`�<�R�l��j���8>1(��@CQZ�<� !���ԑ��mX6���*/FL�<!���`��͠c�ů*&$�kC�A�<Q�
����ͻ�a�0l�N�S`�b�<bO���q�-�`@�Ua��ی�yRdݪ{���z1-T�Ze*iX��
3�y�M�f�  �/خ1��C�
@��y2���_�p�o�,��	[��y�݁1��B�I��nx`�d`��y�.T�Fh�����T���6K�y"��v�x�Ӂ���fI�B��y2DüM������S-ό<�uO�;�y��$��}Sᬀ�o�ڌa4#�y⩈/@g�-�G�mC�ȨP�
1�y"�:޸��&F�d}<]2@�Ǯ�y�N	X��ݢץ�UL�p��=�y(�l��������h3�ژL|C�/;�ؒ�'^�9��t�h\�H�B��8y[P(�����X���X���e�,B�ɗm�T́��QC!v؉p���s�"O��`IӬa�$48F�L�_� ���"OH|*!�?�Qi�4e��Qx!"O�۔�[1�ֽs1�'vq��#�"O^��@�T/X�;$�I�ڤ��"O�#��
5o�##��i��T+T"ONL�4���,��֏!���q�"Oli�M�"+ �3�gX��l��t"O
-c�WjB6����Y'Z��#"O�xK��Ƴ=g�)�EDC�M��"O�ݠ��74��D?JUbq�"O@�����i���6X<��� "O�,:U��� 9e�7����"O���b��N|�`��<<쐑"O��R�ԾX�͙3J��f��yQ1"O�9�EA?A�^<;c��o�
���"O(4���$ij�"�Y�b���"O հ��;WO�L��'� ����"O�pq)J�p�F�7�G��8`Y�"O�d�'� پ�z!D_7J�Z�(�"O�iӤ�1yRx��#��'P�Խ9�"O���JB��Ĉ�$��K�f"OP�	s�G�0�Z�z�[�MI�Pf"O� @�g=	Az S'���9:`䈦"O���&�G/�	S!@ ���ӂ"O|u:Շ_.����Q(
V~��P�"O� ���L�`�(���*q~=�c"O��c�.̋#�T����*�:,��"OZ� � ѝe���;�L9q��E��'��X".��y gd�j*�3s�1%�!��u.��ɗ1h6��PL�aZ!��y]��rg
P�e�ء
V=+!�d�,M �Z��֬����C�	!�Ē-L�Ċ�u7���\�2�!��b}�́%���d�h�	ΰ%�!�z�` ��CV<Z� d�E!7�!�$�5mSXT�E�p�"(1W�ǅ(�!�ĖL� r2m֬Q5��`ǠB�!�I~ -赣С =�qX I��!�D�%Y��Ʀ�_3�����_6X�!�DM/h}�-��*@
4l���B~~!򄗅g	P�1w��+$z<��ɝ�PyB�ڏ=��й������}i2Ŝ"�y�8�z���-9z�-)���yң΢dט�A��پZFNU9�f��y�G�7i��Cd�&~������y2�"�f��R/�)���5�_��y��E3r#xkGL�N��5x�A��y�o�(h�$�V쀐V���zA&H8�y�_�<`�u���|�J!떓�y��_(�TiR��"p�i���W�y��H&D8x��5e�2��h�y��U� �\����D��!I�yB��'r?
ZF#��a7zE� ��6�yA�
0uP���@_�g��d@7ď5�yr�N+ nЇii�M)�%��Py��߿^ft�A��0����&X]�<Å����|�U��4m�EH���W�<)�'C����2��űiQ��u�H�<���?v�-"��*?�T��� i�<q�� .%����& #c
�XS,�_�<�eHJ/&u�=�t�T�^9�L���`�<���3
��H" �=O��e���]�<�s��T���j$�I:_8�S�Rm�<��N$59c���l1k���e�<�(Ӟl�`��6sN�XiA*\�<�DɄ@��H�5a��oin鷭�T�<I�O rH���B��b�q�Q�<�ILD��, �q���8��I�<�E�]&4�Ƭ��,ҕe��8H�lKI�<��I�OR}0�m�KP�=P�Άp�<�nH&2��,�1h�U��Gf�<a���~1RY@���*6D���͒a�<Qfٵ
�I�pc8O���[�aT`�<���ւf�&t5c��q䎜��OY�<Y��E͎$:N�*j�p��HW�<��dX�G���2�b=D��qǓV�<q5��Y؄L!�,?G/�+�B�P�<a ��ti,x�V��8!��d�\s�<�AUܘT���25S����y�<y�\�"W�5��.&��!G�@L�<Y򁍁"�&	�Ꮐ/Jq�!���H�<�G�9a{Z����,7�����h�<9��=v�(�p���I�b9{���P�<��/F�cm�R�_#9j�izv�FG�<����}��̀�Y�<B,"&\@�<iWo�>�l"��@��@��KA�<���ONU����d���pt$�@�<ɥ�^/nH�؂Rn�D���W�x�<�Q�n|�ä(�6��e�V,�h�<� ��y�FEZ~dբ���k:J��"O
�y��	=q�P�&��36~���"O�=�Sj�cA`(�a��<'$��Ba"O|���Y� 604`qI Z>���"O^mymN�+�Z�g/��~X`�"O�Yk�e �~kA�MZJҺ؋A"O��ɲ�K����7
�5`���"O$��R�N��i�/���1"OR1��`1x�<,����4]dN��C"Ov�{5���%n,iG@�rQh�iD"Or���.Ǭ��ʐ�Jd�N���"O��z��[	s�R)�(��I��"Ox�x� u�	�0���:�h0[F"O����W 6��8�#��(���"O�`Jd�גslQ1k�k��m��"O����MU�J��@LHa<�'"Oب��HXh���aG����"Ox��ň���q�/Ϝc�Z�"O4=���;Rt��UΒl���e"O�es�F�.��M*�I�fT(aQ�"O`q��)z���S#��|���+W"O2��v,�~���"8M�2=�v"O��{s�%u��M0v�U�~�*��"O�����WTݫ���D��!�#"OV=Дdö�h��KC�l�na�"O���G�O�rtcc!�Q`@�"O����w�h0�2����)[#"O�5��ڳ?���̆�:�.<�5"OjQ��ב+�>��K�(®Qrd"O�H�K�u@$�b�4O�`�+�"O�e�͓�K��l��J(_(5�"O�e��F0S��.J�|0"OŘ3��>(���^
B�B"O.�Pu�\�n�HP���M RMl�6"Ot���Zy�d���Zi90��"O��#ßQ�T5zw�_�l7D<cR"O<q�Vn�|PdõlD0\8x&"OX�(`l��{�f�0a�)n���W"OR�sfI5MJ@�Xo�5�"O�ô�;)��4� ɟ~N�k�"OȬ��/d�x�(]�j��P�"O�P����~�l��b7Y�p�"ON9a�/�C��
��	2���v"Ol�[t�W�zе-�� �"O��Bw�G&v�$h�˙�6�*�G"O�QP��_�El&��c�P���=�"On�r�ɯ0X���Z�6��l�"O�  r�ĤзFʹW�<!�g"O<�)g��,N�Z�B��J"O��p���*:���ʜ5�D��1"Or�"敤@ana�R�O��e�6"O��r�O�Py�V��]�",��"OFU��N�*P�3B�=9�4m��"O�գ����;�f�+8Y����"OH9�(�[6�ru`>^:�P�"O�`�`�F�.i�l��'���sW"O !��L����VOߴ0ɚ�)F"O�0��\]��Aw�Q�9^x�pg"O\�i���$�LѱF�F���"O��`��6�Q�C��?o)�q�"O�� �$E,_?T�Aq�%<"|�ɤ"O�Lcr�W529^i��T�m�JL��"O�p�UE�F��puhܶQǂ��R"O��a��Aif=��'W01���{&"O� �AÈ&�d}��_�.�"��u"O���*E��T��N>V�B0"O(�㎴R%Z��#�޵cZ:��$"OX�yaB2B�lW!�35NR��"O� c���&p�d,��2O8p��"O@9��Z��	4��q#��Pe"O�q+e(�/Z|X�Ѳ!V�s�� 1�"O�]c��P�qͼe���\4#�X,� "OhkN� u���a��1m�F�"O^�3R�J�7�e�Q˘ R�9�"OtDJ+��7��K2
	����"O$嚧(�][P�Ȕ��aᾑ�"O���
�;kN����P
c��5Y%"Ott�ŀ��F:썘��S|j0�%"O�\�����=����ԇ�J]:-;�"Ov���"�$�nݒ��R#+�=�"O�����M���e-?�I"Ohl�"�NI�¦��L[�`p"O,ŨGI�B�dt���D>F�c"O���N)~uq��W�G���*5"O���G��Q�Ti%ۧe����"O�pD�/������>L��"O��@vl�v Τ���Ĥw����"O|���9Ph��ꅯ�"s����""OL�C��;P�q��"M���)�"O|Ó����s�O�*����A"O�gM��o;>}K�̖�_��6"OD�w��8gI>����*�f�8v"OD�[��	�^�k �TD�H��"O\(T�߫=r��q��� K�P���"O��ug�2�vL�T,��r�1�"OFH����9h�V�i�MJ
J��m�1"O��9cR7A𴠡��Qi�+�"O��PM�-d�,jdσ�@V(��"O�\rƈ�"/�Y���D��%�>�y�`٬��T��/�b�-� ��/�y����{��p�(J�	qp@�
ۦ�y���|�����ҁ�R�Kf�Z�y"*��~���`�-����r�Bΐ�yr��|���T�M� �U����y��I����6{�t´ߟ�y�c�}Y�|!�	�#_�Mp�@��y"c�z�a9 ��B�޴J4��y��UF��2/"p�Lږ���y��f���#E�Q8T�Jts6�Z=�y2K�"��yV�N7H���%Ő�yR��m{�dY4dI>�d�u�ã�y�o�H$��#�O��3��ʴ���y�e}Ii�i�)��ÏB�]Mt��i"7/)6�V�	r��67����i �b&J��$f\�)5��t�P!��_6?'}z07	�^'�x�M�o�<�"�iK��Y����D����rNe�<�Y0��R��d>T8S�`�<Te� 
B�"&�+lQ���!q�<!�N'Y�������4��DQ��w�<�JWI0�(��kTQ�0��CO_t�<��-�L��ҫ]V
��n�<���z��(j"�D�=�T9���i�<QV.�d%���(0�T����K�<��*@?M���4�/]������G�<B$�;<��3N���+��w�<�C<
Q6YSbnٹ͌�k�J�q�<��\�x��5�J1h�B�Cq�l����S�? ��e)� Q�r�P��Y�f�]ʡ"O�`��.ٝQ�,�#D�,�]×�'�"=��\!:�h�ŉ�ie�U��h�<�%a�2=��)AN�x4���q�d2�S�'o� ��(E�%C/�F�R�ȓGdB�b � ;���s�jI�\���&�\��	({֙Pb�"=ˬy8~������0`_�汐�m�&Wo��8�k(D��f	�j�6�W.�(q|��e�"D��U>*�d��7Ņ�B�,D)�&!D�X�F�
^�	˗�B�l�>�[3� D��FЊ1wNMR�' �1;��`� D�P�d�T8�H���"CL��1�!>D��*���5&|�#��#����SE)D��8���*y���0؎�`�'D�|2��آ)�2�K�i��,^���&D��2!��An�;�n�xH}� I$D�LxA�_8I���^�b@b�#D���5�Y1 �v]�6.�&p&��f�!D�dSD�K�(�j�)VX�X�!�!D�|ӤA�1{�S�@���V�Ka� D�$ڰ�5��E)���d�tq���>D���5g��{�jLJv({!R�ԏ=D�L@�Y�t߀DJi��X�J��pM:D����^�)
�l��fإa�����9D�@	6��(��e��+ֺ�̽#� 9D�l�E�Q-�"�#�@O�z\�8��3D�dB�Њ$������'�Ӑ�=D��E��(?����8"�.9�G7D�T��W�qž�+�	��<yf\Q9D���,�!M6.<�ԃҊg�`���-D�x�oO�=�(��2-էph|-3�)�� E{����)���6�P/7����W�Q�B�!��=\�8�����`���DߣBl���>)����\�`WO�l���FL����DU"F ˹lt����A��b\��� �� @��W.�ԉ�h@8B�����})I�R6���.�93y�y�њ�yRL����)�*@�b��m��h׃�y�&ǟ�*F�|����K�p�
ɣd�~7��H!��,��w�l<|��W�.G�	��
��\x��õ'�|�,9�nL�\�P	�&l%�O�ʥ2O �GBE���is�F!\��u"OM�cN�4V�� 4$<&e� �'0�O�tR3���u�#���(�"O��ڴ��QpVIa�B|��|y��OtT�����h������{�0��'��9��P��"Oh�I�ˑ�����7u�`�!��x�e8�O��1��ſx\�M�&���2� ���'�$M��nt���S�5�N��r��6�,C�I�[���X�&�	(WfϷ.�#?9��	?�85Y�e�+��\�C�
A�B�I�m?XX��L��V�
� ��9 ��s琣<E�d�޸~@굛!�A*dhr|@ӥ���y�ě8����͙a�Bp�".т��'��{�@C�5R���F	޹Q���9��T	�y��I*����䀖:�a��"U �y"�
6 0���7Z.l@�IŬ�y�H�2���qU+Y/ќh� +L��y�7"����B��3�`����y⤚�M�(�S��F)g&�2�a��y҆MN��Q�լ1񆀀�i��y�&^�c�4��]1�ۥ�@�y�V?V1�4mO(~E0�jP�I7�y
� գ�Ax(#�$T�h\u �"O.q���B-�̢�e֜:Y�"O��à��f�\e�d��=�(!1S"Oxy�$�H8 Kr(�(���D,b6"O�4)�B�x��x�M��f�K�"O�iۄ���6�!v�B�P��a�S"O҄����-=�E�T�]�G���Q�"O aڔ�Hj�Xe��ƍ/��D`&"Ox�y���$����\�R"O�]+'�!*�hM!��9�||b"O
&��!@�ɣ���
8�$��"O��pW�iŢ$��
�������"O��­w~�I���Pp*��"O.��n��uM��Ǌ%���"Or�RD�B�)�'���-i��2s"O�\�b�U�5	�be�^+Q�dPU"O:���FKAd�
 I�wK�4(�"O%+��T>�sR	#0\(�p�"O<m�gզ>��
s(_�D
�	�"Otq�
 !۪h�4h�@28L�p"O�𕏆&3�����ޑ\B6��G"O�`��[*/%��%h�L:�x"O����r��Q��f�X+f��"O� �L�?� d�֥�� �~�C�"O�j�DZtpd�%Ȓ�l�v"O^�h�V$1��Ē2e�}�ny�"Oيш�5g��p�C��t�p"�"Oz0)#F\�{�`�е�W=�\L��"Op��G�Ǽo
���+7��w"O�1 ��iD�q�W�ރ|*By۳"OȈB�
�1e>��	5��x��� "O`���䅟E���*glE!5u���"OD����3[�p�ϩ.��ا"Or�{eF	��� �$��%�t-t"OJ��$	�0oq�|(�.7x�n��U"O8��Ea�N�48:1�R��MZ�"O�����F6o� A�T)6�uR�"O�|�%N�ht��JǬӀ"Ę�$"O|Q�
ƶ;V�D��jV�8�L��"O�9X�%'>H=9�+���k�"O�8���A���s��D�3P�d7"Oܹ��D׭u� ��F�Z6?�=Hc"O~�4�X�?칀/F=B��H�A"O�`ӕ$�2-x��T�o  X"OY:���@L}Y�@S�҄1�"O�!Y�LWri	C /eɢ���"O$0� Ɩ�r2��#��ױ1��d�c"O|mS�]/	��x��D�f氵��"O��AȠ{�<	8�-^j4��y�"O�9ULG�k��8�M�9;�ju@"OB�yTjOu� #�'�{��ts�"O,�����.�Bp�c�Y�,�Թ:A"Oു&Lζj��ē�C4t��5"OT+����Ht�9kr̒K�V�H�"O�ܨf�F�5(6��2-L�:�~��
Iæ��ݴ_���0�G�gr�'�b�'��֝ݟ�NA��$��$�C�~8(���Th�3��_N�Ѵ-ÚD��h �J�?���]�y��O<3��0O�h�#w��\�� *�HšQJ	CծԸr�"���	;T��S�A�.1r��|���0�S�J��U�
���$@�q�"�b�F�$����ן|�'a�x�P�@�|��jQ��E�ҝ{K��D{��Ĵiz�]I�IO�#=�}а�R�j��񠥇��)�4�����'����+l�}I�A/P���;��� unB$�E�k��d�O�$�O��-FX��'e�5��󳂓837��P�@� VZ8��D6D|��J 	NE����C8iJ��2���A�H\|9Ka#ď`���ŀ��K���2�7;i��r���m,�x�'lӎŋ���<X<��0HP]�WlU�~����H�O@K$զ���Vy2�'��O�3� ���@+[Ҭ�XA�ĸC�M���Ox��$O�MR�i�F�5L$��Lإ8i�$�0��m�oyr��s�x�ݟT��t��ֳQ��I�,����jŭ4q8�W��O��O 0P@͹L5>q@����8�f	;�j��윫�%#ZU����G+1��J��X�_3Q��&�Y:J:0�'aK�uvK��"lV�1�ve�"`0p�bAG�]�`�R%�.9Q�t�c�O�n����'�M�C퀲p6n�a�J#6��X�� �;+����O�s���L͆DsDJX��0���>���4�,Un%�M޴\��yv��- ��)�I:	<�e�}��1�$�i�2�'��S�%�5�IڟLoZ�Akf��f�zx��2'��~4셑ĂK�X?V!9!����r��r� j������&ט c�>Ex��,�x�����x�7��<:\u��,��%�͡3� }��%�%���5�bM�#�4�Ôi����xa��MT����0�4b��("|n�UR��'�����9m�1I��?qH>��d� V��Z�L�?@R���ŕ�3�qOz���z�4����阒v"@�'��f	@\�Ǣ�u�$�$�O�]��C$F!(�d�O����O||�O���:=�J�A�J�<Ar�T�GZz����ɒ8ĖU���7rՆ��"�H��@�//�'� �j�Jڃiu�=��O�n���)Q���(�f� &4$�%'����)�։K>i�j�#=�j�qd�A������/@�����G(B(�O�t�����Ol�ec&FL�3�@y���{M�Y��*]�i��Μ:~*G@�6"�P��"*}���m�\yr�'���O剀����Q"l��T�C�U�p��+�E���P����`�3�����I�ܛ�
��(�ޡ�5��&vn`�bt&�#v��eہ��7M�2�$ »t(�K4R+)���<�`L�,]��9��&^
U��2U��#�����qn(%���W2S	�%@��R�~A&�<�7d��4��CF�S�����=�	"R���d`�O<���?Q�*��%r1���\��5Y7��$&X�#6�O,�Fz�S�e��Y��:}~��:#t6�	�M�1�i��'��'�'T�X�� ��      Ĵ���	��Z��wiD�:\���dC}"�ײK*<ac�ʄ��iZ�Fm��x�G��;�6Y4�8�B ;>��l�{���Q�
2)&�m��M3��_�x�뎄
7#"��	�p�&,�	����toA��ԽA�1!a���ǟ*�@�QY�����x<&�[H���6��/kVAʷ V�*������Q1$*� �P�����>+<��NfqO`�pL�̒u�z�廱/<rAs&��z�6<	�.�~�I�c�HQ�aOj�S� VE�҈Y�1~j%)�,UF4̓GA	��)�O�	��M��.0�O@|I!�,�LQ�Ii��ġ��g��	�H5��5���.3F �g�=1����-1��Sza�M�(�PD
�'Lu���S�����Y�J�P}�L��;c��7�J�OH�cԎ�;��@��Cf ْ2�Ôn:X�x��_�j�THpH>���P�d(�'G�83ၭj�hXڔ��dIЭC��F@���c�	V �-�5�&��P��j��fE�->����:lw2��1�ķ��;ب�0��q�ɖ9��x0�d�n�3�9)���a��.�%J�?�6�'<����ދ����QfN�^�$ŘkxȈbIK	'�0���`��B�R�0����O
��cJL2��'��eC�'��,��]�*���$ ب/�6-'��I���)���OX�e���$Y5%>���f����Zv�Ɩ���'-�ԁ,<��ΈG���(G�|��Ҟw��M��%�1H�D tkl#���owӸ�I�?��j�� �b����g�"�-�)!����/uʹ��^�N��M�Y��A��0%�>`���h�4�Y�$zByA��O� S�ʂO��1:0�5�xdSE[�ࡪ�9���O���&#1Չ'�HY�`S%r�f���Rzx�*bHBP!�M>i䈦`@&U�<)2���hd|�ssM�+��Ȉ$e��E�_X�<	B.� 2  �@����K<	�ԣ%��݋O|�b���MX,�b�-�a+�����.=E�Y�/L�II�~�2���:�'���ҡ�A}�c�68h-�wB߲J�X���_��z�䏑KHjm"��|r�-BJ�L>)$�ډN����'
[y?�TѴ�ڮ ����dT�8���I���+�n�W?�>O>�r��2�?i` �Ft�(�%3d@"�^~�O�+7��(N>�0�O3Z�ȥO���̯;�ʙ��D˿���j�E��Ll�,   �  /  �!  ,  H2  �8  �>  'E  �K  �Q   Ĵ���	����Zv����P��a+zX��M�!r�V�CB�{�`�@-7��!:7�� 2d01G]G��{u�+TR�S�тrF�[BR�l6��Q���q����9tNqZ�� 	��A�;���L�����OT&+�R���VY�ّT)[��f=�r�$ow@y���C��5���О5k��g`�uaL��vL�M����D��( �Hy��s��J�^��Q �?�\THU ��=]�L:�(~Ӹ�㡃�&�|�c�k��9������)$J�E���%��=R�h�1C�_�|�\�x��'�B�'bj�U�	>S�ొa�V$14�S����9�y�?/T��� %��G뤔+����4���I<�҄H n�za�. �3�"��#�J�m(�se�[�G�4t!�ȏ�,&v��OirCcy�L�e�p�A<��EϚ&�:�py@ �	ϟ ��R����4��*�� $�����iz��D1�y�i�r� �y�.�/���%�ċ�M˷�i>��	iy")���<�@�[���*2ʈm��Ȋ4���$�O����O橭;�?�����,RM���@iJ�&�E¥"��$P�ï˔xB�,!�dT,uOV��Q#��d�DyR�KL-:�Y�B�+:�T����A��I��o�$L�Pi�CW�ɠ��М��@�CG�V�'��H��=T�U;��F�X8 � M�Cy��Ӳi"=�����Hw�"�IŰk�a�䠏G2ay"��1�n�#a&˻qĒ��SE1}��L��V�'�i��x�ȼ~j������ڿ(z��0�[�o)�E��2�M[��?���?���(� �qgH&S���͇�V,����&i��)��B,S�����)�%c��GyBL�]��Q��ƽi�0Qp�o�8X��P2EK�;b�a����I(�����Kd�n,�c�W�M,�'�h,���a.��L%�))�*Xxt	ӭEIfah�Цl ���p?��Ie��)2I�+�z�ɔUI�	e���$D0?��m� 6t�I���À���HXB}�I�]<�7-�OP��|�ԍ˱�?��Q�<�yŮCne����R�U�y)w�i�xɉSK� H�������LX4ן�c>�c�
er�U ��R�I"����)e`�W�@Q`Ԣ�j�#��H�P�z�K0T}:�)�E&ZԔrC��OjC��'�"������'�XۢŇd��3�Cӗ+���"�'32���� D�����#]<+/��2��dHN�Ofl ����H�pI�SSĉ��xӀ�d�O`,�B���x�$�OP��O�8���?�C���ݸ`	ţƜ�zŠs��S�P�2�dh�jZ�����X>�ъ��4eh<JRE�z�����e�|0@ �9;T<U�$o\�	$5�*�2��?�*BH5qШ��:��U�q��{y��A#�?��hOl��9�ݹ0eU,iĴ��x�C�; �����^7��ܢ�JĥJ �7��l�����'���DAzdb�bG�(�yjSM�/�Z�pION~����@�I���^w r�'��i
>�`���F�9�0y�K�n� ���Ӻ��թ���'�N�AŬ�k������Ժ�`m�` 	�(n$=j�e*�|	����6������߸l�	�n+N�z���D���2��3J�$1J��
[xsF���x7�@�'�Q�l�e�[�>i0��Q�= ��h��#D��&j�8���P 1�e�¶>�ӺibT�Ty�b	�����O���\}�	��W�~Q�T��F���6-����$�O�Ĝ�.�@KR����h �u�˿] ����ױKg�p���"n�0`�Vh� �`\�i��Y�@�]���jC�V�p���2"�m�H3� 7�������H|�`R�� O�'x
��ƛ�'��Bi��ZE�D�VSrk��g��ꓳp?ѐ�E���Ļ2D/@\ĈDNNX�Ds�O^l��e��̬/e��ఃnq�'��Y�'>��'0�'������HЂNB
y���V�߀<�L���C�"�M�!
��vtk���B��ȖJЙ'��b�J�$��O����E�Ȓ�4Š���S�2�#t�'tV���^�=�ʘ���2k�.U"D��"��}�}"��.ZK���R�еW��E#�e�?����ӟ<jݴD��)�I8��ю#*��Ð�(O�h��OI��yR��pR��cH
�/���E·�HO�YE���)��r�i��Ω�'G@�a7��O��dY��	Qt��O��d�O������{�h�(T�6mέQ��IP,�H�ⱡVO@�2��ځ[�`��.��P��S)\f���x��N�&�H�3��
6
ή�k�@=EĮ�B!(��9���,�%� 2/�,k���w�P�be.�(kBA�K�v�'X��0�y>��8ғ�~2KQqq��IU��[N��R�@��yk�;�D���aH[9, 1`��M���i>���\y�莙]�y���-;�q�Bf �]�*#�Ύ�%��'@�'M&֝��0�Iȟĳ�*U>L|RBA?j�XH2%�U�UQ�B�- 4�LŎ 9�Tx�\�AB(�<	�b̥7R��3�LZ1:�&-�F�2X����7h�+CҺ9��L	]t�� K�:��ǋ���J�:��	�
�Z�`����;8��$%��K$�ȠݴTR�V�'1��ǟ�?�O�=��g�L���M��2��$b޴��Ol�<�$џP�L �тgŚ�6�i}�˅��6-�<Q0�ŵd��O��d�?&�4.����8X6�d"u�}�ld����Oz���O��RS�m�0:�	�F�D�-V�5��� \�>Ե鵯��]�(�����Q���)��	1
-��Ιk38���CJ� �(� Z�`� �VLvk��Q������NV}Y��|�.��?є�iU�b>u3酖-^���2��,��T�>i
��0��Cf"8)�萇%�|�ʱ$��E{�O.��B��Aj��,��$��M�e�>0�''�U��i�����O�˧kt�����?	�bU<,E���R'��M��% AL�402���,94|�Q��'UP�'�J0B>@�hB��'8�1��	E��OLR����ΆY�R9�c��OԥXW�ȡm�"쨧��(Ԡ��s�
8�����+�`i@���ȥTY�@1�IZ
c��fԟ�?���i>�S�SU����33pI��+v ��0����!�$�Qo�Q�R��Z|0-�@�	�DױO$��J���$ꍲ���b�ղe��d��K 82��6m�O��$�I��1f�Od���Or�d������_����@A�G��PC��8`��:�!`a�tsg-±I%���`�:t�哮��1�đxr�D)A �M�%R� J��@I��k'���;0`��8z�,���'o�BN
�"�|� �C�%4&(���m��s[��;r��<�P�O��L������?y�OF܄[�g�4O��{���n����'�5��H�#8�)`��bN�;Ъj��Fz�O"�W�@H� �� 
f�eG��x���F$(����韄�	���I�?��	���ΧoG�)iaf��bmԅ���E�t
8���Ú�un�D*�ė�Wa�1�̈́X?ni "ʓhb��/E�B$C��fGpEb �����t���ҝu�??��H*Q�mP�@��P�ɜlP
��	�R?X��m07cd,"DD�Nd�$lZ����?!���i��)ŧF�3�B�� !��/.���˓�(OR�enXp��mA��7n��dY�|�۴�?+O`a��_�T�'��I÷i��Q�iI.?��њ�B�@q���� �2�'�ID�V�"q�.ߚvy�4,$�:h�R�7��a0M�m��Ea��Ga1�(J���G�X:T`���G�
�`�M�[P��8ZqY�̮6C�\�K-�f�*bF�o�TSH>RFY͟t��w�':,hQp�P��%�L�~e�|3��>���p>�$�;ex�9@��A6`�`e�i�	`����:?1���2v��C*�%VL���\}�*��A�,7��O"��|�0n���?!�
�Voҩ7���s�� KR�\�A�i�d�[��'|1O�3��˴�[E���i;�I�Kǯ�����c�"~�BO��鐥�(6UjDHԈ� �?�t�ߟ��K>E��I������\\�( ��DEY!�dNS����P+],}\)p�Q�3m��`����T(g���7l@0F̭x�Ӑn붴m��	��谁�֟0��؟���!�u��5vJY�`���
"O�R0 {��I�v�x�{����4�,i���DO>@:,�t�0��ē]2t����\�*���=L~h��v%K<��  ���3_��D�� 
D��@�e���'����T� v��&�8$e�iע�<��c���;�k��<r�*	>]>� `M��P�D���:� ��R��?�Ѩ4*
�"-F�nڛ�HO�;���+a�<�㕡�]��Z�&��Ir^�X%���m����O$���Op|�;�?i���䆘�(���%@Z�(�� ,�3S%��Y�X��$h	�O�&���ƀ)P]Ey���)���q�Q?��*&aN Sᬩ֥�N�`��6��Kw2ЁFעZ4d�Dy2#��?yeՌ@z]��%��~wT��#J�\a��/ғ�O0��u��#3�֤)l;.���'`Q�<#�����CiU*p��U҆��>1"�i��_�j�������O��S�p6(q��� 1P9�$��Y�7M˰s����O��d �B�D�J2%4�p{Eo>�M��f������]�[^��a�,A '�G{R(���4��Z�S/�|�JH��&��@A�q: @JS�'J©���қ'"��
c,�̑�n�| ��;����p?�r�Ν	_~,�f�ۥ.T8p����\X���O�mk�+*|L��"��ÞYuF�{4V�`�*Z*�M����?a*� ���G�O���ͯ����e�0B�ћ
Йoڝ`^l�j#e��qht�� ��#IK���ǫ6O�e�|"D+�;n�^�Ce�:+�D�B#���?��Ș� "�����C	Q��H�-Y�\��
�&��+p�qr�#�,;�l��o�
Qd��ɦ;��Ҧ��)O�O���|�<Tqʆ� ıyu�I����ȓ}��X�#��;D�Q�P���;<�0�>���Ss���+^DաG��g����@�\*~���4�?���w@q�P�Ɏ�?Y��?������OL����r& ���g��%�09C�QD�<hp4��ft�M���t��;���bT�Kz6�&�H��?W����K϶pf�Q%*�	?u:FGӽh���S`Ɲa���'M�~Ӳ�Q�#T9C�'w�D@��{J�$Hs.���*O�!q�'�h6m�d�矘�Ih?I��VwJ�YbA3Or��h}2�)§X-��Ȃ䟲e�M�E��@h���iQn7��Ȧ]'����?Q�'���B%��"Ρ���Ͳ7%�dSi!j����'�2�'�-s�A������';�z��G���@�\4"�'� �*���挜>����9�E���,���4�����:FX��뛕qR�У�B�]�
	z���Q�l����6/x)�6.�: gQ��pF�O|�� `iڤ��/$P�-R�) &B�T�kf�i�"=���D�y�D���ȣ_b҈�+E3�ay��� �A�H�y��s1��4|�T�����'��� K*64��4�?�����,� 5��{�ͅ�_c d�VgΉ�M��Ӂ�?����?�AT-ԝX��ߘ���'��/�B�Pr�[<N�6(��
���x����!d}Fy¥�<|�ҌP��N5*�|����̡3t�}B7�Ӹ;������=R���*3+�3jo�5Fy��^��?���SF���&冎Y�DU;#NT�_��C�fE�*TEѾzG�}SDKV�	����dIS~���+�rl��b�&;R���?���@
]�l���	~�t���B�'ڮ��CjU�p;�89&#���Rt�R�h�h���K��P��>X.��B@��1����j&��*T?��KS�Z�8�(�`E@�����I(�`E� nFI�Cn�aJJ:@
�q�̕q0h��!w<(%$r��P�cf�O�(�'��O?�A�e��..�xe�;q���a��E�<	�I��R���o̜u�pYi䬙V��?�Q�i>�s�ӧe�Lc���m���L��M��?��F-s"��A���?����?�b������ ˕���p����$�� {8A��_�,�>�Ov0q��!vߦd��/M&:���P�`�Q'�O*U��
�`�����^�\yj�_�����Oj���	�L�eA�-A[�a��Q�S5,C��O�0����l�jG�R�}�7��Y�����|�/~]2}�Lބw6 �C���B���J_.3�"�'���'�ם�<���|�c�&t����d�A>LK
!3�N<��)^�,�:����R"�έ�p��h�'^tp�G@מ|�!�d��I����C�ĝ|��L�dD�|1��Vk��
�џ�{3��Ob��C�%�~!2�J�4)���6H�˦�	n��h���U�  *	[!�ȡc4���T/�y�CɄB��|2j��$@�GE���LΦy��By�Dͦ<�p꧔?��O���3���2_�%QV��}����ٴ^XX���?���}h���F�07��Z�k��1����t5�J�R���.=�II��X�
�pV�#�J�R���pL\�*ܦ;V^��'=�da�g�[<THkDàr��}E{�%ϸ�?����O�4�ud�.w����%*J�3��0�O^�D,�O6�XdD.\T��2��
5MR���'�d�Uw.da��^>ZB��ÃlpF�'n��K�Jl�(�$�O�ʧ��Ѩ��?�����t��	���$b�V���!ĊL˛�O�8e�T��j�q� A��W��3Sg �~�1�*�;�� �G�L!�%!��|��3E��O�,�̔�H}�Y��M�b��%:E��Gڞ����t��(z��85��<�~�3��*w����?�7�|��I'	�����,6� #��-A��C�ɺs¼"���'XPD��C�!��"=����0����C��
�*P�!�Q	]��(��4�?a�D$p��ĝ��?����?���:��Ok��Qll=U�\�a���`��?)�L���3e=�u�6�ޝ+ Ț�X>II�锾L�'m� ��'K4
m� �1�)4��G`�C�����+�,sB�&��i� d|jI<I�.�/q~��A�GP 9I��by�NW8�?A��'�t�Q ��s�.�j#IC,�Hd0�'d�\�a�݊�$�fIo�I8�4tΑ��J�ɷUUDd����f�ڽ�uOW$C{��h�>? �	�����۟qZwJb�'��iK�?#�� EbU0�h�Z"��

�`r6&Q�YS@di�lJ5BR�`��=g�����T�X7@�hP�FFH��Ǐ5.��UzǊ�3!|�rb�-p����־w�Zd@��DE'�

�,�f}H0`�kT�EL5P�B�I�<��Qz��VFW�	��5i&2C�ɿ>�9�`��9׬���ٛV���t��f�|���-?�6��O����?Nk���m�==V�l�����B��6횆s֪���OT��ލ3Kfi�doW#k7z\�wKU�8}0sb�r�ű�b�;m��A$���@ԅ���	pr�!ƀL" >���&@9��!OR��`�Ovޝ
0�:��̊��	�z<��U�O��@����is~��\$TMKphD�<)�@�j��:g.��9߸PH���IX��Z�O�����8<Dx�q�H���,X���d�2͸�4�?�����)Ј~76���O�h��F
�=Ц�
aǢ�CQ$]��!�'�̩�t��#N�MAL��S�K��t�L-zW1�`Qx%$N��}�u$èq�a:���O쭁g�X+K(�b�P<2�4�y�N�Z��K�7�rt��-?Z�;�/ǖY��G�?�ǐ|����8�T�`��π,�&�Pt���>�C�	+,������d�R��a�T�>�p#=q�S�#?��ӣ�N,�����IzT��4�?���)���+�?9��?���?���Ok�D�y�������oF�rG$^(��ؚ7�R�	6�x�Ɨ�@"��+]>e�cW�h��'L�"���DȮ?�����1�P�����x\Pˀ#����O2�K<Q�^H����Ξo���" KFy��8�?	���� ��� �>�ƨt�I�P�R"O����D��:��DKV.�>�)¼i�h#=�'��."d�J�� �bHC��#P�ꜩtT�ϐ����?A���?��������O����`o.$�FR?/>��@iٓ ����`â���'���2�X1+1K?�x�剑n�x1�!!1 h!��Q��;�EN!��LÃ��6����-�)A>�����)a��&����O�On�"ƭ�_������Jr�ؓ��	#ٴ�?�(O���3�i>U#�L����7��4jX�P%�,����'�Q��+�IX�d�X��I�:2 ��	�>��i~�6ʹ<���A8��F�'�ݟ�h�A2(��$�ƠP��r�ix����'��'>20BS�W+�PRU�z�(��v%F#e�-����/JҜ+�E�YG�U�w&��(Ol,���^6%4(R�,��Y*6��D!��^)>�	���9�\����E�O�G�(��#��O
�E�T�4Ar��E$1Vo`��7L�7�y��&D@���R*D)UT:�𦈛���>�����FA�A�h�a�^�P��|�q��>!�G�'����'��U>��������	yԎ� A��zh����"56yh�4\E��rT��I���Ӏ"�.&(|�rv��.O��h��$����}R⨜$eоuQ#DٯE����<��*e�߆.L}�v�ڛ,>��qNܧ?ݤ)�`�H�:�Mb�O���9K����,�Ɇ��S�Oh�(Ǭ��xs��/0�v"O��a�`��wP��AO�F/������ȟ<�ժS�0���2#��t��%�� �撚�I��[G��^_���埀�����C^wbZc�:(ɖ�X)26�3��KuJ�У�^�dM3r㏾:����G��iD��T�I<��^E�\D�B"j�@�`��Q�˼,i�����	)��\�O�n ��h�]�	��P4Gą&\�Y����?�ʓ�pe��8�0=�V,,$� ��d�r2$i�ńCH<y ������%xx$�#̳2[���=��|O>�P x2�ǏNڰ4"�`A>(0�����?i���?�mM��ON��i>aq��W�7�Z��aTm�)��f
%��٩we^S{���à��jn� �L�M9Q�`�W�R�d�X@��Y~2�:2��R�$$���	&?e.����)or�Q&�QQ���e�O>�x��ؗ�n(�4�ͅyN�P$��k�<y eK�?���!�+ia��tPd�<I�)^4G������1|XZ�y���i}bIyӾ�O�`�����U�	埜�'|o�Ӓ�_�,�\�a��?�Tn��H?z��I�����i����æyy���Ŏ�o$��gɁ.|�r�ް�p)�"M冠�F�0ʓNօ���-��Hf$���lx���\���q�j�&6��	��EϞ�yQ-,���Ʉ�����p�+h�>��gGku�Ĉ�"O~�a+��y0�  �5:m�����'�$��\phB�K�B��@��EM 8�'��P�l���D�O�ʧ��0��?q�A�$>� ��(LǢ2$dD�@��Ʀ)5��Td/T<e�J(H�I
�2 -"f�1��]Q�D@^D8�E+K�n���!#��O����CJ�~��-��R�P��*��Ў�$��\qX1 C��xF�8i�8�b�?�S�|��)΢Q�(83Q��"6-�unǀ�^C䉖O2@|�aj�6?;@�9i��"7#=A���i�U2�\2��wcP�t�D��4�?Y��'h��&��?����?���7�n�Ok�ӰR`�Q�v�@�󥦈��<h����|^9X5˝�ޞY��$
6�	�@:��� �yT���,t�
uvźV�5p���D	}������Rg����g��Z�}x5�,D���5�a�f!�$��1ḄЅ/�Ϧ��4�d�O�Q����n�}H���6
��qDg�ĩ#���O ���O`�ćO���'D(OG�8�`�1��Q�#L8i���:D�D䁡 �9��;bɋePF~��?5(]����	C��Pc�I&u[b1��-��W-@I�M=�ܨ��:^��"=�EG�����6�I Z�F��ė(��I��-�@���9�4�?q-OP���?Q����s��Z/l�S��f.z݀��B�	H!���
W�t$Z6a��e�h�u@�s!�f�'�R6M�˦a��)�Ms�LO�Gi�	�&��vG�!9���ڦQr��8Q4Ղ1�K�-MD����/D����g��Dl���P�o�N��wC.D�`��A�=f2�x��@�"�Р���9D�|�u�O�8��4��B��u|�ps�*%D��b���=,Rk_�M�^��A$D��ӦF�R��vGޢE��=r��!D����9C�D�(B��/)���A� D�h��ۘ>�p����ąg�\1�TE2D�t;Qo�&��P#��(z�t���'1D�8�!+ˋP�x�ǮQ?P��a(�`0D�� V}R�g�5��,ɡ�MW]L �"Oh�u*�B�؃&Ώ�R4P�1"O-jšN�5�hA��
��1�<(�P"O���%�X-|��&l�,J��8�"O����OQ*L!t�i���<:q�͠q"O�q����;����&Elꐐ�"OFe���]�D<
 ̃�W�V��P"O`�`R��R��1���"q��y��"Od�#��L.���ʃLL����"OZ�)������"�h�J��'"O���d�0�_F�����"O���BC�#���;S�L'-:.X�$"O^���EP�� �c6@?h24�"O����a\Vd�Z6g]�c�����"ON�w'O�*�~��X�d��h�"Ox��3�N�)G��,ʌ/y�]��"O
��b��"�
ȣ ��;`�l��"O̐:c�ה4^���ԣO@���"OB�t��=�\a�a�ԑXB� 2"O��r�&J�4���3�����X8��"OV!�DKK�:l�9d��$8��B"OB3$�;�X �Ď2�p9d"O���p���h������B�.��3"O��F@S�,�F\Z��_�tIl���"O~%з!EOd����a�r��"OԄ��C����T� hZ	t2v�%"O�@BP/�<���值*~��p"O�����)�lA�"�Y�r1��"O�ŋu�W�:u%�R�c$�k"Oҝ����,A<��j׼0��-��"O�����n k鞇i.��ـ"O����Q�Yێ��p��Fڱ!�"Of�ơP��2ΙN�J�"O�|ai ��,�zV慣?���;�"O>a���>Q���D�0"O���?��Q�� �K��|��"OXH�D�|��=�uՋtΪ�с"Ov�x�K���lBZɠ@��"O���G�ߡg)�� b�h-�$"O�+���`)
`AO�	aɠ"OZ�+�+=V"0�P� �_:���q"O���i#zTh���d
|��"O�ź���F���B+||��"O��A5�U%�������8Y$�0@�"ORx�'�H�I�TTڧ�̀l�02g"Oh��Ň�LB��0Gb��#�"O�� gZ{/��$
	����"O��cd"z�L؉%	�7G��B"O�X��D�d�0�~���8�"Oڝ��(%M�q�M�/&�#4"O�i��E �p9�禄�3, U��"O�y����JI�)ve �W��I��"OA��.Bx%�u񋒫]Ʃ�"OPd�#8�,2���5�����"O����Ôl9XYCD�M�H:�"Onp��O q��u�SfS�B���"O0L'���L(�e�7w��%"O0�P@ÍM�(��X����� "O�U@/��7�X9p�'��<�\�5"O$͹���C`���7{�'"O���!X�\�X@�F��Ll��`@*O�bbT�G�l���5]+� �'Nx(��5\��p�G�)VE��'��e	�"��m)l0��?�=C��� �5z@ �D@��b4�4`dN1[�"O���f�VR�<�P=cN<-C`"O�ѳ�H��'	���[���"O,��g�  t) �3eE� �"O�� �ӛ8ƶ��AA����s�"O�\�2���A
G9��`C�"On�xfk,�v�=���X�"O��q��,1�A���K��̳�"Of�� `��V9
��N�Q5�(x�"O���V�d���Eʆs6ܡ�"O\I(`@Є>��Y�)Փ?-�h��"O�-2���$�%��	�/)la�Q"O�i�w�B`����(U5t�$��"O������n,���L����%"O�Y����;�T��,���5aw"O�5Rg)�I�0��Ƶ��"Od�@�D8౧�	�����"O�]�q��3M�$�3T �Q�B�a�"O0%G�T�$�6�cV ��m�"O��Yǡ@Y-���D@�zЬњC"O�!�JU�0���;ʛ+I¨ip�"O�y���H����$N|���"O�9��&�pm@p���M::V"O�P���Q52��A��0^"Ѐ�"O�Bfb^�;��d:ĆЮGA�Xs�"O耩��K2j��]�uHPh���XS"O��J��O�)�����ɦ�4=(t"Ot�*���,b�n�p��=񰩪�"O�Eh�N�MGd��C'A����"O&��(N�oO��*�T3B��`KG"O$caQ�G���`�V��Ek�"O4�TH��I���-J���)s*O���W�Ή[�+�5�6]8�MX�<)%�P���jh�!eJ���P�<�!��^|"�+D�*���ҭs�<)P�Q�#� 1`�(�%:�qT@�J�<if&Qr�x ʆ��J�VY1N�F�<A��.yDHY�Gd\�62։�K�W�<� =@6�0���T9YTٳu��P�<9qǜ)NL��uQ0m��	��A�g�<���� �p�uN��v`5Hi�<�R�ڼU�*ڱa&5΄*&&�j�<aG,͹�����/HT� �jF|�<0$��z�2���%;$����1cFt�<Ѡ��iE����`�@�����JN�<9�Di��C���As���b�BM�<!5B_��UqgD8k��T�'��F�<�!�2��9�J�*p��̰Ɓ\g�<�'f��!,0�vi���y(�fl�<�NG�qjV̪���+ ���`��O�<�`茧E�릥�;�={ �q�<��N�-I
R� )[��Hy�%�s�<ǠC� ��U31�ߘ ��Q���s�<Id̃Z�� I�;�2l�"� H�<����5%(��FP=�:�*5n�G�<y!�G<\Z��˕?XQH��siP@�<ym�w�.��e��:X��Z��c�<q��@���Rm�k@�l�4.Uu�<���Ďڢ����������[�<���TJ�S&��"k �tڦ[�<�Ň�[�P,*rh��@�J����U�<�A�%B]xP����Ƕ��n�g�<�`͉1d%��0�	�%mFh�RS��k�<����a��mˤ�N�9M�8k���f�<� �1s.	�z�v��C�$/3���"O>�cp���l�s�Q
����"O�@ۆg�x�pH״P&L��e"O�ꗯՍQz�z�E�J����"O�5�E-7��eG�H�M�C"Ov�A%�X	����M�j:9��'�<�X"	�2C�a��ђ.ބ�	�'�*<�AGN�N�>�E��<&���'Vn���J�)@���a�j�8%�*��'. ���ֹ=�����e\" �z�j�'���(dBZ+7ZU�kEG��M[�'A$}�铠}6U�ɔ3D�4U�	�'����n���=x��#uPy"�'�`��@�����6���;�''�l��G�dG����\*{H���'�����0S+]�T�u�b8s�'�$�t���-�����ό���'�H�d,8C��&� &���)�'���9A���`�"l�)F%X"�P
�'�l둅D9�X,H<}�"Q
�'8�(:�E�aHf0��¨rv���'EF	�&+X;mu�"ƳpE�ȓ?�F�!@�,4��l(s���5� �ȓUI�2$���aW0X��E*9R��ȓt���`�H�.�a��Q#�+"O(��B蚊d7*��GC�^\T�V"Ob�$LD�
�:-yS� "'�Pҡ"O�]�4${���0��\�!�,\a�"O,��\�Qy��A� ��M p"O@�Z�%@V�D���v�I�"O�h������Mcg+(4>��)�"O"5��'M�Vj=(�F0P�2 ��"Ol��"�[_�=��M��-�a!�"O��uꍖI*�U�-߀^&��"O�X`e��
�s�%�m�`���"OP��/�)�J��2Eί,�XLk@"O�H��D�>�� ���L����s"O��R�M� ,� رBo�5:��""OH�[d�ohpIKam�dEj���"O"䘓�$,޲C`G�tH�B�"O�xAL�A�b0�Ӎ�tX��S�"O���̌��N���ķ&c���"O"�����.,d"�r��2^Nm�d"Ox��q(�<G�Dm�WM�,qI�<
�"O.�9u�~P1cI��&�2"O2D��k@�(d���w$�1����"OZ���@�
�h�3mٺf����"O�} �LX<NN�TH#L^#v��q["O�����[{�a��(:~�*1��"O���%#�o�!x�P8F�f�"O�(���	/ĸ��ƠEb!iw"O�ģ�."]��d�Q!	��w"OZUZQ�ЄNZ�6Ŗ/��E5"Oz�!Ɯ�W�<��+��
Ӵ0!�"O�lyt�װ!�d	�H�K�P��"OLQB�݁�6���M���$"O,!Rc \|�epr�E�!�P"O��je`]�V��lU���|q�I;#��4��fϰG�z�u��s��7�cV�qa�[�2�����ˍ-!�F�*�XU3��Z��Pr�ŗ`�!��% D)�G�T�>�>�2s��k�!򤚊$[��r�
T�C�p`�燄;Q!�DY/>���۳%H+QwN5�gY�.E!�d����a���g��uy�%�e3!�� �e n�s@��4���pL��a"O��'���X�P.�Rdf�s"On����>@	�L�`p#%"O���r��Kg0���j7B�@�%"O<����0Zz�dZ����k����"OA��#{���1b�!	�"O֝���P�g��PiQ��_X�`�e"O�ܩ��L){�]�@(Ew�<�b�"O0���`M�`ӜI��DO�}�<�!3"Ot�Qg��mh�8eL�w$��"O�	�������X�ƝUa\IQ"OB�y`Z�	d�A�'%�~8����"O`ْb��(bn�����R�� �"Ol\�]#Q�=��
�*��W"O��al�|,�c�k�&��P"Oz����P���	����D",�c"OZQrF�~{�Y�ȕ>M5���p"O�Djǡ�+
�@��(�<\�n��"O
�H��ה��B'ZU;$�!p"O��H0�D�hh$I���|5�D"O<� �L6��bFϾ8�2��0"O0����#� ���dHV�C"O6���-+C�Ub�Y&PQ ��"O�ั�p/LD����4Q긹�"O�P��Nffp0���*6C�t"O�8K�o)i�N4��c�7�5K�"O��h�W=��㡋V,4�U"O\qt��uw�}*5��i���2"O,�J��;��A�v�M �hن"O��tk�6u(��B�J��Ъ�"O�	�E��'J31D��=�9ZS"O��F��.Nt$�t�Ϲ~���%"O�EIr+�lǶu�ǤН|r$�y�"O"h��I��1xD�A]�!%"O�9��f�*@�F� ��
�PQ`!z7"O���2�ױn_8� ��6E9���v"O��bR��N,�+� ������"O4����-�PQ�7&��uW"O�!j�#����d!�ͥev} �"O��J^!"_HD�F�,>ߢ�KF*O��ӕ"��ve���F�^����',P�dU9)�Z�kĥ��N�2Ũ�'��	:w��u����	q��X�'����`V6���S�f�:c����'L�5[e�Ū1
0�J��]����'�0	"�S�u�8\	ƁO_�t�
�'��q�f.��7���8 䛆P�&�!
�'���(Cc.-� ���+�"fp	�'�K��0g�D�(d�ښO@]Y�'�X1��s5x�2p��f��L��'��� G�ҿY��� b�ZWX�J�'x����AE3 xѶĞW1l�1�'�z�+^�p\4DK&�
)a�8-�'�V^8�$�DjX:���Bn��y���C���V Pn�2����y2i�M��ݢ��C��P�q�O�ycL�m��y����0Q�X���B���yrH��v���ӓCKF����!c�)�y�.��%|y2��R9�B�����y@���&��7yF���y��ŊlL.���m�HJ̈p�㉥�yb�e@t�i��>?�hLA��y�H�46TH'�;;c؈��֍�y�(��fl~�۷�:9���,�y
� .����N����㈏��d�`"O���˛<X��,H�Ȭ�:��"OZ��t,c��E�7R�ܥ1 "Ozl��Ph`I�Dn�S��X#�"O�E遂�,��(a�慡�M�f"O�� �k�+~�8�I#F�!�,X�!"O�yڐ�=cg�M����I�L��w"Ob�B��
nQ�&�Ҝb�T�w�I{����U�{j��R{3����!�	�
C�I��ف�kT�S���G�� %����)�矠:c�������c�O��Pn/D�x�%_
2�J9AE�8*Ҭ0��>��7eB�(C
�/����G��OV���@�
ϠD*��0~��h��Ģ$�����m�J�B�S�v��"+͜@�F��?1���~�L�����L:T0]��O�u�<i�G��6�h���!�	E@�k�<�Q��?m5H�@r �mר�#���e�<	SI2U�P��%9���s��c�<I-;m�&�	ǁ<+�>�K�X�<ك#�7�@ѩa�]"+I�}��iYP�<�b��d2���:;|t�R��N�<�r�aab�:D�C�9�>�6eJH�<�pӲM�^����0� �r�\Z�<�6 �0+�<���1V�>upjA[�<��� :{��B�c�"8�P��#�B�<����]�tH`G��!%�T��J�i�<A�J#Jv��pq@Ѡ/u�E��Nd�<ynAB�*�HdF�"��A�2��`�<aVg�#���{E��<��M���It�<�·1N)��i�,�g�d�5ho�<���O-e�ؠ�ᇪ|P�)#���h�<�!O��E���F��#$���q� e�<���M"A:��`�&L8 $a�/�I�<ᦍD�j�1� E�4 �}�G�YH�<qbIB�k~�˰��)���Pg�\�<��eB')=b7�M�N�]qԤ
&�y� ��H�Y�DźSu$��yB��)|��2/X�-:]�W����y�m˙V!Lq��g.������M�
�'��l'��?4Fl��r�\ۓ��'�>Ҡ�� Gr
��Pکh�x%�	�'�Ё��	!�h�F�˪]�&�؈�d4�S���ƨ]"���?S*��9�+�>�y2�&Cj����R�FL��Q���w�R�T�S��?�T�`�P�14)��5�ZU�W��u�<!O�:�`a��=[�$�b��0��F9a}b�]�`���fA�<%/��`�Eү�p=Q�Ȇ��?ɮOni�'��[�r�:�nܬc�r�;q"O l	Ca	�*�0��w(ư��!z$��V�H������(�f��s�P]�ĬW�	�L  V"O�l`�K֞BN x ���#1��#RR��F{�􉆽,hJ�AaeА�{`�M�S�!��(# �"�6C���6������<��I�xͼ�T#��oY�ٹGS��P��dO�	4i@�q� o?/��qAE�K�$C�	���d�a��DN���:.��㟼����(0������9�?b�<�"O�(!p�Q�~���q�ڞ\��Y�n)��h��d�!9ΆH��!V4���D�!�D�,h�f����'k��4o���b̀J؟���'�<cP���=���@*6�OnO�}C��B�.(�2p�ĺL�RԉQ"O�����Z�+�Z���˅Z�L@�Q"O� Hp6����9��U�k��<R�"OH�����R�ԡ[�+M�L��"O�HR`0p������Z#��0"OPt��Ǔ��`
'�>�p""O��8��$}���$(Ԁ*�UbA"O�tɐ���;�Je�Ȍ'N�TX�"O�XQU� [��� F�~4Ҡ�"OD���ͼ@�n��6#ҿ0$$��"O �8U��8 T=A��H
l>x `$"O�X(�F!�����8"���"O�h{ah�;��
F#B�(>B�"O�� G̵I��`�s��8	j|�"ON��Ǐ[[/6H����+_!� 4"OH@���Ʒ"�ܡa��b~��a"O(a�R&,j�x�.+��4"O���ݑL:hٹ��E�t�p(�g"O�($���T���Ò�XS�\��"O0Հ�+3
��j��`l�a��"O<�r3��^��%�s��Q�R "O�mxH�Yu���� ��+R"O��34M:w��gfG
ڐ8�"O��"�,H ��Ȉ��E�d�3�"O�IK�PF��AA`
w!���QE!��[�_�F	ɀ�L8������#
!�D_��\l�Xu|A�ph[>�!�!h<�iK�L@ �N�Ц���g�!��|�����\�X�!�ً6�!�DG�
!��i���\>ld��F*(�!�%o(��w/�WR��CE��.�!�d�]�l��F"p=�͘���.a�!�V�,��!�,67,��Ѥ�z�!�ߜ4�Б��ɠxb��X�4L!�$�{ ��s3������a�ō�]!�R!^�МI4��3�$$ˢe�!�$ɘ4.��C�5庐�7����!�-��H��*�up�kVl�D!�$β+.�9��
af$֤ɩy�!�DE�n?��R���#]�d���˹X�!�ċ8
�>4W���.P~����Ɖ`�!��1�ɠV(͍]0	����7"�!�ƺ @�� 56�v�V�	�!��]̨U�F)(q`gƠG�!�D_r�lڑ�4TgfL�r��K�!�D�U�H���-' ��Ju�X%�Py�H��9%>�i��� �3��"�'��<��`��>!>�����,��B�'=JAs�M
}��p�ӛ]��y	�'\�} � �A�x�����Q�*0j�'�8l��D V��%(�55W�0�'﬽���h��P�$
�<��H�'���eBF�a|�C��� ����
�'�BlC@�#1����	��J���'o��Iqi2:{����)�'�6e×锚d�F�BV���dC�'�~�YbϮl�X�c���O,U��''�@�e�
��3���>I����'�0I����!X�Сc�$ҝS��qq�'5�����ǒ,���룦�LiF|j�'<F9�EnӞJ���P�GF*���'A� A��& 3��S9m�L�'�JDH��85L� �&�'G�L���'�n�:�ိ�0�`���:����'N�@ ��   8   Ĵ���	��Z�+tI:E���dC}"�ײK*<ac�ʄ��iZ�Fm��xRCc�7�	 >NL�:�$jc$@:��9*�"�$�"B�l�n���M+î�%
��N"G�h���� �����jªҘ29�@z"#L�%���sV+,k�,��RP� �� s&���L���eY�J|b1U)��(�R���	�(PĚ�s��,'��	���M� &Fr�	�6l0i'1g�ɗ��j���N�(N�q��iPr�;s�`$��3b&S"p��ͧP����z`YJ��ҁA�d�開��MU��0�xZ*�'�|c���Z��'��i��LS�����$T�	�qJ�e�΍ҁ�"b�,L�� 	� �֦���I\r��`�^��?mx�	d��)|��U�R`�r$ m���0���[5��u�d�
���X��|�h�$����\	�Ajb���JÀ8x$����=?��ؓ\-H���O��扎B�A1�R�`��Ì02��xz��f>%����7�?I�B�?*�P���@�1���T	L���t�'�@)�f����B��M.Q�3˘�@�n�@�[yb��}a�*�'���ɿT3��C�'a�m[ԯ�s#����m�7{�i��O����ȇb��'Y:�0/X��I��VTp+��"[�(Q��>-o�5�D�}:%��JUI��Xh��O~}{�G�D~P��dN:�|tQs
ܭ\2�N>�E	�^}0E'���NV1yh��[��x�`O۞'��yR�3#M��	�݁�@�F�W;6����&���&7�તj�^5���V�#H��� �7Mr�TS�R��5�� �n?�55O��AR)����E�'�y���q�ʜ`��	@����~�{`*�7���� \��Q!�/ƹ��9�c�P�pLQ%�'a~���랎U����8&��/O�Ő&b�r��'c��9�E���ē_����c�� ����u�C�& ���P)I�Ǝ`%���&A�<�*b���(I-�y��
Jրt�!�F)X��,����y  @�?�l d  �,g�Y�V�}�Hp���7�O�x�Oj̐�`�?i:]�m^֜q4"O�M���ح��놛v��G�'	r�����Q界H�Z	�fM޴5l�P�ȓ�fT�Qrm�h��[1��h&�܅�	:
7�ܓ1cZ3 ���Vk����C≔!�����)5�t�i���N�*��ٴ�Px�Ã�V�"h�G��#;�$ؔJ�y��ėȨ�&�Ѡ��5�͡�eίK��@&"O|����u[~�)1dA0^6���2O~!��Ÿ>��O���*���m #>bȐ)G}8B�&Z8�[Iȕk�uK��'6�6���9�D֮8��	S�,̿��d����<	!�d^
t����T4Di��B���J�O�����~�q ��<��8��#�CF��N:W�OB��S(�~*!�pɈ j��tb�`�BF*-�̣<ً��O���(�wjZ`q��.#F�ҥZEH<�&�]$ ���LM�HN��H�� ֟�ە�'�Jd��G�=�Ddk �S�}.X��>��'7qO�$�H�g��H�b`��^]Ѿ]s�8�'�S���k'��C�e�CP)��-.�>qM<��O�>yA��O:&�ށ���#Kk"�C1m6�I��az҈�%bzr����٦(��Q�N��#�J"<Yw�>AT#�O�6Dy"O:1�N0"�PL�<	��!K�L,:�nηa�eJ�JƟx���'��HaR���T����<Z�S�b?�O�a2"AD�,\�-ٵo�=k�O>�żt�S�֏@��KM�{!�P[Wʱp���@%>dJ��
�'`��2 *j��-N5J���'�N5x�Ϝdr��Wb��Tm 
�'����'�������Ľ9	�'��K#�(Y:��K����!�j�Y�'K`U�0��+%�� PC�^4F�	�'>��q$g jt����,� q�ez
�'s�uRT��fE0�:R�V6G�X�	�'��ƨs��(bQ��h&�p�'��X����R�:�*Kj3��J�'��u'd�RAhu1N��3V�LP��� ���*u����̾W�$��"O�`j�3(g�M+Dn��(�V$"OҸ�r뀥=h����W+G蒝�"O��0Cʄz���Lȏ�&��"O��hǊ�-��
��E,�,���"O��Ô\� i�����:�*4��%Rc�<є�	�U���h[�
���� �y�<���_$x��	�GH�O����x�<�ENBN��h���%`|�� �H|�<�#��:&�i"�&:SF�����I{�<ɀ�Y�2ҙ1d���|�\m��O�w�<9��"���1@��d��9��r�<	e%G4p�4ʔe�8Â���A�k�<1��˖V���yEϔ�;�X!SA�]n�<1"X�I>0����]�lV<�Ǎ�f�<����p�Z�CF(Ⱥ9/^��Jb�<)f��-)e|p�p	�C ��	`��a�<�KM�(7B2�!U����aC�CZ�<Y5i(l,��G��@E�3�J�^�<� ʆ�XV���*B����A�H\�<�F��p�(sKL�s&�~�<�DX�+T乹%�X.��d#f}�<��(��
:
໥�(m�4)�q��z�<1u����$j"��oN�5�	[�<!6C
�m�̹���	4�v<�䢈@�<�a�Ɵ=>� ���QT��[u��y�<���V�Z8��O�|A��s��@�<��*O�FXdDHŋ1G�d+��v�<����U�2퉄��+�6����Y}�<!�%��,`�I҉�<5x~h4M��%T ���\G���Bu���e���'�=O^�0��%D�@�F�Y�)�ddk#��:0�\$��-7D�d��%V
I��Y��;&p�Ȳ  D�� C 
k�L=ȑ� ;)�L�	!D���S�OC�>\���	18���{`k%D�pah��z-���5o�t��t�"D��u�����Y���Vԉ��#D��K�;H���afBvl���	!D�Љ��N�oo��S�A� NdA�>D��{�!н 邭�RI/����{�C�`��#�`�;n�L��u��ʲC�	�s�z��d��#
v�08tfEJ��B䉙�݉1$�$\��̋��1�B�I�y{4�1w���?&!�mO1$�C�	��1�Vg�n�p���ӯ+ͬC�	�X�^	s�*~p���cÈO@JB�I�{N�=(���0ixya�jB6�NB�	:	���9��ZTv�D���4B�I���ҧ�ŀ�z��4�B�	�o"���O�g�jx���C�C�	-�M9b�+QT�뵮-G�C䉷<ݖYڇK�5.x��È�[0H�O,p����Z2J��D<:�]�ƍK���l��c��.�a�ŕ�zq~�2%��K��(*1�YQ�D8�g�U�QV�u��I;,8��3!�G&�h�2*͌���IhⅨ��S�h���%>A����蜍	E����%2��2D�4ʇ#S�.l$I3��X8FY�ᰟ|ACIu�p�QJBPy���ъJ�����ן�"dp���@�!��_�5{�+J.xbH}!1�hM$��'��q5�k�)���On��jJ#G�2ň3����d9�R�'�H��GB)�R-Pt�#.)��2�+��]�h�G�a�y��X����) ���Ƣ	�Q�hhR/����cu�^hⓩ8K��.���Kb#6V2�*"Ob�[��I.&C�`b'>Y<P;��Ov!)2 �,�����<E�� ��S�	�>n�(����0b\8R"O��JFh׮.ib�`QË�TPTY##�lyR�,u\]i��M���΁~.���7'�:�\YC_�,aB�E�V,�ƪ����Jˋ�H�v��k�.������e͏Kl�JօĂX�X�?9@fj�Q�MV�'qd�A
gF�Pq�d�CdUh)�ȓ�8���![�Da�$q��$i������8�zWm�y���_�qXl�'=��&�?}�ɧ(��9�Ej߿�"�Y�J�{����x�$��k��zr�R<�F�:7O4pl6�ʖL0v�h��xBō�7b���[�2p$A��/�,f2M���ԉo7��8�,��p?#G >�������R�XTK=k�l�b08Nj�ӈ2'ɯq,�F�Nɽ¦-�˖(p� �>��O��˧,[��x��Gg,�i��F����f���e�:y?�$V>ybv);�{��I
�j��į�)�x��Ȃ5�D�}�0}!�E�/C�S�Ot�Q���9��M0P�/�3I�أ��ˁ1az���|=�D� �"���sa����!���GOD:l�\�����U)2!*�Oԩgzڠa ȶ'�8��!��~�T����M�v�t�h����#<"t� (C7i��xB����qc6�k�K'�'�I1�-kݮ4�g�#j@��F}RA@�ي��v��z��O��U��"ǝ,�Z��咵:�j��4
3P���%�*!��ҧ���&Lk��5@�/�Q��I[H���'�4�g�O�`u԰� S��}���X7����K֢�"����[}����X��t�Hvx��peI����Q��i�R��5O�I�F#t��h7�z�s��K�.�>r*HE:�oA�'�"qJV/ 4�H�`�/�	{�ar�_�M��r�d����R�	ູ��\/K�O,�;w �'(\����G	 ?y���FB���U��y2-��s!!�Ԩ_,=��5�7���M#%� �ݳ��4}���ibΙ�F�G0NRl�2�4$~Ҡ 	�'��$qcL���T8a鐍'$4�C�O��'ʲC�Ix�ā��X ���N>dr1Q��79�a}�@$k~"���!@-��! r	�>[��u�*&e�T�Ɠ�v%�@�^�]{�d�w���Fz�֏q����5��o�'Hd6y�UǄ�r6�${u��C�ք��a�h�G��c��6�X-q��InZ�ZG�t���]��S��M����*I�a�� *'�4���D`�<tծ:�Z@��:U��SԀt�'��Y�KT�{�az���)u��q�3�ӴZ��4i�&P��0?Q3hWF�L�+���7Y�)��ś��@j��I�<Iw,��k�� &'�?r��R� �J�<)���[}b-���ǳr�d9�7�F�<y�D�vO��$��`z��y@�fqO�4�!`-�3}�I>b�5���A�*�lm���W��x����H}k�.� @��rv��z��q1+ԶG��~2�߶:腛6���,�0 �$DI���O��7�Z�y=��� D3��擢��Mi���>6���I'-�m�<1%�L��ݛ��5>��'�k}���<%���S	�>X��I �� ���t�|�3���t�!��q�v��4�R	g�bE
�M�.9�D]0��OH0�t˒�n�n�yL?㟄���`�2��c6~Bn��D�.�O&A��*S�K�Y���y���&��R�B	�Yd���$V�5;b�/[N�`pd��)wB�E}B埲&
v��%$B�D��O<Ȋ'��;`�^2 �F�B�B�'�lk��d	�8P$�#z�q��'��<�%��%{
�;t�o>�� �Vk{.8���
h���R7!D�`k�H�K��ظ�H�r��UZ���7d̈�I-E�*�Ç�#d�g�=k�'ab��2���+ȮH����)�D��V*d��ʎ�#�ر�f�h)1%¦�p?���'g>��r5b��^�f�1Nw�'�mB�-T&b��ś���¤3�����@�`~��G��	�yB�@9!.��'��i���7aX����>3Q�\�t�8��B�}`� �&�,�)��>��4��8�L��b��3!�
�&�<љ�b
�z��	8�Ά�$���?��+X����>��w J��1^?�;���!z T���%Qe{�d� f.D�� ����*v��էY�SFx*��J�P��	�g nP!�I�c�3�I%%l�"�ه%O��p�(K�d
����I&-x�8��G�I�LB��ƥ5����u"G�vrnT��)�O����LA�bV.��#Bڟ	#�e�4�I��i�`j�lx,��O�~a�v��)w��U���;^�IK�'���V��&C� Գ��-��m�+O�;�oK�	e����E/�銈j�Բ�����"iE�*��j'㚨m6�-��'������&^؂i�����"6�'�ýo��P��m�<������E���Wv��{�k� $�j�y�)J�{�P��w��8��ODh�N�$��<�/O��*�@��q�n��q~�}�G���~�ĠK'���cL,��gZ���=a��j �Y僛3�l�r@BQ?��*ֈ��'�<�b��H�rlK��-P
�T ��.H`�9PfΆ9}���0�T ΘA�'�RI�eFI�|�v0R �Jh<�S�O��h��W�5��l��L��j��<y��Y�Dt1r�IL~���˃zg����
ۋr��	�H
�J��~b2*��1$7m5`�b��Y���1��#G�`��À�.дE�� Y���5bT��w��|�A��Yޔ(Po
� 	������?��m	2���� ɡ�~��-jF�1�G��@��,4��a��B@�p��壠��V�����d�C4���>02��䇧Q�����i�?��	`�*A,}�||��;����N߁5���gݟ����I�q��a����(��F^V8��(Z��Pw��NF:��Sx*���5-/�T�ǀK��:4����d{�4Z�W$y�Lh��c�~�����EM.躄o���exH�T�9����.	l���œ3|�����Ϸ}F��W`Ŷ_�0e��&e���Q��X�[
?��8GԚք�Ғ`	"[����
�xH��H�hC���'@��3���p������&I�!=A0G��z)��@Ҥ�A����AZΟ܍̻h�d�A�eW�y����4;̐��,0��-C>d����D\�x5���"�B�bZ$��.ʾ]��W��/�"�A��|���A�y7���'��M��'C�ntX���&�^��ҁM�`l�KG�#LO�i��&^�4޹��A�+���*	!V<�ĥ��.�p�]1�� B��@�N]>��R���Ð�I`�l���	���󡀦Z�jh�t×�*c�l�DC���&=�Ṕ-9H��hL3tQ ��P�ƃ�gB��j����q�4j9�ya6�'��m+���A:��1p͝�rTx�S��]71�^�S4�[���Y�>E��e��;B<��	m�rV|�s�w�����/ѩg�XX���w���:�'��x�o@�o�2� �o_�."�$Ф��Q� �*̦�����H�r*��%�^E���^�WP| Il�T�kG'4��ZӉ	!f�JQ$)<O�B�)��v��D��]�`���AF�j�A˄5a�QX"���XY�F �Bps�͑�#d��q �F���"ʞ�#�h`p� 4�D�$�hh��H7�T�8$k�/��a��Gs	�$a�D�C��������DSs�IeȊ�P�$
l3�A�@�t��Q�"�BFI�7m�5}2��w!�' X����x�>l�7A��}�q���M��ۇn�8dp�O�ݼ#F���z�裒G� �4l����Th<�5@���>���$Ύ~$xu��kI!�@9����)M���'W&|��,J�ϕ�0��RD�x*dM�ȣ�y��Զ����u��8{�v%���Z	��<�Ej�9x�x�W�[�X�VU���Ć5��9��,�;�-͸��� PL3�_o��{�h��1"�E��O`cӦ�9h3��Z��"�6����|����8��$��40`����C^�0�(<
�͓K�tK��:�z��ł�/e�t�Awe�f��E�3/ǹ�p?���W�d�� �X�q9��x�F�/9nQ��K�f���y'c�Rm��颃חe��&�؜p8��`��Hؼ;Q�˰m�"�;@���B�P��ITh<	��p�a�Aǔ��TxX�l�V�L{ gݤ~X�)̈́���X"5*1v�A���DR3`��-��!�x��ᷠ��=��y�aѬz� ��7��8�2[���7V�В䍁[�&H��f�T�d�1��.L����'B$�!eH�-;PHu�ӭ,+ hL>����..,(�d�W�@�⣥U�<�&t��b����/��s톡⃀�>/�`���=�y�>BB�]Z�e�0�LTA�,^�-D���$�'V$-�A�EW���"䍾��T����w4�y��A�w7J𺐭O8=o ��	�'H�)P� �cw5�f&7���2𤞙���Qin�1��, I��	,�y�'F���ē�p6�R�C�!th�ӓ8�j��a�Q
=��¤�5e����^@�{�(�Cľ�k#�@�N�"�i�%4�O���#H*G�����.C1p;��A�����B�0JD^
G\%�ĭu���1$�~R���<n,Zh�V0�"v�<i��9hȦ�Yk\n ̓� �g�h����
���(鵦�=��a��)�ۼ���T�O���W�s�$#	|�<1fI-ؔ��cP��1A��[�b��Ԃ�-�(>4a0�QF��i�m�'���ˑ(^�%A:�����#@6�R�4�����Wh�����c1ꌱ��9',
 V��*�(!6�.�O���Hؖf�܋��ѱ�̥B��	�����(e�ԛ���qⓓ.�ɓ�֊qİҪӜZ�,B�)� �T�e�R!H�v�p�&��D��̃u�'�(��)Gi��@d]�"~26�5�<��z���+����y"�MvXLPI�-hDe��y2 ބ]�~���kצ	h��+��y�"L�r�$���H5�ޥ �� ��y���b��<�Z�I	2-I����y�Ă��X��M�B����V���y����QUD���ϧ9FԼ�"+[��y��U���Y�%�g�8�páٽ�y�ɝ�Xg����ᖿ`�����%�yB�i�i�C�ìT�r ��H1�y��D�a<$��#\B�@\�fE�6�yLN9\$�E��g�"1WN�*v�A�y�<<\��0 OW�>� 9����=�y���(`C(p����)��je	�y�b�5:D���G:?>���G�ye�"v�^,P��E�4E��:Â��yR�L�s\ȣ�jC
4@\l#��[��y��C9��z@�)��4�P`�
�yR�7_�;���7�$�S���yrҫ%�9SA�F'X��;�,�y2 ӭPoDt�7D�}����6��2�yr��/�D�hr�N�cц貅�g��'�L1�JC�
Y�e���:^�Tp��'ϖ�����Y^��dE�Rq���'�DP��l�B胓*B�O{��	�'OP@� ޱ+f4�0Ê.HrV)[�'ĬU�0.���tڰ�Q$9N���'��K'��1 �iP��2����'��d�J��nb猖/����
�'s�lSf!(�*x����!{����'Ƅ�f��zc������,�����'��qfF�:�$�6F����)�'_fa��[�CPai3b��J����'��5��bCX��b@�#1qDz�'1~�� ��	=����cK6+���'h�!z��6!9R��Q#H#6#~���'�v�Q�m$,)"��уΆ,?݁�'�� SR$��,ov����

�8{�']������)���wO�i#�'��i�R�و�(����üf��3�'fN���k�-�`$q�F�bO`���'p\d�%��UOX-�kI*V	�9�
�'A|1A4k?o�@�����X<�'P"0��P(4�~ �I�/%�9�'�P�C�灲� =��� B���'���`�Z9Sf�ꡣ�T���H�'$Љ��/�x�d
�d�*>>�8��'�y���=t4���ư1)li	�'��<!g�֙K4���J���)�''J�;4�ђT�2�cp��� �'����&��(��Z�ǝ�L�
y�'	��I�|DAvD�irB��'6�P�� :\~ ��/�lf���'�x�E(�K���
1�
�a�<�'��@3F�ё���e�U�.�,�O>�E�չ/�(��^D�#aU�W�b3&]`���m��4��<rT` ���>�+4I\^.:�c0�'��|9��A�7�6�hvJ�n�8�J��dLq��B3�Sd%���M#����q��g*���68	�"OJ�c��-`{IQ���2ux ���Oj�c�E� ���C�<E�ħYQ'���v�P�2	���
��yB�S�6*� ��!�b!�#�'R�>˓6Ո��E �"�F���'ݠ8+�fЈv8
��AꃚLcR�X��.X]�,-� d��#/�0K)xH��+@	�T� ���8�x��ɣ&a�a{%i <.P�@��[>#�Ȣ>yB���Q� �C���' ��zR�*�X��-��	�ȓ)��h��`���1��&~^������|���;#6<��*O�>esV�L�W��Q���[� ��� 'D�Pʰ�5����#E
Y�N��%��D�/j�E �5��3���z��u� 6	�K���tL����	;)��oO�<k�Y��jU�>h�����ܻ������). a3e�nnJ��U��=�G��wN��9�4H"(a;%�S4�j�H "Z�a�!�X+Z����d8~Y�lk�E�B3!�$&).��q�ȝ2q������%�	"v��Q�7*l�)ʧ�<�"a�3n��3�հ�`�ȓ"�-�թ�$�<�R��6o�@�H�|��n��o�:!�J|�>1�⏏(�� &�"�2��i�d��D
s	P
<9�*2��3]8�ܲ$�ê��k֨Щ!��8���"5��`hP$I���8���&���>A�)
���)�4ŉORR���`��
ut��#�&<b���'��`����4E~���ֈJ�?�dPp�'��5��Nִ@X��IS��}�pa�j@��䍮]f��R��x�<Yq�3S2I�Q�-t���c�?���-A(��1ꞌ��gyb�})��qKА�tRW	X�$������p?q���.GO��a����q9ƈ��N)k5a�=��{�{����l�حеᓴ�Q(�gƣkU�r+�m۴�>q�wr��@��ħ2zX4����..�����gK�zʚ�nZ�g2-��_��S��M˕kI�E�p����?7X�q'Lh?��+1FX�������S�Q�xp�!��$����F�SY�.�`
�\���۴�'Z���,�GXa9%G�*�zd���>�R��=W!���v���'�H�m��x�f(!2���KK�a:��	�[�f��0iR؟�Pb$ֽVc���!�~>^P��Z'td�x&�`�G(P����_���?���˙4S��{�"_}u��W' D�<#��J�uVm��X�c�h��~�8Hq�!ϩk���J�"~nڰI�(���.�R"T���%�2�B�I8eF����ؓ5fb��`ȇ�y;��\���Qヌ�@;P���&�Y�(Ń'��f�D@a}�m����q��R=?�����h�ع���	<�̅Ɠe*I�aӷl�<(5���]���Dz�G�6���i�v�'^ߜ���1�(\3t��U�NЄȓ	Tp!�5< #���Rho�
/a�!��&�a��S��M��k���=rX�Q�Ԁ�,@�<�6�H�S.��ID�,R� �ȧ�VybgA��Bi��'Pq#��	r!R`l��m��F��䂠��ώ��h�p� ���g vA��b��E���\
r� �B�E�G٦�� !`�B�(Z�r�hQa���b��1�ȓb�*�`Rjݓ<��w��8R]��9�d��/���?�'�tԀi	/Vv\M2խ�i�d<��'4$�%)ުq���TkiІ���ɯX��* �'v������"T�r�Z$��[�>A{��F�Z��%��"l�'Y��xӥL
�8�H)�$�%N%��ȓq��-Kx����'Ż{ u�'XFЃ�않;#ʍ�C�+�0���	�vg �� I� btx1�"O�`zgO�,0�T�1�˽-n����D�'u����[[�qI��4��3���R�J���-Ҵr[d���� ���d	n�^{���="(��jC<RX1��&f�2���"���0?1F�^%�t��g���^��Xn�'"и��H�s^�)�K�Q�4��= v��sCX";���9�.���ybk�?D!�� O�l��lj1�;�~��}��T'҉��çQZ��*G
H�P�q��Ҁ�ƕ�ȓH�F�ӂ�ųU@��� x�H��*{?��@*K��4�8��B� �>�r���'N����7�4�p?�B�+���p��B$g����5Gϩ }�Y���t(&Tb��'Ɣ�E�1$��(DmL�n8a���D̩Xb�(#b��C���H��DeޜK��b3�����;�"O� ���5�E�zH`\x�Y�e<�z�R��SBC�2=̮0$��DF�f}�Q%>=	�!�3@�x�/L�=M�-�&�!D����*J<�h���3[��u@��<?��0d���۰$;}��c�h1S�!�~���ÌzW�;᜴$+Ь�t�<)��:y���Q����*�fO�A.J��'i��7JX>��ϸ'�B��A�\�.w�ASC I�M*����k�N���JŁy��� �/.�U�t+�=0�@4�߽�0?9J��SH��e�Q���KU�'yD=itK�AHPA(B�?I�s_0>�5AW�ɯ���0&7D��c (�>���w�U�b�����<Y4�_Q���r�΋���'W���w.�~�։\��@0-ޓ@����Sg؟��tS8FJ����!��t~l0x!���Z��C$ښ��Ł5L@��ǎkn�3�	�>��DH�J�kA�2q,�>����B����q��<����<�$�!��ф�	
Tu$iY	S�2�a�k�L���$�h�@\rw�1]R��bG+@�Ge����h����¯:��ěI蠅֫�<_�l`�L=Ѿ]�g6���gCߘ(R�Y�*D��`�/ܰkΊeڵE]5�����(?��K:m%B�Cf�G�K��+&��L���/��1��h>����/0 �Z���K���@�=�O2B��jh��0�E�a� ݃�� 57�h8z&&��
;J<KF��<I+
Xc���f`f�H?�O*|reJ� �B�; �P�#G�<�&�I�5V�j0k�9�1��<����-�=��
��of5�@�O|ih7Q�Zh+ӓU_��J���4}�L�����bNV�5٨�3�bE=`�ҧ��O�*΄�j
KV�ꈨ�c׸{��ψ*@F̣	�'rD$�u�B�.���A�O7��J�L+sBm.�[���b�D��>���k>�3��
Z��X#��hk �ڕ$'�O��(&�D:�x�
4�Ǚ�dyb\�`����(W�D�h��!��V�DPo��?��66Of�� 
�m���c�_�'��4��&�h�"/����ǒq��A��,o�(��W>������"��,LO��c􄘊:�n�8 EQ�z�s�'H�(UF<|����"�+b�P�j�F%/ZeAѡ-D�dy2�HOB�%�1/ےh���-N�c\�-�de�� [��8��3�	м3��֛M���ՌĚUzѹ���G؟�� ��,5Ȉ����O�j%�ʲ�+�i*�,ȎK�����s`��ȀG �^a�̨I� =�>9'�_
x�e�KHS��'^���2���pB��aBX����ȓD�Z�����5#\n����jӄL����9���=u\t�f$*��m$�U�P���&̆�"Ob-!f*�ET��&�L�F��q	�d�`��Đ�mB�EJ���3�����񆡍%K/��ZeKR�l�0��d[�P^H���!dE��F�/j��sd���u�b\x �0?���_�z����ܭ=�R��Z^�'���ha��;e����Y�dǓ�P�T��c+�\�XRC&�3�y���c��驗��R�����+��~r�ϼ��2�e��[����ӫX�zE�����	�AA�(F	{�B�ɹ.>�q��&Wα�T��n4��B����j N&y\h��~�?��Ę�x��u�g�QD/�q��aT؟H�"ɰ%SJY�CK:V5Լ��Ŕ,j�4��w�'=����	���#f�K��I�G* w�?���.#�%�	�b�5X�dZ; C�I�b\<�!�d-T\չ��ښ/I���b'Q1�!��3|������'隨���n!�d�V~��B>o�`y�@R�_!��#�Qi�#����1�8 �!���R�(A��C7���c���!��' o:]`��	_��	Ɔ�S/!�Dא�V`� �^z�yAWeK6�!�ĝ��������,+|@�H�$ߟc�!�$8XJ���N�	z��/���H�'9�Pr�.R7r��TS�������'8����PzL@R��P�*4��'�Y8�(	%=������>x����'�R Q�c°S �A�5����4X�'�����
�{jpAǃ�C3�'3�0����6
���Bu�H�2���c��� ���U;�!3biϮ�l-�r"O�1��#sO"�R3'N�t�@ a�"O2�c���
����0c~A�J��y�צi�`��>M�������yҠ�	:�gc�,�Ҁ�H��y2�V�(�����j�y-+&۠�y�� �T	�F��T��Yu���y�e�4j��s�J!N���Suc�3�y����ef��Ŧ	�4S�ɚ4d�:�y��ٍ_~N�c.�HQ�#�yR�]*&b���g@n�Y���Y��y�N�s���J��VZC��a D��y�Ά1v���e	�$I��H��ܱ�y�ƭL\���G��ab�	��y��>���q�a� �p�!C��yB�,^��*���z�����5�yr��S�BU;�N�
*�q8�!N��y2NQ�1Xu�����$�y"��8�h�'���y%����H$�y�N�=�t� �nşE�82 �6�y*�`i��[��̦8X| �1"@��y"D	3$��`Z�nC�ay&�!�͉�y"%F�0F�Ÿ��UR��g�	�y�j:"���eL�I�~�1B��(�y�	�\'r$��йU'��r7Lյ�y��jc��b���\T�F&�y���%~ ��6��;^�u(v�L��yB���2dलV�̡UR����6�yr�;����1 
�3��[�*C��y�%ܱ{�����L�<UzE�k��y� ��o@P�	�@S� W����) �y"�+>c�u!�g��/-�YA㛭�y���8u��ӥF8���%a�0�y�C�
jtZݨc�˓m���'χ��yl[�K5�M��ѩZ��6HM0�y�%�'��6䏈
ߖ��BF�9�y��d�ze� `�;�p$��N	�y ��3g�]Ȱb��<ʼ��FeT,LI��]�����(&Y��;1O�DW �����vF�k�%��P�H@y��Oa��l@�a̢�Y�Ι�5��8q^��O�ă��O2�M� !�H��Y�g�+A`2Y�y�Gԫ�hO�c�T�j�[�kΒ�P��*g(�$��D{��DeA6UE\��)�����'f�AUў�M`ԈL~%J�J��V�\
}
@	r����<�4��!a$ʡط Ԡ���� wz�� Ӱ]�B���({�	`�W�q2	Ӆ�Xy���)"�4K�K��Rs$Q3��hk�H����	b?a�h�>*��"���8j񰗏,b��eGP?�@��=|E"dC&׭+9�"~���d�T-���3���p��(B�C�o��/p�=K�o� V��z0��q��M�'Vђ!��$�t��S��	'��D+�@U��xI�n�?�?yBMt>�����	U�z�b�].<�L��4m֎j�Xe�Op�w�%i�a�Dj����a��m`Խ��铥�t<��$>�l�΍�L�.�D���ܼA� �u"
?5"^ FDأ@���'kF���0G�����;cH5 ��4�P��ѷK��I�o���`������S�O2���v�O3}I�U
��Q�{���ݴx،�a�	�J �9����Oq�68�W3O���`D�S�zP�H�3{��5�<��O�҄{��
�}�iS��qk�S�-�ɖqj�[�'+�D�'��ݳ4N��p�K�tk蠮�Y���<��jB2X��b>�J n�PR�Dr�N���9�$?��
�5�1c�xʟ��''�(�4+J$e�x-�&@2zlX̓N��@Zƨ�"m� �/O?���
å2 �ȡ��2l����;O�2X"b̜*��$��0|b��ʟh�"Ĺ	��97����������Ĝ���^�@�ÃuE��	 ����&ͮg`� �"HȺ;����4ht9c%�AC�ٕ�h�V}"b`� 0��(a�G)7<�1q"OZ��c *.1)C�CyP@�2"O� pXæ�?+Mh0���ُ9�9�t"O�8�g ��z4�&#0�\}"O���	c����b�R��"O��s�/~:�t��
����W"Ojɣ H�C�ٱ����
���"ONt�֍���`�Ə�pς-إ"O���A��B�^��$U�X��z�"O����1}i����5�P���"O�5�ЬϞR)"0r�����(Hb"OR9be�$E~�x�ŗ��(�HP"O�Ax���$S���sJȁ��s�"O�i �큂7�R!h! p�s"O(�h�>�Ys���gR��u"O�stKO�9���*��[�q���iQ"O���Ձ� 8&NL"}��"O�DX����P$�s�ːC�|!��"O�)W����U�"�}��@"Oҭct�[q�xtC�G�xƂ@�b"O�G!�?&�̤�a��<��Ő3"O�ձ�C7+���Y��ȩw\<��2"O�1�rf^�t��%��.1c��i"O�a`�J�W�D�T�ĳ><��"O�-��/��&�}*�K	AS���"O"T3���� q �UK"O��k	�b�05�����
sr�z�"Ot9���V�������NTD�I�"O�V%݊�:E+7.���!�W`�<��N_��Lu��Ͱ|��en�[�<�dI�6�h����-�H<��E\[�<�@P��H��5��fTo�<1UeE٪r�o]�F3��)� �!�$R7~B�@���ѻ{+��$�܍r�!�$�M���� 	��+rHyeW%!�G�8��dkWZqlQ� [u!�D�L�$�ќL^Zݪ@�A�k!� (n`Hp`�!Lq$	X���3]!�d�
z��@�Ԋ�C���ѣ_�l�!��B� �漚F�R�Ǫ���D��/3!�݃X� !�� J�(A��ޙ0!��F�q���*�)=��U�w.���!�ۑt����^Ju�iK��M%6�!�¹<���M��2i�4�����I�!��S�'j���*�}L����!j!�d�+~
H��bS=D>�� �ņ�,�!�X�COH�G�j����eR�-�!��f�Ԕ�m֏��t��	�!�Յz�!�M��0@��#��e�!�� v�(��/
)�V�փF!���X,��!�{
��i��F�6�!�$V�`pBĂׇ �<�r��j�!��MV,i���q�$�q�¾L�!�R�9Bi�e���(�]@����!�$�0��9�u��-�� 	��p�!�D�(r��2��ȷ�h���!7K!��;]�Ṱ" ,���s�_�!��ߘp�6��f�$�n�P��'_!�$�gޢ݊(N�0����є.�!��|�.8i��f�-u�'j3!�Dԑ{(��C"F�(/&բD�_;b!�$F�v�����^!*	�4�B%6�!��t/�PD�+:#�a���#�!�d%!��H�unؗk�(gӄ6�!��b`^�"�鄮~�[���!@!��ۣw�8����ceF�K!�� ��Y�+�;ަX
DdQ�4�#`"O�h�&ͧ<��Ã�����P"O�I�s��b�H �#h�$.,z��"On���P�3���(Ea�NtU��"O\!���8?-;��G�X���7"Opa����@ݡ�.'��P�"O��"$4���gG�;5�TrU"O
�{$��1~I(<�6�C ~	!�"O��u�Ֆ0̤+5luڱ�5"O9��!T�0H��ƴM,TA3�"O:��"ٸ���c��]4<	̔х"Op}*�pW,�閈�3>�$��"O�i��H��>]��'؞$��{�"O±.��o:e4��y|��j�"Odܡӫ�c���%�P�:^*Q�u"O(�{U�ߥ�����bG����"O����4��M����X��К0"O"�#��W�Mm8<����5�u"O.M�VE� "�����Pp�Ę�"O64aS�˄ t�<��#Ĺm�D�{"O�y�6�F�Z9�I�3�^�A"O�d*��+Q|؂͉;�*-8""OjyGTs�R9�Vl�7{�����"O�\
 �L/������=���:C"O��P�8!N.� A!( ����"OHt�W/��~�e�f�K�y���"Op(0�/�d����V�2r"�h "O������)y�^X�s�s�8�"O�$J��	�\��`rY�P�ڔ#f"O4:� R3���r�����@f"OHu`�c� ��x�7G�))Gd-"O��BF
X������vʶI)�"O EG��@��}৥�!/�r�"O<j��\�p�kR�)�ԕ+�"O�y����}�l����$� "OZ0���]2IoT��� ������"O.�(F�I�^�Ե���I�A�eCv"OLq���h K��:B�Eɥ"O���K�.P�zy�qٻ/� 0""Ov=� C��4�d�*�j|�U�C"O���D�^����oO�Up�Q�"O(%�U�P�9(��dO�6w�z@��*O�ͨ�d��Z̊�� �0w�@z
�'/�L00Z��
����P؁�	�'��1@�	=Z��"B�9}1�'7ΐ�ak�Aߺ��s�^�a<N���'���S��ȴ4�`��� �$K�hB�')���MV.Jΰ4�7Ԭ�Q��''^p�wMߵ��ErF7�&T��'I�@�Ӫ\�l����͉m�8�#�'X�'NG1gӦ yՆ��g����'k�h���?W�yʔ��K��t��'���H�MV#E���"�B��8��`�'�j�z��$��xSP�G�-x���'��!��ل$���9�,��'��h�&/�'�~����^��@k�'ĳta�6b����6l��Sl�i�'�.�� �%B��,�0L�*�:	�'��ݓ�AB�}~�@�io*-k�'�fa�� �:c���g��[/|���3�tm��$38�hm�Ũk~$����i��
��O���3�%o�J]�ȓ^Ӓ(�a�Q?��@����Q]���ȓ+b���娆�&�P[���q^F$��S�? 
9 F��-hF䝠�+�K���d"OX�[q��9b���6
П1�ؐ�W"O6S��~A�Y�bՃU9:ABU"OX<Y`)	-07�]��}�"O2���ǽT^1h$.^1>"O�!	�lݒ��%��M�� xza"O���pÝx� h(7MգD��d8�"OlĹ�#ҁ'�ꙻ���[�tt@�"ONH�枬[h���I܆*���
OR7���A��tqV&ςk��}�E�-we!�8g�t��.dx���%K�8!�Jg
[@��kX��	�i�)mP!�����1��M�{���#n�(C�!�$�$-�.�@�׭a���*�:�!��m�f���^8ʅp�P�7� ��"O��:ׅ'G�L��"c�kpX���"O�y��b�PSθ��l�e^\��'"O�12`�U�f�!��+�tP��sU"On�ʑd¼pE�2���.EE,H�"O��z�#��C9����h�e7@�"O�
���H��KchƏb�6��`"O�}ZGI<Y�m�E�s^¬��"O��ڥ�ކZ�� �_H����"O�W���9C���2�R9=0x��G"O�!Q�Tvu��{�k�5;�A`�"O����?B����(�V��b"O�a�� ~iha�GM�ըx�3"O"-�/E�Y�"� T���"O�!��;�N��g��J�L�X&"OX���
�O���ڲ���}p�M�"O��sd�	CFD��$LE@��R"O��a5�>+�}g�Q,;B80"O�L��$�GR��7(	:E��"O���B�S��u���1� ��%"O�����J�~ݒ���7��LHA"OD*�ޭ?�ny��E�')�v�y2"Ov��4-�`�00����� w��@"O����_P�,z�l�'�|w"O�����ǎs���Kĥ7���)c"O8�E�ML�P�yKõV�	�"O湉�o8Fr�d���e��"Oȸ!cJ�2N�}��ݹT���"O�|0ӌ@;S�B<�=�.%��"Od��(�6f�la��"ɾ��LA�"O, �`
��$�sA���Z�QE"O�Ӄ�L�V%Xf=:�u� "O:����]�M=�\�c嚺dY�٣#"O��"���P|t"��M�(�@�4"Oؘ��"0�l���4.x0�j��<D�@BEʙ&��x��H�Tp,T��(D���a�;[605�2c���K(D����b(r��XF� J��¬ D�Ġa�_�h-"���׹~�a[t/:D�lj6�ǔ���pNT6|r�K��6D��#�� *���Y��NR�֌2D������*P%vm����'J,&U9�`0D���a�?���� ��:X��T���/D�����+�:!����v3�u�e�.D�|	$P*&�vP3ǭ2V�;7�9D���#KE3q�U8����Q�,- �)$D�<#� !g,��Q�LPTL�X�c�!D��
��^&n�"�����Xf�l bf4D��IQ�(u!�1�eዘ"��9��.D��YQ��0f#'���2�����)D�� T�J.ȷ
TA���������"O(�as�Uo+��lW��2��7"OyѬ���0<�kD o-����"OJ��W   ��   l  =  �  ]   ;,  [7  XC  \N  �W  �c   o  Tu  �{  �  D�  ��  Ȕ  �  P�  ��  ׭  �  ^�  ��  ��  )�  l�  2�  �  ��  �  �  V  � � � � �% +, w.  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�I�Q�"~����	����!`��t������S��y¥�#k`a���\�n�x�P�����D/�O�`c�������g��#���@A"O��H"�\D�,�:�HX)l}f����O�n�|X����((t��<�P�Q�W=���e�'�I^�'~�D�U�O �rAl�,c�2�0�!^�g�� 	�"O�0¶���.N �إ��&P����"O�Ya� :�� �Ѡ� .�	��'��XYbh��@�$��b�]֜�#')D���֊�m���g	�=f��1�!%LO��LH��S�Z&>l�W�
/h�z2F�>
�Nٶ��q�� HF���gL�}?<I���T��D(ʅ"�X)p��ħ�
���ȓy)�t�r!V�F4��ѭM�Fy���j��~bMr�0L2VZKr�Qq������=Y�{g�%���5�N�E=f}:t+�4%L��p��ޭ���I�5��(�-�%n1�fF��DC>��$�'s��r1�[�/v*􂒇�$b��2�O�y����]G�Q�C�$Lw�xc"<OH�'�� ��|��@D�M�Na r�Ӆ
���ā�n��ԗ'Q h�$�0P�5��V/�f|Q���%�r<� m�N}ɷ�Y(4�Ԉ��n�OSa�4͏f���҂��m���ܴ�����S�I�ܴ_6��ɰ� �Hz�H��eg\����B~�j�>�M3##�(T(tuZ-�|V���g�O�<�ˋ;���"�	;��+�,�Mܓ���6�Sk��ٸ	!HE[�n�J��[��έ�y�iE#H6jw��~�XŒ����d�<9����O'哝	�)�g���r4���e@>B�C�I�e�����V�	�Ⴔ�Ў%d��	�䓗�퓣l��@ˇ��)�f5�G	;D�C�)� ��8S':@q����bK�)�$>O�=E��g���Q�`C@�\'�L�al���'x��'o�?��u-]H�LQ�0�ښrf}�E�5D�������������.�
�H�H3D� b�)ʓ*����fI�8��q�Շ0D���Ҏ1���0��jG��:�ꯟ��I�4J��*�S�F�j1%��5�C�	F8��1r����Ƃ	z�C�ɖ~�QQ���3[~��v
�)C76�=��'��>��r`�y������-G�>�Sf,D�@[���o�H��4�Oa��Rqw���Fz���ip��Z�+N6Fu��bs	�>-�L!���!�|�μz��I3'n$,���R*X8 �ȓqʅ�CX!}R��X��?���	F~b�W~�pd��t8��jd\��y2�Y)�
I���v���"d+0���O��$p�d�?�����rhř/�	Bpk�_H�T2�"O���\�vA4�"�*VA�`æ�O���$P�(�i��� A���Y$"��8ڑ��F��M� 5Lȴ
�$�K)�M �l���y"O�6G��ۧ��"�b��lѝ�~r�~��y��3U�	PǦ8.�Ѹ���!�y2E��S>�1��z�l���C���$xx�8����au<����"�q	,D�����S��d
\p�@P����<���:@�ȫѢև)*L<z6jD�^M�C�	�� \��ۥV�d���$B�ed#<ٔ�'�\����U>�p��!�Q=����'N0�����F�0�1��&L��$B�'�l9aÂ�N��E!�N��D��@��'�ў�}��@T�{�&`ѣ�ŗN%�@��S�<��,]�]�0(Ҡߏd
-h��Rj�<��	..��Er��N-%�T��H�z�<�`-�
�֌�&
�0��U�פ��<�
,�� 1$A�-��lôz�<a,U.��T F�n��~�<����}�,�֤�󅔦Q�q�Ie�������;0%��ʗX� �ch6D��z$A�3e
���!W������ D���m�(=���SiZ�y�Qv%$�O��M}R����Ҩ�d�8�!�4]���	V������ �
C�R�Z	���:DƑl�2D�|ڤś�7o4\�����{��M���0?��LCJ���&}92��CMu����hO��l�ɒ!D�R��ΛI>qI�$��I9B�ɣi���+�&ּN�4�T��>m�LC�I�D&�t*��ǰ!��{���>@��C䉹O�!���հ �i��;!��C�	aф<C���
��	��0ْC�I�~X�i�u�Y�dݢ�M[�0f����#C�U��
��/�V��p��4V�`#<�	�?��rFDZ���C(X��<i�"��I��Q1d�C����ȓhۜ��l��vC���͍�x. ���Q��́��!Z��%�0#�<A�6��?�v�5�S�� !C\h1��R7�J賐×e��'�ўb?�����F��!Kؚ a� aK�w�<�1�'U��|�Ѐ���i(G/���D{���S�v1���Ka��T���P#�j����I72=b�k
�%� �С��	Df��p<aO>��(ҒuBJ��u�8�,]:E�}�<q�I[-&�H����I�P��/�w̓�M�f[{���S<$!^]����0��Û/�\�<ɄG1��ܨqD�0Ѻ��'h��:i��w"O� DE�qm�.8��w�VP�ͨ��I\�OԌ��V+�7��9 C"Kj0L���'ar��;Z�dA{�(7 ��$
��G���>1�O\5Yb�؜a�>@�T�3�"��3�'d�'޶����w���@�e>"j�4���p=�a,��%���e�4|���]�<y�&��a�@q$�,$�Icd@�Ԧ�F{���i~�@� .��@�d ��.�B`���hO?Qs"ɴX��m�Af�*/J���"+c�<�AIB�vTj��*@("�q��`ܓ��=��\�hİC���@��pk�Ò_x��)/O�D���X�oV ��UE�<� Iۧ�']���_�Or}���&|^�4�V7&��H��|b�)�<y���1|!:�pĩ�? ̈�'��tH��?��@�*]����1�)�C�q@~B�;
$Dr��

��JI9�B�I)!��$rP�Ef�4����7|[|��?Ɋ��?��Qʊ�|cH2�d�8n����8D�<���R< j��cb+!�b|� "B�'��>�	�j�>�� K�-2��#FFD8�jC�n�����[�r����?!��o�m�������?u�A�O�g����d5�p>AK<�W��2a�✱K�#A�J�!���o�{8�hKqA�,p���B'zx��F+!D�b�*�-[Ɔ�p"��k;$H��+D�0@��{�p�;t#@#pk���J(D����ϥ.�t���^�b����%�O��O�,���.(�Mspct����"O���rM�5i�p!�0"�Vmr���Ic���՛#�"�S�ļ;6½uG�8!�$A �v�Z3�4a$|�#f`�b!�dS*�$��'�)Q4�X���8j!�D�-�h�B 2=r p� �G�!򤂖B���(��U�D\ѻ��A��!��R
��%�Ѯ��l�4DzE&[.}^!�>"�\��W��o�����CN�Mb!�	�q�� p#U�"����I�z�!�ˑE�4��u��b"X�j#(�:wx!�D��D0��JAG�/ RGm$=a!��C3��s��O5[�T	p��!�d�|t��!� �<���vZ��!���$c*��3,[�.���j�=u!�$
�x��Ia�5=�\�3�H6e!�D��U �2%��)�@��bN!�C�y�h��B��k�5���~4!��͚IH!'`�|���q�ʯ!�$[�3�����8I�v�2�)��!���p�Ҽ�b���$H�F���!�W��KEIه{+V�TF���!��8�fa`��ُt
�)��A��!�䎕Au*Eʤ��(%�@�8T�!򤃒7����CL!J�="���$~�!��[�u`FAh�Ø�r�Js�͚�!���10��m�%M�:Ȳ�cd�qp!����u�u���)f�xܠ4��!��J7n�X�R�;��mk�D1
!��ص9Rl���LB�'�!з��9�!��j�Z�׎�.����Ⱦ]�!��0G� 0!D��в�+�� �!�D�v��B����Q��s2-N�@�!�HH����
���@uɜ	�!���2kl æ�<xŨ�n�a�!�$�h"Fh �)G�W��`լK�N=!� O<0�G@ �f`��fU\!�� ����i�;
.Z}��	^��Y6"ON�D�<���.��\`"O��E�r-�uGۑJ��y#�"Oj�q��-g_���e�4 �9�"O��
Tû;Ms�i���{��'q��'q�'���'"��'~b�'��g��`)�Q�Qύ�p�`�E�'�'pR�'�"�'��'h��' �1bH�;�� �9U��q���'g��'L2�'���'7R�'oR�'c��y�a�P�xy�b��)d�5�e�'��'&��'�R�'�2�'���'�p���!hą��s���9��'��'���'���'R��'�r�'����_� xTd÷��I�^`���'l�'kB�'���'"��'�"�'o���NW�Nf��$_%T��۰�'���'G2�'�R�' ��'�R�'�����݈R��	k�bIA�9�d�'|��'fB�'z"�'���'�r�'DF�"#.�9t1U�Ad�f�&�'J��'S��'���'���'��'	�p�\7�d"���:@1J9z�'F2�'Z��'���'���'�R�'�Ry�#*�:�@�iU��&:S��	'�'���'�b�'���'�2�'Y��'����OP�t|�1�� \����'��'���'��'j��'Vb�'���:�mT$N�mSC��%bC��'�2�'o�'�b�'���p�����O��="Sv��FE�e�!���AIy��'��)�3?���iҸ}+��X����5���x �[���$N�=�?��<ѽi������ %+HYX�5/訓'jӔ���0%
p7M>?SgT�)�8L�b�(��ҭoI��ǆP�(�h��-���'�]� E��Κ�	�ҙK4B {J�@���k��7mT:N�1O��?�����{�Z?T��E�6.�7v�!�2C��g}���qӀ�	]}��4��>H���7O�5z@A�qI��0p�X,x��9p=O��bD�/��
u�*��|j�T� �`Q�o���p3��?��͓���-���ަ��W�$�	�RH�r�Vc&|�!��f��D�?�"_�H�ڴjǛ�<O��,;P�ȅ�����ъ�iI��'
<�Au�W�?�hڈ��֦'9�n֟ ���a���Zŧ��<<h9Ԃ@ry�[�l�)��<)c�Yr����s{=9"?O1mZ��F�_I�6�4�ƌqV�0�6p8�f��$��{�?ONoڶ�M3��m��Bܴ�����t B�+P�L�O8�
�풺v� �)1L8�l���#���<�|�<�#�a�6 ��//����U��z~r�w��8G��O����Of�?Q�o�� 	^�0ơV(m2�E��#���L���4���|
���?ɓ�>Tp��Bс	�?����F�G�p�(3v�Q
��D������Xj)R�O�ʓ ���7J�1:�܄
3�V"V�|$��	��M�ԍK��?���ܔ%E��AG)�@����R!�?餷i��O��'�.6Ѧ���4m�"�p�,BN-��(&����`�\�=�@Γ�?iBo�� �~�����$ퟴ�b�)��a�R�K}��A(_��"*4x����=z�bt�#���!�U�WE��C��D"K$��/9�đ3C�N&Jh0$��٩bf�apS�<9����E�E�4�mʧ%��%��I��ȪRXn��S�\#v\��@R(�)O�j	�쁮|T�x�a�,Jz��d(�%z�FX.;s�U"��*'y�R�H6z7���^"6�Qa�6o��9��ǌ(}��9���A��8���i�ز��ݛ)품�%
�
ꨙZPċ&a���y��U���sH׼=�D�9ENS� "�ʘ�#���ڴ�?����?���5���O������O��y��P���͐!�;f3b��d����z�(�O���O���]�QH�L�w��U��c��̦9��lZٟde��jy��'a��'�ɧ5�怠
-hͱ�HI={I:�D-���'tM�Od�D�Oz�D�<qE	�pݐҧI(e~�9�2����j��)O���Op�$"�$�Or��RDQQ�B�3�d�t�	����A� �ǟH����P�'B��;C֟*y·`]�Q���v A25� ��i�r�'S��|b�'R2EBW�d ��Rфܠk���ިm��Ɵ����h�'Fr�D]>y�I�=T��օ�xuHM��A"�ڌ��4�?aO>���?	5��t�%��u0ǤV;u[.��⎅d���o����eybÕB�������?5� ,�K:v1��i��Y���p�*����?���o�������1�df�".qv9�v
�d���I��i��I�)�h���џD�I֟��vyZc��#
	�%�5o�h�.��޴�?	�C5�Fx��$�پ�B�E��O�>��D��M;���?����?Y����9O����O��p*$J����7Gݙ�z��idǓp�S�O���i���KK���Ȃ+�X>*6M�O(���O��;s��<����?����~R�6=`���@� .��r!��"��'�ȭ���|2�'�B�'��x����7
�,�ꉺO��	 �j�>�d�W�˓�?���?M>��y ʕ��8D�$a�';p4ވ�'x"4��''�I����П��'��xy0mA$3��0�S�A/f/�A������	�����@'������[��X "�V�UO�S�r��Y�tX@$������|��Ay�Nǵm���ȠL��pʲg��x�t-{p�D˛��']�'/�'\�'ƨ��O x�S�0h
���C�'Bt]���	�����`y�+�W���ة
� �\�F�	�8b�t�6��t`�	ԻiX�|�'Y���qO�h�� X*M=p�A!VD
0��i��'�>G�ؔO��'��Ta5o�6�iN�7C�����A�P��Of��Ol����<��~��B��(��YL�����oC򦍗'pJ1Z��~�$�O��O���J�N� !l_�Z$6��gʡM�`n�ɟ��I���I
���<�*��F��X�0%c��N��`���E��M�bӣ�&�'k"�'F��!�4�k�I	��Їk՟cߌ����ҪN���'���'��Y����DZY���P�{�T;#ҭm���m����џ�9��\$���|j���?�Vʏ(~_h�+�ș7o��Jw�Kzϛv�'���'h���~�'B�'���AC�G�tr��^��8�.�|��7�O���L�H�i>%�	ԟ��'�x �����"�v�X�H�ZΜ����w�p�d �X)H�d�<���?����9E)0"��$��y�Dpᔌ��#�c�	ȟ,����ė'!��'
T�S!4��`x�&L2Z�HtA`���Z�L�	Ɵ���ky�V��@�Ӛm90�ȡ��!La�$2ōB�B��?��?�+O��$�O��s�f�O$`���߉rƈl��G�]B�p��h}R�'�Y���I�?���O��ġH�ᩑ�nu��G�07�?�	�����,J6|�C"*8�D�]Ut!۱��%8�BЃ�S���'	W�`�』��'�?!����@̳�V��8~���馍�'7��'�l���'��Or�\c�СvD� pX��A
�7�����O����	
E����Od���Ot�I�<��Z@�]����-wo��
��j�`�m��T�	�~��A(��'�)��.0�ޔBa�K�	�Q²��66ĿX?�|m䟨�I͟p�#���|�1d�9�q͗8.ʂ��"(���nڶ>�M��ڟ����� ��o��'���ɉT^��±�G�;�IqF��N7��O����OX�i�i>%������׭ڝ/h�"���B~��9�o���M����?Q��;D�1��Y?ݖOA�O2�yB�8�<p�7�ؑ��$ڤ�M��_R",�/O��O��O���B�U�[$.Qa��ӷ:�R5룬M]}��B  c@(J�y��'!�	۟DI��կ���P��ZR:��aH�DVt��'��'H�O��$�O6�[U���L����d`���%��+�4�7�d�Oʓ�?�dW��� �#�Ubb� ������M���?i���'���3= ��ڴ��P�C�i�6��IŅPz(�%����Yy��'6Hq��Y>9�� բ���B��a�n=I�C[�K9NQ۴��'D�S���G�$�P/d��D`@��yԔi�ӷ����'B2_�\�I��ħ�?Y��{����U2��� ��쑷H���y�'�2�'(�'���yZc-L1³�F<|�,�	cL!3D�l�ߴ��$Zt^�m���I�OZ��Y~�nW:V�r�����V�4�K'�_�MC��?q���?����'��s�~��򯕓H�Av�ǦV������i����2�a�(���O��D㟖5$��s�ձ�+N=$�dKp�T)dM��{�<iB�@�O����O�����,��<��Uq�y�"�D��ŉ!	FP�$0I'�i��'9� ��-�6-�O���O��$�O�.����M\��GW0I���'��X�0�)*���?����(�r�ECe��2��8H�	�1�iS�"�+�@7-�O��D�O���h�$�O�@���3w�]�w����`i��Q�$a��e�`�	ğh�Iԟ��IƟD�	���3gu��t�E�=�x0s��M+��?����?1�W?]�'lR��
�~��301�a�%�#�h�yr�'�'"�'��0��m���`�Q?.y�RjS���H@M�ͦ�������ן,�I`y��'��0�O�Z`����v��kUl��%z^��'�q����O����O�D�O�09������'"��2Q��ϒO���e��_>7��O���O@��?13��|B-O6d��i��b�L��V��m%>	cS��ۦ���۟��矬�gѪ�M;���?�����b����8�0���N��hsT�i�U�p��X��Sן�����4��dJ���,YdfZ'~�uoZޟ��I�Z���ܴ�?���?��'�b��C�
�P����?��Y�S
�By#c_����2~�\�'��i>�Ӻs��ײoV��T%]:�r]�%ӦI��o� �M��?Y����'�?9���?9�L�73H�k`�%�h���<9��K�HL"�'�+�~bJ~J��63�1!t�
�wL���T+�t���i�r�'��τ��46��O"���O6�$�O���[҄Q`u�E/RNԭat�܊1�v�'��	����)����?��O�*t�hܾTa���H��%Rva��4�?yB-H�DC���'���'.�i�~��'��!�!�fg&-q�ϻF]qٴ�?�ɇ�<1/O����O>���O���:�=0�N[�ͼx ����=�!�æm�	ʟ��I⟔`�����?��),;�P̊���
�( 릀Q�aҎ�ϓ���O��d�Oh���O"�b$hE����L�X-H��w�ֽq�����M��?	���?Y�����O����5�<��=n���;�h��)�>o� J�O����O\���Ol���6Y�po���8��qJ����n����,a��L:ڴ�?a��?i*O��DL17Y���O$�	��>�B��K�~���U Bz6��O�ķ<�)�
-��O�r�O�>!�� 	1YV�
��\�H��eq��8��O��d��5��+�T?��R&]�.�1�EZ�;�,y�h���dqxiH��i̊꧆?���J�)� ��pG�f,�ԛbٛT� Ҹi���'�x�q��'Cɧ�O:�@��
t1�@�zE�۴R����տiB�'R�ON�O���(�����ɶhL�	 /ּ�*9o�/�P��v�)�'�?��/�ZL�4� W+lYh����lΛV�'��'`"�9�$�O�������ۣbM�x{G��<iK8�cQ�:��1?��&�D�����	.of꠰2g��ZY���R0Ds6��ߴ�?��J�.W0�')�'�ɧ5�@�iW���� Z�4=�	H;����1Oh���ON�ĩ<)�ܚ{~JЁ2l�
u���F�s��yЗxb�'{�|r�'z��Ŷ��A��ٗc�t��rK4D�4+�'����l�	a�ӄ}�>0�OGPd&��g�`Ұ��8.��)�O��$�O�O���O S�-��<�SB�x�<�a��&����O�>���?����E5�d}$>��%H�yq�8�LS1���M�����?����m���h�<�+&�ǻJ�V 0���y�7��O��$�<qSk±�O�"�O�<��S��;<䤩�c��F�L����"�d�O����n7���9�h��S	Mn\(��<XVڥnZmyB�&�7m^j���'H�DO>?�� �q���ؤ�^/Hx��3�+S���֟Ġ��d�|&�b?qۀ��hּZrM.+���3bw����bLOצ��IƟ����?	�J<��O:D��N��� �WF���mU.�MCa
�<9K>E���'��ő�Y�>B:�+&#R�0��,#5Is�,�d�Ob�D�g��d&����ޟ��'��ӑ�LSz.��W,�-"Dn�c�,'�@�L|����?��F�Bݒc"��`���5��*A8����it��E�RF O����O��Ok�% ��i��
>,X&�Y�@R����&2��byr�'�����׏b�p��D/�!tz��������ve7�d�Ox��(�D�Oz�d;-b2%�G' G �H�Ė@�͛2�O�˓�?����?q/O1pE�|�D�Ĩ*g�Ѓpo^	{��|QsIy}R�'�Җ|B�'��B��iRb�wxZ4�� ��T�c�D;����?����?�.OfQʲBLJ�Ӟ�f�� ��x6�b0gƥ8[R���4�?K>����?��OE�c�2YJĢ�R��h@u�L$5m����]y�"M1Cq*������Y!j
�u�3B�UǜD� �L���<�	�t�����w�~"�	���ZV�
'�~H�5H]�%�'vZ��/bӄ��O�"�O$�L����х�4T1�NĽ���'���|&/����ү��Aƶ���9F����id�Iq�'*b�'p��O��\����P��k��C���mp��0R��6ML���S����B0b���X�y��s�0LqN��M[��?a��;@�)F�x�OR�'
��uc��w���F�=n�0��>��6
$c����ӟd���(h-��!z��(r�f�71h:�ߴ�?����?���V��S؟ &�(���Κ-<���ŏ����"�|��'�v�b����d�O��d�O�˓s�^�7�Ǜ&Bj��d��sV�`�P
���'��'�'��'&��D@�`��	�%�Y/9uZa�D� Ϙ'5��'&�^��ksbX���4jE:M6!9.�i�t�[@����D�OF�$?�d�OD���8�	!'D�����m~�i��ݵZO"��?����?q*O��z��RU��>�z��7�/<�`\��C#d���4�?aM>Q���?ɃAV�Gl8#	rM<E���5{��l՟l��gy"k^=������T���-L���M�^<*E�BMP�	۟P�	=�p"<�O�DV�Ӝ';�=�s^n~y��4��d-L�}l���	�O^��G~B��efU9�l�]l���#���Mk��?�j���O4t�WhHr���p�Mx$�J�4;�V�Ħ���Ο��	�?}�H<I��@��,�.x^t�P0A;i��g�i_@�[�����^����ci�!8�rT��M����?�jA`�s(O�˧�?��'����e��~d��r�FܲcV�b�.�I�� M|B��?��Yµ:���� �*,�a�4*�I#�iRbN��O��O��$-}���5?F�P�"�b�h@��L���^�g�1O,��O��$�O�dY�O],��N��*	s���<�R���O��$�ON�$�O(�OL���8��yj9��EC�\��m��Dm�@<8a���I֟��	^y��0����=v�H�wM
���iů�J���?y����?q��C@�`�'�T�:S��]@����I5���ɩOl���O���<ѧ�W5N��O����ш�\�J���O�H˘D�P	f����0���O���X�ұO�99ǒI��L�0�J�c�
���iD�'b�'��Q�R�'���'���O��J@e�v=�aV��F��d2��>��O���4#lV�K5�T?�p�P;n���F�!6Ҭa�h���h$�P餶iy��'�?���2i�I�9XZ�v�:p�J 7�WM;�O���3O4�i>O.�Z2
F1��M��C�&#�Hh)��iؔ�2�'�2�'���O1r�'G�ӂQ ��P�	ny��ⴭD�`(Hb�O��0��)����Qg'ܾ�`���\�A;֤#C��5�M����?1����-{��xB�'d��O� ����BF�c��퐖�	$BI�����$�@�1O$�$�O ����F���3g�;>Q�0��k�j��n�۟�z1舩���?�������H �1}Pp[0�X��	��p}�.Bǘ'B��'�_�8p��h���f� �@#�/P�`x�!�N<���?�H>����?i(�$������3d?H���D�$��P�<���?q����^l{B��'r����֋*z���84��35δ�'�2�'��'�":O��s�O�x����/�(@ �":!9$�� Y�|�I��IEy2��:hV���sԢ��C��� ��<���0���릱��Y������	�vc�(I"
>�����f��a���JB�r���D�O��TTj�I���D�'D�#��^�x�An=Ӽ8�����O����O"MG�~z��C-0��Y �=�}��G�y�'� �[��{�0T�O`��O����8�9��T'"��%�S�0t�\�mZ矜��_d#<�~z������é�*D�:=3'�Ħ!Zt,ޗ�M���?��:��x�'��і�Q���,Ӄk*q0��`�:��q�)§�?	ňA(!z�,�6捕7�0��1A ���'���'="t�Y�X�O\�O<mID@[�L�(I�ҠG�nƥ�� i�'(������O&���XI&��f_���˗>S�Jeo�� `W	��M����?i��?�1V?�F�]���B�-y���A�W?�Z}&��%���ן8����$lc�{7KR�^��*�⋐���a��xy2�'GB�'��'FR�O� ��N�T�u&/~8��i?�$��O����O����O���)V�l��0��4 QL�)2��6���hHsٴ�?���?Y���?!(O>��̓1_�i 	V���pr��	{|�9��!ڿ�8lZ�������	ߟ��	 E���h�4�?��t?�L3r�)#��4a��Û}���°i'b�'�BP���	���������M�p���P���
�@!eDF�oٟ���ԟ��I�B�(A3޴�?���?��'�V�`s�U�b4�A��X�v��I(F�im�S���� ���O�i>7P�Y���as$����H� �(��&�'mB�|d6�Ot���O������� !:�@j�&��;��
,S��'�rFm��'ybS>e��΅�3Ç�S�HY1�ԛ.'�1��i��x�Bav�����O������I�OF���O���F팙�z4��!��FW���撚+��ϟ8%��O����0�,΋h�����:vN��ʳ>�M���?�� �0�i~��'��'Zw]<8h!CBMҩ�&��e��Īܴ�?�)OK]��yʟ �$�O���A8���0�Ϛy\�cP��t��hm���$�0m�&�M���?A��?Y$\?��� �v"2dC�d��
�{���'\�*�'�r�'r�'��'vrO�S�A1�gޞ+�|LQw���X7X��������O<���Ov��O���՟�[�͍�%�V�҂A�:B�	#���/�>�	oy��'ABZ>��������ڴ{K,�A��]�LȖi��˕�d����i2�'>�'�"^���I�\��s��(KѧI�?A�p�*΢6���ֱi+b�'���'���'�ڍY��u�����OD���c�R 9�@[�bA#����)�����Sy��'TP��OM��O��He)��dg�x S��(��P��i���'a�'�J@�rӐ�$�O��d�rY.d�H����u2"@"@OS�G.�Im�П�'�R�[�����'�i>7�Ĝ+wr�h��שs�����K<�f�',�@Ӫ:WV7M�O����Oz�������(��ea�Țv��*�&cy���'F�ҚsX��'��i>a��蜚�
�1
�ބ���b8 ����i}���u�����O��$������Ot�$�OP�t�G�5ln�� �*���&�ݦ����D%��m�埐�F�sSb	���%�h��B���M����?��B+���v�i���'�R�'�Zw�`͡р��U ���C������4�?�/O.Y��1O��֟(����ȡ1�^�)�|³�ُ4�vܩ���M3���m;��ivr�'���'���'�~�B��:�J�05��!,�`R�) 4��D�h��O����Ob�$�O8�'i�L��L���ˠ$�	o�b�Ӏ`
S\�&�'�B�'{b��~�(O��d��u ���M�V6<�@�*[;SOZ�C�2O���?����?a���?���"�!�\�CR	�M"�o�b��7-�O8���O����O�˓�?��,�|�
�R���s��µQ��}�K"}��v�'��'���'����`KX7m�O����? =6qbT��{�rHjc�M�;x
�n�����	ΟH�'�򯗽��D�'���#<'Np�v�G�er�x�pf�j�J�Kp��Z���%��3�A��e�
���y�!�@솂k1
D��f����p'$D�гP���2f*�+a)[!7|������=	0�h��C���)��K�{�Čs��S�<{�+pk�)%Y�Z��7T	+��Wk�+s T�(*H��'��h����s!�s��B$�ck
�jV�Z2: ��%_�:s� Q���&s����t��L���!S��
$��bG�]�u�� hw	��U��E<���S�O�,�	̟����u7�K g��a(U�P	�:�� �U7f�sv.Q�R��}l�y�2�a7N*�3�d��@Gf�6�6!(`cE�������Dd��ش'w�聡�:�3�ˌH����Ŋ3GͺH#��0-��l�&��Ě�+�����?a�ql��� j!��}Ō���'�Xs$)�n��%�u蜯W��p��O&Dz�]>ݖ'�.-RO�@� ��♱HU�	˂��� s��b��'r�'�ro�~������Y�? \9���Eji�mj���mJLx���0uc�,���a��  ��ȟG���*���;rj2ٱ�Mܖ/�<r` ſt���R A��%�%����'0&�@ڤn6s�M ѭQ�?R&�'�H(�m�7!b���BA��PMV�\� ���OP���Ol��?��B�
�v�܍Q�A��w���B_��0>iN>)���d�r�B�2S!T	A�E\`̓,ޛ��'���9 m������Z�!
��W�,C�,�$f�f0���O�����O�>��t�7-n2��Ub_�?"Ai!�=5����,0 �*U�X�x���,��CFD;n����t� 0r�Jʵ��>Įm�D�¥����	+�Z�$���]��O~EJ �R� �ڹ�wF�'*z��@'��O��󤍋D�NɋV醲�ح��H<f�!�DR��=YG��H����a�����R���D�<�c�ނ6]�F�'i�U>I�d�Qџ���4o�5af R/�~\�1*�ϟ��I�Ei����ˏ/�"l� ���\"�H�&^���X�O�8�Ӓ�'k�PS#o.(��`�J�4�e�҂z1v�F�Y?@3.��4��X	���C[5��Nȼ�
٤9	�����9�ĦO413�'�O�6I5�Oh�¹�կӼ*�@��"O��B�FQ2*(�0�X�f��G�(��|�c�ɬ�jB��im�T3��΀	�j�b�Ot�D�O�H��Ɔ4R�d�Oj���O�nX:jvЫ���
T��\"�l`U��/��I�� �� ��O�e9���<a��E��J�ïB
� EY�A�a��҃,	��*Ԩ�/^�7v��!�*�8���!��(b�y��i�k�����(�?ATx���ٟ��Iߟ� D��>˓�?�4�X�@�J��u`˷g��S������x���B�"��rٮd�ޱ���A��y��'�n"=I���?�-Op��e�/z�T�L�4H�be�c`	i�%br��O����O����o�D�'���Β�t�pE�ͷ~�X�& �9�����ϖpK��eG��ke�v���C�}k��	#&�Y�ċ�?#��%c2F����hA���6z��C@��cZ7�[��嚵�ӢLf��:M>����52�!��ަUE����"[D��	����	ʟT�'���$Ov�PX��V�����Bka|�|ҏ�<=��Qc_��D��B��' �6-�O˓mJ���]�P�	� �&�T%�KNl�ub� 	j��Iʟ��QB�ş8�	�|:�Î�%��V�#?N ���:=
����P��!qdǼqZt���~�֣<q�� ��)XR�˼G6F<ӳ!�_ӲE+��0�!���x�����W)F���<iT̟���Ο��I�� �yD-��J�l:Ն�#�ll�'2�ᓐ �85��≻l�@Ķl�NB�I/�M�#ǆ��H{A`^�Bt(���?i*OT a�Nߦ�Ɵ��Os8Y���'xޱbBHu�R����Z7:� �{W�'�rM_$7�pŢb�εT:%sQ�u��U�����}��5��Q�]��� �ߏ
��T^@�dG�,52y`�	�� �� �	�$YP��D�Nu�H������!� �	��M�%��?M��^Yo����!6�D
���wh<R���1��3�Q <Dx��2,QQ�pr��͠i�Cg�	mr��R�〲[^�t�'|��'%"�A�/ �R�'R�'h8�?W:�(�)�yx�i7kO���t3��PV����+n���F�?�3�D�7B}:�X���"�.�ڀ�6|�$X
�!ޑb��D�+��]
��L>y�G��N�*,[v�Qc���P�kݙs{�V�<�ԧǟ�S�?%�?�'��-��Bd�<���X2�P�<A���d����KM6��	6#�E~Ҏ(�	��	ky"$� ��-d�2�T��K�v(��H��I�Gg2�'���'����ڟ���柤�0�@�fJ2��EJ%�����A_���	h�"W$x>L����' �BQ�b�>{\��r� �����=��|��f�R�z/$*5r���p��L`�&R�N-6����U>���	x�.��ฑ��\�Y2c$B�C�p��<ٔ˝N�� ��[-�fd�7�0�z	1S!��@�_z�6�'�S?jG�ګ����"{��\Cf�ՈhkЈ[qV�m��D�OP�e��Oz��}>ZE�ثiFZ0M��Z�x�#�OV!ּm���-i���;Wh�'M��G��W0�|IZ��X4��dȉ�/�����M�"��!*�� 2�I�7I.���O8�r�"���b
�H�����
�VM�<Q���<�Ԡ��y:�<pc.1:�vL�P�\u<i#�i�f$�SaZ�v���e�B"�h�k�'H�	�$Rؐ��4�?�����B����@0Vk�L#��Ô]�\(4B\�|����Ol���ͅt����)a����c�|/��IqM��؃��,��i�>q⁚�Y^h��� ��{LF͒ G�	�mQN|���C��ּ����,1v��(�O�ćYJ��'��O�O����$@լ1N����0�
M��y�'��ybd		��e"�nn�� �f��0<���[�!�KM�%]xE8p�*c
nH�O2��Op�p�� ��
���O���O��N:�6D �,��/�f�����{�2<ґm�y�5�⭘oH�d�w�.��X)f�ٔ;O� ��1t�B�a����5)�Fc�q�1�S7�@��]�ƕZ$\�Ͳx@� �e�4�]J�λrZ��yp'�?,���!')�%��h�������)K�O"�d�)�>1��N4:g�
�f�J+!���IG��Pu���3Q,EKwfM��$�O�DzBoz�.�d�<�T(P�s0ҔP����bG*�2�ŀ�=�j��#� ��?���?Y��p1�L6M�O|��?`��<����L�L���DT)gXY��$!h�Z)��"����@��U�V���*r&T@�2S�2\�g��>		AGF3-yp�i`�դ!`�铋���q�1_��'���qj9SA�
;i� �Y�Ҭ.k2k��'lҔ|�'b2�$\-Yz�H��C��W�!SrV�V�a|�|b�H�8�tY ��O�h$��+�3��'�T7��O�]ٶ%�Z�(�	�dg��s�Si�fͨ�b\9mL�d�I���#���ϟ��I�|�T��"H��%����V"��3UA�H�6y��?K���� �!W ~���DQp����ō�����C��wml���`K��-4jʆ-O����@+�-P���I�����ß,BG�<&nREC\�i@X[��GSyb�'Q�O>�:gn��<UJ��g�[�Wz�ɫ4�%�t�ش
~�hC!Ҡ �h��@�.9��=̓���ƹ�̘�'%2U>1�K�ʟ�c��T�3���X�»`$kᡞ��D���t��
���2{(Y*1X �,Qq��&TK��O��"�Mg6� �i�$J�P;N�d� ޢ~�r؈ej�B&�IA�.��!�	�/�]�b��;k���k����v���h�.Y��Oz��'��6��`�O���G_,E���P�\+������&(����A�{�(�En�)��@f &4��=ͧu|�� T��7���hӢ]BF�P���M�����>YW��N��8���Z�>�6�Cэ��<��-8� �kS�[����`�q�<��֐tM�M�4g�3�ĔJb�Pj�<�FɆ�P1���0g�tu�f[b�<95� [28�6�\�\ ��Z�<a�-�	_0A�л적`(�A�<��-�%W�앙��\�3�l�1M[@�<�g%W
0��U�a�X���C���|�<��G�
ũ��^���MkW�u�<��ΐpD��+C�Ņ;^F-c Kr�<���2~IX�y��j�<5����l�<��AX�m%X<����Nyƕ�dFVO�<���\�Ta*��t�v���oNA�<	��\i�� �]햬ˀ�~�<)&�D;h�T�����&e�<�e^~.�(��ѿ�K�*	Y�B�	�*8�LK�-F�{��K�Œ$H�B�	5"ȴ����5�a�F�R=hUtB�	�-�S�ӼF��ؔG?B��B�ɣY��=
������c#^8�LB�	6/��xi�JMʌAx\>+C�	/0w��;3)ƞn���4ۺ%��B�	=�(���B�b��T� ჭTc�B䉘w�Lu����!,��;��W.�jB䉸ih��#
�p:������`�"C�ɐ$�(h���#򬜈��=y�C�ILp�����վ�� JZ�a`�B�I= /ܩ���U���Q$�X���B�	�W�nc�ꛫ;�T�p�+�&J,����J� G|}�Ff+���'�O6P`�H�>�2�W>i�X�E#U�Gܞ���m	j��K͂Z)J=��$�/�PH�#�/Pd�A�	�6,u����.���$
�eG��(7�C��`�%��Q��FBU�t�K�$�#���d)�TT�G�>5%�gc���ʱjK>����Zw4�ܒ' ��vDI`�OR>hȘ��F��9�RD}bO�$6}$䁂��	����ꜶgO�	�G��i������*(�hy�� ?�,����	搘�⍔#��׽<���+�y�퐘_P$ԣT�W�[!�}+CI�ޘ'��|)GA�Y��MR
�z$��t��'��m@Bbz�e�Q���p�8�a�/� ,@���K���Н<���Z�����M���]�����8Q恒��W5�,Y�M�ahi�xT�Ƃa^��$o>�������$18���H�<��$�e�"0A�P��MK��Q3V�J�>1��5k��Â͘�FVJ��CΟ�S����O���B^Z���B'%��s�HH�P}�g 6	����\,��(�%�(�a�ԣ�!Zn���;6�^x��$ lK���$)�!*�X�'��,�2�'�則K�� �'�T����+��+1�&� A�կ��}� ��yҧ��Q�����̑R�n�cv$���� �����ЄR�D�
'd	y�8��I�ha�=80��Q9�[J�E��I/-5�H�w
Px��)rw�߬_���VK��=' ԃCG�7g���$R�!>|s��7BR�K�ǚ59v�K�7�pA$,����X�g/B��O���_M�N,�G͋��H��"O���
S^�tQ��[������gڽn)04��D�yѾT�fO��͎H�x��K�2�ƹ�6�I?n��}2�Y.s��*����yc��3f��C����nqOP��LK$w���������|"���,,
�×�.�>]a�'���0<aU��L.�q3��#~Q$��ACT�~� "� �q�݊ujGҺ��C� f�0�S��ˍ'v��%���>��! ��?��'��Q��N'R��0��"ؙ}���1I�dc��U�s{z�+g���uJ2��@ �	gT�����)j�>P�S,�-X��0sB@�8N������w8����pt(rUN�vL�x�g�Z~T1I�exbìL��(O�%8o��DJ��@�Ѻ1DȆDs(�	Am�3fX�'�̣��'hθ!E��c4n�Q��'`Oh��΃>Ř�⅊*`��@���>��0,.�a���%O��0!��5@&��@m<{�,H6O�|�����\�28��M�c��D�t�W:,�xҧ���g�l�!��>��y�$ؘPGȡ��C�'�T���]0�I��8^�(�(tJ[�L��a�y>���3��ɸ��$�3��2|m,��X�I�h�b��O��W�� tƜD�	V��%�7��8�@c��;^�����?K>��7�^�4,@��'X��[��>���2�B�y���C���ÂH�k�l�6I�+{��p%m�,lD���ц(�Y���;O��ō&F��E� �a�Kbj+kp��R�'���0�ď�V��{yʟLpY����Y[r$��ᑟj����`6ړܖ��ghƶ\I�x���#n�P���&?��a��0�`�	79hI�GX�H�O�xhlZ�w`�#�H��%�U$_��^�d�N:��d PGqӊ�I�Iȋ@L�Kè�<�{�I�L��)H³�d�	5HM
y��S�nǓEH��he�'�Ą�GIH21efmZ<]-���b��Pz(K"��W�[�n�-mD`,�̌!V�^t��O�q�	�D7^�z�O��!s�ԨU��uW�n�q&i�>8dB@F�ǗB�ȱ�� V�G.$�CH���V���  �!��?t �7���(a��O�����\?� Gg��\�'�?%��O��|z�j���!pt.F;,��]0p�v�'д�[1@��=x98��z.���tM��o����\re������Ӣ�Y�'Ӝs\X���OΘ�g�S��_�4��Qb@��U؎(�G�C��M�v��2s����1ept���������8�=�Q�E��R5mOpț�ӗg�*��=E��4g�j�IgEԥIXj�):(@&�sң�4�D]����^�'C"�C��yǨ[�p#HmZ&�U���K"����d���#?!�LT�a�t)�N�9-�,C(�$��ಇ��s��;f���Z�[�,@�}�qO
	h%J������9of�z`�ɊG
j!B�?9����/�6���R��]�)�o�d�Q��S/A ,��Ea�%1���R@=%�8�����s�%���;5bU�X���R�N|7`�Yf̟�V���'ў@r��;r���p�e�6) 4c��W�B��#~ 4%��ЪU�����P�&��<�H�O
�=ͧi|n�BЩ��y��F�p� Ã��_����	_$�0>�q��x"(�`��!���	�_�% ��]���&�$�	�W������.���щNA������?Q�e.X���(��'
�h9���H�'B\9�d�*0rl�Uh�	���p���yRE��z����Ǝ X�q����]]��7�'��	`��+� ��QM��:;��	��D�7l�� �҂�d�pv���y�2��o����TI�)'�����'�ў�`�[�X�VɀCӼIL>ؠ  HƸt�f�H�4̙�8B��%�'B1�"�#��;���q�+ā�M���ԟ����o���ճwP=*$�\.>0��a �oa}2�� *_���ɯG��I��BhL��"c҂��x�h�<1�{�-wЙJ�MքE�>�ͻg��L��8��r4H>?��`DzR�NNx��O�`8 �?��� �Y�N�Yb��&���5a��N��'�L}C�c�B0�ϩpkB���}�cI*gv �*V#��96�M`d��"�MK�� Ej���Il�X ��ryE�|�3Ѷe�`ǳ�)�1CW��̅3eK&NFp=ID'�Z�t��DM"ky�qq��##���*�k^3V^�%���
w?1��O)���uף�Oy���=}ƺ�� M:<�JdjX$ka}��Đ^��1��*�A`�)�,F��B������=A����~��S8�p�E#w��0Q������y$(T.�`�C1�K�}x>IEz�A�&M�=�	7�Ԡ��-��M�F��{6��CLF�*��)���i��Y�ed�
���2z/�@��㋕ƶ��E@^�j���2l
q;H		�!oxళ�%jӆ�C%f��?9�<6��E$�i�D�#(T8G<���O�@S�AǧQ(f�0b�MQ]�T%5�t}�j�/cv��	�m��x��X�'�d�cFN
<D����f�'N�dz�M/$$A�E CI~�OL�H��ߟk�G"N{�L��ܘW4���]�!�dN"l�d��6��%H�cu�J�Bhf%-g���
c��=�P��}���u�ʼ& �22�ͱJ��λ;�|� U �)���P��U��0��H'�� ��ѭ7�ƵpQ��!�,p�� ռ~+pp�1(A7��<Cs��,�R��
�]�3���p?�q��}
� �#�jJ{ϊ�R���&�����ɶa?:0�C�դh64�#HW��l�'.��Am�T�
�Y�B�B���%��[\���ѿQ�����I\�V��G Q\�,ԩ$�A)?y��'	*���G7}����5�~��C�N���o_�?�cq�R���P��,�'.�;4mX��3�Mu�#=�;���[�GL07��Ǒ�.x ���@)�,��Ú�>�h��p?9daI�y��b�@S'��9O�xRS�x�u#�ڪl���A��C�7άu�sK5�I�wN�t�wCE20����8d�<�'�:��ӡH�F�p̫GD��N6 �2�٬tu�*BϬZ��O�5hQ��5	����v!��֟`�JׅZY��3�^>��)x��1O!t\������S���s�N�F.�@��מ��	�� ��x�	�����#A�_�2�Юg����J(����������d�X�<@�E(��z�$�D���'������0jb�Ăw��tKM/D�^�е�3���2����[�@c���AM�yS-(�e=��?	��K� ㌝λ7@�y6���Rq��AR'|�@y�HM�<R�&?q��IB|��z�P�!���Rd�$T|���"ѬXS*<�=i�`F�i�3�NV�bk$���v}�OSZh�����Pǔ%
P��UM���6�����'+�yI#eJ25�−��H?��%�S�E�@Xc`�N0�&�C�Njӄ}�@(+������3��HÃC�?Yaf�V~�I�: � c�;y_"�� �+�jU��h�J�F���-��MP�����&FxcӘ%�PTH�Eďk	z��b*�	S�6�[�U��D�����-�O��Ý�@[w���gD$1�ʒGNF��7��57XYxB�Q2@џ8��Ϩ�y��<:�ԕ�F.ˡ:��Tx!a�/�O$m�A�|R���J��D!8�l��6�"ɪD��	*��#R�I5�@��@�]�2*��r��$-q���O���fQSQ0(1��
n�V�c��ɯ]��0���U3�2|���`_����	*��pm� .@&01/@�����"܀M djN�$�\<�%A��0��O$��$�ڸ/@��'�ǋF���$O�O�������(��$͚_���P
�BǔĲL��ҭ�AC�O��)p���O�)�a�,X��杚^ڙqS.�l�p	K�)	�K�l�9wer����'�byk#C�!<�����ڥZ9�������䓚?���F�4�gg�Z�\��~2��kO4������&���R�ԟ��'Ԋ��W`V�MV�i��A/��4�'��$L*s��-�fBX2K����P�g�¥0sbȂ/��$��Á�.A�ϸ'2<��qr����?�"��[�~5Z#o�Mo���5&�)A��S�OX�=a�ˋ�:;���q��*u�����P*�?��k�O��Ԣ|�:�|(i�?戅����d���6O6�Ez��	�)o�\�5A��.T�q�@�'���b�ի���F�W�����1�^�]+-��3�\�V 8Arw�ِH' ��3S�B��'�JI��#=vd�81��B�(��Ҫ�O�@��bQ�G�ٓ�Ԕ
���d
#��6���sj��y�&`1�?@K�F�OΫqn�4��̀�| ,�S�]!9u^��cɇ"&��GM�?:]�Ճb�ջ|)`6�ޡ;T����MO,nN������~*E����� ��
�i��Xy�NI0��(��]2Z�J�aGb�!#e�%��X�Q[�Iv��#<}�1�E�Z�<�$X5� /qO�}�ɁE��Jq�Њx�t��aTLZ �T�����^�\c��S	���P3�w�h�@N�58U���cS�X8!��'������]x����CA%b��Q[�P3;4H㵢)h�ֽ�>iAʉ5��(CeY4����$��|��@����I�j��(�r�D�rC~|G�Ϝ"E��ɦ��)S����WP&h�ȓ�.�
�I0�K:G�� ȣ�Ư|���� �DӾ�q ��|:���~r�́=�� 8��ձx�[��qy��RO�pdg�6F0qd u��`cq�D7�;D��aQ)z�:ٙ%�'�V�a��D�(��$Ӊ1z�qCe.[\ �U�1�2�w��9wԶ����azR��B����2N�E�����n���+ !:nc�|R�j���k4A�9aK�m�:?����g�$�x2I�!��TX�&)x��5iwa��O�:�8��d��\,���Ҭͥa�> ��ęp����DZ>yP���X7,`>���5O��q�J��E�`���X-t`&E����J#���))� ���d]�'�&�(���/FĚ�`�

(g �9U���
�<�t���w�1��x���H\�X@�)��#L�*h��L�D���4��f
�B�I6�8!x$
Ӣ�hɃ��2o��Ubׅ�"0,(D��OH-�B�+擶|��!�aKGn�>T�&%ёk��]��-��a%`��ҴTN.��ELT���y{0��9�*LI��9DDI��Gs����ޯ8g�L��*AĐGC�&�ax�$��U&(�x��5k`�G�s�u��$w�y�T�Nbʀ�"��Aw(<I�	�j�����,	TEpuJY�D6k�����
r	2��W��3!u4c?��m��
����eǊC� |�F)D���4�RL{�ME�z�@h�$$#D�t�p�Y�E�Z���FE�Y�F͠e�!D�h�ᬒ|���q��Omh�x���1D�(D���$��iB�?Lt���*O� t�Ԣ_Z݌�y��:YX���"O�T�/�*��Ш���KTpL"�"O0����
gb�z�Lʵk6$��"Of)C�&=����d\"O"T{�"O6 ��*��t\|��da�3o!H��"O���l�W�fE����'Rj� 0"O��c)O�(x m:�ݛ
�v���"O�pb� ײ �
y	B��js���"OХ���t�m�Q#�;kx*\;"O&�������t9�AU�F�B蒱"O�TIqd��(?��IP��?>�>�A"O��:����0Y���U��J�"O���bF)$��D"#����z�#"O���'�>2n:=(�ˀqf���"O����'L�\`�K�mf|C�"O�EctϘ0�шG�A= NI;�"O��yg '���b�`R#�6!��"O@� ��N4�h�τB��"O�݊C�ҭ0�FQ�%�� �<�K�"O�H��"� c���Yf���$e7"O��� ����Q7���`p"�"O]��ه1~���æG(9�R�ru"Ob�)�ې�jD�S�\�[�>9�"O�ʒj��/0�'�F�`�yʃ"O��M��a� �C0���	3�"O�Q��^�[(V�"A@�A��z�"O�ęv��7~�J: �� w�x
�"O�\���:�� BS&ߴ�ц"O� �ګb�>Xq��F�'��"O���!d�K>m�E������"O�1bPc�=5K��iW���b� "OUp̌-.�c�%��0�)�"O19��8}�Պ��ܩ^Q� "O�5�Ň�>@�d�1��lG��a"OƠ:�b�Y3�3�-�=e��P�a"O��4*�?H�nt�!���Bh
`�"O��D��U�m�#�4P���	�"OPH�SG^�d���G��K�<쑀"O����͠E�ҵ:�c(Cؐਲ"O�-тD�C�������.M�N]�"O0���g��?o�[c�F�b��P"O����O	�-^�ĩ7(ciB�r4"O�q뚁PZ0=RE�&L6H��"O^� ���k�Ls�o��#(h "O��j�
 �6�l ��tx���"O2�ba�l�,��땖z�|1�"O@0#��̓4$�R"+�2�n�!�"Op዆���k'����'J�2�ڥ"O:�j�읔bK�L���IJ�@8W"O�%����!$��	�o�vF&���"O��1�_�^[>D�#O�9��v"Ol��'`�L�De�N$Q����"O�9JQ�Z:�j`��K6	����e"O�dl�	-=R��*��|����"O~���<x��W���nw���'��as%�',nL�asi ;�����'�@���h#[����B?a�aPN<i�+$nY��k�h����ԪP�B���wyB��>�0��6�r*���B�yR���-���S��
z=�(;�ɚĨO2#� �IaT���꘿)0�A��I�<�S��x�������I�6�I�����eD{���i�
񓢬�7b�24��&��SEZ:�'���t�1�$հ>�x�j�-�y
� ��S�ƕ0@  �RlD�Js0S�"Ov�qbK�I�ɑ`�
eU���g"O*����0�ܡ���h/���&"O�lz�/A�.��1�!#�9 E�5"O"��C��l��)�a��;�V�"O�Ph�&%��R��x䜤�E"OT�FM�$����1��&D�<�05"O�ґ��j��3�>^L`�"OB���{�,�T���GI�5	4"O��t�^�X,����e�WN���G"O^����	SFt���Ј%?t}�"O-� ��g�����H� �8(��"Op!�AQ�-V�4��"/ti�����H������H�9\0�+�+ש�ԙJDn]��yRCA7C�H���&�7���y`���y�f׸l'��q�[4s�~\�V�Χ�ya\>X9���M��b���ƿ�y�ވb��%��#	�̩�v�3�y�EQ4�TˀɎ �d���yV"e�\��g!�% ɜ���'���y�㕚i��U��#�`�
���Ҙ���/�O�����R�D[N����'-A3�'��'�����I..�f jqFZ�\*�'w �	�c�($ƨX:��c�- �'�Ee yPIx��)R�\X
�'5�S�$�K'|qk�Q<�̝b	�'�ؔiӊ��h!)��Q�>�Q
�'��� W�O,80Hw��)(��
�'��H�s�F�(w��5*�Y1�'����Ҥѭ}�6��LU��
� 
�'`���G�� =(��E�O�RGf���'k��G� v~fuE&ڶD%�|��'=��p�l��Q	7��3Tn�y�'chD!�P!�Ì΅+�4�`�'@����h[D����c �3R��Y�
�'&��@������g��>�N�
��HO��'iך"s�|�#�^�ص�%"O|Uil6L�� ��C�j��G"O��`w�2H�ؠ��FH"2)bB"O"�1��=;�$�D��"b0��(5"OĨ�$�է`�땉��.�;�"Or|���[�$��)� ���k�"O�h�b�˼T��8H��=��!�"O�I*��6:�Q��3�^��"O0黗�!|jj�)I���	���O���D�	����v�c�y2�,�!��^�;�.���.�'~��j��'5!�$�j�����76^(�,�P!!���9t`<zvb�!)�ĥE����!�d�_��Gc��0��*� �0�!�*d�)	7�H�Ŝi���'.�!򤃽��}�bQ��:���#�'�!򄕾Ϡ|�`�Zu�t�2��\u!�\A��X��̪&���(�a�		!�$J�.g�	�½^����O���!��qf��d������C2�j�!�d��^�fUrӯ�x}�̙rj�K�!��E��`]�Ү����|�!�d=5K���Rf�_v
Di0�!��"�^m#Q`�WY���H
� 4!�$�3	@������ ��,ıf(!�7BHhi��T�PVJ�t�!򤂌Lô��&aG��
P�6�"h�!�K��P9�g�4��q�R�&h!�� |�r%�K2TPf!zGS�apF�y�"O�ݑ$�	��>EHC�/_`�Y�D"O�D+q�F�0�zwdQ�O��3"Oj��s$R�h4���C(qI�A�#"O2d��C�Z���'�'V@d"O�@1fk��B��E��ۨ`-Ԁ9@"OشBVi ��dH�ğ�V�eKw"O���I��&`��8$�"#"OV��B�
��(4��_^pJ "O��'G�!-AȰ(A"#K����"O��$g�����V2<��"O�����B+��]��iZ\1
Ћ�"O�=P�$R�I7�x�G&D�"
U��"OQ8�O�<f5����Z�~] �"O�]��lu��BTg<cKLu4"O�!a��$3�݈vŜ-=���E"O��6f�L�����W����"O�a!�>�ybw@����"O�T��Ʉ��pQH5�ӛ��9�"O(�pp�	�h{�IYu�3(�X�[��,�S��yRj�;�j��"�� �:��!���y���$��t���|=�M��͉��yb-6x��Hμp�x�tm�2�~�'�.e�B��I���6(נl
I �'�L��G� z`v��cW�T;l�S�'��qpaĞ�a��!�BP8;��'i���4�*<��5�A�;|k�'yd���( B�@�%��%�T��'�f��(9�l��4��1/60��'#b�����7h~�"��ɵ	�c�'k��#�@�)�D�ʥ+��
0��8	�'���� #�(��:�r���'�Z��C�BɃÉٴ9����'�����Y ݎi#��z)��;�'��P��%-.�Vqr��U�(u
�'_ ���c�+?��a6$��F1S
�'m|�2�F[Qq�L���C GE��Ó�hO �@�߰z���e�[v�MjR�'��IP�����]E*,(
����B�	�HA��4��_b�Uc�J	��B�I�Z�2m���$H�=���
��B�I��<�����ı �	Ex�B�	��25��OI!� ��J�uԚB��B��PD̐o�6���H8h��C�ɑw�lY+���9)0�F��%X�B��($����CL8e ��A�ް+��F{J?�Y�mոzz�!+��,Z)�0;D� (a
O��� EY8'�"s�>D�<QC����8��Ri�;����M D��3�c�@q�(r ��xY�-(P�?D��y�l��U��thAL��qXch>D�X ���>�H��KL�`I�o(D��prA�`�`��1W	@9��.�<	
�)�M;�"���tm�(ۥ5"Jx��pCȡ��A�3?���j�D��ȓ{��b��͕R�Y�4�LPb8�ȓS��s�iZ�/��"P-��>�ȓz0"-�QL�.*}��(�E��Yi8�ȓ����Sh���q�D���͇�D����k�xŒ�0�	+IR���F�V)�PH�#�[�eR�V���ȓB	D�+ �����Acć�0���e/�ueFz�VE��K
6H�
 ��F
�E�Θ'J����M5(d�-��S�? j�aQ��>����#��3<*�I�$"OҐ;T����l���	�M P)z"O��0+���\��Q''�A�R"O�h1�#N�N���͝9}{"!��"O�Q�V�����X��g�Qp�"O�Std���"�X#n�2
�y�"O�`�%O���+э
 ���s"O2\pU	�kYʵR�L�?�J�0q"O�iq���fx�(t�Q�.�*t�"O�٣���I:�P�KՆ��`"O�.<��x�l�-��IЕ[�yB�T�/L�!�)�%[,*b���yB'ri�ъ��K�A�ApQ�4�yBR�|�Hh�,_.L�ִ!ݸ�y�/�6�f��)Ε?�� a%�O��y"$)$0�1[ch^�?L�d����yk�H��.e<���e˟�yb��<1��0˱nKtŦ���]�yҎént��%o�J0�T��y�H���0���,~]b=��O6�yb柀�"��@��f ����O.�yB�۾@ ���bL
�\�����	��y��:^��F�Z��*&I��yR�^�z�p�BJ��D�X��y�nM8�p#���B�ص���y�o��^�M���K4������yB���b�d ��T-��iP���y��4�p�r4�Z+"䐩�V����y"�Oհ�5��e[r젴���y��-�b@�_�]w�����R�y��S�|�(�̃$Y�r��rɜ�y� ߬&�Q�` �0CSڡ�dß)�y'Ԕ�80S�@��3�Zi���$�yb*�C������% Z��I^�y�@�P�cȚ}�r�'���y�aV�O�xʲ�M�E����y����#�ޡ؀LZ*y��j�!��y�ֲO�`I�)�}�$���R
�y�L�kߚ��'i�5n큰ˈ��y2���,p|as�`ܕ�%��yBTr/\��(ڴVx���^��y���YN��uk�M�H\k'O�y�F�0�����a>T���� ���y��V��Ҙ{ei�L�1�2��0�y��1k:�q"��b�R|i"���y�#���d�A���i��p�A̽�yBI3z[f'�'�xysЄM#�y�M4/Y2��V�Hwt�k!
S�y������FƖ�nF���s�S�y���?H�p�B��w�� �����y2lr�lD�Ū�<�Q*R�Q/�yh� /<� kvIґ%{�Q u��yR!̫Y��� ��(��8t.ֻ�y�CN#/�lq���KY
���葔�y2 �~���kh��D�6�����,�yN�.�@��MXp�i�e���y�j�Wvi��H�A�D#bќ�ymĂ�2|�I�55(ٛҦ�y"�v�l�F�V���b��)�y2�[:� �:���<}zH���N �y�
$7
�D��f�w�ډ �eڥ�y��IX��{�D'g�]���G��y⬙Q�4I�r�J�M����1j�3�y"+;˸�R��N>L�F�d�y
� ^Q ��	L�IQC\�%40��"O4T`,��_8�����
A��,��"O��c��^13R<�J%g��T"O:�
$��q�<Y�٥G	f��"O�D�$FȌ���	�kZP�l�2�"Oh�8�#\.m�4L�Rʞ�ꄓF"Ob �F�3����I��;�t4i�"O���e���J���K)W|��|��"O����6<�H=��͘3r_xu��"Op1������KbM�WB��X"O2`�� T!$`�7�n#�3�"O����M?$��!+ I�2$>�)q4"OlT�`��~�։K��F�$.>1��*O�Y���bq��-h��'�~�"��$q@�� 8ƙ�'�� O�8��X����	�>��'$��R� ʂN6��c����T����
�':#���V��87 W�W���'���@�A��Y]�0PoJ�U����'S���.+Gxub2n�Kf�uC�'Y�,�֪�-	��)��R�l!H�'UV���	(��YF+
�\]��'��0٧�P�FΜ���Fذ �'*n���A��	5�Q!�<�J�'*֜�$�5�f�R��÷}�4�#�'�jY2���6`�`cp*�r�N��'�l���݄kmV�r�I*kE6�C�'IԐ�',<��A��J 3�&1��'�|< �g@�����胳% P��'�R��$�Mg����EF�)p�`�'��<{��<H1p�b2���,��y)�'�ԡ� ��6N"F<�4��j�'������>���t(Q �إi�']
	�f_�X5�q���`m"��'28K� ���@�wC	V��X�'�
� �H�Kg�Ɂ��D�Q̤Z�'������ X��C���: �lIH�'#px���ēE\6=�s�פ 3@�'�ڝ��a�����#g�9E��@�'�^�kG�ę^��â/��t��I��'c�Q��ݷe
D��fҽ8lLk�'�L\�
�y�H%00���H���'������_8_�a��oUzY��'/. �fFF�d�(��w����(�	�')���M�^����'V9��mB	�'�\0i�	M�'z���#I�[�L�`�'Rڴ4M�F�\�Y�MH<	,�K�'��KEL@�"E$Ĳ��H���'�,��3D��eF��aAR/v�0Q�'�~ah�:��x�aD1m|J�3
�'��k�g�)]���$L�e:�S	�'�V0�G��;3l �� F?^�$<;�'E�0���BҴ8K�曥^T�
�'%t5�!G�6]ΐ��I(.L���'�0���=�@�re�%6p�X�'u��c�H�b,��Id���'Gh�kA?�z��B��A��*�'���A k��)p��
U�����'��E`>dm65
�'�3)�� �'��`o�,���JŹZ�@�j	�'IZà$�%0O2�y���Y��ĺ�'r&	u��T�h�r���N����'�x�b�� v(,@"Z,4⪭��'6ހ4�U�0B���mO�t������ �8d"�7.��&�E%f���C"O��	'O�`=r� RZ wz��cP"O���!I=f>`�B�:Nnb���"Oĭ�#�_�^3�Ll�Y9c"O�QCmxN�䛀�Ji|�"O���C+���\
�i�b���"Ous�[8���� 
�mFTs�"O��B�>mp� JT^$�7"O���:� ��C:�["O�T�d�U�]��=y��FQ���"O�]3��C�7�\���s�PR�"OP8傎)�L��E�P����"OTE���y*��X��"OL,��PB�Er�c�T�����"O� ��P�<b	 �k�0\0#"OTpAS��6|5;��\�:�b�#3"O
�'��o�� ��_@o<ۡ"O(i#�!˧Jh.4�c�9]_h%��"OJ�� �R	'عFD�1B��S6"O
��ɕ]�E�TL�zML���"Oɘ��\�
q�іY���@��]��yRCbA�4�Re�:Xh��c���9�yJ�q�%����K���X�.O��y2 E3"�jq��JD,Hx1(�	�yB��"��@�By*�+�6�y2!�?h�\ب��P�1d|9��S,�yRe!-��M� ���V L��7����y��ʦ�ҩ2�V�����%�y�G�����"�¦>��sgkȌ�y�CܶL9��H�̕�|�|'�A��yB8T�>1$K��~m��e��y��M�+ qZ5�%b�tr�D�yRM̗mc,ipvcX���lSU�ک�y2��.]��|���S�3��=�En��y��,��GM( �[u�9�y�D��&C�PkQ(ڼg���������y��_�wA��{a�YZ��A�DS$�yba�i+�epE	(h� ���D�yr�
p^����L���6DV�yh�(��,
G��!�I�B��y�*�
�t�*B�v�D����y���f�m�b7�R1J���y�nA�#��0c�$O�)��8q$���y�-�a�r�A / �j�L���yJ@:/��}	���7 تp�@�y2�DZ`�8��Eo���FMG��y��B7;�%�e���R%�y)�?Ӕ�+P�.
�����y�
�_�dpH��-RW���3oج�y2!�.���f$�T��б����y2_�M�N4iҋ�+IL��I�'�y�,(��̹��<H�4{�J��yrb֡|������G@V%��O��y����܊�lЌ\���׀_�yr��	�v{fo��|6�""� )�yb=T�"<��oƤ�I�,ي�y���d6ЍrF��y�2E��a�9�y2#���#��3m9D!i��T7�yR��7'��qUNa:�$���ף�yR!�1CHYՏ�	�<a2��y�O�E��;�Iӝ	�&=�p�̝�yҧ|>�[�l�3 x�`*UQ�<abO����`K��ac�]����e�<���8T9�@���QC�AH��`�<� �U3�U����2'Wwf�w"Oƹ���%X�8)�fJ�85��3G"Oh��c�:7~B1Sp�ͨ&X�rv"Ob4B���}EB����ߴN0�0F"O���s�ߟd���`b۝I���"O�i��#����&�?Y���f"O��PiG��\��;1Ő��"O�b�*�2?����@�ق\ Z�"O�)Ge�!n�|�Z��\�lN-jq"O�Uh2��e��a�H�P8.�F"O6M��K�b�T��F��X&�U�"Opi"-�<�I24/�#"��5"O�I��*d���iSn�;&��C�"O�q�D.��Z*9q�����Q)�"O�1*�/ŰQ�P�RM�@LԬ��"O�}r��j�L5��"���P�"O�|�UCWM��Y8E �}qrEJ�"O���q�["XI����8 ^���"O0��5+�+�����X(|pIA`"Oe�2)�+"Ff�6&V����"O�ف��
fɌ��$��Y(��"O�li�f	2pvR ��D�(u8��!"O(x�C��p�YCV�,p��|��"O<P����9@Z�y��P����V"O���T��Ԁ)X�Pd�<y�"OȘ� �GTb$# �ɹg2�-�R"O.hѦ�<pC��r�`ɗQp�C�"O|�K#�وwg�ЀB<�8r"O�0�čB�r�fir��B�x�!!"O"�k"	�b�B� !.R�k�|�y�"O�|��L_"	�b);��9)B�@"OH�Q�̫$�T��U��(~0��F"O�A3���3f�P�k�4��"O�����JCW��h5�F&t����"Ot��E�V6v߀�a�EۚK��� �"O��cڬJU�����b�����"OLe���܏>G��77��	#���y҇מ�v�ba$�*Kp��b����yN؃N\u�fd�& �eCCN�=�y��nTLP�v�$@]�SN��y���/b��0���#�`$C�I��y£�����@D�\ DO�D�K��y�V�64�a2���pȤ��a�G��y2-���7�c��{���2�yRC�.�mJӭ[
V�Z�pԩA��y��'XΈ��r���V �c'��yB�ŌE�uꄩ8�p��"׏�y����}itQإ���i(�擘�yrJ�"s�F��W��w8��dԟ�yҬ�:]�ū�H
�sz�}�L���y�@�1-�rk��[���&�y"Ý "]l�1�^S&�����
�y��D.BS��r��^ZEB�ځ$ï�y"%�)i����YI��2a���y�Kǩ9���0���D�r��Q��yBɃ!	����X.��e ��2�y��/#]p!�F�>"?��r	]�yb���4�,�JT
�%&L4sw��%�y��8��#O�IS&��6N���yR,F�JD襠��ȬFS܉#�L��y2�N� �&xɁ��G;�B��B�y��.fex��d'���{�%Ż�y��ȩZ�ܸ���	˨H��E5�y�i�e���yw#ĴS������y
� ��NZ�Qq�$�q�ʬ��<�"O�̀E�#�|�"V�+|��"O��
���	��!%I,���B"Op��b|E@��iv:��K��<�c@7%%�h��ω�ր����R�<����^%�D���[���⅃F�<q���?=���
`�4-���d�i�<y�* Y*N8���S60@1b��h�<��_�_
�h�<5��P%e�c�<�殃Z��I�� ��`s��]�<���eG�o�D�0�[�<�Sn�;,T��!�S[d�z��V�<��B�$k}�ixS`E�H��%D�y�<yA(/��xѡ�@�[`"Ồi^y�<A�%80� ���h�"!l�0��u�<��Zx��8�%F���|J��[�<y��M�0ΈEd�9UZ8�i��<���S_�t��5=�D��Ěy�<a��R)0��80n�:Dp큢J�@�<�s�ť. ���,�zC��a��~�<a�":~�p��@��)���s�<1�*�!,tͻ4 �0 $ViP�NSm�<!��Z���
�/W�\m���C�<qF-˵wl p�䛨;�(1����<ᣂ�([Ul��� Y%���*��T�<Ѥ�V��s�l��؝��cJF�<I$@+RԒa��R9z��bKP[�<A����6��h@$�ڽ.t�<���Js�<i@� 7�4�kļRI�� D{�<�w�[4��t�ͬ�LQ���@x�<9F�D�U��xP�@.LdP��dq�<1�' & F���)F�*�X0l�o�<Y!k�"T����r�+@��0�i�g�<�� ��}l�U�C�Ěcy@퐐 b�<��M���UN�-َp ��Z�<	�dW���ӣK�$��r�[B�<�3�P5���0�c��B�$�u�<1��s(<pg#�Bb�R�n�<!��Α3�J���d4jD��s�<��l��@���PQ��H�RC�s�<)���r8������&R��9s'�w�<!���,�C!CB�<� 3�l�<�a昉kN���(ɵ<�zd;S��k�<���20m�x��gF(t*�@�<9b�%*�f=��OS�%�lz&��}�<)d�ȋ2%Z���ަ��h��d|�<���	6�|���� d �I�1��t�<)s����PEm��0;.��j_X�<��+�l�p��?���ì�R�<QR�Z�(�i�FhK�U��(��ZP�<�A�Ƚ�|��d-ؒCd��#�K�<1�^#,�Z1T�3똅���I�<)�@�61pt�#LV4��\���AZ�<��MU�JT��6nVQO����E�<�� ���y�G�@:\)b���y�<��=T	��H&�N�$q�i����l�<�6_�A|��m��𽀦/�k�<�@��p�d�DanX,	��k�A�<���'h8�8@G=Z. ��G�Az�<y�-�'�,�JPT�{�� ��`_�<A���erT���^��Y0��^�<y���/��ɑ"�� �lQxR�P�<1�P�?q(H`@݅����פ�N�<1�` �J��g�
��2���@�_�<� �E�л&�%#��
jjt=xC"O��yv E;02�4sD�͹3e� h�"O�y�O�YX��R �.���S4"OD�R��, ��@�b��v�*���y�T��i)����Dq����ybN��~�,��T��J��x#WcS��yJ�6Ǭu[1�A���b��֦�y"b�����Ӫ>52%�Ǥ���yB ��]LFA8�l��.�,�pwb¸�y�eѵ$~�h�1�F�(�X��C1�y�(r�JESTH���pF�C��y�$�k�tmc�_"rs<s���#�Py�@�M��l  M�2 ���p��{�<�p�<Z��A��C.R�25�$�PQ�<�EN�7H��u����s9H5��gOs�<)aI�+M�^*6-
#u�&U� �l�<	��ת0y͛��W5
/0Y��a�<���V��e�3πq��`�<���!	��s����hs��ڡ�Y�<�F�E�4�hş,R}L�Ѧ/a�<�C
�8G\�����O-�ı	�]�<����6dL`�񂐿Tr
Q��I�Y�<i���eP1ò�ѹv�X�6��Y�<yB��O�y��� ���k&�W�<�ь[4Q������>����D��U�<��ħ,'t���=rc^�S�'XS�<�K�ne��ŷg�~\�b�N�<I�h>�1Kdl��d����Rd�<��`��h�D���T"�D�A�`�<����2x\*mH���f�%C`$�_�<!�ė�z1
�At+;���ց�W�<Q��X��D�B��U�P%�R�<y��7	����*X�z�$�΃w�<0a�J�d � R%W�p��^J�<�		([��If��<Y��_�<��*۲��� Lb`��8!#Z�<1�瓿
dm�@���lx$bFX�<a���_D>�93�#q�T �RL�<���9~A�4q���;�pd���<9�瓚M�v
�O �=؞l��ʍx�<a��T�%���cp-�7�)R'ɏv�<�����	�L�s�g�dE.�)r��H�<y�OM�P���SRB��&�İ�W��O�<�sۜr8��Hb��I$��f"L�<I�,��P����"�Z�i6�u���_K�<AO,$ze���C;���aUo�<Q$�&^ڨ��-8#������j�<A�'W�t��G�J2Q�:���Ne�<��C50P�,��d$(�V�ʦIAl�<�U���9{(l�&I��*�ln�<)w��"h�L�9����`O4���F�f�<鷦�� 0L�jˮ��͎f�<iC%�)6x*m���_t��bd��g�<v�H%i�]��?װ\R3�x�<�@"�������\&u��ls���x�<)ah��(��%�_'B��ӅBs�<��A�v����m��= �v�<y�
�\�H@�V��	Ku` xh�x�<Y�mˢb�A�fN�"�����~�<��f��a��C�H�£}�<�w��<6�.�2�b�k�L���)u�<��f�w�Lh��f��s+���`@f�<�dᑍ$�Ƅ�QfE ���0��d�<����#��X( �N��T�X�#�^�<� &S���Ae�����].)�%��"Oxy2�M9����j���<�"Ov�iV@>`�����	A��$8`"O&t�S��[����f�K�va"Or����/f@��jI7_� @�"O��j�O�0oB� !��&".���"O:�r)�n ���D)L
_e���"O6��eKN���31�1�`�v"O0Ek�畫K�Jy9@�1'�5H�"O��@!��I�E+��[��E"O֡��'3.�	3��׭~��a"O���J�!>KnY;e��4ʔ�t"O�@b�_�+Kr�ʖ�>g
��f"OF���Fӱc�8 ՄY1P!��#�"O���cb꼳$D?U8���"O���	�;�9��A�26U�,R�"OB�A��"_|�Dዊh?l���"O*a����m��P5~, ��"Obȑ+! �^��Do�15'���"Oڹ�w̆0�-C'�[�)潱F"O�h�j��c"6��"�پxqp��"O4��tL	�~Έ`�wN�62x���"O|��S.ƹ
�\u����z��T"O�Cp@�Arf��<OyB���"Oj��P�U�ckF!4 U#2�@EK"O\1�,��L�=����:y�&��A"O|��ӯďZD��`B�y�����"O�A�o˗S����l����X�"O@T{�� Z蘔�n��/^�a�"O 쪰H+%st����Ғa�	�d"O�E8���&/-�������R0�"Ol�a���LA�$SX��>��b"On�9�d�?Z�|#b�a����"O��H$�عe���t��S�Btp"O�ػ"Mݏxez5���kUق�"O8���N��Q��副w7P���"O����?y�3��B'_���"Of���ڴ-Z2M�CS�6�x��"O^d��J��9C��Ȟ]��8�"O�`��%v
|���9�Hr"O�\	�'���2)ٰտT����D"O,��iV�{~	����v�ݹ�"Ox�V�����"9LW����"O��X�~x$���@ޔG���"O�P#Bd��*�XH���}����"O�4J��"w�:��2�ª��t�f"O���E�"Fæ��oY�'���"O&U��g8
O|��!�X��9�"OZݠ�BQ+(5���B<s��)�"OX@�AL^{n�b1�W�U  a�"O���5*R�q3�9x�c�-�C"O:P�3$Þ9%��K$݇\��+�"O�T+&,�Zg@����·R��"O�8���-:jD�'סG����"Ox��N�:<�@���Ѹ��"O��(g�tf"��v�D!p���%"O��w�O:.lb�� <n}t"O�IÖ ��:7�G�f7��+�"O�m����;���Taٰ ��h��"O�=iS�Xk�z�fm��C�����"O!��I�B���ڲ��=%��s�"O`
' @*[�������cD\���"O ĳ5*�#\�$|�ϓ�� ,�4"O>}q�`�UN����`��m��x�s"O� ���%��;iT������ا"O�E��-�u��P�l�v���Q�"O(�	�C\^�Z`��P�-��ݓa"O&�Q"��|R�)��(W~dP�"OFU@ �,e��D�7��eDs"O�pq�D��R��Z<���5Ζ�y��۹+6���2N�/U�P�C��yRñS���4CZ�"o��KT�C�y�/5d�n��V�т�3W䟌�y��	#�^P���|�㑑�y�͈pud�Q�A�UDQ�bY��y2�Ȱc[���b��.��偢*���yB�Ռy򈒣��!���bE&�yr�
*t$��v��/�0��;�y2�7D�,(�c�"*��%S���7�y�#�AX����1l�1��Mޤ�y2'��`Q�ѧѹd!�x�J�y�cD�*�B=j�� �bm���D̈�yBiK 
��;d���\z����'�y�/��$�3QK��=��ɰ!����yre��ѐ�T�5�Bi	��W8�y���GX�Ѱs#�:|zdbCm��y��_=����we׈"�*(��d��yr(�� �-b�M#JЩudE��yr�Q�@V�۷F�K�bd؄�B-�yBɟ%meF�В��%= x��6a�?�y��ޕuA3�/
�� �q��y��� m���S>ch�<�p��$�y�Y���|�6�ϴaCu�A	<�y��ӊq$Fc��R]������yb`��!S&@i�@�%�+�-
��y�K�?�� iw�V���i�r���y�
�Lr�l���C�h"�ۚ�y�C�|�$�qREW�G����ؾ�yb��j#����mߌs	
���U��y"�K(���H����h����M�yb��5`{tiٔ�:m��`!��yrCY ^�)��T�b׶YR��	�y"&�9dl�RWB.�f%��yr$&+�0%BfO ~<���en +�y��7�怐��Y)��D:����'�x�Jd���Ab�,2��� nD*T
�'~�Q�	�!K��0.��[��E��'7�%;#X�[�<�S�.�-N��$0�'����M�c��=2�98�L��'�
Ո��z	�y�ɤEЬ��	�'�xH��$S�0 �� G@�8&��8�'�����F?5H��3��,�b���'l�K4c�7$�r�@�
1����'���0�!�,B~4!Z�!ݸ�J�@�'�>\s��7y�5���5���#�'�d�	B�X�Ĩ��kC�}�^8�'fA�
cA�]#�:A9���'%��I/�>��m�/�<��
�'��:S�"mH�׎�)y����	�'���jg+Pe8��H�pi�1�
�'զ|�E	�fM1��A�?�}�	�'t|Ѡ#@!5�@yBꎄ;>"��
�'�H ��$U Hd(k�dͅ&iZS
�'���HaF�!�J!oT��UX�'&�<�v�J����3v���(��'�Hik'�ʀS�f(Z����A	ج�
�'4��c��`%�P���<GD��'�
���^ ����$ :��� p�(�.*3�yVH�)�x��%"O�LS,��_D��kq�]�R��!"O���C ŀP��y���:�<�3"OԵ��Z� 
1C�QSh"�!"O�]��h�;d���!�N%Sc��b%"O�S��B#v�� �N�t_LęC"O��kĠA"� 	���-hIds�"Oұ+L 6�3pH��/P �Y�"O�`R5fא�&��&*�;M�@2"OL�Z�g�b��"��Q�)K�8�"O.q��\+.-�s"Ĝ2���"O���
�-|��f���-�J$"O IqRf߄t��Ѫ�퍑;X0*u"O�QbR�(���*8f$�uB�"O�h���R 2Ӗ�;���#���"Ob݂�%�W��aƤ��K
d�3e"Ot��P�S2U5>�!��8^eх"O��ٷ�@1|������r �"Oi(��"�t���ǔ�]欥�!"O�� A�&��M�A�j:��b"O09��	 E<�㵥R�z�[P"O2l�4�R�L�ZxYu�	-ܴ�cr"O�#@��o6ƨ�`g��a�*��"O����4�1æZ�RɌ�"O�􈆭�3��iCf�9຀e"O�	P"�C;Xy�E�&#Ɗ���x"O�I���ѯ
�v���,T�llN�"OX�;�
��[_J���H�U3B ��"O�p0�B�X��!ѪE�e����"O����FMH��[ �b�B��B"O�U2�Iߒkrv���+]�h�x��""O2Y�B
!W6��,G#u�Bm��"O�M����M�쭛�
�F��=	@"O"	��"-O����j�(R�� "OV}��lM���B0*�7b>8�&"O�Q��V�U�.�9�gW���"O�h2�H�<e*�G���T��"O��z�	���hG �\t�U"O�ir���hڤ�Qg&ܷ`nE�"OX@z�'�6*{�m0�ʗI:e�"O !7�[p��*V��}X��R"O�e!F#�<�\�Ra�)��h�"O48��4�L=
������*w"OU�&��4,s�Y���e~|,"Ort��aN�')\�[5m�&m��s"O&�*eΊ�DO�9*�,��8a�{�"O�aY�I��ȸ̂�e�&���2�"OP�����+n��	�S�� �2u��"O�t���*Z��x�,��9���h�"O��Z���%JV�K��=�0ʰ"O$x���P5,uTXp��S�ĈTS�"O�	�er�����is$�H�"O��p���wԚ�i�&���x�A"O�8
����X��Ƹmٌ�Qr"O@TPe�Ǫ(t.<�!�P�+���J@"O��+E�I$=3d遰��+��1r�"O�Y��P�\jW���|Jg"O< �k�"8���A�.\W�V��e"O��2DIy d)� (�>df����"O�xq@N6ok�)��R:Hd$I�"O�*'	�0 $��Y.�ð"Orx��M�����E��u"O�\)�o�H7�=����-x��p�1"OZK�Ή+p�`���h�"lR�"O� �T��f��if�i"$��1$���Ɂ"O� 6ݵ'G�	���%v�`�"Ohu87� �f��z G>Dc\l�!"O���U�F�)C��� ` �7H�|��"O�i��fW5�z��p(C�0H@�a�"O6��w)@	Ux��a2��3C���1"O`ܓ)M�D"��Iل�J�"OdIs6E� ׺����8�PL�q"O6�I1�O>t{�d�@��9��p��"O���&!�23��,@�Q�4b!�"O<}����"[��j�Ȓ��! b"O���&�Ձt�[&䗝7d��"OleZ���V�|�ELY9PY"OL���:c���1��p��0�"OD4��Ö2N����>$8q[�"O����-@�{�@����Fy��{�"Oi��|�	� �:ir��B�"O �zE��$7JT9p�8yax��"Od�����aCTX���{Dv���"O���G�H{�{&O�V"h�f"Ox�ط�ֵW�X$`DK�Xi�"O4 j ����A���ɂ w"�;�"O��"'���@0;��Y(>hʘ3�"O�8T�C�0�B倆	<����"O0i��	�>���I�d��"O�f,�1��u,Θ6CT��"O,�BF�˾h�>u���
|�C"ORd�k�lf@�
Ӫۿ�U�"Oؽ���Q�|= A,�!(��I"O�V�W�ix�)J�$�8;�m��"O��Ѝ�!pa
� �cE4-�d}a�"O�M�S�V�&�@r�A��+�$Q��"O�\A윺r�:�Y4���&X`ܛR"O����/��w'��Ѧ��#M��A1"O`�0JN�O.�a�`��=I�@W"O���DɌ�� s`��PAP85"O��s��;��M��`[	"9d��"O�{�����6Ղ�n�k�%8%"O$��`č	1�t*�n���(*"O��Cτ�Z��ƭ�(i��"O�q�!N�B����U�G�$�6"O��q�M�$���+��څs�vT҇"O��R��>���aC��lB�P�c"O.��R1n�F�q�*��t;m�r"Oze2�G�Di	p�h'"��a"O�T҆ƎB�]IT�>X�"O��3�I���I�b�X3u�2U�0"O>E�v���&�)B@j�����K�"O��@�&�<D���KҲ�"-h�"O:�*RF�	8P�X"gk�RmxMT"OvQ#����h��`*�)],�"�"O�5�W7F�l0���K-���"O5� ��h�,Ȑ���N`!"O�B��H�h����¼"�
�bb"O�((��ɉ6j�y�Bwޱ �"O -���>E����D��pV�zR"Oڄ��iO5B���Q"���C_�!ȇ"O��Y����l!�ڙg�b@�"O�����?}��P�N!o����"O��q,S�
y����)�`�`�"OB]��L�+g������A">�d}9"O��z��Ն �VQ��˅��,C"O����B�o����K�%D�X��P"Ob�ja�A�	��I�H$�"O� �8熛NЮ}�@�.I��3"O��j��ח?8Nػc�(1�:��1"O�\�CL@+-���S�ȽK�h9�`"O(��F�Ye����$�x�F�C6"O��h��J3%�=��o�	)u�!	!"O��d��#D6����U͎ɺU"O0�A�F�
��e
dMۤl�Ia�"OVH)��ו��0����2Y��:�"O<1�-�t/n��_�p�H��q"O�T#en�=L�2���8А\�W"O���qc�?�`Dؖ�nǔ���"O���c�þ|~T���	SI*��R"O<4�ת#]^�#q u.���7"OBY3�F�(X��Q�bj�$4���P�"O҅r��8{���(�6N�.�X�"O��A��jY�gĵz~��"OIi��S#@t8u��"'`]S�"O���@h�3Fu@�	�@DR�h�"ODQ��o�8�|���K+R,$�C�"OJ!d�K�@"��Q>&�{s"O�P*���r�@��еA ���"Ob}�f(����a <)0�Ic"O@!�n!c�p��b�]�<��\��"O���b�3�r��WG[9!�F���"Oڌ�+�Fs�ѻ��R-,�"���"O:|�nڌ.��B��6��Y�A"O�1C�E"��8�ġ�7w�r�˃"O���B&S���)�%.�� Q"O�x�Qß�l�$uyD��
�nq!�"OJ���&o��%�F]�o�����"O��+��F�n�	�R�X��"O��`2$K8�2����J,H���(�"O�0�����h�|��.μ����"O����/Hi�LӸ
�2i
Q"O�L�k�3��
tB�($��+R"O��%�cqQR�,���2�"O�5`��ØU���@� _#>A�q"O�1c�\7�){0�,|±q&"O�b��"ќI�v)���t9�"Oȼ(�jW�?},�d)��:���"O*����z6�Ad�\+?T#�"O�A#�؞D 1�ƒ3J���"O@��E]�m�x�j�B�̉�"O�dpcB�7�x���!k� ��P"O���/�k�d�1C�45�
0Z�"ODei��$M|�����
^�"O,yP�cнi*L!D덅jҸ0�"OZ����;/�r�GJ+wa�%("O�(�`�Z�5�|\�o�+xgT `"O���R��~��CΜm�A�"O�E(��G�	��h����CZ�)�@"O~��4�@P��1�hٽ}�h�8"O���w�@�8k ��b؂Y�b"O�]�F+[�z�0@��Ɛ%#���r"O|��Jďb�p!��_�(��"Oh 
 EA^��š�AJ`u�"O~U��h��Z����"|>n�HP"O�H������8*���Q�j�jD"On�9���<LȔ뀂`�=9�'��q��·?xl��M�^u�Y	�'�-ѓ!���0��ݼR#V%��'1�%U�F9�4mW�}�8IP�'��wE�*��BU�³x��t��'D��r�K<�<Y!�,w|P�#��� l�3�ءsDL�E�G�X�R"O�}ᲈ�?ke8ɺ�j�%Jƌ���"Ov`��=�v�8VI�z���r"O�}2�!����(r�G�'���"Or��%Jա6��-h���P�Y�"OB4p�
B� `��,Nl���4"OzɈ�+�WBd�d"�8b� R�"O�����>p1>�������dH�"O�P:�ɛ��<R3.A�LC&%p"O�y`.P(}�
t�"�W�'n��"OT���ۜ3�JԀ7M��!�U��"O`�I�c�!C��H.�*Ph��"O�8�"S)4�8剑�˓^Qd��"OH����hѠ�kwm�0H.2<��"Oܑ�&GԵC����Q*5&�)��"O
�Bvđ3}��)�'K=��)"�"O���e�t� �sF'*���PE"Om�I<Z&�\�K��$v��(3"O�ܛA�ь24�5b��	x"���"O�c�G<5�:�K�+�Aa��"O\�P�T�VU�t���+6R|��"O��E�7��5K�+��U�p�"Ok�g�x��1q�	9uf���"O���dT	"/�Ir��$}�``"OPBa���|�'$�+�����"Ox|!��OL��� &]�+�lm�P"O�p{���#=��C��Y��@Ř"OzDy�ǃ#(@J�������8H�"O�X��M�/h�3�ſO���ZE"O`�¶�ԮWRV�B��Q1����"O�ܰt��>:�X Aɐ@P2�3"O��f�
m��P_�
9�W"Oԛ�+���+���Nt %�B"O2%ѠS�lw����MX�n,�u"O�jC�\,d�}I%�:r�T��"O����]r^���m�u^�8y�"O9:1�ֺ+ ��.Rn4:�"On�2���9�&U�D͊sGP��"O(�c@�O$}�����N6��8r"On��$'�X��(�Un�GT�;�"ODm�VăA��R�YHmV�ȱ"O�T�D�� vXq&v]`u��"O<):��&,�� ,	����"Ov=��1
�s�ΰ8.�-�""O��SB(.X�5��Ȭ�ijC"O6Ac�\7@m*)��^wd�ٕ"O�DZ�B&�����?Q$T-8�"O:���	S���#�!6� {F"O2��ЧP`0��B�2���"O��)�A×>�qRԪ�ZD�qF"OL���
u	V�̃?���QS"O�Lr�XMN�!��ɘ.gT���"O�$��%!8q)q�F�PM��ѣ"O�t�CDăy@l���+�LS"Oڬ�c(�0P����[�ʍ�g"O�p
���<�� c*|�2!�"O�x��(��ol�4P�65N<��$"O����#�-	�� �"II�y�B�X7"O޽Y�D��z�$ki+ �d���"O�IB�H�}Db�8�n˗^����4"O���MȾ���`�L�+�LI�"O8�aU`-"�lI����}��)�P"ODĂ$�Pӌ<��a_O�d��"O��H0��
��\2a�:"Oj���"O� ���B>K �kp.O�-ce21"O�h٥`D.$�� Ad��N��w"O���cGui�X0tk��d�H�G"O^��,�R�Zj�Cד ��i�"O���On7 h�C��-3�z4"O�p��/p*�`W,�7T��"O`���D�>�sQޅ���K�"O����e�>��8뵪�/�~��"O�IiB/
��)��I�'r�D�Ѵ"O��g{^�R���2$ov(��"Oz�R�˷ ��ˡ��kcd;�"O(��$�~b�z�3��1"Oz��D�:���3&�G���A�"O�Y�P�}#��I�.A11���"O��/�~��*e����y "Ov�!�^�+�9�G�̩z�x��"O�0z�B�(6k��� )^(k���"O$З�E�5�XJ�(�}d����"O��	��F�;�v���^h`�E"O��[�`���nq�a�ǭ�ȕ�d"O�[��J'��d��	�q���`"O�%cA�ȧ]���h��]�j]{�"O�ydJ@@w��)pU#P��Y*�"O�E,��S���e"T��� "O�m�*I7S��O�|"\�X"O�I�"�b�����
�%�XU1"O^麷c1{I�=�eϳk.\!�"O�(���#����p�����"O�(��a��_���W���P}X�K�"O��f���K.��`ݗ,�8��&"O�����0i^��R�ֺ ƞ���"Ot�	s/�$al�42�E�Y
�i@�"O� q%�&�ʅ�dN�'"����"O�q� Ȋjj��8J�"ObbF��,X� ��=3(��"ODzj�G:���IDĴr�"O:9��Mq��h���-m>~���"O���G��m���&r,ȕ2"OF�s�c�a�)"���
�
Ƶ�yBD�8/r~m�����=�$e�<�y�e֊uEr�zDg��(@�ء�'�1�y�"� �:�!�h_�*L<����yB&�;H
��"�ᄑy��a���Τ�y�M]� �<�aFFntfL�5EP��y�bҕ@�:�� J�s�(��*���y��D���x�o֍i�(�#�?�y"� 	�p(��8񞨳���y�ݓR���ʙ2�, �-�-�y� <,��p��#4�yХ/>�y"�s/L@��A��ha�����Q��y��Y32�����8��r3��-�y�� NU����;-s��*���/�yB$ϟ|4B噃��w�݀�ă�y�d_��X0�jԟr������?�y��T6a�Ͳ�	dU����/�	�y���:���HԶl�к�����y"���Q��2	��Ί8zr���y�Y00X�x
���:c���i�M��yB.B�xg�YI��j�443��
�yR*�`�`�v�c� u���y"�H*Y���o�0S�0A�E��yrE-c~ꌩ�M�R�,H�q���y�I���	��\�F�RL�a���yRn�U�ȘQ�L�C�
Y���y
� `x���	��R��aŖ�,�ۄ"OL��0JC7C�(�:��մK���*V"O(9��ݵNP�#��	�Y䲙�%"O`�HI��J"���;*�څ"O��S�+��m�<�Â]���x�"O�<���&_�谓� �\s6��"O�x�u��\0:�	� c���!"O�x��<O�9B�ռC����"OFQ����+��MS�}�4T�"O~�Q�!��EA�� R��)_����"O�DD�9Y��t:�,N bM��b�"O��А����+��0ir�x�"O�M���m�m�U���0-��]�l�t�'�vI BBH�hl0��&@ 
�;��~��O��i���	��4j�)q"O���bj��p��Ɵe�FAy���nx�?����_�T�P���@�NӖM�2L=D�� �$�{^ ܒ�����,�#�B?9�{��9O�1Y�P&�B�/\=Y�%��"O����؛}����GmɉwQ��c"O����G��H�q�	����x	��'҉'��I�?�pu��lէ/�ЁYf�Pv��B�	7��@�Pk���Uo	��,B�IQl� Y ��Ұ�R6'Eh�B��%�"�;"��)�b�Q�A�r�C�I�ev�P��B�N��4$@�8��D{*��"<���z�` ��U<W.��Cc�<�@�Ԩl����ӋF�I2�m_}�d$����dq�^����J5S~�2bG�Vo 4�uOu�B��7�v��w�K�R�X�`�>����?9����� S!E�Ju�"�fź�T��(O��=�O~R��1@мvv8�$�?�2��	�'���:dJ
�*X�!O�=�:��4@� �<E�ܴ2h���+_�W�}0s�
�+K���S�d�8�����1E��
F��=��~b�/�(?YAiI������La<(kb*Cy�<��E�#���i҅N��``�C{�<����h銉�@�?��lc��v�<ٳ
^����#�2"$�@'������)���CB��%� �h�BW��=��D8���I�?��R��Ս6~`-�f�ֺ*�rC�{��U3"�yg^���rf��>�K�p��"���I����ԨS%@evp#��!��C�	vz��AA \�LP�fD���IR�$"}��i��Hf��AJ�%�p/�-�!��]�z��fJ�δ2	E�`ڥ�g���Ox�?�'��z�C�jƂ��ɑv0��M>э����	s]��f�F�=���jԮ��_�!���,u}������{PX��-�>!��\�2;F��dn9}x\�Ps�E-�!�d-�( k@Ğ"�*����.L�!�D�p�z�kX8}�)�ۅ]��}"��8i���3n�"�Rt@&3�XJ3�2D��s�">��P��j�}ƶų�;D���w��uV�*�`�cg��p�:D�`yp�D;�V���䒅O�����8D�`���A{(�"��7d��	�Q�"D��R� TQ��xbti�����b"3D�� �������Q̄�fX5`6D��F�^����!	,H�>1���9D�����h����?HRAg=D���$�ŤGRLU� �3&ꌪ��(D� 9B䘾964��SjR;.��h�a%D��Itg��4�	��0�� %�L�)� D�'�+I�|�Ò&�D8peS�"Ob�K�� {ӠY�g9!F<��"O��I@�5[�e�Ɛ�1�;1�xB�'|�X�$�fc$,1G��n��ۓ��'0PC�`(7������&�xq�'�܄zGT$o�qQC��l\H<����$�<)!�ӻ��IB�N�m�����J�.Etȅ�[���Pr�]�y�I{�l/
L9�>
דz;tዡ����⧖�-�K$D��K�G	�b��.�9WR�Y�L�t�Q��Gb]�l/�I�7�C;O���H�=Ɍ{BG.4�0�a��?G:Yx�,A��yr��
z��`�Gܫ60�x(s��-�O��=�Oh�h�E��^����*����'�p�����
��y�
��)�<���'�	��h��<���I$�=&����'�\���̌����(=�+�'Xp-sF�Wid��7�V=%�v�q��D$�'$�#0�Q�z2��o³"� P �'�֩���Z������I�DU���ēvځ��l�.'d)��%�GT��ȓ.���E�D_
$��S8��F|R�_t�O���2TB�F�����0 �dX��'�<m��C�_�6��T ��!g��H�'Rx)P���@I%K��M�D��~��ؓh��3���=���� �՗�y�Dύ� sc�U 1?���c����Ol�~rR [�����x�b��v�Z�<�NW$:���ebi2Ȱ��UY�<��K:����`�zn��B�	Q��d��5�v�lВQY|�'�~��0�"`���L��dC%��?���)�S�O`~ч��5��ّBA���c�"O���¯K�9�h����l�4@Y�'t�6�Z~R�O�#=)���,*�XR�C 03R���痧t�&
O$�:��'v��p�ᛗqW���bEBu?	�2s�4a1C�h�APrؚB��l��5b�daR�@*m�p{�D�<l<6%��.��$����zNlxV�D9[v����d�"��%�P��@��;a�H1��Ŷl�GB�1\�	���Y�ڔ�ȓj009TIF �H�f͚�6g���ȓxvL�3Dś�gd�}�cǉUj\�'�ў"|��&C��I(dǟ?H�������q�<��˓^�@���4v+΀�t�Qp���=��T�a�z�k�.T7Nd�Y�B�ɣk��}���^�>�nQp#�^K&�!s�OqZsn~;�X�h�͂�R�8��t�|��'-�Oq��y�"�I�[�E�5̊8'lT��"Of��D�r��iF��ql�i+��e��;��@�N؝�eI��`k�DA%�/D�`0� Y*"�h ��� z<�(�+�>���p>��9�Ĕ���Ƭ>0�%�mL{���'u���}REN�1��bk�#.{�8��Ė}�<�& �?	�A�Uc�9T\�ae��p�'Ҹ�9S]��>�=��� �X���\�b[N���	���Q�n:��d�u��n�r|���M3%i݆E\b�z�$׮s�XrV�<�$���xt�!P*ۤM��P� Ah�'���D�����j\���ƣ<�V�`T�	�~B�'f�O�>mCu�:2}D ���I�Ty�f�`�*�� PBQ��|2r���cH�ӑ/D����b
�~��0�O�a0ū���y���4&P(�ĝ|B̝s؞��vE�Y�����tI�P��_;�y"��S<�M� ��c��Gd����jZ	2p� $�t�����w� ���ƞ�ch����ӗn��*?�M<Q��I(o_�a���"Wvܫ��ݼ�4�S��)���)�뎐q���V��|����O�>�۴�O�>@!W-?ޙ�D�ǳz���C�/D��ir��!�"ex'�P1~���B�-��S���=�cD�$r3f��"̬D)�� r��x[#�i���aG#O@���]�>ͻ
�'���X΃� ��,���܈l��ә'�������̐��"L&��86�T�y��
�~�2��E��1L�!C��/�y2�ݨG]�ɚSNə,i��B��-�y"�Z�z&,哢���'�0�'���y���peDa��<,�QB��!�y��wF�Y[�a�?w��Rd�C��y�+F�UO~��#�	s�z4I ��y���]+>\�#���D�	�y��`?\,�d��C{48�S�
��yB�I�}VJ<RL4�d�5&�4�yb�P�����^ (�^%�
��yO���H!΢,��"�$�yr#P��:�
�*��0@F�@KT��y�c�C?l!��d�e��yrM��9���S���,Ad,ҍ�y"j������3T6�����y��F�7��!�e#G�L]<��B�X�y��U�T��i�2���.�Qr���=�y��уo�"�SC�P�{u�eq�)Z��y�JG�zK��ic�U:||b�&��<�y�B�-v`P�$-G��.ٸ��7�y"�F�Hm �ُR�4�7Ç�y�M�m�*9
�g {_�)Hw�N�<�bF�����
!]F�)k�OK[�<�W�>�H�I��e��ʧ@V�<�d�4u"HHp�lQ =D	����w�<!d�,��i�ѩǽ�%h���C��9�>ɀ�E�0�a�X��fB�I?t���prd�1O��#�c r�*B�	-K��e�Ӵv⾹��産��C�ɴ�m17��=l���/SJƪC�I(nA����'zF�`�@ŇݒC�I�.���r��ߧ+���X�z�pC�� {�6�G
)�(�����'ܜB�ɰ��)����9�lТ�@�_RxB�	-L\![#k@�ܜ�%e�2B䉙kɚq`�a�.SF�+��;]�BC�	��gh�.O�`c�I��2HtC䉦k�$��e�1L����+@~1C�	�"U�P$�:erA�=��B�I�@6�5�F�B�Q����,>��r���#V�pRD�ц}�����2�i�,��De�TJ ��3!�Ĕ��R,��(��vGو��t!�D�Z����Աv2N� ãN�]l!�$�[��䱶��[����ͳxR!��P0q���`��Q
��
M!�䞑J�H!J@�7�6MAB�
2�!�d��h����;`��APrC� -�!�D=%����ɱ�Ȭwș�!�ԄP��H�$iI�(�1�� �+�!��|ƪa �H�Ŗ�G�vd!�C�T��Y�E�h�|+�L�#
6!�d)q��\0�,X�*�P�kD���!�	8���p�Fݻ��Y��`3!�Q+h�n`� -̈�r���?!�� &�r�K(>��	
V�N�8�Ό#'"O)�F��K$�11��C@�"O@T*�G�lofİīW�2��X�"O�����\��� _�P��"Ot�!�+[<��H��� ]0e�"O�`��Rsv�]�B��-Cn�yg"O�ԛ��Y�	X��;V� �"O��!�IG�`��B���E�lrR��c�p,v�|B��8ed�,`��	R��ɥR�J�RDo'D�4kS�v.����P ^�(&�e�ȵ1�nE���h�!sp�b��O�$ǺD��
�p_�E�뉱/,�:�e��m�5�N���[l\|Q#���,t��C��RP�|S�  >2�%�Ӆ	�����ɢ��Q肸�eB�Ona��lޠ!�����#�2�;
�'���(�CX=*|�%�B ����ʡo��0����'�<ac�'�gy"�)b���0$|V��-T��yb�-
J
	�"���p[`m��vD͚ $Q#)-��3�M7lO؁б/U���iBcv,�1�'�Z�� Mb�I'�i��p1^8/��p��O���	�'zňT�)k�2��}˾Mi�{"�G�aղ��(ǥ@�>���F�{H����	����0D��9u�£l�z$$f�6ۀ�Z��P�$ �v	�2��D͆�(��I�J����a�(�v� n�)Z&B䉙F�i�U�ӗ`J�MF�=B�:6�2O��i�B̉1��=�v�	;�hd�'�M�V�^�j#H���z�ŭ7 ��̓D���6�&;+*Ճ�/�(Q����h��(�	ې:�ܘ{R�A�4>����l-�7�[O�X��&aFh�b5�?a#�ݬg:l�R��	T3prܪÁ�)�l���k�H� �Rm6�g}"*��(Y����P"����=^��8I!)�)z�{��>�%PDp��*��=�Z0#7�ÁQ�yZ"��\�����	�k��y�'$�l�d)�e�"=�P�f(�}E̜�V����'�����@~��
�|]2��9.�-��J�p=�N˩@����F�
�M��_ M]�%s��ߔ2�|a�D�~ܓs��q���?�$����Q}���a㋏Aӎ)X����!j�����͆�"}�c̗�EPR��a��D���ʆ�;�r5�=��)�gy��&���"��oDIX�,Ľ$���b�@�-Hʓ�|�'i�7F�(�:`�)D�
B�a���rd���
�L^h� ��q�����oGVI�}R�DE���y׬̝�qO��KF�9��C[`��s��y�Ε��ݛc㞵�뉱qc�,)W�Y�c�em�/��zc+ҘSh��	%e�POҠ��͓I̞�X���2Iw��As(�,\��z�� Q�qOn5���@){`�Q��,.ҧj��ă�i� ;y0��Խؽ�g۷}�ɥOڭI�KOt�g�	-k`����+���g��{�fQ��Ɵm�޹�O8�F��'ij�h���V``�ȣe�n�����)s�F�9u��Hx�����Os�̺�&�>6�X@8��O��QGO�Zi�b���c�W�+�̤J!Q�Y�� �P����AmŵwSZ�G� D����M���5�G���cFlq��*��H�͔�r������@�M0G�l�+gG��!k�"O�M#4* <(�de��Ɨ� � ��0^�A��'C](7�#�3��X�f<���
Zj��q��}!�Dֺ8�b8�n��|�s�����������8�8܁	�@3��S�\&f@��R�y����剦&�\�Іդx��I�*�ޕ���I�9�,�爈b��B�I��`�	2��K�>|+q"Chf�O�u�6�1��hC��I��L�<�#��U�8��13�[*<!�dW�%̝�$��a�1҆ʉ+!|�A�|����$��U#�u�P#��^su��B�9<���7��=Ys�[�tGR�w$�#h,�x��X�4U���$��\� )��ؑS���Y��2�!�I-os�����(|�B5�e�1y�!��\t)�0QuF����z^~�!��r��*��/�)�YC��n���͝�@�*�0
�'YЙ�u
��gtZأ �&U�Lik�OF4��b^��4��� 8�@r'�$B0 CS�H*�b�` �'�|���֌�4�PbgG�>G�ك1�7Z�n�C��+Z	!�$��
�F�0d"��x;MR�#$/�O�(Si˽ P>x[QBI�O�`5�s
��$�j�)1f�5���'�"0�R�IjhDkab�䖼���²+����&��~���}����<p0 �KL1h���wAN:!��_I���ꊢIn<<�S��h����(���$��caz��W)q��W�M*�|�bC��p=aCg�>"S������\ �����V
6}�#����`H�E8D�$���]�8s�u��%���zЁwb<��V:��C�n�*�ݹ��S* ���� �V%k����$�zC䉤:Ȳa�#��_d�A��R>2'�`�C��$9� %��e�����<ـ�� 3����cZ�;�^JU+S_�<�'I�U`�e9FD/0(b~����Fݔg2�a�"#\O>0b`>'���$n�|`�1�'�19�g�6�tD�иi��9	��,JP��1�O<����'52�D�-zujMcQ@A��( I<��� �/*9xP"�&�ħ�M�� ����ʔ9]L�#8���Q��R'!�ЇS��At�ʢ5(�xIH�$u(�\t}R�G3I@8�H��d�	�O�x"q2��@�7+׷#7D��π�
��}ˆ�'9�L�gkư>p � �,X��h`VHʿ�h�#g1F<ݒ�_�(�aOJ�6%?�	-D)\���\kF��t�ϴ`��"?A�ʄt��DrD '2~�˧
x����5�Ykq'��!7L��I�/0Ƞ���q
���ɶpgZ\�цG_fU��|���7?z������  �Ӵ$;�)�BC �'�H4sb^���T�5u�� �3�3-D�|�''�k�QS@�.�s1#וyw����,��2
Ѳ3xA�ק�#h��E�H䀝w#
,I�->�I��U�a#��!�~vB�h d̟)�� 穔)l���2
>&?���b�Ns�X���F�<1B��<�a�J[��'�
 �4eט{�̨�&j�G�Z�>9���Yi�-[s��%� 1�u>y��m�83� 5𱣘�	J�@e�'�R�3O�1�9����U���I�&�q�B��37T�чSu�8�I�#��a�L�b����e�Вy���*5��}Ҏ֦EH�1$d?�l�!����k�J��gJ	BG��3�6�On��e��V*��ƃ�0���౯�[�<��@�­o9-#шJ��d��5��
S&��棑3����?���c�����H�"k$Dh6�'���$��\HX�)ĨE�;��R�MYB�U�ěF�@<��+�.����0YDN�yHD�>�����"-
�,��E��>1� aF ���O��겈X�;���۱��l
�I�O�(��̏kQ��/�$
�~Lۇ/���ɞKL��v��|"��2=�Jp�f�,Q1`�"���4Yj��r��Iд�^�O���!��_�C��R���x>)hp��
G��uiDN�h��l���
���bT�C�>{0�r��E:�ȉ�k�|�Ǐ'Z�p��'����`:?{8����`�-D�
%�3 HsP���	
�Ȑ�o�<}e<�!.O5P�T}AC#Q,|���fP��LC�T02ͦO���}�aL	="5N�gZ�J������m��Q�P=�L\b������6"a��
��+`c���#'��}3�>��爿Mr�>�O�U����)[.�����3Vv��ґx��M�f�2��=�|�˅ `�e���/R�Dʱ��иH R�ޖ�p?I�h��i�F��AȾt���ؔ&��%�a�&()O铝�锧@��M<�dꊰ	>dY0OB�t�F` d�r�<�mD�wV>�;��V�<�~��N����n��}�Ȃѧ�O���3 ��*k!�͑A�����b2\O�h[D�P(k�8��Do ڸ�@�ˍ�s�4H!�2R�(Y�'�����Ӏ[sE�a��S�P!+�{��H(h�����%�5��F���J�#:|�'�A���X��ɧ�y˕?l���!���B�ո�'�8�Dɣ��42�H1�'ˢ�E�,O�8��� f.l�bh^���C"OB�s��$�j���v��q*)3@|`0"����}A�'M&��ç,%�f,���؈35F��דNd�P�b͏Wwn��&�cB8�[d�{r*]�w!ܙa�B䉾�4b�	,-+̘��'��o������CQ�~D�pp��:Nr>M�g�:>��г��
_���"D����Z�/�*Y rg�\IAA�Mj֢}�"M� UR�I
;jQ>˓a��(HS@��f��CЫ�7Ȱ �ȓ��x[o ���kc"�3 Y0aono���T�qiH ��	#~�%gŃ2����#){T����3F������M� l�!1gD�32��I�N�G�蕉2"O��3&ӭZ��QIp�R�;sl �"O4Lj�*�>�JӃ{lX(�"O:��6��~��)K4�$AWB{"O�1᫞�|�
�b���E���G"O��Sp�X�3V��fIN|J��P"O]9S�ٱ?ؐ��C>=*�"O� � �9'&���Ug! zD�'}���i�C ���¹7�PI	�'��	�M��@X �!�ā�Bb���y����L�+�cYr\r�_�HO8��R�\�, ���p��5ӣD�!��wҌ��M�1�:��"���"�!��2*Nq�i1���C�d�
j�!�P���RQi�� Uf���㎄[�!���{`"� {}�,�)X�
g!�O{�X5H��U�hX�| "�.n!��E�Q�� �� @�a�СcM!�$ĹQ���z��P�y �=���@�R9!��NF�@�Ɠ�j:���@ګj!�$F/|�r,9����4��3��4S!��ދq2،���a��yy���!�H�I1�YX��d�դ��!�$�2��ea�*�$i�$!q�+, !��	�n[��	H�,���#�Aе0�!��T!z"�Tˀ����kҢI0�!�ė���ypd�Z	V��T���M'.�!�d�#�5� 
�%��o�H�!�[/��Y��O�;�@�QOE;�!�d�	R��h��+��� 3��5t�!��ůg���b�R�3�J��#�!Z!���Jŀ��I�9D︨"�F�3 !�D��e1���eN�r����P%�z!�3��%2V�F�0C��[e�$l�!�+La�Az�`U)G �تD@ϰTU!�D��DUU�t��^�`�%�rA!�d��GV�y��n��y�<Z@���X!�d� ��3�A%>H0E��ÚL�!�ʝEmT`�J�N=b� �c�b�!򄙛 ���YT�ަn�,<0/�b�!򄒖�hL��HK?`�k%��!�C-6p�|�U.@4 2�}����2Mi!��^�z��0�A�G> �0���U�a!��GT!^�FW'C�����טq�!�ā(-{�8�%�P%#����e߿|6!�x����ϔ>G���1b��o7!��Л0]��ѡ]� ��I���[I�!�D�\��0��#��]�2`�f��!{!�dM&R���jC~��scQ=7h!���?�,��2U�Y;����t@!�$Y�.e�� Bϟ�nm1�ŗS!�Z�%�V�r'%,&�g�U�M!�_�����A��O7<Q�P�ڴ>�!��A�vB�Л �F+5���aύ�%�!�$�(S�$�#�\7T����E � :!��&*,��R3�_���4 ��� !�ܤsg$p����b����t��E�!��-l�脨M�0Y����!��!��Z:{�xx��!�<B�hA�<`�!�$C�W�I������x� �!��R�_�=��kM�Ks����C	�2q!���"���zq$�R�B�2]�!��>�>�0�$ԫ�<��d%͙tf!� {uZ� s�رj�@8p�W'i@!�� ��I&'O�t�)����D�2�"O4��C#_-�
y��"�6^�H��"O��S�}��QಁZ�e�	�P"O����F�>l \a䦑�
^��"O�i��-��x�@$�^�x��'���UO�c���V�M����
�'����'ɂ_/��%���r�hiR
�'8�iH�����i��͕�bH�#�'�jt��E�@�~t:D��f��L1�'�h|��lE31A�x���f�P%��'��؂���(�Ȭ�nۛZ����'l;�KEOt�D4�@�T���s����P��L>y���Or�k�탨 Є̘�BS?t�p�K3"O��I7)[
]x� ��B;�*A["�i�"uc��"?^��I�?�Dhb�U>x�D`�!�7_���$^�z�I�-�G��6MЦ7N�,�B��/�x0y�!K)p[!��
nd��q �B�e�ʙZ�c2qOH����3\�P��,�'�\��ᖈ&�Hs-ճ;L�a��/�j����$x$���#�$(e��+��XvhP�gR��8��<��KݎE������/K�H0r�e�N�<QV �6$i�@.�`�t�Ѭ�e
�1��
��<"&�'�\@��N�2��M�S�6$�0R	�q��<!s���1�Z b�4X�8uI�C��+s@] �ʕb�f4�ȓ8�T��a
Ⱦ�>�5J�K\$c���ÓLW�<Պi�O�ՙ�\�:��\�WMY4�l	��'D@�Z����4�����?�ڤi%�D-����j�<a�5�gyB
�2!���,��$���cd��y¡�`.�a
ec��]��U��M#LŵN����@,6|O��˗hN�5Ȯɓ��o8=)��'�Ε�F�S����. Ò�i����q�G��!��^?&riY$�&B����po�Z�!�$�2�Dc@�\(m�����ڭs��O�T�Un�d<""~����	JP��R0��H�� 0o�`�<����M`G�_j!�p�#�%>��ī�w��K~�>��B�%�ǳf���,A� qԩ��Gm��bK�<��1�ր }m��p��_�)�J��[��'#$L�w��QVH0�CQ5-�x�ד�� t̉(�"��ش��i@�kǆJb�e�T^�$��ȓ�\!ӆU-@�l� �:�l�=��̟��8F��7�H�����&-h����mze#�"O�4�� �֠�#��E%)�ZH�IK���i��xy��g����J���`"Ǽ���M�.X��J����p?���'z��-�DX�5$`@QG���$l�+فiM�9rc��@�$��!#*?q0O�T<�3�Geb�O�`�����F9*���CHA��e���i�Q��]��X�/�$��)�24�ь����e��"�k ��C�V�S�B ���E)Q'i�B��3F"}�^7[/�Lc�E5f�&�3�5f�e�M�DY����V E C��y[@�1�^�PBU��2q՘O�� ��9OQׄoGڥ�e+	�3..,���sG0ܙ�D��>i��w��iK���l8H���#ҟL`W��Eʎ�>�֍�%L���&�<q��=�ƕ�t� (� i�S�<��SVZ���rH@><8��J�e�	 ~6@���T�I��?�`chdQΤy���� ;� 'D��󡆑�!&-�	�	��1jF:m��Oz=���O�g≵6���p'��k/��@��\k�C�I�j)�5�Q�ܽqDpX`�D�9w���bY)��3g�'P~	�΅)vi܄���<D&��
�R�ޘY���z�HʓD�ȍ"���
j�\�t� 5~�0�ȓm`(xp�G/KS�')yJ�$�42Ə��3��С��is^�@���"�v�jW�^ k�C�I!S���B�G�E�x-��,�4L�P0e?�4N��?�'��J���g��h�U�@a[�@�
�'j�Zt�H�O��ѥ��
�z����D5�@��	
F�V��WÂ����сOS��B�)� j��%�Pdt����"O����$Ush�u�R��< ���'NVm �G�S�OOʈae�J+��]��cЊ'��];7"O>m��OD�%��D�P!��r��2�W�(96�E����I=t��]�`���8��F����d��b�bܰ�a̼v�����T$mZNk�H�&x��'D����&y�m��c�i����C%�I�r���`A�N��p�!��E�k�Ҡ�R�Kn��(�&~!���0�jA�(��2W �Zc@D�<�0S�"��e S�O����Y����n{2��(���y��� D��
��&5��W�G�o+��#Q�ߩq�$H#.�w�d���8LO���H����$(�DN:%P@�r�'�9�S�UK�,��Т�؀*q凞
w��qҩ��+�=�ȓ4����Eԃ}�f9(��>V�j]�=�$��)o�6��� �',�"|Z5G��e�v�Q�f%T��b���e�<��˘.�%�"�JBh��P�9���ِ"ٳ,`R�ɻ�Q>�H��M���@&b�n�A0��qb����P'���F�?M��DǓ�~|Ne UىT`�ՓT�INv>��D�]P9[S�ϙO�B��K���zb�S��J�b��(|�V���D��1�w��҄��eZ �yb�]R�FX�� �w�����E���'g�xyщ��vP�'��H��B�>Z��n_j�$@'�2�4��ӄ�0~H!�/0$��Cn�ZRa�u��6W��c"�k≫.h� �U&�!Vz1����9ڢ YSR�C��E(�)E�d�TC��::A��;�� M�����J��H#褋s$�=`���t��<����O��7�+y�t}��g9!�A��"O2	�S��~˜<*W'_�!"q)G�'����H�w�m8��'%P%���93Gn5ۑ#�45z�(ߓ<d3S!�T/^1�%m^�[м�7�	�"�b U��y�R*M�p�`�0�>U����&�$��T-'}"M� H3q2e��1�O?�n+_�t�1��;b���'�23'!�]�6-qw��l+\��f�-u�$�uj��s��t�R�`��]�>9Y',����Ovq�t��
����p`D<�6�B��'~6(a��N����}�r`r�
��4��@��_-&�h���.�&E��p�o�`���r�ɖ�?�>ɢO@�R̂ꓣp0K4#k�9���1�T~�ʓG�x戆�U_��B]d4��QI�5{.��2��9)��i��H�� "�戼U����H5c�R��ƞ Dc��c�).?97N�F�������R�6�*s����;:�R���.W�p@qb/N=6m���ȓN;R�3��^����B�9A�����<'.�ɫ��@X#�S�	I�N9X�c�B�[�쥟�	��5�����c��-�����p=ip'صu����x��q��ےZ�z���J
�1�nMѴ	��4��'a���b�w�g����Y)�=C��a��H9,/l�8������0�哏C�Nqؓ�ӈE��Kg�0h���:5(� q�'�L����P!<P�р.��-iM��/T�)�K� ��ݟ
���������O*@�î�w���"3�Y�C�Dѕ"Oʌ %��&k��IeLB,:�i��`ʄ��4?���S��A�FC��'|P�>��b#�~p�UZe�ֱD�-$I=|Ona\"��D��{=�U�jR:e�rj�G��x]�Ǔ>9������>�O�y��Ý|��D�����x��O�,�$�ۜ6�yJp�»~����/E0M����@�;�O���U �$��Ѧ�J��ಂ�_F@Q��Q�$�|�U�64��O�� ��Sl�	�A�K'w/�lY "O��r %�D��,�!�16�
�i�TH��QG:N(@%�'+zb�F�Jq�A֥�R��u�x�m��E�+q��q���K>��	7I�SSb�*A�пi��C�	"3�4�H�͐�(��H��%�vi��H��˹1� ���ǃn�>=��
�[���+� �%t��P��:D��unE�X�N�
 ˟	V(@�P�9W�N���h�-���	 (�Q>˓�&�B�M�.&ڲ�J@'��n"���E�4��2$I�f�"T���+H\pS�S:(O�T;��C�
� ����4�͛C�C������9W!����E9&����NT�3j��V��� �< �gL��Aqq�Z
�y�͙�vrm2��̺M6;Î!��'���!��hĘ��#�a�O`̠�7/
�E��&.�zC
��� \��%��z�<r4��_�ɱa�\����"F��d��(���9S�L��bO:_#Hݳ��~oLB��X�k��_(C�Z%j��C'�P6�vH��+5�F������V@���bLՂk�Z,9u)_�q��{��E�R��m
���Ŧ�����T9��a��Q>٪�d#D�`�QlJ�iU�5����"Ñd-D��٣�����u�bI�VV�4�..D����E�~��]�H>)����4�:D����@
q�=�q�x󜔺�i5D��Äo�����o�/$�X�(1D��ؗ&��{��@d�N�- ����;T�� �,N�
dn�ч��
L{*"O��q���'�h%AC��*8 a�"O6e G	 Q���6G�K�"O��K�B�}h��t�] "Ș�&"O��@E�3a̼X��_�o�}�"O���`R�K�����?�QY�"Ov|[CE�����G�F��Y��"O�����̴]�xX�^.r��q"OV\���/�$���*φ'�8� "Ox� ��炜��H��X�v\;U"O!pC�ٱ:v�b�AI�_`�M"D"O��s!�,/�$a� �>k[�d�C"O��6K( ؚ���[�Q_�̋�"O�&m[��ĸ2�)P?2��"O�ѳs�m�y���
�C"O8Mȁ�U	2u*<�VZ�*�C"ON�krdPy�pu�Bb[�	�` �""Oh�%��-� �`��*�����"O�P��Z��Z����^%��"O�q`���bO|2шG�`����"OB��<h0�р��-����"O��-W�'�Ԥ84�V�>�T�S"O�I�cV3y�x��/˽� "O�U�O�4P�	��''���u"O���/lQ�{�l�:i�="B"O�s�T�KF�#����^�l=y!"O�}��e�.�p�Ɵ��(�"O8�`g��F�պ�l�|}�}hW"O��8�(�P��@ʖ�R��Ik�"OD��I޸�C�-$�Dm��"O�Qx��]�ql�I3)-���W"O>�kPC�2,�"@ȕ7)!��iG"Oz(�ӪnRE�@�\?`�Ա[�"O�8� �.@���u���GVR"O*��D�W��kW��,H^�l�E"OZ����݁���/��ON����"O�h��]���� �4N"ODI��c��}C���� -@#��K�"O����*�#E���nC)2����"O�x��/IR��4B�L]��\ �&"O��"�չbpv(�l]���qô"O:Y����6>V��h5;)��)�#"O:=P!��d���3ß/=��|��"O
v.��w�m��#U&4�T"O���.Ǩ\O���3�Q�*f"��#"O�RWAT[8\W	k�8B"/D��2Fmޘ����⮓���!J�`�/d���],�&1��M??i ^:�?i��~~��@�4�Ԓal��4�*p0�]�y��'�TC�y��i���e��Q��Y4�M�h��d�.X��"~��ъ\�u*��]�]2<�*v�O+Z\�Dx���'*��qQ�A�ΐ-@%��2����Ic>� t��-S�0�CMOh ��-?9���?m�O�X5���h�E��!o%���8Ox�#��ሟ� ����i< ;Jъ��P�ѫ��������i�&+Thpt%%�:��%=�4��Ɇ�?YÑ_*ZY���O����O\�;%ď�)��!��Z4C����P�|j��2k���SN ����e�ܥ3|l��6DE`y~�EP���aʚ�<���I<E��� z����Jim����yүJ�����.����A�ʏ#P����?�6<h�N��T��0J<��)Ρ`��	�L(2f�\8	���J �\:��p҅���O�(ȁeo�6PB�Q3 �;(������#�HO�� T��dIĄC�\nڬJ1�(kGVc����O��~*g��.h�sD0��b�P�ɠ����<qH?�{���;�	.�"�@����z��;�Q�t9�g��'�"}z��;Z4L��"	:� 0Z0i����{�O��O�t'�Eh�P>m�5,A�ѣa)X�.�,�d"D��e��G
��p&�(_&�{��>D�<�Ш�
U�zC��yɦ�*'C>�V
�>�$�[ I�y��S�%p��AY\�'��ӧ<1S!����i�/��Ai��&.�j�(\{1ZY�~Q؄���K#8���<����R~���=#\��e*�/Q4�� ��V1:�T�#�<����"Z�j��*G%b���
7�$Axa	א���ē�,S��Hp�Q�dI!cp�Y��Q*$�kG�
'5T91�(�i��Є�PB$���)Y`��x�a[�kn��\�p��7L KIb89�L�)m \B�	�8�X��ϡ-�X��,C�	4T��=Sq�.ris�n�C䉮C����0$B!@ )��k��B�	�D|YN��#� MS�@�k�B�I�\��̃�kY((��lj�Y! �(C䉏"����7��!���Q$k��B�� nw�Q�d/#C X �a��-�B䉉U����MŪi���s ��1|B�	8(JCgD�.T"�AY� �!fB��V'>QRT`�0ܘ��8e��B�ɑu%��&KP�//v��a 
�P��B�	<`vhb���l�0�+pP�B䉫DC��{@oA�!�	jv���B�N��8�i�1YT�Y��	/g��B�Ɏyˈ��぀�/z�h�P��'%̆C�ɼY.>y@�e�/�
0t�CT��B�I�}�T��;>����ߓ��B�	"4�t�d��9n�&`2šP"C��
k��9���L��@�H�Mpg�B�	
P��9����'�@�bL���NC�I�?���&άt:0a$N�d�C�I8���j�%G�9X��[4���!1 C�CL�9��B<kDQ��8b�C���`qJ䫅&d/��ҥ�@��B�	%��W��<C�q��(Y�B�$Y��� ?�)��hG��B�ɾV�u�$"�9aŐ��G�"L��B�ɑe�֙i�"-�Xq �'�[��B�I�p ��r���'~<�1u�U�%�B�	'.Nyz �P5tI�DÓ�O�B�I4�~�¤ESs�$�ؔ�_�R��B䉦 �Xe ��ǚ0,��S�ޕb��B䉍kJp����ܻ O�Ӏ�%)(hB�I�� ��@�(o�
Y�v'GTv6B�I$ >Q��תOA,�A��% mB�I]�� I��L�?�PQ*���R(B�I�T��f�G,�w� T�PB�ɗT�>P��B�4Qrbg+)�<B��&�J��0|��ґ�8��B�	�x�T���ƭd�\��`��B�I%b�X��d���$�B�2��w	�B�)� p�0��x��9#ÀL4s�)A�"O1f�N�PW����6��`��"Ot1Q�af���E!ҁb ��5"O�0:�W�&$x����;$d�B�"O��5��  �� �a�@}���u"O���1�Pg!�ň�Ó�L�8�b"O �1v��Q� !�$��
�Li3e"O�<��GV�`���N�9p�r��c"Oh�x�A�<E@ R6'�t�jAI�"OΕ8�a
^��(b��ݳ�"O�ܱ�AԑZӐ��a�
]kP"O�a{Q��`k�0���ь~.�0"O��qA�Ē�������u�\���"O\�&�P�s�̩ូ>��U!�"O�p��Q2�MK��@(?sf4�P"O��d�37uX]+4��7]<<h'"O�F�C6,Ҽ$YV�K� F ��"OR����Y�p��.��a��P�"O����O�/��JL� ļ��"O�'�:>��0�K7���Sr"O:��׈q���xwZU�^�qs"O�3���&YT���I�!co>�3�"O�@E��	F:�b� V�D�� "O*�qu)�y��<��A�F"O��W�̞g�d�jd&A,e��Z"OrI㡏ҧn9�6���F���c"O���e߻7���%�5���X�"OHi(f�4C}$ 1��I��؃V"OX}b@G?zK�P�C���[p"O���ۆga@` e�K�`x��W"O�I�1j_/r�
5����kH�=�"O>5AB	�F��jԧšI:����"O��	E��0t��װa�#�"O2�j�O�$'�6@�5lZ�]�d�W"O��)s�5@n9���ƍ1g"���"OH����J�L�����ncP��A"O�8��!��Z �g�jj�"O��*�//\� Cg��~�b"O:$`�OE
H�U��?8��#"O�qc���f�	2v�����S"O���E׎�X�͞0��(�"O����ڞI�� �rJU����"O�i�gŗ:Kv�{Vi�`�&�P�"OiSBbԞO6T��'K Sy�#"On(`@�N�>\ ���<��3T"O({%�>_��[�F��q�>�KA"Od�YPbS0Ay��(a�	g���"O�]�SÕ���8�%�͗Z�Ha�T"O:�mɏV���͘��B�*�"O@���\,IHq1�&8��Qc"O�����ō2���S�CآC��h�"O
Q��L�pϴ`�eC<!���u"O0�3��,sJ�&"YCܔ��s"O�=��.܅)t�狕N�t�9Q"O��k3_��ؕ��_���{5"O��"�*y
��S$zf����"O�dˡ%��!K0���ܷs^.�q�"Oxd�]��jDSeCޤhR`�S"O�1S%�	b�@]XBiG�d�"OX��n�I|1� �%�E"Oj�a*�'|;Z!�b�% ���("OR�Ifd�O��#��C�~���"Or��3Ƅ-)��@����,�`�"O  Q�`�?$�9�u��Ka����"O� @�3c�= ��Y��K�&{V:43�"O�	s������U�0j�����"O�y����;Q|I�i�����)�"O��n�)&]�c"�D�I���"O�*�,�A�D�S
�c��uq""OL���#�.To��{E��+'�%"�"O|���8L��욌����"On$�thY�U�|��
K6��
�"Od�Y�M,�EP0���`��=1g"O��QaF�h	b]녫M$m���Z"Oٸ�M���*����Ƌk��x%"O*��Ѹ�H�����$8��-$!��&@���1�ЦP�����0hH!�[Հ�p��$vb���T(H0!�D�3�bl)b�)� ���a�RB�IH��$�������)���PB䉕q��b �����A�C�	�}@����L|�9��1vC��.}��lБBܗm�J�J���dFC�	��4]j'��*/�@�s�ˎ�B C�ɽ��\"t�8Q$+��Y�g?C��0�ʰ
ץT�-A�-=��B�+ct|��gӰ]� ����ЮY��B��\�
lw�Un$��MP�mHFB�IF8>p�bf�Q0h�A��VjC�I��Υ�T�N %���#��͏0�ZC�ɟ�����g�3�-kvč5e�nB�I4P ��)�79�j|j��Y�B�!��-�p�76W8���
�$�,B�ɳA���V(9�d�'�D�
}jC��$h��{eE��i��+,�ZC��<;��`�tOׅ<��{��/;�C�ɘ����R�0��JINa�C�	8vL3��GO�;N�B�I�(�(02·	�-[�K4�C�	�g���(�.	�~��� +�C�I*�P�9R�ː ���²cX Q�B䉣`�V��1�ȧ�L�S%ԊC�B�	X}j@�J
�`�0\q���Z��C�	�\�rq��@@�h�HP��.��C�I�o�Y!Sm,_�N٪��N�n%ZB䉊[I���oI�M���BL�.�>B�I�\� �s�ΘI���CE�$�(B�	
�`�z�Ĉ
���j�G#O��C�Il� X�B,drp���B䉉b�ȹ��ޜ%"h���5dy�B�I�X��j'�_xI�4c��&PjB��t*@1�O�)��/pB�I�}�\����']��V�<Y�B�I*k��ȷΏ�1�����˛/�6C䉎d�d�D�:z$�cDK�+��C�	�i\� `��]�@ r�"E�[��B䉝9(��A��D6>��ѫ�g-�B�ɃaM&a;��ڃ[ĐJDM�([��B���^<ЅY��� [��,9nC䉕x�J�*�@/>o4�ҡ �Gp�B�!�pA�̉� WE��A�sFB䉯��\S'�R'�6u�D;f#�B䉣Xe|���;�, ��!fMvC�.I7`��3=4첨h��"tC�ɐ6z��a�AL�(A��5�7
0>C䉣v������H�'$�:b'C�	~=~@�TG��eX�C��M 	�C�I�ݚLr�'(���VhC�)� hik��N��p�c�˘s4�!�"O4����ø+�z�a�� 5sx(�"O���!�-��) BED�s_��`#"Oʌ҄ Ą/�x��0䖴<��P"O��%�Z$���*����"O.h��k��r�*9J���Y�Vr�"O��qG�9\4���ܒ>���)"OqS5F��a����@��	���y�"OhM쓂rp���+Z+�<LZ�"O(�xT��:5B� )����~i�D"O�����T3?vQj�T�R�D�9q"O L�ū	^1�-�� �_꩘�"O� �%'�Z9B=i�8/�Ε`�"O����,]� =a�l��
�J��"OZ(I�hI���!A�Lbd��"OB0�tIG�a�᠚	K@��"O<<���Y�i=j�pӎ�00���f"O�xK@H�Ad�����[<$�^!K�"OV(��ho��Y6�V(3���r�"Oxi���C|�Y�hհ-!ZyY�"O������h� &,˒E��)�"O�����U��1Z�D
�H��!�"OX�tE�*;O:h��ȉ��c�"O�H92   ��   M    �  ~   ,  K8  �C  6O  �Z  Ud  �o  �{  ��  �  l�  ��  ��  >�  ~�  ��  �  H�  ��  ��  �  W�  ��  ��  l�  `�  '�  a�  � � m b =( �/ �5 7< �@  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!��	y̓0�ƙ"�/�o:�="�I�1���G|"�S�r:�HT��"��cS�pC�ɩ#��c�ٶfv��j/*�t��hO>Qz�C=H�䈊�I�(���@9D�<x����������G1����3�I��hO�O�tͪ�B�1�6���<Xf�D��'����焘C|%[dP�D-h���'�e�4'K/@
�Dce�Qjzġ
ד��'�,����KZ����.�Kx�(O����T�okzѫo�����aE��=hayI"��}��(���(f���ɒ-�g�&��5}��'�a{b�A�&��d�i�7;b�D�Wu�9J�-�'�u'mm�rQ�L)b�.�Ո��	͊%�a"O����.�g���J�Tl���C�>�K>���H�xС��>,�n �$�?t�|�O�ѱ�B��,����g<���Ɇ��X�O<�*Od�O��O
��)�.5���A���܀m&�y��	*�TFi�9�u��ˣ���y4�'%|5H�ȃ:#J�q���Y�B�<]��'&�1�D�̄(��ń�<ZF�:`�+$� ���X%E�Lk `�3+�Xa��=��'fq�*"eBQ%�p��h�6KB\��&"O��%+�m'ĵ�ph��EH)r���w��8��/��a�f�Ɇ_��3 j9D�䱲 �4f�\���	�6U ��<����a�>){Ej��c`���`�(����)}��M<>J����(�^���G��y'Ǜ+94|���܋��-��i��(O��=�O��l@6g	)*�V-r�L�2B\��'�(�����6�T�Gf��<��8�'tB)R���>�Hx�D�d�zh���� ��HQ&��(�%O��Ax�"O��Dh�:�q�.Vy�Q���x��'U�;�Zg.�`�!� V:���'�@�"d�ʨ=f4���!�~-��'��-¥�ΠT6t؉͊���`�'D�1Z��ȣNʂ%s�N�#���S�'��� H�L<t�����
Z���q�'�6pK''NA\���+�%�,�[��x���$8�����C禠3q��<�y�S��}���Ւ?��tk��V��yi�|�����֒!s$��4KB��hO����V����ʷe_FU�E).?�!��&0��2E��6�.d㢧����4��7�D���ŊI"R �� �0ȄȓU�4���#y��9��,z�b��=S�OV�?�񭆲v�5�����z�e�1-]b��X�?i�n�c��M��cI��4�(���[�<1�)��Rz%
�c�* �$�7�CZ̓�hO1��l�,D�;������
U��H��'�I<5�*M �\�f��4����"}r�.?E�T)��[�i9��9*j��H�QV!��CG���a$gȄqW��@�F1pO!�d�G9�ܪ'��6%�U��j��b���uӦ�)��*P��JC�R� ��k�"O������/�*a����P�ġ��"OL��6#Fz,�C�w��Y��"O�dx��ˬo�R����vÒy���5�S�'+�>t2�
�B��E�m�.I�EGxR�)*��E8��a��D��Ms�'�q��p=9B�W3*��@C`Pl��A�v�<��狫j�l�8�OG/d���QdNX�<I��J�?�z����wN�B$�X�<%ă�;z�R�yz��qV��P�<y�����u��� L����ƕI�<i�%�:1%��B�� �d�s���A�<1a�lS�"MC�U�aK����<i�!-���*a��e��X3�I^g����>9���5	�x�&nO�sS:���Ób�<�& Ȕi��Tе��&hgNA)d�u�IO���D��<;�(Z�i"�Lt�ÐP�n�aQ�+D�t�&�ox(D���ߋ<�T�SpOL�(O��~��
����C��@~�S����JRC�	&-̜%�V"�+A1j\��$�<$0�D=�S�O΢�	S�E�v�V|���VL�t�P 7O��'{�S�'�MP'�(1גUc�+
�Gı)���q5��&�O�x0F�d,�ڗL�K�zj傀P���OW���W�������bȮ�AŠ��W����ĥ��'BF4��Nq��AҌ�^��q�{��)�i�1-h,#�!	�J�Qa*\�I����?+��dB�B%[@88֋I9��T��i�~������Q%n� ����0T�R���-�"ۈO:��c	��Z ���4���r���k�<�7�$b���B���dx���k�<y�d��%̻�'��g��|s���gx���''�hID�DKz캔�^%HȘ�L<Ɉ���:y�Ε��I�C�Y�yl���'N:�;G��6pZ-�7b�Y�txb�'BF)�V��&k��"�i�G�ܭ�~��)ڧs��1Cl�49R1�2g�0�ȓ���0" ��I o�K}}�Or����]]$`��"�6x�I���57%!���}�^PebR���0�F�I�?v!򄂔bY�PS�EC�fR@b��T!���9��y d�+AN伲AV�#�	i��� X�iҝQ�4��0���%���*P�$)�S�I� l�1��.L#}�b��VHS�3��{b�D[�D���hT�;�x�����)��Ɂ�Q�"|ڵ �!Z0����d�9hs��hO�LV��
X�#ۆ\��ؒ|��I��x"�'��h���.�(��eJ�-�tM`���.�M����'�~¥�C�aqZ,¨IA�^6�y���Sv���MJ
Y���8����y�^�Z��́Q���V��E�`��6�y�ː�>�j�#F*]p:�xE�]��d0}��>%>˓pOZ�`a.P�;GؒQLQ�@����	T̓\�:�YdDP�ZA$D+a=�q�ȓ=�n�4f�2*�Yi jY�̑��NΤݡ*��=O���CjژI^�U����ē�0>�K?�H))�BI�7A��"�D�o�4d���$���L<���'0�)#Pe� F�0TQ��C\��C�'��A�%Ċ�Y`� ���&]��ZM�mZ��zu�M>ͧ��'5O�8�"%������*J�����O�'�����b�`��B��80�L�P��"��xr��/6��� �Q�
q
Uo��~��)ғ���$���Ϙd�A�"оy�Jarp�FF�<qb!��8��" FJd�8BΐE~2��d8���bK�n�v9	��ʆS�:Dr�.D��ص�)#��m��?3p��'}B�'�<<*v�/�������Hb	�'���t�/L�ر8�$��,�CJ�8c1�=|O8k��]#F��ر�l��gڰb��'n�>	�S�B*!�6I�Ji�!�Ğ�lDp����k�dQ�Ɩ�)����)���0E՘bz�RS���H��I��?D��`�M��AR^}�$G�&�`�p`
=D��;�i��=@��wM�IT3��-D�� ��Шh�0+U�d(��A*?���"�O ��WDO�O0}��I�<.(�bg"O��
ᬐ�{�ވZ����R;�� @"O(�
WMK���e�E�eB0q�"O�傄�.���Q�Ň�
�ڤ"�"O��[a��R1
���T�*�ꄐ"Ol!C�+B�*�C��:Cq�	1"O`y�$l��.�f�#¶7ˌ�	�*OTq�#��
[��7dU8g�F4b	�'a�Y��"��	wv�3�bI"��
�'����	C'T���/��
�'xT�,�Vf:��6��%`��S	�'�z&�� e��a	�E?C�d=�	�'��q�"�Ƴn:콙��AE���'3.�	'C�$8@qW�S>�!��'�H�s�nٿ����9 L��c	�'�r���+B�e�t;ce�&m���	�'�P��@b%H��Y�3�hG�L��'_*�A�!X�*Ҕ<8�l�$s�>I�'�t�k���2�d��a�i��ȉ�'�䫄bX&h�B8Y�d�p��J�'��8��a�n�[w��J��;
�'7th
sυ��>ĩc��4p�	�'k��Sd��'0�AC$2I�*أ�'hL`�� ���I��C�
���ȓH�-�AN�3��0p]v(��,D��A3�
D�-���K��vp�4�(D�$��̜P�[b�J�W늤�u�$D�8�a���!Q��"��7�*v�"D� B�CB�3�U����% �!�&D�cGg�f^-��CƓx6���9D�H����m���2�!��l�(mS�!D�� t�j��աA"TBѱ+��H�g"O"�#����T�����6)����"O��+���k��`ʉ���5#�"Ox � N�.Nl~��h^�Ee:��"O8�в�ߙ@JF��c�)�r	+F�'!�'�'���'���'R"�'���A�KƇW��p�%B>lF�`Q�'���'K��'q��'r�'�R�'/dt�&���?�X�� yqA��'y��'BB�'���'���'�"�'��p�P�m� 17*�Z�4��'�"�'��'�B�''b�'���'�18�DJ-'D�V.,����w�''�'�R�'[��'b�'���'7ɻb#U;s��QZ(Z/�`Q���'��'��'��'��'���';��S�!�ʨp��\DyV�r��'<��'��'���'4��'v��'3��P'��u�v͐Ǖ�n&*���'�B�'Ub�'t��'�"�'9��'�&�{ �B+1���s�mFV� 	u�'��'���'`R�'���'���'d��!�JS8pc�ЎO�m+�����'�r�'��'���'���'�r�',�# �ϭ3:���`W"2��f�'���'k�'�2�'���'�r�'g��r��c�.�H'���r�'�2�'���'`B�'�B�'���'�0d-�1T��Ġ̦f�"��W�'���'w2�'���'�2�lӬ���O�:b�	^\X	�q�4C���ay2�'��)�3?�u�i-Q��ę1	�M�t��4!���A����D@Ѧ��?��<鶸iN���EU?U&��d�!��H��(xӞ���;6���#Ԙ��Qե��ԁ�W�~�S,P��#Cjҡ"��@7��l��?I/OP�}Ϫ&xx��O�� "e�Z�x����1��'���=nz���� ����P)Gk̃�2q�c]��MS��iA�>�|Bu��>i�b0͓y:��+�G�>U�q��,tK(�͓g|��*�%�~���J��4����ްU��T��kP&?lHL:��V�-���<)I>1R�i�2p�y�`H$J�~ ѕlN�.�F�A�B�G
�O��'$|6-�ܦ�ϓ���7o�0�� ���IM�=���P����5'3�Ae��3cF�b>���\2`���I	D�Q��H��8:eڔTt␔':�ԟ"~Γ9�X,��V�;���	�̴n�n��R�vD����������?ͧ,|� �)��UpJ�Q�#�;[�l(�`������������IЧAe~R'G�p�p��E��9+��C?��)+��g8d�ן|�V�b>c�\he�Y
�5 Ӫd`�ȅ�>?��i`4�R���IB�'H&��	L�wxv`Ul��Z�D8*�W���۴1Ûv+>�4���)���)�+K��r<pZd$�"z���
s�
��䕑h�ظ#��L�)(b�O���T�'O�J�z���Ş���I��M�Q���?Y��Z=����\�����E��<iG�iz�Op��'�F7�צ%�ܴ0F(,ن�/O����c��B�����G��
�@a��?!4��<}P|�����/�������U6 ��r_�DЋ&4�$?�O4�2�
�1Q5�<�0�ߕ|�"M��"�<!�eg�jZ������9'�pgaԄ+�Eѧ�ܛ~��p���ēW��ƍ|�~���d�8��64O8��8k��(��	��i�i�Ccr<����l�����4�d�<1����_}:����ſ[�Q���Oȸl�2Mv��'U>q��*�Jk�rS"�: �a�!?�wS� ��4N��f�2�4����@��Rh�O��D�s Y9 �Q���Q�r ��<�'#��#��\
���ui/��QF�7v�
s��"��K$�"��Gx��O$l��� C�.��؇	G��c%�we��[���,��	�����Z0K��+�x�ii��V䲩��@[��|�B
՝?���;�n����p���(�t�As�B�.�Qac
�j&!b�n�*;6A��mT��	��%H��� ��n�����f�^w��#wh�Cơ0���/W����&�rp���T-}��|Q3�ϰ6EZ!�G�ضrx�r7�Ɍ��js�Bb���X�I��D��`�(�, 8����-�&q:�b2}��&�X���@%�\���h���-D1��R�X�4��d��?X����	���ҟ����D��ោӠdX���X�hg��{s���)� �`�.qѺֳic�I���'���	���aB
a�\6M�>G�ƍ"'�"H֜�5��
��	ş�I�P����R�)�џ��Iğ4Va&U�5��g��+���
���M����䓅?��6$���D��d≴x�$<31n	o�@t��-W��7M�O��D�O��$D�f˧�?Y���
%!	�m��ܺ#�]��D��隐+�'<��'x�aF��,�����R&&H^D!'��:ޞ�J�H����'���L)].��'H�'!��S�֘�et�ȢdoګJ��	����:��7��O�����%����i��*�5��F�<�2]8Pj�Jʿ�R�'^R�'<�t�'��U>uQW�"���Ӌ�&ivIpbo����1��NBvb�"|��g\��7�By�t�Q�T�W�����i�r_����a�xy2_�H��|?�'�[:�4�P���e��eМ �1O�Qyc�c������	؟|k��OL2��3a�1N���	�'��M���`��9(/OT�$�O���8���px20��9\y�hï8&�k�W�ɣ��� �'6"�'V�T�ȊuÜt,
�J��3/Ej�-�<�*@�'�2�'�|"�'�g9� 2)�#?�!Y�eEFL�cp�Ԟ���?9���?�+Op8c��?��i��I�e�%ˌ5���ӣl�0���O���9���O��$U�|r�	�G�������8`��[V������?1��?�,O�yIЬ�|��JJ��� J�l)j}�0d>?�*<yưix��|��'y���&qO,��ۚ\3���9'��<a��i�2�'#�	�&�`L�O'��'|���A���a,�Hl"�J��UO��$�Oh$��*8��~B���<���q#�q��{7a�ЦY�'��9�c�'�"�'�R�O��i��ÀO4+�c%jB�n�A�&f�����Oy�d/�)�S�>����(0�Ƀ��9$6m��b6,�d�O>���O����<���?�F��ф܃�JI�^���% �1�����O>I���h�<���l!4���
ʣC�tcߴ�?��?�U�@����OT�D�O���bpA��Y*.+�1�2JO�t��c��3��}��Ɵ��I��Y@M͊n&���%�Y�mV�`pp
�Ms�y�S(OZ�D�O"�D%����\��#�BĔ���.V�<
g[�@Xd!#�����I�\�'���:���U�(Л��W04�˵��o�	������<%�����J�Ώ�T �q��J̡��*� �s�tb�P�I֟(�Igy�L�v�I�7S.^h��+��Qx��*u˛6�'�"�'O�'�2�'��9���O�M�GO������ь+��XZ�[�\����T��Ry2	��f��ӟܣWe]�T��X��o.(�00Ë՞�M�����?���hk̠�>�W��A�ơ���D>B1RK��������X�'��E�Sa#��O���Ơ�*#W"u|Z��u�R�P�x�s�id��쟀��/�-��q��?�MQ�`y�ǯ�`@I��H��6�<�C�֛FK�~b����V���tNց�R�ሗ'�z�+�t�����O�̣���O�&>u��p��4;����t*J�}�,���].}��in�8vT�3�4�?I���?��'剧�$�������3S�\��B��7�B�=�����OR���OH�)�|Γ�?	�挱/"H����*380hjV��}p���'`"�'��4a.�4���$�O��(�����|�c�d�05�����nզ������I'[�U����D�Oz���O<�AL�H�C�T"�̙0V��Ҧ��	<�r0I<ͧ�?q����d�_���CQ#[$�Ȳ���"�mZ��d��D�ϟX�'��'rU��i�
؍-�h�B�H�Ec�,3�G��%D�}�J<y���?������O<���,e4�X*DUz�y��+��l¢��O�˓�?!��|b/O�+�|�2��=r4
 {��SH���`t��v}�'�2�'��	��x��/9A��I�{�4!�$�ʃq6��;7%�,�,t�O�d�O���<Ѵ�[1�O�4m�%HL�H��<�d�\�.�^Za+vӆ���O.ʓ�?�D�*������%R�u���U������/�P7��O���?��&������O��D�k�+�����N�?��5�����'~2�'���6�^�혧��Ѩ8��RGN�
_��8y7e�(A��������h�����ڟ����?���u'�W�;��r1��>�Exk���M�����'������ )S������M�D�b��io�a�1�'*�'���Ob�)�� ؉?p�Uf�=C����5���M�"<�|R��^��'ې_�赁�b
�i��ݙķi���'�r��={�O���O�����(k�IiFe[ n���gA.�Eo���h��ty.�~�'"b�'Ĥ̪��Y��=zG�j�X�2U�w�T�Dڷ2��$����x�	by��r�����7E
��!ի`7�O&K�"�Ot��|�����D�O
���#GD`����o1 �#Ϙ/AL˓�?I����'�b�'t����nC
�0�����ބ�a�"&�Y+�Ov�$�OP���<iqfQw���.ݦ�P��C��Y��(
[�������ߟT�'�"�'6�ˤ�'�ٛpm3�~������#���
�>���?	���D��'�$>M[ѭсZ��5*�Q@���M3��?�.O����OJ���*�O.˧"���� R ? i�2"�3lªa���i���'Y剹!3�QPH|����1o���R�
�1��٠��l�AmVyb�'�B��Twҙ����5��Q���s�h�1/ǘl�dՎ�M�*O�XiD���驟����$D�'��4��>��Ju�;-R��4�?��P�6� ��58�O���^>7�[�6�q�Y�:BLH�c"�'8����6�7m�O���O^��`�i>��� ʌ�%���˃L[���g#�"�M��d�-�?���?Q���B,��$�O̤�3�[�}(ƭ��M�v`�˶L���e������	�x3��cO<ͧ�?�L]����L�Ф�(�:�i���'�"�8��g~��'P�mK/�:6�_��]���>Ǣ7��O���!�b�i>��	͟ �'.@K�$��Tp��RBb��^z�0R�vӐ��\L$��<Y��?�����[�Z��a$ꍺ��,��5+�Re�r��Y�	����	ş��'���'n�6m͖1�x��b�%@s���Sg��K�2\���Iϟ��'7b�C29t�ɛ�h��a�e�S�L���ҟ���'���$�O����dn����iLȈ6(�HtrU���B ©OR���O,�$�<�CT�:��O1�UKQd<ׄ����]
wt�����f����O�ʓ�?)��Q�������3� HX��L!��A(�'��A���iE��')剀�6�zN|j���1 ��S���x���A�#�.�l�ry�' ¯݇�rY>��	�?�X>`(1�j�P�4��D&�7-�<A���+Y$�6'�~B���r�����K*XiM�tL_1@��j�>��O}1��O(\%>�@��43���馆�� �ݺ@M�C�Tm�4t6�ȩ�4�?Q��?9�'����?��#j�����<dL�iЌ���|;S�i�֘���'ɧ������'�P�5��cH��0�LY3�65��hӆ��O���IS��m����I��	��]wJX!�ć6&VE�$���%�J���?u�i>}�	ğ���V�lm���D+oHE����ei,��ش�?iE�P�tw���'���'���~��'n
q�q���C��+�H��3��ҮOjIIQ5O��$�OL�$�O����O � �-� �a#�cޘH�#�,���ۦA�����͟�a�����?�s(ް#���h0�F8��k �ӯ�`���?���?�����i�O2��#��A�	I�S���D�Ʃ/��=y%I]��M���?1���?A�����O~���;����ȑ�'�"���$8}�$�Je}b�'��'V��'{re��i�:���O92��G&5������HF�����˦y�������Gy��'B�`i�O��O��3��W�
J�,U�Ʀ9�ְi^R�'(��'5@�	f�^��OL�d��̐��mh-�T���(����L�զ���Ryr�'@Tx�OJb]��sӌ(C����^z�����	
 �7�i���'O��j��'�b�'����O�r#G�=�� Tό#i�b�3�T�0�*��?��?�M>�'���1�0�x��ǁvC �A�#7��Av�g��d�OP�D�~�i�O��D�O�a��a^sp&X�M~���������ğ��I۟���$��|�dU]?��Z4Kм:<T�p�ٶ(���oZϟ(����Ȣ+S��M���?Y��?��Ӻ�l]�\�P��dm��&l���	������jy҆��yʟ��d�O>�D]�,z�-s��2,���Ht��}1pDoZ���P0���M#���?���?��S?���_��X��Ԉw�l�8a�C)�~M�'(�*�'�I����ߟ`���l�7 `)�vHW�h�$	��,�:<޴�?����?���O���iy�'4�h��̖�R,�f�AJ��%-�1�yB�'���'���'��S�2�v��4\dʔy���v���" �!��ò�iZr�'e"�'YRZ����L#��ө-6N�8-=hR�������X(Zݴ�?i��?���E��)��H�ٴ�?�gVp�bI�-�<Il�	.@�趹iO��'c�^�8�	%{�����p�V]L�华zԀ����Q^<9n�ПD�I�0��G����4�?I��?9�'6H��M�(1Z�[��S Z`t��i��Z��ɻW2��?�禍zPa�	�:5cS�f�6ldlm�(��6���i���'���O�6�Ӻ�3O�p�.�H)d&dPx������ş���!n��'���}��g��h}C��\���݋�G�y��l�M��?�����'�?����?Y"��� �`
�a������q��f� 3b�'��i>a$?i��I0� 'L3KW�M
G�*[Zz���4�?)���?�B#,����'3"�'=��u�4��%z"�4@B�:C��M����V	~��?�������I4n2�ӱ��1cM�h#�IC�^�� ܴ�?�a�TG�F�'���'Z"�~b�'kR8��b؝Dt1IA��*[N���۴�?1b`M�<��?���?!���?)�	�:�d�(u��x��Y8i������2B��'���'��C�~*)Of���iwN�p�[� �=$����7O����Or���O���O����H)|�m��T�0і�ѹ%?�-q��ӷG�ʑ��4�?q��?y���?)*OV�d��J��Ɉ�3�Ұ�ǎ�nO�$�)tc^��'�"�'���'h�D�!��7�OL�+i�r�i�wȈ-AЪ��KXN\oZ�,�I�ȗ'�"�����'&""�L�t��V�ܽy'd0��O�"(�7-�O����O�����T���n៸������(]�x�(�i�I�Q�P�C&�"D
�4�?	/O@�DK(?l�	�O��d�|nںQK)�K�?�T8%Ƥ�`7M�Or���"j�lZ��I�@��?��	-,�xJ#��J�2,�%��?��O��D˦ ����O>��|K?m�-�uHE{��b/l�-t��,�w��馭��ɟD�	�?����D�	���K����#�j�{G!�#`p +�m�M�(ݾ�?a����4�򓟲�D�M�(��2G���[b�)5�B���i^"�'C�	�2Y��7��O�D�O����O��(T՚�o��	�PMs�I:;9��'R�I?	��)R��?��O�z��%�kZN���e�>}�B���4�?�E%��*��'�r�'�Rd�~R�'Ĩ���G�H��CȒ:zנq��4�?9W�<���?y���?������<�u&�/�HEr�
V9jj���$�Nq�����	Y����Iocf��D��P�5����'��Gk�L�'���'="U�q�/N4�����|Zi�	;d���Δ����OR��2���OP���m��ɟ3,���E�M��#rʁ�?x���?���?�+O�	���Y�
A��B�c�O�\H%g�� ��ݴ�?QJ>9��?i����?	M�TQ'g�/�P�Ce*&)��9��sӐ�d�O�ʓA�~������'?�$f8nPtY{Ď�8�D��фHD.��?����?�B������kN���e	]�Dux�/�)]��oPy�M��~R�7M�|���'f��
=?�7�� Ȯ��fL�s���#!�ަ���՟hR gY���$�b?� �x�H�Zc���6M��
�j,"�i�F���l����O��D�č�>Y󈎞+��mj�GB>Lư�ȴ��%cD�V"�
�y��|b�i�O�ˀ.��l����D��/?�H@J���Ц�������	&^��} J<����?y�'7(@�C>1�d�+���$vj�4�����Ԕ���'}��'и�T;��ӆǝ�"*A	��f���G
� �'���I֟@&��*I�8a� �	Ʋ�� �B� �O �͓��$�OV���O�ʓu��Y��B�s�`�� ��Xfȅy�f�9�'���'b�'���'��T�
�rB�0��A%	Zҝ�FP*T�T�p�	��P�	PybU�k�	t�@�!�6tO>���+�`&���?q��䓌?y�`�2�ϓa T:h�=V5���ō�(�A�T���I�p�IBy�/y�����*�~Icq�ؽ(�&0ڦJ�̦1��k��؟4�I��ID�D�jEK�*Y7�uҁ
T�(�v�'8�V��Ȃ"�<��'�?��'�81�[�o�� y㉐�ghB#Аx��'�B�زQ"��|��H�*7D�6;a�@0�u j�7�i���a�$��4Z�ܟ���1����&a6�HQDV�ku���q@ϒ�6�'��DN�36���)�R�ر���j���f і"��fA��0�^6��O����O��iK�	џ�r�͒nd���$�=���J�a�'�M{"b�?�O>E���'(��#����Aɐ�x�ݠ	�Xy��wӚ��O���1^�l�&�0�	��8�V��a�L��h�P��//���nJ�	����M|z��?Y����3�$C(K̾���18�>;��iG"�-3\�O�i$�mh�%J �E0�^���1l�2)nZ��lc"��ޟ�'���']RP� ��b�2D�>�c�m��t��q�XL<����hO��	 D޼2A!�49X�I`g���_UN7M�OH�$�O�$�O
���<�)��^��i��A�d-c���K窡���C}�I�XG{r]�`�	/e�(��a��qp���2z��z�4�?	��?9����P���%>ט<⦘#��g��@@�G>n��6m4�����O2��?-	Ċߗ.���0���+� aJn�f�d�O����OL�ň������������?���A�m#�Hr��z.���seȂ�M�������OH�2�ޒO�iM�$�U�]�~���-Ѭ	?d���4�?���,2`�is2�'0R�O��$�'6h�rL�����̚�.�����)�>�����)�����|�O?)��M�-��p&�YK�話� c��@�r"���e��� ���?������I���gF0*TYIjX
`� �3҈6�M����?i���4�������	�@��r7�j:���a�X��o����I�����E�=�M����?y��?1�Ӻ��D�ujn�@'Vkd�������Imyb��yʟ$�$�O��$D#m2�A�*��W�Tq�ցO/QdLn����p@����M����?i��?�Q?�����"�7E(�B�BB-@��'� �'�'�B�'�Q>A `�03ЕY���[���`��k, ɔ'��'"�|��' ��I:w?�� �]�#�b�b�_q��q�������O����O����O*L��nK���P=�����,P.�}ᇈǮ�M���?����?эZ��ON��FO&
�(�J�J���Ё�^�t�I������L�	:�z��O���&.Ez�y!��&��[.Ȋ����'?�'��'i,�RW�A��ē5S������.蠙�3+�a�nTlZ� �I������V��(��ݟP�'���(e�<��hߕ���۰f��e�O&�D�O���!+�<X1O�)\n��p�"��!˾��w���Mx+O�� !
������:�$��P��'3���ǀ��֘i��Z"o=��bH<1+"����L<y5�O� I����BL�<Q����B���	K��Hğl�I��<���?��֟��O?b��LH	.<)@��W�����bi�^8#�a:X�1O>���&!�*�K�+�m����\+6�{ٴ�?i��?���ۢ,�'(�'�d�-h2�
�LG;R���q3F��O�@���OJ���Of��5���6��Ғ���]�N�0�Ō����I4~�(��H<���?�M>��8z咅k_�D�!�vH	3����'�
iʊy��'�2�'��I`FF��'��Ht���7��V�2������?y����?q�C��
��;z.P���둷
��� jQk̓�?����?�/O�)�qB]�|��)S�~t�z� ֮o<a"�-�\}��'���|��'� �=����$Φ1�1��P���p�˒Tr�	ݟ��ʟ��Iҟ$[��蟼�I�0qv�A%���6�H�5�sDG����	]���� �I0?���@�l?��[�d(��\4fKTU`3M_3VΛ�'��\����&���'�?���S��=;����N����������i��O�	à�s�.0fJY�?D"�Y��v�挛A�i���'�нp�'wr�'|��O�b��5�C��v�h�2���3%'0�q�M{���?����L���<�~�A�D2^0�&(S
ִ���HIצJp���M����?	�����'�?!���?���
)��U��I+_ڙ ����t\�F��d=r�|�O=�O�r���h����G
���p��`۬6��O����O��lDզ5��៰������i�����o�X�ۑj47����ac�4��<yt"\�<�O���'R�=� 
[嬌*h 1�����-k�i��@ݚ`�6M�Ov�D�O��dB_�D�O��)d�Ӭ5�~�h���
�(Q�i2+��y��''��'�R�'b�'L]��fA	!y�$H��I�P}$Q8�� �<�6�O����OT��B�$P���	=bp��Q!M8sZ}�V)۽-�����(v���I矈������I��p�ɧqY������̸7"׈�2%Pv��$��i�޴�?1��?�K>9����Ԉ1����ْr  ��Ou�Pj�U����OT�d�O��J���i�����\�Sg�9��V�O�m�$CψR��6��O~�d>�	 >"�c?�+��޺u��1H��] %xP�gv�0�$�O���O�-p�@�O���<��',��d��E�H����;.BL���x��'v�	�a�4#<��	��p7$R�S!f��%���n�}y���7ג7�m�$�'T��B9?���X�Q���"\�0��T�Y�9�I��h!/;�S�L+&T�P&�+ulL�i�$�3K^�9n�+6��Lc�4�?���?���O��DJ�R= �C�KO�;3�%��#��@�D|n���#<E���'��iK��5;�(�6��f��W�^�X�ħ<�bM���D�<����~�(�#�p7��yGΰ��� nt,"<�7��4�'���'�\sb��af��6i�;`�T�%,dӢ�DB�t۶�oZ؟P��џH����Y�\�Rm�=���PLڱ���C�"��9���OP�d�O0���OR����h�I�ьۋ#j�4�ՅM�NAx���O����O��%���O�ɍ[t�l3�dl�Vظf˱2�
6m�,��	ȟ��I��<����t���(�%M�~аp�����x����M�(On��$���OlʓS�Z�mZ?
���؄D\�p$i>>���?a���?�/OT��G�^kⓏ#z��"A�~��=�D�=@�^��޴�?���'Fl������W��i2PBǐD����6"�9�M���?���?�"@4���<9�'�f��1!J_ ,M��L�Q˔`Ѧ�xb�'��I0v��#<��Y��p����di���h��$l]y�`���.6MCB���'���"?I���;����(_�2�&�	��ԦU��Пl��G5�S�'*E���㓴B�h"B�_'��l�|Yh��޴�?���?��'M҉'r��j^Z�i�� d���5�6-�gI�"|�%-6�����2]H��Q7J"s��E �iA��'��g
<O��d�OX�IU:Hqg.ٚ�B�[�&��/��c�Pa�D&�;k�n��@C	<Gg�-��D��m@���P�F�s���*y<�ł�2����'>`lq(잰���#ME��#���t ����+����a���<P���ɴ�J�#V�L�4���PK8'��[Q,�1t����S�� �l���̾#����ԍG� � ��M�L��0b�ϝs�(Sb�T�VD@&��=��taq$�?��ݢ� �Y:� p�J>$-Pd��4g��Ɂ��|�ĩ����TS&`�&�&�����?�g�6�?���4�=JJ��CEf	���0��h��6@�ȤI �	pf���63$m�!�����6|8|9׎��I�4j0���`x}H�@�u=��ӮJ#P���1��`o��Fz���:�?�����D0y�Ic�G3nX��� T1O��D"<O���g�$VFs�D��g��WORynZHT��G_�V��L��H�|�`��ey"�^�mW6=�
�d�|��NB�?��lݽ(���9�+ŏVq�43�(]��?���+�4��D�f%��*U�IXB���/�0�uZ>�â���z�����3>B�t���.}"�[P\,�G��M9p�*!d^�.��Y�U�EA�$�گF�n�z�'���܍q2����L3�������������c��D<��s"�:|����m!4���E��:�G&�6K�R� :O�1Gz�"\�k��p��,��B�?'�7��O��$�Ov��e�{�&���O��d�O^8��G~)2�N"Y<���ƌ0M P�1b"[~�V� �!���y���
>�
�+עL
�Z�����)T���H��YF�Ih<q��'[�����_4�|�B�͇P�t�Q�'��6��O@����O���|���O�D�OĜ[ ��79c�P��ۻ4퀘�i�<A����<镭��<y����O~s��}���s0�>j��E�E3O��d�@}R_��'?��'�z�n�:O���D@�bX,;���J��$���'��'~�n|�e�	ßd�',����h�\6���k[�#��M��o�8����fA�p�d= A�Q�z�D� n"ʓ$��[d�(�(�ÀS�=���1QjB�fAj�r�3<`�� ,R ��"�bK
����H>�b��g�:l*�%W=^̈́��%{���I�G{r�ē	_O��CE�#.)��*��ʼ`a|�|���"Rs8�'d�^�$�C���'�7��O��lۚ�0��i��'��Ÿ�gZ�A.m8 �ܘ!aUS��'h�GJ	��'�󉒎/�(�'А �US��!Xΐxbƈ�i�up�� �\�)�B�^�����h��q�O �i`���%�6�b���U�H�%-�P��D�_�7뾜)���o���O��)��'
�'c6\�`'�;�$8{��[�L��'������-�$Ș�@FJL�ˎ��)��|�i�2��!�Z�X��m.ӌ@7�|���'ێꓦ?�*���yS��O؀A�L�Q��(K��A>��w��O
�dM�b����L�N�\ɂ5O��'��� 8t\J�h�����^�=���>YUcZ�w���z��M��F4£O�H2x��O|J�,;�� �Dd��:�]c�E���&O4�Fi�
�m�ݟ|��b)� 'axq�C�o@u0��D̓�?���=�v�WXf-�Ѫh�<���	�Mc�������O[[����B��yi�LkѸi�R�'
��X/�܊��'�2�'j��wD��!�O�}^��u����|�p���q�Y�t1[!�\�`iG
0E1�<��#N��y��ҿDK�Gȍe9L:�@�?fS�}s��MFdYF���c>���T�\�1v&��A�@�Z��q(�3��� =�IIB�F��J+O�	�!�����O��O��[קR��Pͱŕ�#�SF"O���LɃ=>���"�>\	:�4�������ЦA��~y�I�_��l��e��?��K�*	`�n�;�iV�]TR�'���'���֟����|"s�V�9�j�hP�ܸe�V�����@N��l�5�f1�ulA��Rh�d���*�<a��L 'P��@K�&6�qۀJ���iX2%DW@XӁ#:��1�ɔ<��<)�㉇N@Va�.P��a��%>}�I⟔��[���O/z��6�^��Fu��ĝe��'��0m �/����u�����<!��i�P��*I�����O���ܴL2�Y[A��5	�z���O�����"	v�$�O�� }@&iI����%@J�ҭ�g���D�Q9}d��K��Oa^�C)R{�'�2Yx@�@�'�~�X��L9|��Ѫ���Py��mO�?�D��l���0<�S�ϟl��Qy����d�JpjpJ@�Ă@ 
8��'�'<tX�D�:60���O,Xd�#
�'Ê6 ,>֜��c�=A�`]ReD��f;��<	�i+��OP>��!�Fß��*V��I!"��b�R|I祏���SN�5(W^;"��@��'�		��V��x�O�h��B�Հi� ��Ba�9Y<ȸJ�H�T�ϖ�(���M4bxSjU�K;�HX�!�.>FM�;+"\��b! b��E���޾O&�O���R�'Ì6M�J�ON�%�����k�"$ �� q��Ĝ�b�ve�g(0)Dl�`��]*���=�'"摞P��_����%�F���px�$��M[��?��5>\�V��<�?����?����!I��7�̀�G&�M�R�x�-L
+�N|
0�ȜJ���'mƍ~�\��I~�$���D��͓XN`�jd� ��H ����Io��)��
�V���BLI�n
���Iܧ,	�̫��Ot0�'��#�
IQ��59Ti��@Ц�i޴�?aS�D��?�'�r���?q���?9Cj �[&^UEB��8���C)����?�����P�RW�ɒJ
�E�qh\�^�DI���s۴��|�q����<�Q�W����Hr)U)2<��;k�<剠�C
�?��?1�����O���t>�ga�>2D��g��f�.�j4G�	,"���CP/I:�(�I�2r �fc*l��<��g0��!�B�D��E)4 �=:��83�����{j��;�m�*����@TM� H�I࣍�lJ���6��7	|��ަ��4��'�Fb?���g¢/[�i0+kݸh�-D�S���@ *H��عy��0 �)�	����<IS���	��ع���=k���:�Y�/�5�DeRʟ����#.�5�	��$ͧB�@D[!dܸ=�����	�1��5:�)3R�?H�KQ�Q��P�4ʓ(6��H���1�r�E��!?2�Kw����Kg��B�d�a��R��M#����J�P�) �|���?������٬5*nQ�*ԇ^ L)�c̞�1O`��><O�`�S�!U/2�
@��&ņ�JV�IQ�����l��ɳ�l̐�p����{�X�V��Ov�o�xs���D�'��ӒB����I�CZ�A0��K1�b�Q��K|��	ܟ� ���:���%p?A!GfF1��̐�#Ph����X�\ �A,�	y.�i��b�Đ�$�t8Ѥßu���	[rM�]8b�H�mT��o�uI4�CZJ�� 0�f@�`�$}"a�?�a�i�#}*�'	+$ez�@R>���!Ai�Ae`�'fR�� ��.�r�-�hH� �i>u�����'H�ް0p-��Hm��������'���'$J	з�?ib��'�B�'����4�-�6�ӸT��-��dZT�cϚ�\��1�f+٤B��$b���t�'u���+eCq�l�c'D�j��mS<x
6\��B	
V�R�H �6abv [.l1�Ƀ��iT�48�Q�w'��Qdc�/�2lT�O<<����x���'{����|�'��'���"Hr)�C�7���
�'��KQ)�%�q�(�9��(�'�O%����'R�	$\�N`�TNӜ,�@��^S�"A��8�.���ȟ��	��@�\wr��'X�)&5�d�	���.w�*�R��$	�E8d�ˇ0�flJ�/߳#��9��I>��a��(9� � Ï_)ZE�}hV��)���ꏗ���˓6Ql��L�P��&=q��ҩ��� �4RǛ�D�q�j�u��O�bYZR���\tL����Bj�o���Q�i�&"�Ρ�<�DU���'� )Q��>Y���X�qW+@42RxX�4��+�n���?Ad��?�����tύ�ax���F����e	��X�Ƙr֧�1=����P�(M�=	ۼc�(�A���j_�[<�h��
�P�q�@6� <�����2 �a�-J8�hҤ��=������I);n`�$�֦mʬO4q2�ˉ^ꖹ��kTS��õ�d�O����\�6�S�h�2X���H���%>���D{�O 7MB	�*�g�P+y˔q�`�Ƈt'&�D�<!��;��'��\>M��H�ǟ\�d�C�j�:�A6hخ?�ଓu�֟T��B�Zq�*�'c+�陖h���'��靲V���D�T,A�9�ĥ�"l��~�Z�s׭G���=C$�:�'-ƞ�� XT��Ӕ�OZ.��OU��'v�6MV���h��3�@�P��T#)d� �@����<����<���]��LP�ǌv�N��b�_E��c���C���	d阃{Dd`��@��E��'x��'x|Q��awR�'R��'� ֝o���ÝnZX�����2��1�5c 1f�ܡC �tb:� ��H�'F�I�
z����Ȼ6%�P��EْH�"Hp�S�K 
 ������)B� 2�I��1�ڬ�'��pA�oU�0�ڼ	�j\8M
�ie+k�b��'�<�a��|Z����'��E3fo����9h�(*�+
�'k���F�=LgL=Sq,��*e`�'��)+ғ3��f�'��ɺ]L>�K�D���.[�^0ɲE��%�z�C&�B���Iߟ�I>�uW�'��1�0{��/AI�]��SHK�({rYY��W�.�ɓ���~#рO������P��P,9A���6�
8qRg�U�t�y���4{@I[�Lu�y[��g���8��d��;����i�q!)U�f�:�'�H7m���?�D�I2e�4�rb�dA�Qj��8�a|B�|�ጽQ�J-��=z8h���,�(��'Ǽ6��O�ʓ<�	z�T�0�ɱz��(�AE�d��Z��ӺF�ƥ��ɟ렀�韘�I�|JQ���Yf!�׭S��)Y<@��x�]�(2��Z�gؠ#��I���j��EyB��lH 0���S����$O��?W842di�Qj@i1N�-x���͸w���d��!�H�$���d#�O�l��MS��д�J��_�_�u"�n��ƭ�)O���!�)�'
/�!� m^�jtiBU��71��Fx��i>���41�� ��'�UJ~��ml@�]���DY�	��v9����|ꖦ�?�G�I�"����ƣ]�Dз$_��?��#�����'FJ-�q�$��KK���gxd��/��
e��3A��fS�Gfda�>�@�^�Lp��,�s�n	�G%Wc��͌��a2_wO�� �J��
9y�/F+v��܂K�j�f�O�mڅ�H���)����#!�C�tj�@ӆ�ޱM{�C�	<c�,��C,I��|I$��/yE{�O��"=#!�,�J����@}�x!� 5���'�2�'8�T����9!T��'���'b
��\���Q�3̞=Z�(E�}j�:pҢ����3]�ZI�EJ�O�̭SBn_�yB	�
�0��gH��� ��ާnDx���OO�qH$b��,z}�F��>>���'at�owޡ��e��rP��C3���F(f�
�h��4�?�#׈�?AÝ�,O��� �RS�q;�#��B�]�����CnHB�	\���a��H���'�b���Iٟ�1�4F��6�|��O��4[�T��'<ɖ� d�^ 
�@�qg�#, Ys�H˟@���|�	��u�'�2�'��)�-�/&���Rp�ˏJ���b0f+m���o04�fL��C�<l	�e��6�(ON��p��+4�ą
�n�v�;R	�h��Q��}|r���lǡ3����U�0�(O�cꀱD0�E�<Y�9Ywf�=[���'��6M�O�ʓ�?y���)��t����&-�p�*�Ą7�y��'��T�`L�)�t	1OS��ܡ	q�|��q�(�o�H�	ßT�i�!��K�1jI�)a�i��:k�H6D� ���$-��R�@!�p�;A�2D��iSA�����F�A��h��,/D��je�� 9��4e�<�v�yR:D��Z��O.3�����$IO>U�� 8D��x��ShQ�WĐ^��$�):D���=.*�E��	ݒ�i��:D�KQ
��Zd�PY���
�pE��6D��QC��|ݖTvE�h���o0D���́cxD���E�%BjA��/D���ꊵ$W��"SO��B�6j.D�,� O='D��I������b"8D�X�4��;��c� k��U#�-6D�x$�6 ��sp���;M��ta5D��P���e�V�0�Ŀ3N�A#��2D���D��,�)��+����Y�"c-D� �C��n����%��B�p=yP�=D�;f�f��;6�3z��)U.��yR�G5v5� �N�������� �yrһ:[�D(�l�[B0;�	�y
� ��fD:%�p���A���� "OF9YѬ��n^m�C#\�K�X]"S"O�h�w�@�@�*�/�&K��%�e"OB@W�ܓ6n�	���N����"O��SӋ�;&���)/�~�f"O�!y`��   
[�)bܓ�"Oh�DQ
�XDA�*C4 �/�y��Pc�L5
���?�(�ş��ya�#���D��o]>T��Y�E�&�3v�OQ�M�*O���U�yw���W0ǒ��!�=	\�s�k!a~�/�
L¼a�*¼]2-#$`��MS�A�,�ZD�3�[�%�)�:x��Ć�e|�㠮H�o��G{B�'&���b	?1D8�)��K�~�^$Qy���k�� ����Թp��D��h�x�ᱩ�1�2�8&�����)̡4M>����T�&Z���cS�!����٧R���H��P�?:~mH0,G�����\c�� *]�ʶ��חX�*XB�	L!M ��ִ���K%����'�T�!$�[�tU�qf XP��s�DE>����SD��P�D搤|��U�̤kq�X1��I7a�Hȳf ���xb͈�f]���0Ȁ�g�F�Qpp⴮E�W�j��;�B�$���z���p��}IP�F(������T6f�<�B�$!�g��%�s+����}jp"f��'�d�A�?�<�+�.#k�P���䂬1�(��h��9���`@h�=j�󤕮R����
ܰ,�Q�ElN�;9�V�BzcZ�R�U
6��Kr/W��O a�g�5�>�ɀ.SF�P�!��S��ÑP�0a�1 �?�_�����=L�R���(IRD�-^a��y��V��$H� ؋ܸ :te�l
had]��p>)Ш��1�p����#D!!͜xlry�"�w��̋�.��o�q��(ިL}8 \�k\\-!�'͟A	��d�g �Dh�\��b�|��HgD�~��Ŋ��Ɛe.�i���
	OD����P�H�Ĉ��ְ%��k���*I��ɭ�� ��F�#]�8�w��'�F�e�=����<I3�F�@�|QF+ѱnԜѹa�m}¢T�v@D"	��a��H���0G,J�iS	T`�8�e@�D�Z	q��I�q�2��6M�wdY��A��7-O�7]ơ���.o�(�Ch��jc�OP�UېQ[��]����@�NZX'�uS�	�uN�4��)@�	#K ��!�R�lxry0�I��T����o�.ـ'�W��	K���'�(IYc�zոI�"��À��+�m��«��\��u!�<~���K�$Y+�
�[�ߦy(l`���ڂ�B��ߟl���!�8ݰ!-YPx
�Y��?	��-)I� ��A�^�g����(��>4�"H`�=1VJ�SD��Y���Ã��$,���_�j�P1kN:=���)�̱-��Ż!��#Q������ra���N��hO6AI�)� �(�#�%F6ܭ�c��zf���C8IHVG�N�|�ߴ��<�<P�$�@��Q�i05h)�W�x���>	�&�:5� Q�>���GG�"�MX�o��I ��#�d��+�`�:yK�lBp�;a{Fy٧+2ҧ֦%�6�n֮�1�+�}m`��>I0NO;X�Y���ˬO��X����_�J�.-�S�ڿkaf(s�nW�F��e� �� :���n��}�
����ע@�<���E/B��Rjk��q��K\~�R�*D0`�*�����ߘ���yWL:V�Ңm�?)�
X�_�;E�%�k�
-�����M�-��
�bH�t&�$��Ã4V�%�N�KPo�'{��ݶ	�JrM|B_w�k��C�	�s�ՙ.�L��bjU��PX�5���w^�G|ҍ��0�L��t�i�	�6) j�g��n]��9��*� �'*�t���*��D�P�Wbl����t/JiG,@p��Q�*`��u@	���'�xR�jÝh��������K����A-I�28za��(6$˧+Q�-Ր0%��WV\aZ�jS�<:�)�S��.��|��t@��x�p��hX�>>J��c]'d�`���:>
�����O�J睙Z\]�B�G9n�أ*E�R�:�5��5j��T�J@�d�7W��Fy�"�-f�깪��Ӑ�Q�piE�.��I�U�}24�J���t��L��qQ��R����)J�m�2�@���Gq��"!琪�E��!3�Ӻk�]r�ͻI��x�"_�V�82�M�y�P����!��jA�#sn�u�c�O�C��OV0�'�ԋ�`�I�JR�@�( a�}� @ J�XLZ�Ď�^���/��~�O|�h;��W%R�r9������J8��o��SxT � �IVȩzL��IQ,C��	H)g��.�-*O
�9R  �^M!X�ؠ��P�c� ���4��Q�S�'<\p%��]���f�Ӆ(���9"@�7Q.�O���wL�/��]ȳ��}Yly���A�D,j��(4�5�U׆7�ui�'*�3C�V�~5�my�P�BT�}rF�	O��و��
w^lK�A�'dܑ�У��h�Ρr�ӼK$�#Gń�1�� &a
�xc�ݸd"n83�L��M� H�8/L�M~&���� �Pa ��21��}q$��H�ax�9o,��c��9E<A���e�
H[J&���� �Z�N��#���1᤬h�mٛ�'a��j�eɻ?����Q�ę~2�i�fԅ G��vi$'�@x���Z�����:��������l�ҍ����!���b�8/��Y��@�JAX3(E�%�(E
c���P�����u�Bd޼�,q�#Yؔ��f@��(O� l�p��҇(v�i�Rp8�����V/7.|n�.T-�y)�
��x��'�P�B���"�`ha�ݟt�x�e�*P
���g͑SJH�c�EW�G�� ��@��p>��-�a�X�$���R"`9�Ə�?�pz�O,���%^d|y���|�c�h���wN���siM��x�[�t�\�	�f���Ҭ�id9��v��9(2�F�~Jd�`D�	@���a�-��+���ON�	�()�q/_K�2p2���Ëu�|��#j�CQԩ�
_-�M��!��L�ć?~b�!9I�
N1 ��N�>!�ˏqqX��%�36���E�RR���)Q�Rp8gK� �\e���fL)�ե�*�	�G���c�Ʉ��*i���0��ap�,�<����"0��"͟)B��D�쀃��I8Y	ZJP,��M���=��>��Q#7���(K0;a̡�&璙;њ�'�l�0����k&�Ol�p���o�nEh��*H�#Q�2�MY�C�'$
�P���-YO�-˥�2E�(�B$��!�E;� �.S�n����$;��MX�SI�	%I~�=p� ��'���ab̍#�2Q�`��!�����D�;Ä���"��_�����Ty̓k�����D��L�7D�j����K>���G��-5��9���S�d�1��8t��0C\ ����uʖŧ�/�,Gx���ī4��%��	0LF�e��ä�Z�
#*��W�@���'�J����Q��^->�HK��[���aP�8U��ՠ���phh��$�&��=2���!�S���L��{��<�zɊ�#�Avb�$D9ɼH�B.�:}�t�2��'�$|#K�;�l��c�`ER�ŉ3r���0	�0C��S�n:|�����7&dse&*zᆁ���X
<2&`�w�L$�@�I���j��UJ����*�TH�n�;'�EP�D�${1Of ��ˠ$eḧ)ͽ|l����hfg�,
�.�;���î˪(�f "�ۀd�����`�i�^p�F¨	*��%��6����P�$����Py�'���8�Ĩ�%뎼`�mZ�
		q!��F��:��I��'����C��8F�`
�a��D������߬��$�O�=�'�y7 >j�9i4�K�v�����b���p<����oQ��a��O��z���_�`��0�̉j��T�n[�U�=a�l�D=q�
zĥ�үV5F݂���څn� Q��ۦt=�<r�m�����їiz={�&�$�@�ԭ*��O�R@�(��(�gBɤE����`,�O��䙒?��MX��[�LF�PD�BQ�Jm�$V|��3�D�;nZ�|8����4P�H`���d⟀Gx��M� m
����M8�@�Q�^z�ޥ֮�;M܅��Ӽ� I�&||d�����kOfU�,�R���@P�A�q����'�"&Т(�,N��O$���f�ܑ�G��6M:�=O��-�8T�_�3l!B�Z�o2Iy��$�>��'C�Y6 @�ؗE��=)͙��尒�F�.����R�6�{%�N.�?��A�)| �E�O��I�x���g��k)����,�=]؅��O�\IU�4'���ƶ�H�#��^+��'�5Y���i�������'����EI��H���(OZ|�<�������ā�FS�\�ɚc���H���c]<h�4dˉ��O��Ș/O�� � �4�%�4�� ��\���>H  �#\��?f�dJ�����l�$n�lH���!G� 3������,0,�İM>����.4$���'^[$A��S)M���@���2rTx�?EN�j?A��C	=��B��g>y�-Q� ������D�Cِ%@0��2DGV����&����GW� ���Ӂ,H!S�p��'rm�=�v՜E8���c�H6�ahV��#/G@� K�:yN��"�	
���t$ړQpĐ{q�&7��i��_�5��[�G�O\`p��y���Z��ۑ���}�i�7N�q7�=���9������_��q{e���Ol����*k������I-\^X�#Z�pJ��J�)�R�����}¼��g�	�4��e�&!��i����[z��P#�[�mR���	�v��<�Uqs�.�6�3�o�8H�܁�=�#N,n����ݺln��~Z�y�gQ��n���@��z�������%	�����!�J�(�v�O�"�㉑Q��u��u� X�_h�1K�	�f��`��c^�ʸ���6L�i�A�I�tؾ�S�0G{�$��:������DpO�����Ԏ9`B�'�Le��=;^�؃&��z�������[?Ȕ�ԣW�:\�D����R��Io����]� 3�Ưe � :��^�sc��g�ȉ�ΓS��483�/��?�c�ة?k�X�#��eR���;qƆ\�t��0ˌ�&�\��Py�A�o�ΟJ�%C7?L< ��ۗR��ek2�ƚ#�hc�di6�ֺcBht����#2�|+G,�	�@��U�����l�H9p�\O��0���~N� *:@�-O��p�'`�4�S�+e�vi9�,��n�j��A�q��P�e��cMb9��'���"�+X/��`�(W��U�G2>�t����*b"���I`ܨÆ �-0�^�Ⓩ��yRU����n� ���B:!V����1E�܌:%b�A؞8z"@��/T{�o�,N9 m3�&J>��� ���|����� q��A��F0-j��[�X ��o�76�}��,�%X�Cs#{�Ak���A�ΜI����sMC�,`L4ݭl��٤ώ8��IH�!�}�^�E%��c剅46�xQ������'�2��x
�KH�w�楙W
�!��p�T�,���1#gO�=��!YV�ޣNwL�Ȗ�I7z椛S�a���L>����Rr�%�Ͷd	½�S��Lޞ�z$-���M	(�i�����h��z�A��V.~oZ����O���!��1xŢw�C�'P�]:4� \D*6'�r͚ТF�Y��h��'TXi( �t貘��d$:�*�����[� �nj��D~�-Q3j7�}Z1Hϊo��uQ�2]P�%���!5�&XH�epcF�	��̺U�	K��g���d)Q����U.��0�p����φM�xs���L�����Zy�� `20�ӢG3w�%��i^E������A)ٸ1� �[S�Ȼ��T�l�AZ����P��%���L[@���غ5���1Ov�0g��tԴ�!7X%�m�,3��HCEK!>�BQ1�'�%��j\�}�NX���!�Vt�q	M��ՙ��J.`��ɏO`��Q� ��j� ĉ�ݦ ���%
FE�$AW�A,��$�����I@��0]��j�FJ)���;EV�t�	zyB�L�@���eߏv褕p41�(���fז����@.j����t�'yxQA�m��+�rh{���l��p²G�%�j��NN	���>)��	�U �y��dx)ˇqQ�D1��\?)���V@�#�xU�G�9jyh9�f˹>�t4���(� �'g�y�D�v��	k��]�y���,H�gJ�j����p>1�iC< �B�k��w��`��*,C6���i(p,��?�\�a�O��i�����<OQ�#��u.�WKޜ�yr��(�L�tJ�(�[58�p��"h(L�pB��?�Q�Ӯ��O�g��ִ`P����o�M�BYhh��dJhN��ɔV2�Q��oD�C4:MB���`�#7��>|F:@�#,O�� pJW�D�X�gE+1�|)�"OV5p��8eU<Q�Ag߸g�:V"ObiS�FQ9�l��ϛ�n�M��"O�8�d���s��,J���'"O��
�H ?�\��k	���Y�"O���ꓛ
�L,��=��$i
�'dҨ[䉗*P$
-i��D"B�d��'T2)x4
�h��r�g���(�'j���@��H2��	bT*3l�H�'�4M�A+Rj��dKBB3s��@��'P��
U��9v�J@K�/�|Äy;�'b���`�'Px�P�$l��y3z�2�'�`�z n�J[Љ�Ԯ@v�c�'�J1a�Np��uk!�"pr���'��S�n�-=H�h!�+�3_վ�;
�'��P5���ud�A�'�KQ�@a	�'��!�e#-r��HB�9����'*�����!c��҈΢:&`�Z
�'���'l�=!���ir�6�:]I�')����+_��	K2aP&+�L���' ����#pzH�0"�� @N	��'�$Պ�X6�Zձ&i��B�����'��@�S>Z>%K���e�:���'T0�C��?a����OY#'O���'0(0hGM�v�y�ρ�L!�y��EN�b�p�nExC��Qa���yR�ں���+�u��l�����y�B�&`�RU��*Gh�=r�-��'*�A�d �=3�mc&�H�fB:9#�'r~��C������g�'��X�'�r��`��h��QaQ)9#@�8�'@�� f���fj�"_���P�'<�|��N��c{�dB�'�` &�
�'�ܻ�K����*Zs���	�'�$:�o�n 5��m�R�^��	�'D0����C?��Hfi��OC�\��'�kd/��k9ʁiS�>�VX	�'jN؋d+ҳs-^�{�́�֞$��'����j�{ת�J���S�)s	�'=<�J�� -�l��W
�'�~���d�,��%
d��!&ɡ�'��ee���$�@���D�	��1b�'N�p��R��PMCpy)�"O�����>�V��G�Ɂb��8s"OReT�BA?�(+�`��k����'
�����?N�jXB �S�y,����� <q*�O�$}�p�J��B�P�T$v"O��rfŘ�t�<l���f���x�"O��K�o�/}QB�r�T�N� k�"O���҂���I@�o4v�ac%"O� �	Q1]�(��(ס"��"ON���.�	 >��q�b ���"O�P�(�􃦣M�2�z"OF�y�L�,$Y�a2�G��R1$4�%"O���􎝃&Z��jTi�/YNp:A"Ol�H�Ӕ���+���9��P"O�9����.-\��h�R�.�Jk�"O��XV*�w�$9����#�M�6"O4UC5"�;6֨��Q��jha�"ON�P�)�&vJ@����h�5`"O�س֠� H�HYR��h�r"OV��rM�x�1 �	چ"4��q"O�tZ��<�\�"�'L$��q"O,4!'��2����G��ĵ�$"OНjUP����ɒ��Ȩ'"O�ҧ��i�~���>N����2"O*��c��3b9١���M�&1I$"O0��S� ���{��J�L����"O4�����<��ٲ�C���!0�"O���Q�I����m�L��UJT"O��HFiY�_$����(��"O^d1�K�	��@����m�l���"O��Y���B�!�5��%��a`"O����D�_Č`VHÈGØ�Q�"O|A���
2�� p����`�F�w"O̩���b���M��8�PE"ON��GD�^b���Â��n	[ "O���烑:`;V�p����or���%"Oq pÏ�&t���fC�y��ɓ"O�e��-�0<sT��doؾ��a�5"O��(�b�!��x���Θ!���xd"O�<Q�� UD���
	�eO�m�7"O�����9{�@1����0`=lU��"OB����1�vu˦��\���P$;�S��y�ήs�8pSf�=n�B)	5����yB�J�9�h�v��c�,|�$F��y���Cr��A��F��@�s�Y.�y�ܙ"� ��6 5U(C�Ɖ��y��8O@�R��T�m0mQ�!H?�y�L�/(�p*3/C��dY�#���y��6N��� ��#Bf��e��y��R(ψU�ϫ"�ji9��	��yB	�"nږ�:E!%z.���0�y�2y��k�"�4f��ĩc���y�ψfM���E�R�+r����
I�y2N؛S�΅�b��N�� j%+��y"��;�`�+�L�Xi�O��O"~��R:Q"��J'/�4R:]ꐀO�<9E��!Jbm�Q���z��y��a�<A$�ݰ �N$`e ��g�@�+l�Z�<9U�@1$^jT��̀�#�E;�lBS�<�D��I7v�i��^	3l�m�6"�P�<��GaH�LI�"_����Xe�<����6�`PP�F	i ը !�^�<i��� J2���2�Tz��$e�Z�<!7��+a�6���ˀ�  � ��^R�<���O<!@�
�*W���(�F�L�<�,u~ի1�D�.�u  NB�<!Q�ڃL�H ��bE�elщ���F�<q�Ó�7�@qKtA�!�	�~�<� �4��L��vI0�B*wf!`'"Or��O���!�S�D�@�t�ѣ�IBX����Z�G�E� �&~WzEq�@1D��H֏X5(�ɕ;5�b*�-D��;ƃL�IFh�I�S�#*L�5D�rB�'9{ �(��]�E^љ�h5D�t��-�s`����@��u3�=D�d���<��$�3C��8�̉�(9D��#1�˶�^@�tAH,B�	��7D���BGI~���GFcRA�V�#D���!M��b7L)�@�b�CN&D�,�7�S^���R�`��2�pva.D�8�G�,s�tH���]�9��Á'2D�d����i֊xI�&O�[N�a�+<�O�O�a{Ƃ
�8��L�\��}��"O4�dmjF@C�K0 �����IS���i\U�m8�� �E��u1�&�@'!��
"Y�}{$�H�Ha�!@
J ��)�'`�t�Q��ޛF;fq��EK�e`��8�'L*Q �������0|�	�'�\ u�K�BJ����F�w�j����Ɋtcd�!p$�=P�|�8�k�>8�B�"��M ����R8�eh4�����=�çK�y�dƻv�4
���ȓjN�q�KN��Ћ0k��&N�y�ȓ'wb)�� _�S��s��Q�@���R���� l�=�2�̇�M�����+��h0#�]	1$�}���al��Fu��b�x�L8�ȓ	zn���M�J���c��q�ꘆȓW}�ē��ȭI<<�Y$� =JQh!F}��S$=�$����oD���d�"O�B�	8DQZ;1l�l=����`��C�ɒr�%j���6C���&iW�~�B䉡U+�9��3heQ���1SJC�I����U�O%=U���O8tVC䉰9)2��E��V������&+�C�	 ���R��@	k����'H;B��*z�b!8��щp���R`ΰ���鉑iT��X5cz��
1��B�I2^I2�óLT0��j���B^C��>)�\y#��]!}jH��+�e��B�I�;ĸպ�b$Db�e '�$����d??�@`ԼN<�w�Ͷ\q"Ar��\t�<�d^7#��U��d])4�h�)3$�J�<!�Ǖ]<,��Vk(:�~9w��I��M����k$LU�k#�R�]�66<�ȓ��e
��iE`	12�(�ȓr�Ψ�a΍8�,�1�]b�"I'��F{��ςX+xH���F<d���1P Ē�yR�� V9�|���'h���rB�M��'a{rQ=4S���F�[��jcJ3�y�H�8g��%r^�2]zSlɗ��ȓ
 <���f��4]�Pa�s�]F��T	H����9J�$@��6!�2C�ɋG�%SbA =]���U"˓�hOQ>m Tl<#۞�j$�C=o����m.��m���'&zJ���ė�J
�ݢa�	&Z ����֤)$��)�n���������Q��1#��Sp���V�$H�"3�Pp��
R�Y��|AΉ�ǔs+h�ȓz<���H3BՈ���qT�)�ȓc� 	B��Er@���+uL�Dx��):Pΐ�qyj���冤N��"�@�D�'��}� �a @�L"f#��ӷj
@�.��E"O��Y�^<<��������2W"O�Q��J��,��0����z�9�"O���&Z1@���bG�ѱ%`x���>O^���д#�`�����[�x��� �!��{�T��6��
*ju1EQ	�!��"}NL�b�X/,|�a�䉎O�!�Dϫ9,���2�#D�N�B�)��	��DK�Nв6�	��~��'��l����B�cCX*��y��'iX�Ǜ�Sr�	+s�B+$��
�'�ݓ��D�t��`2-�9��\��'���g�^�B|�<�1�>�^q[	�'w��5�4zNŘ���.,���'�|�!�C
Ip�����-�>�#�'8����j_�{�TQ�P�ʖ|�X��'X:�2A�^�yÐ�̪q��S�'��P�0�F�*K��a�&N\^H�y�'Ҿ�'AH!( 6�+��Z
�T���'ӌ�@_jf�iA��v��!����z�<A�!@�ֽ���U8t�d��S΄R�<ů�	LT�Sע'4Ā;3`�C�<���^? �n$0�C0R�ܠ�G_|�<���9ʹ�P��/lΞP�rI[w�<�q'��7�z�z���(>Kd]92b�u�<aũC�Gh�.��*Xx�����g�<��זp�"�F��<>5��3��f�<�֮Z�tb���1
��);ab�d�<耢)����.��7`��S�F]�<�#�'RPC���w�p���'�Y�<����������6�H�(@�<!P&�%�}�	�VZ�I	⍕a�<������ۦī6�6Y�D�UY�<�1�$��)h'�p�B�e�@�<I�$��R�U�/��&9A��z�<�+��;����1CB2H�ʹ@���r�<�!��� [A��(1����o�p�<��
.Y"�̡�	�M��@��o�l�<1b凾;*t���Z#�I�F�B�<�"`^���� "�v�� �v�<Q0-C8;�n�9P�(B�JG�h�<�vjteX���σ�=����(g�<��ň�N��q��� "�b���WJ�<�ֱ`�r��D�#�xeI��|�<Y�%Ye_t0e#_^���G�|�<i0lV�d)Z����:�:�G�p�<���*1��� B��:@F�Ԑ7�k�<�S�(e��i���6���S�H�}�<��A�1o��u�L�{O�D�'��]�<�"�߱r��X
ѬO�5%��Yt�[�<�5lF�Fg)���V�܅�RN^�<)�)�7	3�XU�΄>L堅��V�<y��Վ�⹛��I�1��$��iT�<�#Dډ����rmY<g��D���BL�<��'�"���)5H/J���[w��r�<����=A�0I��I�s)J�k��w�<�Al�8"��7�H��B�z�<���ȸ\@X�M͟J�޸JFO�<���,���G�`�*!�fG�<9�A¼p*��Yv��Kw،�t�X�<)0ア
C.ͨ�C�F*a%k�<�$*��'38|)�i�X̐)��B�<a���+c���800�YB�<qF�Ǹr(8Ȋaj\����i~�<� �r���jM�Љ�Q%��{�"OTmk Iv���I�`�7C4��g"O<5�ċ�;J|��d�F�G B.6D����D�7K`�1׎_���=��5D�lx%�+�lqb�[�X�p���f2D���*��=Ω�� F%,�)��*D�8��> u�QÊ��$��Q-)D�@UG�4`'$��b�.���E�9D� s���2RHR����yܠx+�;D�x�������eE��*�D�9��9D� ї��7WlqC�� 1��6D��z�b�)*L�ّY��u9�ƜW�!��]7Z�$���<]�鳷��'|�!���J���VᒽX%\x�#j?!��TP(zĂr�����zmB
�'��{�[�c����b�'
�^e9
�'P8R�-A�+��5i�M���'�h2��6O&�=�G@ȳ �l���'^�Hy L�7$ٴ�hW�Rzz<*�'>��S�Kڜ�R�a����	�6d�'
�q�R,�!K|�qa�6v����'���`�nXK��s0/L e8J�'O4Q�T&$@�H��4�Rf�Ŋ�'&RA$��9>�4L d�@4`����'fn�yq �<�ؼ��m8Z�tD��'K~Y���<� �l_�[�L���'@��goN,U ���ʊ.���'H��E�;A�B��G�S),A�� �'�&����^��٩ǏZD�L�'���x�D)�4�p�H��vt��'3D� C���*Fej1d�e�Z]�	�'�h�R$n��,������޶loT�{�'��z$.1��S�PELЂ�'5�8�(��6c%ҐF$�Ш�'���PW���C�6�qƐ%9"R,��'�X���"��=��*��!��'W���ҫ�^�01�eIR!$��M2�'��(���D��"e�����'C,:���3`V^�b�:8H|�h
�'�F���@�+?�`�t��) W�]�	�'Ux`�����"q�m����'�TҖ�H?"@�R�P�.����'N��cƞ�8�84;�ܵ)]��Q�'{*�����)��#wዪ4��U��'�r@a���/h��Ѫ�`����'����é�|- 8�����`/I��'�`9�ݶi�b�9���!��5��'�t4p�ΨX���[�$wd(�'���7H�Q���(1�W<��!z�'�j1
�+�+�f蒐@�@a�@
�'f�0��#&w��k	N�	��,��'�L {��f�\ڇ��+���	�',��[�k��Mh�,[w�7X.��'��E�B �=��t�U���r�'/jm�PO_fr�(��բR,�a�'@�4��ʯM�8L�����K
���'�����o_*V��h��[�GhY�'���rg�[�t�H�i��_(7��<
�'��TZ�D)7���`-��D��}��'��m둄CTB�0'^�H�6!+�'!�Q��R@�l �nΉIę��'J�i�D,���(p�ɳl ©�	�'Y�}S�b�]̊ p��>X����	�'�>�)a�TgY���n@��	��� &�[�!�@�B	�����Pkq"OX��.Ķ8i ��A�*<X`��"O>E+�l�%t���ï���с�"O$( ���)��Hp�N�C�� �"O�h0F�" 
`r�M޿;vp8À"Oh%YBF�6^�6��3̛�M��(�"OJ��BH�,����DJZ�(���ڂ"O�ps�׋.�t�i���*3$���"O~A�'�
w\B��N�8q6�� "O��2��;
I�U#ծL����"O�a����$�P;с�|��=��"O��x�ڲ��z��*�v�P�"O��r��O�]ӱ������u"O�Lj�M[�Q�xA6��`��)ْ"O�8�	��(���۴R��|Y��"Od��3ؠ"m�����K�K�D$R�"O�ء��Ɍ4
��AL�=v�x�c"O8q`�A�gY�X�O�CJ�a5"O<��p���rZJ0s֌�*ִ�X�"Oj]��
�V8��0��l��IA"O��"�1^Y$c��)`�!#e"Ovm�@
�~Ә�q���gS�g"O�hXCH�*z�V�	3d��7V%PF"O�:�lL�=Da
�)���@�;c"O�,���"t&���ɉ:{���Z�"Ol���� �N/f��fB�tٮ��f"O�Xa,�#���u�>ZeZp[@"OBXoC�^֎�n�	IL���"O<A/�-�\Y�͕�U�@�1"O&�I�� !+���l|��ڀ"O�1LڳfZ�cW�N�3N�$1"O�Űs��9|�Y���H���T��"On0"##�Ҍ���:,����"O�L[E�׀h��a�v22�Fq��"O~���-0���I�h��P3"O�bv�:�6UB�*�e*���B"O(���Bޡ�%C�J��i�"O.atD�}N�0����� ��"O��).���9�n��R|J #�"O�L��m!Ev��B�_�c�U"O�b[���(%�?=��!�p"OP᠆k�,E�,8pA�%�V �%"O��	b�5hi����c��!�DZ�S�eӱ��bD���!�$�ME��b �ʟN�-ِ���F�!򤐹nN:�f��N<�Y��<2�!��ğ.KHA��� ����2'B�@!�d�?FJp,ޡRh�EH�!�!��9QPV���.S>X���']�fY!�8q��Cu%�6*H�q�g��bZ!�D�<@�x�pk��� �p,�(M�!�$݄>"0��Y�vT�8��H�!��\dTY� ���g٢PX䋬$�!�X�|��8��MӲ<^%�ƣS!�!�H�l��L�/K&r_.�A�`D1�!��C,.��
�oI�sT(���:8�!��\�D��:R��g��3�!��>�@��V*�����XEn!��z��|�EՆY b��N�UR!�$I
(����r��h*���⃁�; !�d�<j<����o" <y���#*!�D��!�&a�˗�T<�� ��#B!�	!S`�Õ��;E0~{PLұ?!�$ʹm��M�u@<ҹ9G��e,!�� @IC' ُX�|��#LGd���"O<�w遡:�H��b�<Z��C�"O�e
� �3�9{�B�FS���f*OL��%,�t�6p�L%�&��
�'_�)J�AO�k8�83M�	���'�|�c��A�YiM¦V��%`�'�.�	�`��}:]`Rm���)�'r*���2r����d��xK�'����*]2[�p �F�f���'p�����ο��$�� �(fEb���'����hQ[�ڴ�Ċt��a��'�.�9QH[�6n$)��x���	�'߼�[棇3�
�k2d���^��'�8@a�6�ܱ3�K���1��'.>MS0&V1;��V��}ۢE"�'İ��p̈m�p���"��+	�'���q���F"��T�0Lnʈ	�'�<�Ivo��^Ԋ� w"�<"n�*�'�lRa��څ�(QѬx`�'��(����m�.���<�h<R
�'ў� ���P���%_E�@��'{��y�$�5�xYˇJ^�Qgx�X�'�~`�혍|o�� O�F�d�h
�'�� ��a�4)`���l<Q�}�	�'D�q�%E"�\�	$��$/��(�'$�\�D0��HY'��+���'a�d����6���q�٪w����
�'9�DA��J���5��.sm*��	�'f��!�D�"l��S�G֋n.��')\��p�'Ma��p�hX�s�T@�'U��{�j) ��M� e^�\z�'w��CΖ�5 n+u�ǤR�V�B�'@��Z���&%܉'�HR�u9	�'��P��eQ�g�]�ʊ�@-b�	�'����e�Ͻ&�L� �
�6@�]	�']��� D�8If��R͙�'�J���'|���.@"F���¯{�|
�'՚�C`�
~�f�:�* C�$�S	�'�n-��ɢ?֒ar�ݧ4n]��'�T�Z A�'�T�9V*�K�"OZ��&��2�<9�c^�^��-��"O6���@ͷF9�y	�I҈���A�"O�KF��"%�y����"xa�"OF��`�ٌ`1���NE8~�E�W"O���%�.@��a6mR����1�*O������I0p��eGH z~��x�'��ycǌ��*[H5���5n���X�'���q�CT���f��<y/�j�'4XI�h
��*�Q�Y�e�M9�'����ǂ�vy�d)��K�b|��'��<cB��#t�-:wb��حc�'Nt�@D�A�S���L�Ő%[�'��l��,��Y��kO_�]�p�
�'XV) S]0��!C�Vfɸ�'.�s J,��<ءb�4<�D���'��@xe��M���A8-v.6"O�
c�+��xryD��-�!�D�+���5�I�n��Z��!���Y�L����k~$����~p!�H�4���A�*#aƝ��+�-|!��:��*���@� �	���b!�[_~^��eѫ0��T:�fIyJ!�]JM.��D½/��đ�ɔ4�!��0����Y�k�p�"��!�� X\Q��.KiP�`�_.��m�"O<�Ń�2N�L��FcˑX�Ĵ�@"OD��c��5�nQ±_2s�Ƙ2�"O0��f=K��+��@�H�8��d"O�͝dq��J`&[%z
�y"O$�j#A�i�.@��$�,cd$�1a"O��a�@�'O�d`�3!�1Ĵ�"O�-*����"�h(���2"O� 0FiN�;��h'�Q�q09d"OB1���K�1���0�	4j���"O�P��䋆:�ր�M��XQ��xr"O�D��@�;aXQ��,�<یe+"O��:��
fF���*\�0��x1%"O��1�ˑv�:qz�j�2�� "O� FK�nb���2�>U��"Oȝ��^�w�P��1! 54Q�?�yb � f�V�bvbgZ���߫�y�+*HY��h�}�@�1�k���y��D�<B�5���$B	eӐOR-�y��܎Y^^U�f�� =�P����\(�y2ML�_継0��^�<���S����y�BK��dL���E34"䪦�׿�yBf�V~�:d��!$
�"�yr��Q��iI�+���!�,V��y���*E����c��+�b�*s�@��yB�U+`)J)����/-������!�yr�ȡ����#閺Sh�Q1d� �y7F�m��g�N\fA�Cś��yb&��]��i�uE̖U�lI���;�yB�����}�x���^>!��Q���
��88��X���77!�D��<�|�Gϛ(��1��]!1!�LHUzb��� �J�>s!��ig�d+�ǡh%.��  W�+X!�DL�4�4��;����5mJ!���u0�.e!VD�/E�>7!���;;��*$��0����u�!��&*\z�R�M�	��wĒ,�!��L+�.<����E���{��++~!�D��a�؅� '�'>�:�cr�-b!�S�?�<@(���_�(��R��!�$��%���2EZx�z4 %E�7:�!�D�>d�$��Ɔ�[Ҕ������w�!��\����Tc�$�����`O�w!��+�0�!��H3�֑���C�!�ĄY�b���L�,�x����ɓ�!�D,mj�苕�E�%�t�H�m�<9!���F��2%I�Ow��Вg���!�D����0��3�Dl�F�]t!�*C `$���Ml�051�Dk!�Ĝ�+�`��W-�
^�x8y�ޚ~�!��T/
�596���g�\d0v+ծ2Q!�����ᒪ/�<�F��|[!򄟠%�J��w�ޝ2�F�g�X[!�$�+�2�b�ѕl�L  �7Th!�R�O�)(�/-m�2���(^�!��� 1��p��({W��"fCP<a�!�d��)��9�n���X3t!C= �!�$	0OR�Q�w�N���0��%U�!�DG.$ڄm��H��v`�(@S�S,K:!��/pU̍�f,��u0HH�'Y<\8!�dE�z8&���c�X9Q!��44!��MH :���2'ab�� ��?U!��Y�{8��خo�|�a/�!!�� �!҆��l 
���i�YuZ%��"Ob���`�\��i(ɔ�n6�E"O|�#$�)3�d:��=Z�# "On�fNˢ<#61 B��,`���"O� ��-/;E"�$3m⨙"O�� �@�<��hw$W�6]B�{C"Ol�@ԪAl���c�өNQ �95"O�l	b�R�0��RC-!Qn���"O����V(6�|
#JJ42��"O�&D/s�V�Rǫ�3N��<�F"O���"H/��*E��8|��0�"O	�����.���*�ň�*�"O����[�$����hʹ	
�H3"O�ɘ�!�=:p�=S@H�����!�d�6d�p�B%�Q�Ӑ��%��7�!�V1M���V/N^*�@A��!�D@��rԲ��''���1AeN�#�!�-����k�'vԾ8p!$���!�$
92��� m=+1\��Q�D.z7!�D�1zЈ��1.�����b!��)#!�d �p�r�gӅ,S�X���\�!�$Ж"�q@ݤzDЩ�r;�!��D�5���$�R5޶���gO�O�!�N-R��6�U-!�f5&,�!��A=Ƭ�C�xI�Y �"ZC!�D��4�d�(12̸�b�Z�!�)@pqPeL�"��w*�-~!��&#7^1k5��O��HuiU�$m!��Yhd��d��Z��86#��$X!�ѿ9tQA�F%+�.����Y�<O!�D��n*�P��ޅt�r��/��N!��Uo��S�O0w�� �4)�"k�!��R9jcl�l��� J��F�!��X�wʹ�#JXV����Y�j�!���L�6�B� U6Mvj���ނJ�!�$\�!@5#H�[[�1�Z��!�\=[�@�&ϐ�9Z$@!a!��!�L?�4�R� �l��̞3y!�,g��4��AG�^�nU)��T�T}!�D� ig��6�M��Mq�H̿zw!�D�`
�h�+�7�L�  gض%!��PM��y���F�Jy����E9)�!��+f2Ti��hYF@�c&;!��*�$�Ѯ��B�
9�RL�)h�!�dɆw8*�I�aT#be`U��+�(�!�>DWR9 �(Ӱj~�%K�26Y!���##�\��N�Sh�B��M	5E!���N�s#΋�.�t��HS�!4!�M wob�xU/]�%�J��'��,!�ݼ�`]�b��pk�]��H�
q!��N�_�L|�օ�m ������,he!�$	P`�����h�QXr+#b�!�DB=)�e@Kܖaz��ȧp�!� m��{2-H4{�IS�Nz�!���(7�t%Q��R[O,��%.�{�!�\�V�Z,sf[�9�(X�";l!���8���%��e���\8rY!��;X�*q�	�����D�OK!��/C�y��!d�@��cH(�!�$ڟP|�0H��ur(iA6ʛE�!�d��t��l��J�go����M��p�!��RZ�Ҭ��N]5V���KO��!��^=n}a4H�%
J��)!�[!�� edrYS�R�a� �EIV3?!�� ^`����
9z��
̝��ݺ�"O܄Bp��`J@�ʗ6����v"O���"�{�B�8*M!!j({W"OȰIQ��73'x��aɂ]U��!""O,U�ov)�6�n�6Yّi^��y2�� �lX�R&�(UAȜ��W1�y�LՑ3G��F短5+�(;���yBm��zt����< . �`�Ԙ�y
9*��k�ɘ��f����ٲ�yr��VV8�!��U�Π�PFL��y��F
h�m���K���R�IE��y�)D�a�89�  �03�dj�i��y҆*05
�2�.��4��遲���y �n��0��%��ς��y2/�$��"���,�(d�����y��Hc�2 q1���T!2�MP��y�����J�e	�b9����y�%Z>7Tz�����Eu��8����y�N�3��a�ˉp�n ��@0�Py��Vv
�$��
܋��,sU��M�<y
Y�jʊY�%Z��`�U��b�<I'X�15� ˇ)P��!Y�Ha�<i���>`�2����E^.q�6MY[�<Ӡa��]�����.�#d��S�<	g��LF<#1�؇�Z����K�<�MP
D������%sB0"���G�<eX.r)��0�\�1)&�B�<��.�\�����Ɉ�&�����A�<�vn�)X�����>|m&��v�<�H^���Ћ�-�|��!��[�<9�g��Xl��C��.��E;`[�<�
Z4b �p1q�CC�T��`Nn�<�B��^�:�t	�6�F�\d�<�G#�ft8q�|�xX�&�u�<��g�!{�ZӠ6Z�Y� eU�<�L��Er��dN��R�;�v�<A�I������P�T/̤s�e�p�<M�C����c�&<�i�u�[S�<q��Ϝ|�!�#-�$�`���R�<��EW��\ase+��-��Gc�<1�.�����̗)$9�]�b�^�<���#w/θ(� �<<|�� ��<�`knOj��`����m��/|�<�"DY�=5v<�@�_P��eO{�<�T�j�B�	!ݎd=���NIm�<Q�i��Z�����eB�&
r�8c#�f�<閁U4��8���Ӡ6
h� Me�<YV���D!|���$MN�	kTU^�<�Wj[)���`���LM�2��@f�<B̚�;���A�F^�B����`�<�2I�@���!*��A����F�<����>���h�b�SRZ|ѵ-D�<!�^�<�}�gk�Wv&Ue�W{�<iF��. T�AG[�8))rd[N�<��ŋV��(
r)��0��!����L�<A�q��˅��X�`�@�lO�<!5/�2E�]����8�\�ʕc�S�<�d�P��DX L@�:�h�r�g�i�<�CJ�:\z�$�wl�9�F��iFf�<�F�I�)a�����mW^Y�"�|�<9C�?cW0=�i�<H�%�c	d�<�v�ZoV�h{���e:�s!�x�<	ӄW�=�����gQZ$���\o�<�	K�,� Dc��Z��˷�a�<� B9���>/�Ԝ�"&M�g��-ȕ"Ob�Aq�P%{EJ��eN?C��A�d"O0��<B�p R��P�:V"O�9�
�gʝ	V���,v"OX*�OF+V���C'�z��"O�b7�W|�֔�'p����"O8�ASn�;�i�A��N(<g"O���fH7��	�&R�S'Tm�Q"OF�F��.J0J�)���~Ը�"O|����!"���( P=�Q�'"O�H�F�H8Js�d��/&ؼ�A"O�-j�*�v��-ڄ)ʸ	�`"O��IŅ��x4�QRB/�'�aC4"O���aB�2?����b���ex�@@6"ON�񁒻rfu��+F�#ybx	�"O|�jE�D�%�J�'���rJ@4"O*)i��p��M,#K��"OPg!�>&x�I�ܹH0���T"O��d�ۛp'���UkS 0���g"O������
��T��O���"O�X����(nq�qb�:$1�sc"O���)}&͓��N �U1C"OD��gM�>��h'�R��v1��"O��#ƊB-{�!���\��xw"O:@s!�`6��ۦ�[���"O��ʖ�]�L����G��K���"O��1��	&���8���m��"OVZaJ���B�PQ�%� �� "O����T�m� s�!/�X<�%"O^��K�)������R�0yA"Ol���.F,M���y�� }϶\�"O���,?!�Ĝ�'���S��ɰF"OfQXg��5�]!���sYj�H"O��:1��-qD���F�ÂtA�L�"O�a��E@~tZ��R=F<>|q"Oa��X��aB��5d�T5��"Ob)��f�, � �h$ɝ@,�5�C"O�M��nIN�ڕGS.2s�e�g"Or��&���}�T"R'�$c���"O��[c�)d�����s�t�kj�<���t��e���6l���ۃnA�<a�ҙI�Jp*�@�4���#S��|�<�H����D��-�P�5s%�z�<A䨄�}f��x��58�1�!�k�<A�@Y9�XY뵅լ?~��:� �R�<􌐁xQv݀s.@"7����1πO�<�Ŏ=%��MR�C�/.$����c�<� ��h1��)�*��J� #�b�<��e�V4ʡ���/�xuce�S�<!��_0uS.TC��ȋ'�. rȖN�<�ROKj�0��A��Ⱥa�FI�<�ë�/!M����o���v����
a�<�G�7���E� ^�0����QZ�<�3,T'c��
EI]���a����V�<�ꐬo�f@x��X��DI6CUP�<�&4*�e��@� ���f��B�<�$�ɰ8.�u�@+,P�"�JuJ�{�<� O��"�윻�%Ϫ�^}"�r�<��&ޅ>��BV�k��5��El�<��EN���=��cٔJ���aaN�s�<�7�ȊAB��j��z�.١�h�e�<у�*`ڷ  �2O�k��k�<ɀh[�b�dÀn��J���� Gj�<i�� #���f���A�a2UJWd�<� �Y�6L� I��X��],mz��b"O&��U!ߢn��a��Ϩ:�Ȼ�"OHq�!��P����P?h�`�"O@�*�:1!�p�c���n�p2�"O8���98���o�
�Z�"O#�܏i�^�I�,k��|��"OBa�@�7!�$���@z��`D"O�̂=xX�`+Q1W�ĉU"Or�7h֌;�4d◩
^E(m�U"Op�B=H剓hS !�8(ф"O��v�ʵ!t���'��%_�t��"Oh��g�� wܸ�E�]P��"O�I0�M�	K]���KE���"O0�d#bl"5[�GG66ı�"Of����\|$��E`.f �"O���A �>�pL�4d��3
E+C"O� C%`W�:`L�y6�F���I"ODU`�)<���)�ӽ��H��"O�$�'�k�Ĩ�]���A"O��`G��i�r�m��o�b��Q"O�X;d-Y0h�+��!���
U"O䌃�'����j��kkv��"O��2҈B�yH��$�:7Q8@pV"O�F%M�x��"�Î
lX]�"Ov :�#q�}�@�K"\�>�3�"OBt�T6�Kש�<%�< �'"O
�1D�
<ـ�IK�H���"O0L�� ͣ?S0��F*ͻ}�(h�D"O�pïP�AaR 31`�n��'"O�ݳ͑�w��B�,��Ȇ�J"O �i�����@�]8\4*u"O>i5b\�g��qEI2XVfPW"O�<rDD�E��5���$hF���"O�s*��z��!��Q�gpB)�G"OrH���#1X�`0fT<9b��A"O��Fߑ_��a�e��?K8̳U"OI���x�`P�E"R�Z�"O<Y��,݄g=�]���T`<���"O��� N����Ά�Smޱ�a"O� �2�K�0��,�d.A-'>��"O��cc�<%1���m�Bdi�"O���vBJ�P��E��H��"O�����TC�ͩwK<�\�"OR@0�ˇU�^�*��93~���"O9�@j� JּH�'�1Xn^ո�"O @�``ԧR<�9�)G.Xm¥��"O��_�v�1��oM`epR"O>�0���'Cg����i'J�P8e"O�8�F$�8o���#' ���"OL�ɠFF�.���гcFI��;�"O��C�'?�,�Q��4x>��w"On92�I�uJ(���krr�@"OƁɗ�R8H�0Je��>&E^IP"O�p�Sg@_��ʗѿGR��@"O����`N�+���,�� F���"O��� ф_"�]�pJH�xu:a"O��:�h��Z�H����Jg�TЂ"O�q���K�ܓq��9�>Ay�"O�)QF�_4NH� �#̸��"Oh�8�"��}eh@���ɸ^�^Dk�"O�$k��M5,�:�#H����"O��ȥ@K�ooܙVI�.N�&0�"O�x	��M{O�a����u "OF ���V��T�fF\-��ɻ�"O� �{ Ό�,�kP�Q�v(\y��"O�y8��kYJ��r)H�<ɓ"O�	$������"(R�N����!"O�]��a� GXTs��
#J�|a�#"OP:��O��*8�5@ɏ�B�#�"O�YC�B��E#�0�f�D!N�^ic"OM���1� �ThU�d��]��"O:!��a��<8�S�^�>�"a�A"OF���l��,@4l#�+�"f&��@"O���'�ԾO �rs�
�Ěp��"O@�4DU7Xv�Z�f8Q]�0"O� @mZ�6%��S�W�<�\8��"O��B��;%� �0̙9e��0�Q"O>�`+��O������v��1"ON���o��>�y쎮\j�t��"O<�A�͐xr~�C�A>7��=`�"O<4��ݡ�vE�%���sX���"OF�"�/���(D͉>R�s"OԘ�у݅Fr	���<KAj��R"O�����L-S�i��z�*�8�"O�ABa��V�����B�b�PlQ""O|�Js�I�NS��Y�gT'Q�F�"O\�ڶɎ�I�i�A��3A��d
�"O�p���$�43��H��]��"Ol4�7"�4]�J]��;1o���"OX�)G�@�tr����G� MEH�"O���G�"I���ATf߆�����"Ove��AR�t��*�F�q�"OT]�so���NyS)/C�zm�G"O��4�Y|V|9���Fn���"O��ɒ�(<ّܸw��hQ�B�"O�x�S�,���S�$I`ZX|�T"OHDq/)<tB@�õ1`t:"Ol�)��fԦ|��I�C�0��"O����ݑW��a�0hԄy"O� +��Һ�3��E�A��V"O��r���%XP����Q$5�^e�d"O|�fL�F��|2�&��2���" "O,æ��:@�PtN�u���"O<��h�2K���TeI�u����"O\d�a�)�6I��� JB�k2"O> �(i\|(���m:�Ѐc"O:��FAKHx�㠄��\5��I�"O�S���jm��D&kX!�C"ON!����ZT"�8IF"O�K�+H☝�"a�-yv��B"OH��Ǘ1L ��%��{���"O��)��Q6k5����-(`�)$"O�p0�g
�/�����QbUr1"OJ��c�Z7da���cD�
lHH�"O,���۫	f�A��M$l����"O��J�HԮz] ,8'���7�r�"O����n�G�*��������҇"O �q�
H7�����.�3{��!�"O�M���	��p젱��3g���"O��zOذ&��\�􆞚^c,2"ON�j��/<��%KՅU�
a�@k�"Oht
AƖ�e}<)��D@8c����"Oظ��&��;1����gǸY�!"O��ӡ@�{$�59 \<H`"Oc�ȗT0Y!�jL�ē�"O����@A7�~(�eZ�*���A"OЈ�"S�5%h�hc.���ؠ�"O
�;2��)�RE(Ѭ1-�*г"O� Ltʓǁ�9�c�*)Z�"O���.	�?����j�3�X�"Ob�i��ֹ}%�HBƨ�����"O􈋓)�����G''m᠉��"O�����bWT��fz�*�"Oi��^<>;��i3#�6r���"O��C���x�Ѱ��E�4���Y�"O�U��nA�����['G Lՠ�"O200b�	3ڔ8��L�<"��4T"O��`����
BZ���R	_�j���"O��C�lH�M;��Č�5�dea�"O\�
b���z��U��n@\dA"O�8�U�^ >��9	bbJM\h��"O�T�4�-��8�#��P�d�٦"O2\K�� ��@��E�q�R|ؒ"O�M�v��=�Q�*�{�ԍ�"OH��`	�������@��!H�"Of�Y���H��$���ʝ��"OD�Ѓ\�.k(e�堐 �f\��"O��� 	Ȋ�5���{O�
�"O���ӕH���:V3�Ȳ�"O����f�W����EC2T$v1;"O��	w
������%IUY�"O 9r���J\��%�8#����"Od�K��ʶN�<�Za�S��0ջ�"O��ؤ�� <��IgDU|ۇ"OfȰ#�+PB`��mH��ʤ�P"O�ӂ��/c�B�Vγn�����"Oz]�3կu���I��B9Vh�p1"OЄ��eר{���B�
�=JN~88�"Oj�h�����iKw)��c1 ���"O&$
$�.Qꄝx�(��q�.d��"O����Y����Y!��y�̬��"O�%r���!=���	�vaH#"O�TA�MG9L\B��D���ZB���$"O,YE #b��*J�K7�A��"O�l�0Ɠ1-�:x�tH��2�8)�"O����阠k�V�)�͞K
� �"O�ى�̎�u�pU� �� �"O(�#�(ĵ'�\��?O�	�"OV��c�ܰe#���GOn��9�"O,��A�J;�ju����]�W"OΑ"0	���T2(W����f"O$ �wg�r��Ű(^$8Z5٦"O��A�K�&h�:WƏ�"RU"U"OP�T��:����U� �T�V�ˁ"O�D�+��[E�� �G�9����"O��J�L�>�v0a�-"����"O��c�O0h�`�إ!�BЬ�'"O  (���3�dE��A^�BDdX�"OL��w�ݚ/J!�# #T���"OnP����,)'���)K(;��"ORy��f\a�(�9�'I��e�D"O:TH�m�UC�t�w���4�@"O Mq��P�u�,EY�$]�
��Rt"O��J��N'	n� ��W�R]b�"O.pZ���
X谐�� {ި�P�"O���6�T�x��)@�ڵN�<SB"O�A���X�8k�Y�]��L"O�e(V�#Pxt����n���A�"O> aï�E'��9�D�n�I@�"O84�Ռ%G���1G�E<����"O,���G6���w���fV 5y"O��I�͜xI0tQ�FC����"O� ��U�F"/�n%��RUB��g"O�@`��8[
����ل0�%ʴ"OT|��蓟3�� �H@4}�PH��"O�$�t�ҵ^aZk�A��g�H�!�"O��ƋH- 'l����S~�hY�"O4E����'X�<� �X�P�`Q3�"O0`!��+[�"H�T���J��6"O�$�3쎰[v�ۗA
�K�XJ1"O�"�Gܯ4nJq؃�Ν^_����"O�m���6*d���h�&N�ƨ��"O��!#ǊUg�r#�D*Q�J �"O��r��Ll�����[ wVu�"OH�bc�	q(<�ǕP�A"O��X$���/w�x����%�"O���ޙ;�N@RG�@4K��]y�"OL�PSDL9�ڔa1��+��A��"O��CPL�!+L�:`��y�&T*�"O��cƪf�ع۳� #��{�"ObpSC�� O���I��Z+����"O�4aq��4
vHY��f�MM!�d��+ߊE��Ɋ%@Jp�$��;!�dX:lΥ�a+	 7DXڐ�Q�*!򤜓R�,�ӣM1)(.Y9U#@*�!�dҵ0���p*^E��C��!�$M7/#�q�Cr���1T]�!�D%[0Ax���(!�Mò�K�!��4>^���#X�%��s��l�!� <�$Ah3�ǌ-�.��dӘ'�!�Y�D֎9*gB��bT�dW�!��v�h;�iI����S���XB!�����E2�D?G��1��/@� .!򄆢$i��̀[���9լ<?�!�h�1�UF0P��a� �!�d[)X�P$�����!���ՃJj!�d�$q!� 0�,q�H�?f�!����Tpz�,������3`}!�@�dX��3�W� ��8�`)o!�J�3OH5�g��g}�Aj�o��f!򤌍3�YX��ޭu���C�(hL!��D*j1.a`�勂)����H PJ!�d�C.�����C�@=��E�c3!��@2}��1�5�ݥ �Q��Z
!�d���%��h
�H
�+Sj��t�!�	HE𔨟�	��6)���!�P�p�D@pe[G� }`#cS��!�@ ���X�#I�m�Gk�!�0)�#4 ��W��PBj\�8'!��ŽT�rtK�*8��Ԃ�w�!�z/����U82��*��Ո�!��&���r��B�@���aT5!�d�Kn����ݤ:�(�� 
VF!�DH%�
��/Mf�v�B�ʷ>6!�N�7��}��R;y A���œ>,!�䃛�ʵ+t��:\�HH��C��-*!�$@3UBr\8�&g��ԏ�6r !�$%��T !�û���@�/ӷ(6!�D��~�z� `)��]�U��DZ,(0!�d��%�����k��m�(�Ӂ��?3!��83���g��r|YBʟ�!��"EF��KD�L�l�/A+_K!��_/B.蔥�;�
)�EM6[.!�P#�R���m��L���p���9F!�$ d�����W¼
Wk��*�!�$�IjeF�)�����[�j�!�� M���ҏx{����m�li�!"O,\��34zׇ �.�L��"O ���-��%�����2h �"O�!�dʞ�qUn��E�ٔ�B�"�"O��'@{{ � �(I�}�Z��c"O�;��B�Y���A%�j�)S"O���`�Q��BhhB,�qZpS�"O ��WLG,A(���`,74h�C'"O�1P�-ٹg\�$p�dGP �!�"O�D�#<&�*�P�#^�MD�S'"O�@5)�{���	��Ԭ��� "Oz�SvF4ME��zW��) f���"OTh���y=d9����*��C"OLU#$��s���x�K�9��v"O��"l��t8���KW�Nʐ�a"O�L�v�+S��` ��͙Z�A"O�`�H�7�����M��,Sb"Oj�;��J25�Lb#�ӣk�N��c"O^��5�N'�� ������"O�$����?�R�{��wlj-�T"O�[4D�m+����=AQ|�X�"O�AYa[D\",�#`^�ID�C"O��
T�*���Q,�-�#"O���ցn���Q"��}�t ��"O���s`�>ޑh����}�6��"O� ���=D8j��.��p�b"OL�!�����ܹd�=�(�1"OhK���1������2Y)!"On�d`���rU��k,Tn躆"O@�WA1y�8���}d��"OJ�`7�)X
��i��~(�Z�"O� K�,̶9����f�[
Ց'"O�$��\�0��u���,9?�ٓf"O� ����/'����ac�I� ���"OND�t��|���RŢ��fh�9�"O�I�j��v}�rִWq�+D"Oe��a	�w��'JP�>^���r"OH��	�h���bbcA�h�T�"O�����]M˜�S�A^6A�6%��"O2��ѫU/"�Fh;���gD<:�"O���C�C��ZhBe��&G_�)��"O<i���Y8nAmڕ`��U�\<�s"OX��TD�}��/��`�� "O��JD�K�q�|
���J��@�"O�(��E42ۚ��P'%N��v"O�D�����ylȜ;���,C�`(�"OH�)�gɿ+��5��Au��v"OLd�������R,|i���Q"OD!���<1i�Y	�f}|	�"OrE���/<hHQr��>}��"O �3�!�~���{�-ͨ����"O���W�`�$�(��T�+�4��p"O2�0$g�%Q�~�S��:9��`cs"O���r(T�X�8-�$C4+ȐZ�"O��R�'�As6�6�f��P"O�%���H�.�����V��`"O�9���R���'aY$d��)h�"Ob�2B�.g��,�U�ڳ:��Q�'"O:��2�P�
�"Nٴ��"O��hVA�e���C�^	]q��x�"Opźa��=f��s�J�o~�Q"O��F��r ڌg��*:Q�=�U"OT�ۄw�T��#��B�U�h3D��"i����9����`����	5D�� �yCL�"ve:��ٱ�&�f"OP܀tↂh�ݨR�H�v��l�V"Ol8��3W�5�CJC#=٤Ps"O�B��0C6��9&��&�p��t"OD!i`�M�oGr9��_�DTޔ��"O�hj��
{"��B��>9RR�"O2���a�%d"�M���-3� "O&�`�.������ k�s?�1#�"O�@j1 �
i �2��T���"O�d��h�)C�	ҢK�
�=*�"Ot�@p�F>\;>p�F:8��"O�$K�	I'\�}� 5W����U"Ovu�I�&��`�g�{lP��"O$X��؂<HrPYv)[$_:�"O|�B Z�T����%
~֥f"O6�D�\+o������zx��"O�諰kH bm�v�]4Ti�6"OT�)p�ߧn�dU1s-�3]��ZB"O,�s)�n��IԬT�+�"O@�C��?nߠq��� Ȋ}"O��u��I8ysw)�Z
L��"O��SU��23�j|�fY=�رJv"O��- 9r���V�i����q"O����}ʀ���!��c�"OА:A�߉e�h It��88"O�)�UG��$�A���P��,�2"O�PB  �#lz�y�Fۤ>�R]ʗ"O���7���:��MiæK�9�,��T"O k��.��e���Z"O�U��i�7�$x�6�c��ܢ�"O��Ѷ �zTeu��:\ꚥ
e"O@D��L-N�!ʀ��H6�ii�"O`����*�iS�`H9�q÷"O֕JW.�:'�^���ߦfeT|�"O�dxw�͹U:`-*��#b�s "O(��.͈5�SĬ�*��	q�"O��BKU�hҀDئ�۠���@�"Oք"`��c���Ak̆n�� v"O"P�2c
�@�䡹
	H���"O(+d�'�]�"�]�A�H@�v"O2t	0�̚jB=�`��T��d`�"OJ�g���i�v��ĥ3S�ƐZQ"Opm�犩{�NśTO�c�d��"Ol�S7��11L�qƮ� %S����"OD���7�䰁�$�9e`��R"O�H�T��5x�V$^#1 �f�'h\0����X"�q	��ߎ5c�iX��y@���>Q��C�F�'.�S��/'n��%ȷ4
j<�	�'D$Q�gj�`�h�� W]��"��$�O��������jJ�pBT��%��yᤋ8S�џ������k��D��14��A�̓E�B�		Wt��RϏ�5�=��I@7���Mˏ2C{�$Vt�k�kN�J8�|�� ��X�BɅȓfڼB�	O:�P�AF%B#���$��@��$5��"Ck2 ����0^����
��2�hC�I���|2sG��=V�p��P�)���'��$��(O�-�OLA�eL�Yl.�P��9q����������~���"Ȋ�M���!X�!���j�
��5Uf�`��6]�!�D�/B�.%��/D�	aE�����!��~��8G�V�}KpH�F����qO���D�&1��� I�:!��=!���b�!�D
�}:�D22$r�hgo�X��kT�$D�H+�e� pJ1��G $2p�[�`(,OF�<� Kօ�P�<4j��Wc��M�$��k�����茓=����Ҭ�)el`���͝��d(�S�O�B5�J; ����V�H��;
�'s
� �G�x�F��	��h�	�'�N|��B��xw5�E�KR���9�'�X�Yq�T&������4F��p�}�)�IT�W=F��@�4u�ЍS��HZ�}����*t���J���D�
JR	h��<��p<�V�X됨rF_$&����q�Iv�<�U՘t���i#ކH�%�fO;D��
�ED}��-���\� z��BC�7lOv�ti1�2����rj�>q'��j��'D�P�&ԑ<�@EǊ�Z����w'GO���|�O�����/S�S��r��.u

=j	�'�|	0�Z�o�<�2��!z��%�H��'�0E���Q'r-L�Y�Mܱ�,���և�y�ʕ�ޖ9�d�x�i�VFō+���$0��<��　fc�Go@�{W�}�qB�V�<�f�G>�@��0��H��1*`�RR�<1qB;fV%Ք̪���VK�<��)?<�"�3�Q�i�~e���DD�<��<_�Xĉ��,Y�S��Y?������h�^`B�N?*D�v��,I�ܸ�T"O�5#�8F�p<�4閵B�<��"O|���&U�꘣hV:D{bH3�'��O��D�I�)%u�Q��L�y�ѪC��"!��R�а�GA+MtB1C�	�b�!򤓭LIL �a�U��Z��)Q'�!�v�,�;m�H]�Ta�H[>`1O.�=�|���O2��z���b5��9��y�<��й�P ����]@��{�<y1���t�賂F�%����f��w��hO�O��y8tKDN0��Q� ���AU"O\-[� �0Q�􄂒`��<�0��IR�O�1�˟9�L�P�OƊq�f �'�zՀ�#�@"���Y�d}!I�����0|Z�'̽h�Jɰ�,G�4�ƀ�U�' ��|��I�_4q-{g�C�D�2�!����Oh�kӅ��^��%��R�0�R�	O���)�f��m./�ᩢ'�b��K��0?!׋U�:WI���<а�DhRJ�<�i^-�B@ W�</���@"HH<��Y5�D��v���.��Ѫ���g���X����\�p1S�,H�H1���7Y�C�Is!�5襌B2rcv0¶&�5IX�B�IG^��c�D��-�D�`������2�S�O��������r�!��>�{uS���	�|��R�];0@��Q�C0t��>�94ȕ���-�
lb�nB�G�@i��K�R2FEx����rI�4JJ���4.�q����2��$92��G��">�I#!^��0<�����	E?��T�cl% ��D��%'
	"�|��p?��?ez
1^�(\��4h]m8�@%�d8f@I%��@����#�D��5�>$�PR�l�C�,�#B�Q�m;|i�͞�yR�&"�<���IB�4`�"��̰<Y��D[Ar�@PVa�rz �W��[qO��=%?�� �8�(�1��n��S�*D��8��ҝ�>Q��Nm�,�9&�'�d7�Ol����"7���WD�� ������Or�=�~R�'��x(b�Ŧq��1��1i�N-��'�X���]�p��� +���ɯO��sO���'�Z�R� ��(2�5�v�_�uV�����>D��с/��_6�������<}�0�z�7-+}R�'���3� &��0Fؑq�`PQ�mډ1�^��"O^�6[�&a}��~���3�i��	�<�g!��LG}�h��,�aq���E�%�t(��p>��q��I�pŉ�Ě�E��M�u�V�87m�O
t�W�4)��`�G��Xa�	��ȓ(�.�ȡ%��NlU���͍ab����9�t9�A�s�N(�%�	�X��`%����	)�b��/�nE�C���������'�����[Xі��dKV���aR	�'ц)��,�1���iD+�o��@�oXa�e}�|ʟ���BŦQk��GZs��x��K.n�az��Hq?9(OLQ�a���7�@�1��\d��#"O���Ĉ˱X��㤅P�� CW"O\��� ZU"	�ЦˍM�L���EtH<!�͗
���R���d  �Q	
`�'a�$�{��mȊ`w�3H��d-�On��%:B[�H�kd������؟���	V�ɏ4�剩GEδ���[hnB�c
08
�B�	�	;"D����:x��Fl�Y�V���'mў֝�_~ ఏ��p8����'G<�����)�4�L�iACA�aJ�y��'W���D�g�'h���P&s�"�(�`
�@Er͑��3��O
�g����W�Kfnq�,[�F_z�'�T��I#N$�� �׀d� �׍*4j�dY��p>�'i�Y��
+t~訲h�7U�2������W�dU�샺2��%�ٵ{�O��=L��J��qV��vhE�2���"�b2�hO�9
;dH��c�'w�2dC� �����ɓj$�8i�aֆr����&Q�B��lq�6�׷#��u��3~
rB�q,�=4���6�ia$��Q�<��ҡO<����N��hIv,GY�<16){��������6�,FE�P�<I��7摩��E%H���c6E�C�<Q�(U4Eh�ȷ��~AN���ǀ��iF{���i����S̖�p.h-�P��5v��
�'������8d�5b��.y��i�
�'^+U��"N0��;�B� p���
�'L�Z��Ҩk�l!�稔�ot��c
�'O�����"`��h*DÜ#>��	�'�����d��t��O�M^��	�'�<�GF�@]�l��� {y�=��'P,T��#=T�|�pn�@HZ�h�'��(�4�	4;�z��wM�"��H��'XJaЅH^�0��9ⱁ�?E�I��'f��(գ�,u���Nø;�L�'w^�
2���5	�/�v�2�'l��r�D<[
V� ���|Gؼ��'�Ji2@˄�`��3�����1�y��֨|n$�ɰ��+"|����yN��~��(���t�d`��5�yR`G��BՈ؝C^ZuzJ:�y��K$���XR��)C��[aiǚ�y"O�F�.����
a8��P��y���*P��a���,
�v�@��y���/�P ��Z�Z���:%g��y2�Ş�L�Y�
R�v�0��Ӝ�y��� I8)MΏD�u�֭���y��>fC��R'
�JT��!���yR�\�.w��H]�A4`a�$�y�)��~�pK�I�6<e`q`�?�y"
�)~#>�4��]E �q�	�yBc�?�@YJ�!܎jT�|� �ɐ�y�jst�`�d$�S2�� ��7�y
� dU�#�M>|��K1*��G�vñ"O���r�Ьwf	s�(Q~E���"Ox��O��Eb�P[�Je&�K�"Ob�����%�`���k91��LH"O�A�d[�j�fc&��Y�n\��"O☫�#�e���S�d�]!�"OR�{���uD�%S�D���"��!"O�D󓠈�p�|j3C�h����b�'o ��Qb�7Bnd@���[��T�'	Qip��(Z�K
��
�'�I4+I�e�;R�_$GŌ({
�'��+�A��=Pa��-Ïmf�	�'�4�V��#XL�G�@����	�'�x0a� :z�xg�֠T� PA	�'ߢ�c�o�E�b(鶃��C�~��	�'��	��B+�4y�iAjg(M�'��4X5��{m�E�e/�g��p�'�R�s2��i�D���JAT'��8�'�zɰ���0�@�$iRJ�N�i	�'�&Ժ�f�Һ%BJ��N(�ݰ�'�l�%D�
+7 �F��H�:���'P�J!��Iw��%ƃ)V?���	�'$����e����g�MC��
�'Z
U��AT]1���ؾOA�	�'Ѷ�2��F�\�0q� �;b¤z	�'����tAw*X���ի9�0��'T�$9��E�j�HDI�56��
�'
�Pk��[>] =���,�4<��')���C��u�����t���'~����&ڼ)�J�m�n��P��'8��K�'a��\*S� ^m:,9�'��4�����G�����`ٿ]Vza�
�'OR�x4�m�*8�� H#��!�'B�i��WSm�rdE��K���'�(z�)WNFM�[�
g(X��'�R͒'o� �t���Ҳd	C	�':�xg��d�Nu�r��
|�����'�<I8�#B�e{�@���·�h��'�����K�	�l,1�O^����
�'�e�t��/5�f\c���QN�2�'׮�����u��H_��~��
�'8T�h��<s���s�ċ���A�'�3!"����{��ׁ�d��	�'��a�a�kR"�(�L�vy��'�()�W�D�4��1�O5pw� ��?b��cM<?!0�/d������̶h�����x�<Bń5G&��v���>��(s�dN̓?�4K��V�蟀�Ɖ 7ZP��I���{G"O��ʤ#4&�������q p��@O�I=�I�O4T��G �3}���ڈ�qB)�6�l�Ka$��x�a��l�lq��Y&[���0c�e�ȑ�v�ׄOk�i���0�9x2�B/w��%�&�e�#h9<O"�*�iݐm�L���O�0{$ �i%0PXB-ï:�F,�F"O���ƆG�*S�����
&�Ȁ�W�xR���C�Y�ϕ��~eJ�{�1��(�EȈAw<�c��� (��"O� ��M'OD���E�2��5JdG��N��<�Y���!A|q�J�Qd^��Ӏ��+�s��I,e����,�`�3	Y��˰o �w%lm�
�*jv��0�[����a�l��'��&�P5����'-;. 2�$�o:<Ї������@HY����VJ���6�E8���S��Ȫ[" ÔΎ�hDR��$�"3=�ٸDc��kIR�17�O/��6Ҝ� ���X6�K�'�fD*�͉J��,?��)ڝH�xt��g@?q�"B�ii��g�>�Y�!Z�;��exԠ��Kz���A��c�]�Aq����^�(A�%,|w�0���"!(ԑ�m ���r��/Bcjm�4�[7	��R��?'��r��W4J��=��4�)	�S�? @-y�fӱ�:�%�TH�H8U�'�NP�w�|\53Q���P!�1:����T�	�W�`�Ơ7D�|��-;l��Cq�X� \v���8�Ć�b������1�蟶z��AI��ꇧl�tZ7"O����� �lR�	>9c�sq-�}��'b�cQ��>���Q���FK���qs%�j�<�M�&meꨙ����6�Ad�<�� 5T�!'�����I��h�<m�L�L�,u�c"(����+�R�<y��+%�B�O��T�%�"�ȓG%�}qC�sa�
��5V#p���9�DjU�x��'-�|��Ň�}�B��G�.XȤ2��M
@<�ȓJ�.�2o�r3DusN]�h�n���P�"pC_�A[�l3A��s%�&���F� 5�qO�����LN5"m��!�F۰O��!��"OD!���"�tU�%837�u
����	0qdh�� j4�3�	?3��D1c6zn�y��)=Lz�����2��(`�C؎02����JƯҒ�aȃt9���8�O�:q�a�n�u0E�#��OL	�&w<���I�O�S  �ĸ�`MTT�x� ��C�ɑq�B0�EK�K��<Cf��*z9��[��@ʵ�0o�X��nH8���j��S��C|`Ъ���&�8!v"O|}�A�V9U�n	#��L��	���cb�C���0sn�耱�"���*V���{�yr���(��E�"K�[Qt���p?q��R>϶�Z���-5��!@��<@Մ�Rs%��s���� �R�+n���Xc>]jB�%�� f�P�x
jȫ��7�W#N��bM�f���g >9�~瓸X欭����N[`��#[�X��M��*� �<D���&?�((D�P��Ѱ�͙0{긍B�K���.dfx�&�Y�s�R�]X	+�	��aHP�x���fuDAr��1By�B�L�SIq�q�]q�*X��X#�)�+y	��!Ї�r��M���ȴq����G@H�?UY�jY��P3)�)���J1�\(��ݎ*}�-�1)�5�H��DͯP�P<"kL���4A�^2q����^�U��عЪ�P3���'��]��Qz�˭���a�O̧pX���k߹T����lR%.��F}�e�:-��+�!�Z�(I�M�|�g T5V�f\1� �	�R���xLMKEIf�(��aI"3�*%?㞄��&��cH�J�-���>!�-HF�2`��A�dUJyӍ�IJ)m�J�I,\O����qɘ{	H���E
�a��M�D,�5�|�.��hF̰Є�#��y��P�z%��Fd�, r��M���'jLԈ�d'��a�(Q�<� F	:#�8A��I�%�< �P ���?���pL`R"�*�䰴a�1#=�� C�"!dƍ��l�I�	rQ�8z9���!Y���;c������D�,�$!�I�4N����*
�H!I?*���y�,*&E�� �DÖaP�4� ��^� �`Z7�q��'](K`�B�,�z�!M�""b�H�'�����U�oZ�O�>����V�I���{��SUCY�zu�@@X>��|�M��2�Ե�G�!M�|������	A�zɪ�� ��I�:�.Ů;#���$f�� �$S5KU�`��I�ņ����x9ΰq#[�$�. ��*R:u����T` �^�l�p�>�|�։�P���S7��@C���L�'�Bm[��:p�4I�|�!�ܦa*%7��� �OX�\�y�M:}R*߱�����e@��� RN6^8�'���3���I���X�Q��>{.�S�O�B1��١�����L2B�%�j��	�qi;�O0)�#�=H^���,�%o��)���>��c�9H��	{ M#�$G�r���.Opi3�Bʝ`��q�gI���=j��'L��6.������Ԣ� -K5тiN�.���
ON�Ѣ�A͘�QFg�?Vv�x��	�~=s��)��(ir�Z���d��d��O�!�$Ԃ��`��\�W��d Þ=�F%���W��'��>�I6�E�2)B�H�KCxC䉺�
�CD�T����oX7�֡|�B���a����=���ݱ����`�;-�~� ��g��0���K'9�K�	��)"bZ�ob���أ�������<q�/�>a�z��K>E�ħ��cҺ}�R�O�f��IYp ����'��4x �;w����S>��3���
#�؀�O�;��]�D7x�%>c�pKeE�{L�8Bv��6c�Z��䦊�RZ���g$�"����(�"����U��� �s�)�<�9���m������J14��e��II��J��ơ@��z�˓�O�j��� ]��v J�D����D�w�^�!h�>��O�.��D�� �����S�.>�(	ד=*6	�T#�4D@�ܴw�0�c��.:d��U	܄�=!~�A3HѮ0��\�.O�>s0�;"JٲB�2\D��?�,�f%�f/�]Y�E�ċ�U�B�H"�B%3��[�`H�Ͱ<� )�# �Nx2
=���'��e!�54��E�\0��I��r�˓s�b��&��m$>�3fc� 3B(����B���U 4s�9g ���ɩ�pb"��fQ�T	��N�a��6��CK���
��� ���ScX P��n��ߥ{
����&���P`�':��-���@p5O�!/�29�~��Vl�(4����T�O��ɖ�E6dg\�Yį�<�'ޞ�I��1�J	{�F�ڣ��,M��`��(^]��0��Ǌ�+!"q+�$�>kz��&i�&��q��r��ᇉk��}� �[;�"�?Y�ɍ/Pt(]q�[ 2$�ye	�k�'���Z�g�<)��BU�X�J�/g����K4s�
�ct"2�`F@N|���t�����
��Q]�!�\a2���q�����m�O�� �AO�J����SUp�2�K�2bvj���E�ΒOh�а�����>I��!*p Xd���R�7w��Ӵ����$��e���yR��4`+�	�d�5��ũ��tsa�ޛ���z�ic���=5	(Q�~&�����¼-�a��M�9^�u���O(��p���j��u W8��� �'Ǵ%��K��x<�0���DQ��L�
����蓡�:3Jt
H����`�1��lx�j�<G�<�	�5���Csa�)n��q��1�jX�\�ZdIT��0H�Y�?F�1��5���1 ��h$�0닌1[
y��dD�U�p@��x�/	��^��⥌M�O�9�R�M$��`Y2+ǩz\��E!��.��9���'��)�g?�Pȁ<H�5�Q�=I�F����I�,W̟,����]��u�ޗiϲL��E�?4f����-^R�a�V��~R��S�E�m	�9�l��V��ED���p�Q�g�i��6��2@�C/�A��m:"���#pӯA�-7FaqI���p<	��̽ ��� �E�<	��	�����gD��-�v�f%t�'W6U3B�������,F�Txp��B
�H$zѕ%>��8�D�jkJ,��ʔ˘�%4�2D.G�H"q��m�3�$V���(�>E��4%PY��KX7:p�� �Ge%�0�5���F���L<�G!�D�4�"�d�?@�n�Ȣ��e}�IW%D�*'�VX�D:4�N� �.; -9���B�:d��Nx�()A%�*@�>`p�ь�9#��L��7�H��X$ˇ�T'�`Q�ݨ�g��j�R�a�˅�	�h)G|lJ���(G�t��3�]cg@�#yt��g"Y%�y��C�t*z�ڕO��w�<���mV/�y��V�*q��ϔb��`a��y���	���yq���,�"�k��\��y2H�j
Hz����~���kb/թ�PybaM�$��Y 	ˎO~��H��o�<ٲ+���&����Ԟg̎�xB�Jd�<����A�b�j +�v�ԡ5%�`�<QD��*5(y0GHL�s�b�v�<�Cꋺ���
Vlܮ_���)�Cq�<i�NN�+� ���&�@I�P�<�T�J���!�,�����E�Z�<�׎8R��Ma��R�k�U�<ف͚/Sw�xq4�)�b1��A_�<	���'m�Ń5�N"����&�Z�<�2��(����`�-��*�#W�<�vE��uҙ`!J���&�d�<��lסeX"��k4���.OZ�<!�E�A�X�Ó��0K�N����L�<A�/R9OgꄸF��,	[BE��bHJ�<9@��0�����eX�
k����YF�<�PG�'�z�����!�v�C�z�<�E�K�W���VL�	#�N�U�Tt�<I(S#=������Ά5�tM"�,�i�<ys�J~�g�� YJ�(�ED�<�ҧhc�Bb+��q�|̹���<�scѦoc�����"��͢PM�v�<� 6�C�ND?L@J{�oI������"Ou)��ׇt�AXd�� �>l�u"O��*b	�6j�n��,�Yc"O�m7�H�_z8����8ߖ��"O4�aS��&��D��ڡ<Ȯts�"ORe�0�ɃGH�����		WLt"O45#�e�Sl~����M�d��"OL�@a��1y���b��+����"OV���� ��c��ww���"O�|���}�>4�t���(��\�"OV��7+��AP�pǕ�{v渉�"O�K��af�� %8TA�C�"O>Lr2�ݠ5���*%��/n�ȩI�"O|�Äi˿�|i�P �5>&d�Af"O���ӂ~朰�E�_�Gx�g"OCC,�#D�� �+Fc��k�"OЬ�e%�$\xd�����.�j�)�"O81A�a@G���0U��(s����"O��zQNߪR.t1 �E������"O6�R�gS�]Īp�dڹ��]
�"O���C�u��aA6�qb�"O��9l�@%z9��� .@��rD"OD�I��-pBpx�͟�r��h�"O. ����R��r�"> '��`w"OB�Bb[$Z����� E����	b"O@�X�H�(9�}�� U�@�v�xW"Ot=:$�S�)>��8nŘK�<�R"O�iR��M�,��f��4~�rb"O
� �Ǜ�np��i�v�Mk%"O@ [#�tj ;2�K:4
-RC"O�L	V���N�Z���HΛ1؄xa"O���m�@���Eے��貀"Ota��g�)f@�Q�bΕWѰT{�"O�A�\$�6T�!קz�^��@"O@�C�%p)���ŀ�"��y�"O�9s�nI�},p����O�) �R!"O�ep��@!��r2iѲ��J�"O.�����y�T`K��G�h�"�	"O�@����DDR���"�8���"Oj�x@�ˑ<�����<�(s"Oᇢ�U ��y�ΏF���"O���" Y-"'�����.A^�YC"O�hc�W�r�i2��M�,i�"O�1ʔ�@�n{�q3@I&o�5Y'"Of=ҒNF5Sp�2�_�^JX� "O�)�2'ރ`y�e���,h)����"Ote� 唙A����A�Z/�{�"OD�����9���7�b.�G$_W���w`Z
 �	�ȴ�'m�.L�X���TdB��Wz�ب�l:O��rm�8.\b��Zr��-V�E��gS-#	�	�b�Z*����ݼ�yr�� �hQ@d˘ �nIZ#�J����P/}��B?���DƑR��̇c��q��U+̾�ƓSܠ ΚuƤ|� j82\�#��̈7*��	,*�O��#�@'(�2ق��( o���'�<����I�d�''u2���;UI��!�N�0\���'6��ꃵV)aW/:5 L<Y�N�2PX�(F]�Ocz��h��/��`�[ #	���'גD��kX.3R���F�mQ ��m����˓��Yѐ+6�3�$�&SN@hJM�1;�μb$kg�q
O0�B�c]R�1sȪt��z�̵9gdave��02����^D�v ҥ�<w�ec��**��xr ��[�ĝ;T�ȝ��	�C����#� Eٌ݈AL� ��C�� F1 t(��'`�	ʕ��f���'M�tCT��>�Bi��3� ����ߪ8[�c6�_�+��=b�"OhDk%�eژ��a� :#"Li�G�SVhI�'>���%Tm�g�I6z~�d��HJ��� E`�C�==l (Y$��\�x`�4���J<:�!e
�@h>�e�vX�h�����:�4q�gċm"J��"5O���^�,i�� �>)���hU2�3Ή�\Yj�en�_�<	��U /\�6� 	�Ĝ�4�T��!A*���� )��?m+҈\�jA#al��B�e/ZC�	�s�:e�jJ�-?��p�"�9*�3��"��?�'1�AK� .���D'����'����5�Q�h�P��Q�SZV���'�v1�&��3�l��)�Bx5�
�'td�5Hһ �>�I���C�}�	�'K�(J�/[�I��3��0PV��'��0QF�\]�<�1�����'Yf��F�-Q���;W����H@�'�6e
�V��
L�CEuhD��'i�a��ٱx,�����!jNB=i�'c�m��>JȎAJ��f����'M�-0\5x"���W+fk�)�R�+D���t�j8�8�7�"zAf$D�#�j��:����΢E@9�� D������2
��L�(�*m�� D�X@E�L'YqM�c�ʊ\ޢ��;|O����m�*��$͢;8t��ϰ3�u�Q�hk!�$��W�u��ˏ�U���B$D/R�O�)�+��*�\�~�D��5
g�D�����~l��J�<y�╨>� I�F ��O˜Pq����-P��cO�d�Dϓ��$O�k6|�<A�̖@���AW��j�F516�[k�<ᥥ۟4����Q�N�0XjwF^X��	CN����@�%�����|���#(^ؑ�&f�$�(q8�|qgj�B����#r��ɡ�s�׮�N���vc��O�"�Eõ.�̒�qODMR��ʵe���G�1k�޽���$��/Z�a��Q�*J���?M1UI���F��M��t���탸W��a9�i��[�ab��&EbP)R��O[i[�G1 �4-��F��?���7v{*	;�''@lxI� LL\ys�W�0y'�A8I����5�աv��8@����u��kgc�a�X1��.�-�@A��R�s<�qP��^�^��HյK�"�)��O��ZW�%� ^����-A�h�tHE�u눢?�S�*I@����ܥ+�O�� -� v�n�"�f�Y渹`�@	�׶�lH�����gܓq���H�o�Y��Ѐb�W( cp��'�l%�㋆Z�����ܧ��؝�D��g�R�x@�'yК�Gi5��(�.��R�d�'�'FnZ�hY�*��Ty�#��8�Mh6�F�D���I�&��1�(��?)R�l��e~����Ν@�6��"nd̙Q��
BJrp�"��f�v1���.g�ĸc�JVd�%��!Զw�� d@��S��P~�4���B���43u�ʗ�~���S� �P���	v@��0�^iQ��yQ�˄Z�=�0GTn�S��,�0��C�� �cό�T�`�S���ɀyb�PW��|r�B=h��S6n�%P��3S(���~�.�u�:��b���퓨.�|�S9�( ��gt$��˄fW$����'$�1)W��H���ϙ2��1�N�$R'o�0hp�K��`������r?	U�*Zt���#ؾ)fV`Y5n�J���s�bU�z.�i�I�7�,9i㌣P^,�$��$��IE��pZ�I�&1J�S�'|&�0$	I��d!�Ҍ��D}�� Oʡ����V̧Ur~ԛ�ԗu�x@�$.
�,�`U�<+N�'>L`���z ��莍�f�K����C���`l]762�@
ǟ>E���\a�0�KBO�6��HI'��(G\�M0����&�F��� 6KPm����))���t,Ц"��QX0k�	�!OG&O��p�Ɠ0��d��6�Ti�J\�.䜴'k��o�a�Mэ&fx���i�>Q��_%t��I#@��h��4w���y��J�p�P�Ye�џؚ��M=����IҬ&>� ��O;c��\ "Oʍ;��T�}�U�bB[�D^�-�P�\�kNm��|B�d��c� 1��!S�O�8�c$<D����ҶG �yP2Ð��u�A�p��U�����O�h
�E�iHSd�H#Reѳ�8� �뉈U\�0ز���Il:� 2��-V .�4�sږ	z��TX�X &LiY* $��|r���H�ʣ�ȆL�Hܣ�m�e�Y ����8��hP��iF�n�<��(�c�[�L�$�d�'�(��N�/L2��O�HX({v𶏆 �(��銇�:����WAy�� g�O�d�R��!�d��7I���F����]�f�YA�
~�aR�#N�ȽSF�Նk�j�1�C���$��	8c�FE�f�<yӨ�%q�K���x�=pAq��(pY\�Bi� nx���D�T��p���}�:6��J+H�s+�W�k#�C����X�.�"�%ٙ��S�O��*��3-�:y�W�H(&Q��{�
�%�<�C�� ��>���CYxx�ԁݥBM��P�	�����u�	���#��3�I�_N����Фv�EB	.gV}đ=\�E"(O�=p�򩙂T�f	)4iN����K&�I�2��`�/�0��,Q��=�O���ϊo��	�%^0٬��v�i���q�풷]���'�$��CZ'j�T�7���s ��)gmV*Iiz@A�E�.��=���e_��
�'L�p��	-%��&W%^�j)�'�L|�3�&��FS��}��e��so�+����>@�6�D�<��BP-'Q�U!B��".%
�̓�yEݥ ��
A#B�4a؎��E&7��d�LZT��&k�a|��Z�6�bH��b�V���T�
o���å(yL�D���0<q�U8y,�'�,�[�&s (�F��#�̵`�bDָ+�E�͵�(�`\a�o��i����D��b����|��`��	���OK~��C�t~`�֝R���x�$�: �q������!�g?��I:[���k�
��
�!�$*Ɛ��M�@�E������-��Y�m�s�Ф�]7V%�	|�<Q���N��MxǓoPP1ˤ�@���m�fj�\|Rm[���IpT��9�R&^̂c�Z���U�CA�(2m�pq�@��V�2�A�@H�x�e��BY�p�MBy�Ś/y�t�0*V�I���z��W���'��:��6Y�25�p!4���q��d��&pl��A�u�^e%���'GX�Sh����*f�����O/6 �ŧ��^��"!G_��]��b}��Hr��m+�3I^��&(!�c��$��1�OYh���g�g�I�V�h�B䂍�x�r&�C�2��6(B �H�
�/b4��Ʉ!�@"Pa
$+����F�J��	ad� ��\���I*�;�d�2��8���3u��G�<%iص��JMO8���������I�^�P��*Gr�;2�ރ�ƨKT�+�DG�LS3)	�/@x��� �*9�ژ�G��H��%A��Xf�	!z���"
@�N��?ӥ�L��L�3�(옸�!�rӐ��u��r�n`M�"~nZ63!���� $s2Ur�;>yCZ{�Č�>x`�~&���"�3<5�X�1HD�rעx��˴>�1gBB%���6�;,O�q�V+� O����k�� �Fh�7o��- ��<<O�(���6m��I�.L&�ԝY�� 8Ċ� 1LO�$Ar�����;�r�Hch�=Q����ŋF��">qA'�k�|�*�2R���`eX�;������U�<����F%���oG�]�*8�!�D�<��l	M��H+�	͞����k�<i���(/.�s��<�H��Ig�<��BPy��![�ЕJ����fi�<y�oH�1�vX��%���t��NM�<٤���0���9�nH��%XC��l�<Q�/����x�O".X���J@�<i��W80���"���[��]W�<� G����14�G����N�<a`�ʀq�,# fn��k���s�<Q�nP�f,l��&��Z^��ch�D�<�	LU<�K�� 5�
ik1f�~�<!��+K�C�ڞ@�VE�P��@�<A��:,���gɈ�E5�t۔�L~�<�w�2m�0(�"�s��d`0�v�<ar� 8�<��V#�<5�p���e�<��\�&p\�!��&q�rMB�Au�<�կ�ly��K�[�42EI�<�4GL�[\��W(�<�r�"D�$���I ������X���+R'!D��BE#
�Uj@2��Ch� j�f%D���g,	�z�x�� V'����t�%D�� A�! ��$Qo��`$��X"O6�ȧM�i�ܙ��%ӟ ��8�"O
�	�0L�>��7d|H�5"OP�Y��2E�t�#GBQ�@�b�P�"OTxAu^>t����ôH���8�"O�a@�O3F@�)�樚6vf\�C"O�� �j���d�f
��7"O<y ʃZ�X�DE�J7H�"O�x��Sn	����"��a"O�h��M��R��vEV%2*�axb"O:p +ΎT�����Ҥl
N��0"O欩�C.nE���W�^S�p�1"O�,�A�\�ws�ẓ"�I_N�	u"O6d�����Jpx�p�Z�>��l<D��UK�
#[����$Eq���1D�* �_c$ �P/b�|�g=LO��h�2U���`N�~�i�N�%KF��$�]FP�<Qg�ڦ^��!P�DԈI��S�?��,e����>4P(-hA���ElfEÊ���l>�K��ղd�d�u�� M��o2�	�����=��ߟ�I� PlH;�Ý���T ����O�A�H�DE�T�N�BL���a�����1�~:��my��,O��W'�+~�~1�@�6OĴ1D�
zt��Fz�SЦ��u�ۨn�&/@�ؚl����[f�Or7�)��	�$�V�H��ϸS��6�_ǉ'�`�U�'ɧ�O��ٛ3 �G�>��灑�10nm�M>����	˴Z,�=�F��-���"
ͥY��	�Y_�|S�}��:_���R��RE��%�"�o�/��Q���j�)��B�*��ΫgHذr���zHD�T-2��OJ@��SD�<�0%��L�>�p#LH��*�H��|2l-�(����	Ԫ�J6'�<%3�C�B�}�'Kd�S���H�S�'6�t�� I]�:¶(ńjx=�DT���$OI6E(�O"#<�A��ug�ɉ! J Q���C՟lE{���*:�L�R-��T�`F��7��O>��k?���J\�?�('�K�S����4���t+1N!��[�'������r�>:d�ݚ����__��'�|����I�� �I��?P�h�f߶�	�0|�#iƺK�%�� �
������G0?�d��<���p>[wgΒ��9Y5&в�_�H�1O$Ժ�''H�a����|�,xr�Ƙz �����K��=��w4����V?��𩐥�u���w�:`X�댬h���c�ʅh��ap�C��̂���<'�X���O�xز�d�(�XAG��%�.�iĭǭ+H������t��S��?!%gS�E�Le�UgO59 ��O a�<���W?�5{��J�C�����_�<C�āC�`�cbJ�V���/X�t��n{,K"�p�������#"3�	�ȓ{>���f�#��,:g��)��Մ�b�|����� �C`�m�݇��HT�!IH�5����dN
"Adj؇ȓA%��)���=,�3u��K$��JO�!y�$	
H������<���%��p�7!� @��F3$�9��n�*��F���JX�Q��T����*P%��
#�^�:�1�ȓ3���T�+�R��ƪ�+wSvx��%�l���͋I 1�� }�L�ȓ'�"���dݮk�4��3̜\��Uٺe���A�Z�J�bO\�|���:}��1 b����:1��"⢘�ȓ7-z�9�iχ,��9�t	� \���Ě��G�Q=.+�;�J��Pt��9m&0���:3���:�E-�ȓ%��e��M�j�H}��OJ ^t�l�ȓO�!�盵Ie��J�%�7@���[
M�ç޶M�����ϫD�h���S�? �UI�A�/r�.�c�		?�j�Bw"O^�L:U�%�VH�-N��
"O�`Ռn�����ӼNg�0"O�Is%R:b�~M� nŻ�E�g"O,���+tN<�E�C�*�@��S"O�yw��7^��� H6��� �"On��f���&�ybo	��L�s"OB�*���0���^l3�)�0"O(��fN>)���0�g�z�HP�"O��7MC ?]"��B.j�"Oh8��`F'{��xQ�>>
h	#c"O�ū *s���"2�&�����"Od�+�F]:i�޹�a�φv����T"O����� �hdad�+&R8Y�"O8ld�#�k1)\���)T"O4 Ȣ�GXX �kG�Q��h��"O���@�I=$�ޤ��/��M�R��"Oʕ����b|aW�ϓW�"O�U��U�x�l��%S�R�,�r�"ORx��γ	�u���M�F�)�@"O��q�YH����u��!r�Ιi"Oʙ���<i�.)�� 0���"O��X���b[�""BU�p��T"OX1QR�ٽ
� +�O>k�ʨ"O|���O��:G@|1/"O�X�R"O����c�;W�z�HP
ȎJB"O��q*�� K�L�l^�<8p"On�� 'I(91�=���2w�����"O�+�bS�VrĠD"u֕�f"O�E
u�٘w_\P�T��xj�QU"O�!�W�4a4m�UoB#�zD1�"OLhq���1S��{�m�+OZ�Q"O
��ŉ�%/���a�.2,K��"OLE������Q�N�&]i���3"O��d��k�Z�H�MC>L�l{�"O��SFO�d�pdM��
��0*e"O��Cb*� ���ҫ�gm0(c�"O�YIU��d(�`�
�,5OXy�"Of��D.�>UL��̗S(��;s"O�%P8
��� ����|g"OX�ʢ�	V͞|�%��S#����"O�9a�̮m9t�	��D�J@ٲ�"Ol(&�[*<a�8�R�lZR���"OP�����ż��&ÝYQv��"Ot�В�N:�|\���C�@Q�=�1"O|�)7�Y	o���D�/'�<�c"O�@�/�x�L��'b
%���"O")
ǂG�a��혳�c�����"O�`:��Ѥl�Y
c.�Y���8�"OD��X'Pp�Q��G(|�~� R"O^� �*ݢث�R"7��=S"O8H���<XR�m��OӠ�4y"O�Q��͊�T�R!�)�"�I "O��3��I�_!�����64�\T!"O&���+��&��1�L'{���2"O�*6�	�J�r�8Í�$Ds�0a"O���N58��8�S�^oZ���"O�`�G���bU"`c�9UB�q��"O��*ы�Y ��0`��;^�5"O:�㠃(BzxrF��G)�8��"O-"�o?r��3��J�4K�"O�C��
�X�sҮ] B��9�"OTU� /ә7#t=A��P��b"O���Ǐ>,z�q�R��:9d:�a�"O� ���͢}�EӷѷꌤqC"O"Q�G��,XqCcMM�	�P��"O�ػK�=:���rk� F�ܡ"O��P����(�H��#��f,��"OlI�$h�9`dԩ��X3U��=8f"O���!Ďo�$hJ��܋F�*��"O��֠A�$��K��V�P���Zu"O����G��;�@���hU9a�`Ud"O�4)4�L!Pq�fH+bv�H&"O��c�IG7#���#�ۑܑ"O<�cCQ?G�da� ��\W~ū"Of%"�-HgL�h��<OWz D"O�-*�� ]蕀a�Pi�p�#"O�qx2ɜ;@gzI����h�~ȁc"O�0�`ȋ V?,	0!,���j�"O�{eC�8y̸�
;F�(`��"O����ȍ��t�!6d�Z��q!"OX��c�K	0f����,I��K`"O�}�k�#��T `h�V�$<˷"O� hboٷp���PP[�4��|�"O!Z6O�J��d[��J�i��U�""O,�C�z<���%cߚ|�"O��JBdcBe��(E� ���"Ot�q�69'�ݡ�������"O�����O��<��X�����'�t�!�R,l ���M��@Vp��'�Z�[�m��3T6�vLC�<`"1��'��L�A
S�M��1�v�F#^��
�'��i�F�5#���hC��	E���k
�'�������,=
h�K�4+��t�	�'�\��ĕG�R��A�Q�Y���	�'�x���c�rd (A��.T#�	��'�<����Y��(�Z�����'��X��g�01����5��0Y'f��'�`d	ģv����A(H^Y�
�'g
E-Ƚ:̣���?�� 
�'O�� 7�L9B�,��S Z� h���'#$ım�+.��0�Ӆ�?m#�Ջ�'���3��
8�0	8��f��t��'M�	��� Rbia����-|��'?~) Af�5PpD��@�ݫ<-����'Xz|
3�Ȉ.`����,x��a�'�i9��ɐ,T�9rE��m�de��'3&��%�=JQdl�&�F�` \LA	�'��	�1��I���2v�Wh����'R���Q��/���r��Ls�:�'+�`�eѴ�0��F�C���y�'rP�s���s��=(��M(]>���'��� �e�ext���A�oI
�'�(�Q��:s� �p�I�-g�X�	�'�� #��1TB$�.��dO����'LSaH^�A{�u�4lRR�� ��':��:�|DʐÈ�X�$	�ȓ<Ƕ�z���@<�d���&|�bi��r�di�I
�a�R%ȤO�'�8e�ȓ*L���ΐ3 h(�F�� р���?L�I!f60���0aZ�J���ȓ ��i%�_sĢab��79�9����	����A�UF���j�:����h��D�V�[���M
�ـ1�ȓ	�v{<��%I�3l���J��yRMJE`j��"m�-�@43R��'�y⯗�.�왋��,+:z��R�
��y2���?���cF�q1���֮�	�y
� >Y���׭7���h�K
?dϮ��"O&��)�
��H0k	�sw"O�	��Q�zZ���D'w���9�"OF$B��	r�<|�Z�4���K7"O�����!G�*H�Ջ]C���3"O�IcÇdA2���c,��Q"O�Mq��Q�X]� ��5EV��"O�d2DOR�GB~�q��q��DX"O�p㖃Tr��+��I?`���
"OL��aŸY�^�N2s���1b"O�!��_�}b��֌ͥ�|Y�"O�H��C
{�v���K�m+�L"O�A����&��`u���U0V"O�-AX�oD�� &D<PB���y���$���P�lؘ�^%�v��?�y"-�\�m�֦�4:��h�!Z�y�A�T��eэ�	d�
�m�yb��Wfvl���ڵږlhӠ܄�y�E�5cd��ˍ���bS���y��W��7Kч
=5"&E��y�i~Lhz��l7��� �yB�Zi�9�3IZ��&ؠ�&B��y"��b�fi�QKN���6����y��]�I���:�dY�	�Di���yrk#<dp���B�z��ēbOJ �yr���"s�U8s�ɻy��]�%bW�y� C��ĉ(ׅ�$m� 8��B�2�y�CԌK2p�qb��`�6d�� "�y�Ida����k��1R�H�0I(�Z�'����@J�D�������
��R�'�l��Bc��i��Ti5�!
=V5��'�֩g 3"rԽ�程$b��Q�'��4S�hW/5��|����"�zA��'E0}����C �a���&	C��a
�'tf-k��ٹVf+/.�"�C4D�t��Gٸ9R	zr���1D������c�
�x~�`�'J
C��Aʜi����!�@�Y��_�AC�	�D@�{m��<���Β�r6�B�S�@��҂Y�T;,��O�Y��B�ɉh�d��`�ͳrQ(y������vB�	 [u�m+�F�ak�`p]�2��"O<�q���ߢ�CG�'+�i�5"O������w5�Ϛ(6'�Iі"O�0��+c�́1�˯W��a0g"O�|�   ��   ?    �  Z   #+  6  �@  �I  ~U  [^  �d  k  Qq  �w  �}  �  \�  ��  �  %�  f�  ��  �  0�  t�  ��  t�  "�  {�  ��  ��  ��  ��  ��  �  = � � �  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��'rLa1����%�H����U�ZnL1O@�=�|jE�L(��Y� �<<H��Q�<��@�-Jn �u�J�BB.��r�J�<�R�K�{Q�Y"�[8r_^I[�GG�<����WݾX��E�/q���"�G�<���ҠJ	\8��İ~��X�JJ��1O��g�	~8d�`�Ԃ[`lA���v� B䉌6�j�Y��M�Y�xx!���#`�'��	E�)�'V@�!!���|<(�?T�}z
�'��e��^p�V����@O�
��H<	
���`ìT�W���C��P�B��ȓ2�NM��@��;Y�4��e� D��!g$��i�P!D���x�T�e�2D��
ƠJ�D!�&(I���qxa�0�O�\|򉹕H	�2B��� �H*�ڌ��0�g?iGf�(V�*hp�h]�D����*�C�<���̔mBT)�c#� Y2�4��@�<�h�8�|�����n����� ��hO�nχ�~�f�� �IS�LS��sa�	��y�"Ԧ-,j���!:�:ĩ�ٌ�y�>���"~*�MղQ��� ���i�젊�(WO�<�Rʘ+]��ś&�Y"�I�5�G�<�vi6?�ӓ�� ���2>#���3d�g^����	$m�N}�n�7g[��&�Ϙ(KL���A� �~r�'�z�9���XT`JCe��n�~��H<�Ó��$	�U�%&ۏV�eQ�P�a"�O��kw��*dq��J@�+u�ʼK��	w>}��;V�]X��_�W����!O��=!��M�*�B�F��~�.AK���X�<����a�V�rx�׬ �<щ�ԟ���=� ���u�]\V�,ڃK�9}�9��TC�,�t�5�ߤg�n�"��ݶL@�e�O|7��HO���?i��Ϻq  ᗢ��,j����u<I�(�p�Af�Q�1^6�FCP*����R�'��*7�Z5U�
���Nu,��	�'0B�K͚�4n�-���8t�
0��}B<O"�}�&��bzA�a
�"eD��ȓ�0���.G�4�
p$��04��z`O�5�7�J�J���-��\N����'���<)`N���^(� ��/[�20���	x�<�h	����A*9x��4%J��hO�O�(��
C�n�H�L
V ���'M�����a��S�,�8	���#���4O=	���b�E�&D\���D{"O�nÀ!B5o��u2 ��3-�*�]�H0�O,���2Xo��K#�D���q"O�d����$S#
��L�=Q̚໵"O��� �D������Է+f�� "ObiT��^��Tz��O��A"Of)�񭛔r\X�dљ�I�p�	V8�$[�B�X;X���CG�n�t�`$$�8����cg���wJ���Ȑb���M��'�aKj��O���G�� %Z�'�L<�q�A�]m��x���=�b�'G���2�	}��<�&lՓS����'J����0uO�鑦
�l� i��'*T�un��)�jP�P�]�Dy�'��a��"��B��R.�,Y�m�yr��
�&0H��5����E7�y��0^JL��D*'�� 9����y(�/V�Q$Ƅ��k.�y��S�F�,h�vX?�|�ᡊ��y"b�:j�Υ� `�_�ɫ��U��yr�_+�$D9�"W�^2:��Pb�y�`Ni��mQe�?O)���Lޠ�yr��!toF��D�RW���Z
�y�, �S�O$����ᝯ�^R�N!�&���'Y�Y`"���DA�].���'FrU[E\K	�p���
c�4O>��1}��)8= H�R�њI�W�0=I��n@>ip���Eş4	�V(��G�-�O��Gzʟ֐�DJJ�0��0 r�Z�L񖝈E�>�S�'D�vP�DܪC̦�SQ�1�i��E�>���.t9˧ g�%�p�<Is%��,��r�;`(� wh�ly2�%�O�� ���iq�D2���&� ԩ�<�����t_�@�D.�#5��q �K">���U�1D���5�(y��!�%�$ϲ1�Jo�����&i��4bfKO�;�tD���WR#?����t>}@�E�7l��)��P�&n-Sn*D���7�=R�̉AT�N�]\�Ek��#4��w���|Y�y�� �Q���r2�z�<���߭iI�VM�rB�iB���<���'�ax��>	Ҏ�-Y�Bb��]>թ�i��&�h8�cޛ%�L�2�G�MBb��G%6�IE��l"�d-k�e0�C�L^!ٷ�9D�l��(<#����'B�]2���k�X�=E�ܴ�i vlǓ;o�$��N�;�~l��f���p��5 ��,k��Ք}�F ��p?i"%�.^���� �.(S�M���	C��r��R ��!;'^Aq5CJ6-�U��b�\�`��0���?H Z��1�,�:D�Ȥn��!��0|�c��VƮ�@#�)Q�t���Z؞�=�*��3o�h��ƣ\�H�&��M�<� $�20�YL:ђ���<�p���'��d3�I2P�>�Sc�Bd�*�l�B�	��$Ÿ��4��q��3��������yb��]��]�XD��*JM��t�Ӡ��=�����d��#EB�@��K��*��!�^�	w!�Ă/�R��A�I-0T(6
��%i��OV�"~rf.��A�̘�4�׾{��lxt��yr["-(��J%c5u}p� ��P���'�4�D,�S�4�R�-L���1�S_*����Č���?Y4�f�H��ϕ�$�f��j����&�x�W��$��g}��D�]z��Ɵ�>����p����x���? @Ƙ��π$bd�1Dnɺ#��D0�O:4ô���b�օ����
C��"OR�:gA^�@����I��h�z�"O��['M�'rĀ;�J{��A��"O z�)Ր	M*���I@�1$�8W"Oީk79jK�E��A(w(��3"OLѢ��uDQ�wG_�>��#��'��D�|W���3�.sjfe3�@Q�!�ğ7 �*�����2�`Yc[�/qO�'m?�C�i҇1�a��-ԈH���L/D���7*��{��q�g�D���Ԫ:D��� %W�'ּ�SvF_J�^4(c�7D�0I`돛.[��0veˣ>S\�1��)��;�"5qO2YZ��%�,����$A(�#P"O,5�3�&����!�ضf�����(�Ş"�`A*t뼉��k�"N�E��P=(�KF�n�v��gG��dD{2�'�T@���9b�ơ�!ǉ!#!Yj�yb�)擬qօ��I/ �F<,J  I�B�	�R�@�(��.a�Z��aj<|��B�ɐ[^�颠�F�B��dG�@zB�ɟ`$����>��#(�ritB�I�g�d=VO��f	x����4QJbB�əa�,����Q�L��քB>TB��%c�~�(@h�?Q���$��,�NB�J�-zE���ȋsg�{�nB�	=q��Y� .���4
p�ƌ?'$C�+Xꑠ��.Z�J��C��	p�C�	1?�%��)Z\؉�:!C�	�%��C"˸�B0HfÃ��B䉧fy`bhZ8=M�˷h�9a�C�I :���N3#}��D$S��lB�	�\)()"Ƌfo왱p��_��B��2y����e�Ѻu��Y�R
]�l��B�I"n�B��J{�08�'$2^tB�	�C����d�' �2�����(B�	�_,b�ҋ��%K�Y���_�yFC��4RYVH���1w��Dϝ�g�\C䉈 ��`��S;�ƍ!G(8m�B䉻m�L� �-J5�������S�B�I�a8d�K��k���Q���y]�B��?j���v*;Z;ت� K#I��B�	r�pՉ�O�18��iS%
(��C��/�y�3J��#��{��B�ɫb�1�&eӫHUd�e	Q=�B�	�1u���/9F����mivB�2|�^���
!2�[��rb�B��%��:6��T�*�ӄ��K��C�I8��иa�G�-�� @@
ڼj�VC�:��\	�&H5����$�7"C�	v�v3��Nfг�o
�[C�IMD�(�t"��,�`|���Ȧ�B�IP� q%��;�fP⬌�)o�B�)� z�h��¸`/��3w*�)G����"O���!k�� �T 2
�H�"OΜ{C�ڂc��QKvdEP����v"O�1
V��1m���Z�K�Z��S"O�Ge�J�*���&��]���'R��'{B�'��'���'�B�'��4Ğ�`�BV#�$�R3�'y��'���'=��'2��'��' �!I��K,GG���]Kb� ��'h��'=��'X��'A�'n��'���D���BU���H7�A��'d"�'a�'5r�'��'?��'z%uB
�R�q1$�u(LJ��'E2�'U�'K��'�r�'?��'�ك�g�LE�F���0k�J�O���O^���O&�D�O�$�O��D�O졻��Y?;d�9�-�AĲ���m�O��D�O����O���O����O����OL�YѮB�6�Y�,\go�Z+�O����O���O�$�O��$�O����O��iE�/�l�"�`��5�D����O����O���Op��OH�d�O~���O��a� ?!-�9��*R���j�O>��O\���OX�D�O��d�O��$�O"l����i;�$GcM���1�ON�d�O��O�D�O����O��D�ORU���R���@��ʊ
�0�8���O���O����O����O���O$���O]b7Lϛ+,����ƃ#��!�!��O
���O����Of��Oj�$�æa�I��c���=n(Bw�H#-���	'
\���$�O��S�g~�f�R��섏tz�2(٢-B�l{$S�2��	�M+�����|Γ,������h��d�2p�,��戟w�J7M�OZ��Ń�V�	0{��@����.�8�����t#�Q�1BCA�P��<�����D,�'l�d����,.��bK�><qu�Ӳi�^��y��)�¦�s��m���;G0BM��(�
Zz�:ߴM���?Ot�ŞiFP�3U[�T��F��r�C���TTj�@i��!�%! ,I��Oe���D�'����%nS1j�z0��tr���'��Ip�	)�M�׋�`�C"
��@X$*��V�C�|8��Ż>� �i�"6�x�p�'�}*'\�*P����|n���O�T���y$�ЃA�>�'=\`�g��R�DI_�5��HN�cH�'��5��ʓ���O?�ɲi)��l�8Z����9���)�M�F��t~"u�N��S6X�!���q��D�2��(�	�Mc#�i�m�77VbO\|$�Nr��B­�1Qx�Ի��̢�z��BO�W}������!�3�ڽ"���
�a&�R �G49��-��M�CU� zG㉴�,T)� �&�ܑ�7O�f�
�)�K$i+�eϢ8y�� &:����c��6�`9���Q�L��E�+,);~���'c�R�h��Y��2�b¤'�(����R�X���р)"5T 7·-�fl����2Z���K@SN��y���->��}����
�A�ő��B2��8N��)�TR�x|�d�κ��w���x�#�:c����#ᄣ@�t�@5f�/�M����?a������bVC�4:d�|��+^N���u�hʓ���Fx�OK���5&�):�"0L�*o�ģ�d�5�M3��
����'�R�':�� ���Ot1�`�g�`LX��E�K���RώŦ͸��ZL��|�<	��L@e �V�ME"�	�AۿV�|Dk��i,��'����o��f���'��$B�X�n�`�`��
@�,���9�<����"d<�O(��'���z�d�@ꄫ	ض����B6-�O���v���`�	L�i����)�'ވ��(�bd.�:�ɯj�c���������Fy"o@�{�@W�[��]g����m�w�1�	ޟ�$���'��=��%7����EV>	�������'�"�'hr�'Y�FR6�I���у^3��pAf�Jʛ&�'3��'��'2��'xF ���F��Mc���>K�sAΩr4�F�Ul}2�'9��'��I;[0h"M|ⶏ�ld�)zG�ѱ,��e�"[��?�������¡J˱OZ���Y�MW(�[�F�'�kG�i��'
��'~��T���'/��OB8��2	��^֒t�����Cx^E ��=�D�O��$�� ؼ'�T?	�5�a�~-�$��-��U��$iӄ˓v޸��ix���?	��T�����r���Bӷ@�y�I<*�B6��<!���z���O��1c0�� e�ػ�IA+���aش/�������?A��?��'��|���%4��Iz��+,�i�w�޹l�6D��gP ��y��i�O��2�Y�a�$"���0hm&�s�/����I֟<�ɩ����ߴ�?a���?1���?�����s1g��#�ȹ�G-̎;���o����Ɇ(Vܛ1x���j���?�W.b�r|�D��E6\���Șzޛ��'����!�f���d�O���O���O����$&r@]ri�. Ortrbc��n&���\���Iҟp�Iݟ���˟ �O�p��"�v�&�: �T�F���+*�$7-�O(��O|��d��V���	�vy�����A$1X�d��I=OصYR*f�H�	֟���ן,��d� M�q��6-�����E��Y��p�j1��m�L��ɟ��ԟ,�''����U38+���B�K�PH`�k�S�i*��'2��'+^�'DN�H��i�2�'#��h��;>U�,���>l����#�v����O���<Y�N��̧��ɍ�Uc�cK_��ٚ����!V�6m�O�D�O��dƗ"4n�ϟ(�	��<��=G��q(7e��ˠkTe���ڴ�?)O*��ת-{�)$�4��� �Is�<���P���Lǐx�ÿia2�'��)+`�x�z�$�O�d������O>]A�̑rv��"�C9*):�
���V}��'؆u���'k"V��G���B��ŨW�R���Iul��{�$J#E7��OB���O���������O�����sW����_=����g�	݈�oZ�V���	Z�i>�'?��I�<�V�����*GG�}�U���Ph�4�?���?���vΛ��'U��'u���u�k�Y�rP��jN\�|��S�޻�MI>Y��Y�<�O6��'���� P�Br�c��tΐ�[E�P���F�'�~�)�9�$�O�$ ��Ɗ����&^�&���5F�9"[�L+�N2����	ڟ4�'0r@��0b��uN 걤 �\R����0���O��$+��<�Q�j����u*��yJ݉��'�@�<����?����򤛽\�,4�'m�ԥJd'"_g�脣^!-{�h�'���'��'���t�<�<$b��1+�����>�R��'���'d�Z���b�D��'�lE@���­�`8�T5�Z_m���' �'��	�DB�c�p3�d:^� F��}�j�z��i����O
�IP% �����'.��fK��lq'�H��\�S3�m�O˓q_j�Gx����B2C$81�0s�#D�L����iI��U<�Xݴ���ܟ,��=����%e_�D3�J0L96ac������\�0�S�0�S�7UX\
$�� Y����"jNO%^�nZ�H��` ܴ�?����?I�'h��'����-��Y���C?���%�?<����O>�I+t�h@6a��%��,:�(�'_Ɓ�4�?���?��a;4��Of���K0��*b�I���Ĩp{\��R�-����b�d�	՟|���P����ɑGf��dF���޴�?Y�HBuA�O��D9����Ȼ���+mvY)Ճ�>Hؙ��Z�� ��/���������Ԕ'[:��I�r��a�uf�k�|8�憂~Y�b���I^�ly�떸C�`�r��լY'(���}� ���y��'�r�'}�	,#K�]��O��qJGM�\&�C-��&���(L<1�����A���I��}
��ݘ&�1���-����?	���?A-O��i@"D�S"c�����l�4!�*���-��� ��۴�?�O>�/O���� 6ߊ]���K5v�~�P7�	�pp��'8�^� ���!�ħ�?��'&������.QQ�G4��ꠕx�\��h�K �S�t��._�R�� 4q������M�-Oĸ�p����J��������'�|��U ��c�!�O�6v�D���4����H��b?e#�@�	�Xhq���߆ܩ�j�����˦�����<�	�?ab�}@��>(��Nݘ9*�"���X��6m����"|R��J���J�G]�*�@�8�z�S�i���'҈��x�O���O�����b��1�u� =6�e'߫/@��>i�a�D��?I��?���֜v���+��ȱ0�%�E�ن=���'Y<�@�*=��O��$�Of����˽k�����Ȁ8��P���K}�F܈Θ'C��'bW���Ӄk<ԍ	�K��k�@�w��WS���N<���?!���D�<��l wP�2�/E"��ٵL݁qMJ��<)���?������XB8�'HBrT�ɖX*�`P燙?���'���'B]�Ж'�6蒫����C͏�)�B4ȇ S>&��� S�4�I����IFy����6mM�싓j�tu�@��\��M����?q(O˓�@A����Z#����<M�t�1��E�&�'3�Y��K��ħ�?��'J# y�����W��c�MA(6�@]���x�V����0�S�BP�IA6���J�,�J��U@���MC)O����O�!H������l��'�j=���B2�ơ�Wȑ�U���4��D� Y��b?)jK%f �x���8B�v�hӄu�P�Ħ!�	ß����?�H<��_[$��F3s�n��SMK
c��Td��%m�r���:��4r�h���-��x;bmR�Y��lZ�`��ӟ��ё�ē�?y���~�!Ga�Rp)!a�=d*"ũ`����'���y��'T�'h��"��'���@ �
��3Kn�b�DJ2t��&�������'��|���#��&3�V5QsO
�����D�<���?A���@7/�.	xp� �r�F�B#
_��p�Q�K@�I�����_�	y�*5o����M0/��Y�(�_�|,��y��'�b�'�剽s*`}�OZ�]ӕ ���&������O����O.�O�����'[�)uA�y,,�!�E쀑"�Of�d�O����<yCGH�11�OqJ} ���b2z<s�$Q0(&���jӴ�D"�$�<�k�x�$1:4h- s;^��S<n�2�lZȟl��KyR��	����$��z4hSdP�V�2�SC%�'c���J�e�q�	py��O��"R��$��Qi��h/Ցp�6m�<�a犸�����~J���ڗ���g��$͘�z�J� �j����ԝFx�����pl^,�@��A"�˄���M۴� ?�V�'���'w�dk"�ɽp.|���W!�dP2��5=�<=k	��?��� 2�Ǝ�I��01�A�'�,J#�i�"�''2��G�Bb���I`?��#��d�mzծoY�髤�BC؞��	��8�	$܀��Q ާ{�i���D�yHda@ݴ�?���Q4ix�'j2�'�ɧ5֩M�{���� :b#,�ڣ"����O~���O��$�<��K*HM���5)^~�xM��ðM� ���x��'��|�Q�@_0c��\����b���"�FLc��I՟L��Ey�`2�&擥ڞ��ׅ+8�x���"�6~*ꓯ?y������$���� I|��eBٺe�SUcF�t�듂?i���?�(O� 
D��b�܌8��� �2�bQ�!��4�?�I>I*On��Q��E	6n�Q��̈́^��@bh�
9��'�[��eD��ħ�?��'&n^0�bI^n@�
P��wh�h��xP�ܐ� 9�S���W�{S��b��9�\���kŁ�M�,O�eK���	٨�X�$�N��'m��D�]J�p0�.�8eYVp)�4�?9��k��q������b��d�Hr,����)O5��o��U��8Xڴ�?����?��'{H�'S2�/I#�4Xa�H�H8�d�=!r7�E,k�"��3�I̟�!�����!�oξs�`�Я�'j���'E2�'�\�Ă4���O���O�,�W �� �.��VO,DA8�;$$�`�B&��<	��?��$���hDaX�kP��ѓ'_�{\p(3��i�2b�9��O�D�O$�ľ<��0/���Ս��pT|�1��5���'�0C�y��'���'��Iq�>L�� �-jT��  �%d0�W
�p�֟���t��Vy2��%Q�Ș�(�=w7ȅ�AB�s��m���|B�'���'��	�6�С�����x���6@r�M%>�H��'��'��'��	(f�b��P��5�/���F}hR,��TB�'|R�'nR�T���ħh����KN='$*Ǌ�.��S5�iV��|��'WR�K��y�> X�H0I��΄�[%����S˦]�I����'w��y��3�i�O��	Z�m���"R>WH����Fm$���	ߟ�!e��P&��I�L�R�ϕ-������N�-�  l�IyҢ��Zؼ6�	@���'���+?�1���D���65a  ���5����ܪ�.���%�b?I��@��0"yi1�_Ă(�v|6� > In�ʟ���ݟ�����'��J�j]']1��8��^�J���j!�g�չ3�O��OT�?����u�lD{��Ț�� �k�Z�\8�ٴ�?Q��?A�_{;�'���'��$G�a �<��ۿ;�p����бO4��#&�D�Or�d�O�g$�.�P���#-W;U����!�	�n���}R�'pɧ5&`�~�y���	h*-)�$M���$J�7��<	��?����A�?>�!d��@�  ��J6i:���Z�՟���[��՟��	P�Pͨ��Ã/7Ȩ���)QX�䭐̟8�'�B�'q�OJ���r>)�QU�F��;`杜4B-B�>!���?!I>)��?����<��X�d�����9Iy�c�<G��	ԟ���۟<�'*��[�G/�I��E��7ꚔG' UZ�X�x��tnZ�'���	�̂1&L���O�����7��	6g����t�i�r�'_剹C��O|B��
�ðc��SgBC:[��t�FG 6��'��'�F�V�T?��C)  �
YW��t���(�!~�*�6��c3�iV���?��'J`�I��*I %k���I�6�(���4�?���"�����$*ʧF<��q#�� �ǔ9X��lډm����۴�?����?���x�'z�e�'`��\��h������B"[�N%N6�@�,q�d�<!q��ȟ�K�0C�R%��0<)|����$�M��?��:�T�@�x�'��O"�$��@�<�C�X�
u>y���i��'�h♧���O����O$�	!�X�Df���J�k~�P1F���I�X{F� J<!��?�I>��M�*@��"O.���f*�F8�'jU��'���w)�D��'86<��~H��#�\S��J��ׂh��7"O���s�ǹ+p '��-w��3���?�~6� d�8�5ñp7pU��&^4_A*<�1&�]W��A`R:h~R�ST'ĞO�Yp5䃺�#��W>s�\x�#�i?�X��f_ T�U�� B��5R%"��r�`0׿�v A@��e�
���ʄ������	���ޟW�rC&Fb���ۨR7�iI��)pO�� �*XAb�7Ϗfs"�'�"GY6C�"�T>�h�<N%�0�7��:�*`�'�$��<i�+4uL�Q��$+e�n�A2o�;m�MQ�和�(O*�ȁ�'@h7������R�T߸���	��Ԃ.J����9 ����s�@9���E��*�(�k��0��$�Ov�$��k�(լlr\a���4~��X�t�b�C����$�O��'*�>����?9��sw$h��$�
V�rL�V(�hn��w��n&�)f)�\�0�S����'�0(! �?I�HSi�$J̝�w���(k���b������ק��A+���;ćH�#�����
m���r�'NҘ���r�O޵¤O_Y"	&"���"O� �͘�UT4w��5p���0�	�HO�3� HY�U]�DQQ���):D/�O�����)��D�R,�O���O��D����?ك@��]�"�C,B�`����`���
o��� ��$r%�+<z��g�': ���fRVLH�:&N��g���@C��O�	�Vbɵs����ˁ�����)xH�P�t��1��M�^\�dR�[��'�ў@�'ЅJ �@$V6���Ai�
�	
�'�|��'m�� �F�X��	KPn9�HO�NyR��.�7-QC0�� ���S��Y�1�Q�v2���O���OP�Pd�O���m>�r/�r6��0�ǃ6{�[�ψ�vخa�'�Cv���J�Q��`L�kT�OQ������A� HKc�E�(�������[��ō`������)���:h�!B�Q� :t/�O��D�� `+*�O�D���L<z�2�� ��ei����� n���B���1�A��f�'��R�(K4)��X.�6	}��'vL7M�O�˓-В(�cR?��K���Q�!���!�kШN��-:CT�!8��'���'�r�׃��3�69a�L�3z ̓D*��s T�Iq�� fvF xcEV��i�&I��(Od���mv��81cZ�;�,izuO\EÊ��M�R���ShR� q0ȣ�뒢�(O %���'�r���,;MF\��0T�ܵS�EV<q�$�OtAɄ�z���3KŬI�`�X���$F{�O՘O:��D�r��9�(����65Or\c7���a��П,�Oj�sT�'b��'`����/�*�1TE�E�D)�G		CNpȱO��s'<�QJ�]������1�g��Z|���ekT*9϶����L#\&�|�v�Y�o��q���W�:gȠ�&��'jU����;Q3qȃf^�l7 Q	�����4�E��?I�i���S�S�?ٔ'@�i�JO���Щ�'[ɖ@��'2�u���K�0�0ℭU9��Q���Xj�'9T��^)��fɘ(J\8���S�y�X����?���6c������?���?IԿ�����O0�Iv�����8`�O��J�;{X-�Æ�=Gճ�D۝�vm�'X�=pAn3��">N` ���R# ��]�f�D5��㳂+g4UJ���>=a�h�ť?yH�/�R�1OL4!P�܈M��#JY�um�c�ONd¤�'��|��'�"[��C���W�`�毆 d�pa֪-D��0�,K4H.�;�LF�q�"֠���HO<�	�O�˓V4l�:q�i��#��	d$�H�`Q��NEJ��'��'�!�&���';�	�<1v�Psjp�l����@�
5�$�dJ��Q�� 6�')�E�t�k�&o��bI�D,ԋE�J͠�-��p>	������6�^�!�� #}
�@�7o���$�l�I����?�OMn%�UH��X\�@0s��v���C�'�$钅�Y2:�\	���/?��i��'�d����
Ԗ�l���I|�4"�V�����#��D�(���)��'l��'��q��� %iVd�����3��:p�^�-�Z�X2h�>�Y���C' �P�b퐯�(O�EkBnS�/��OI&�3am�5"���R�oŌ-��&՝r8�KRϗ��(Ox�[��'?b�'92_>ź2�	?0������U��բ��|�?E��' �!�PjD|��s���+I��R�:�'��5���4lьY�'�`K�(�'�9�vQ��?����򉌾v���D�Ob��Lc���ė0 C�58r�ك���X�aV��&�ʧߘ�?)�gH&[�)%�G�Xt��u\�r*\��F��"m7ɧ��r%2tDx�+��K>��<IeC�+WF$CG�'�r�'4���O�!х�A`�Y��Q���>O�D/�O���JH�9>��(0���+�(�Ru��:�HO���\A�&ù@Ohh�E�#I��y�	ǟܻ�` �@�f��Ο��� �]w�b�'H(s��0+�N�� ��ky� 3�%�H���I�#Oq�����0��ĩՍw����<!�I_s�ݹ�#E�lE:�KF����AV$؝g>�x
�S�tp��'�,캒 >�	��iA��ӢX��UJ��^�8x�	e{8��������?��?�)O�i��Y�cBRMq7 RQ,�r�O��d�="oƉ�U��!���s5�-+uX$Dz�O�U�Tcu�ǳ�M��)F�*ǔ���E�4t���C�?���?	��0a�T���?A�O^�qРB<�"�b'؍�l�k���j�@U���	H1BHؿM�����n�'�X%�ADʁ,|M���!;� �`Ȗ�8hRM�̓?;�����7�M+�Xo�'����g�6�+��=�� N%_����j>�61�Ɋ�H��4P�0��>���C����6O<�=��*YaG���oǨX�|�[�<鑾i<bV�D:r�Ĉ����O4ʧ{�>=��φ�m�z�1��3I�Y%)��?���?A�\b�*����1]Ӝ����ɮ &ڭ���R�'<đ!�N,q���94�'uR�Ey�]PY�H�=G�p%lڱy���;��J#��1A��U�8���R�؜v���ӊ��9-��u�60�~�#�]5f���D������^�<�����>�%�ӣ2V�p�Œ�yM��K�@H�0�M<≏�PqFX:��<LK^���Ay��b�2��-<O� ��p��Ts�<)��.�Ԩ83�"O��z���=JS�M���r"O�����
Xq��p�E�'S(b"O���`�d�A�q��/?�$�g"O���4)p�$�a���=D��I"O��Q7,�0Z�Pp��4s�^�j�"O�u ��Ђ+2rtc���E��Ea"O�M �B��%p'�O/�F��"O��`7 �h/��9�GҺ�� �"O$���Ŋ=�AgE"P�2hr�"O���f��4o�H�tF
	B�A�"O~�J���|��MB��"PN�K�"O^D���(rW�%��B�v�N�A"O��ƄR:�0A:r�!(�� �"On#�Nޟ=o�-9!��;Mq��r"O~T:ׁ�3�2<�"W[E*y�'�,�k�ȴx`K�wĀLb�*�p�<��Κ'�b�Ʌ��L�A`�b�<���7I�MHt�C�H`��Z[�<AGŖ+�=�7d7K.I:���R�<1c�*�Z�c$�$T�v����L�<i-��Wk<�����ޒ��el�|�<�B��/;(% P��??�j���]�<Q��J��:���@K�H@LR6�G]�<��E֏N�2���d�5!��<���Ht�<#��6��R&��D����F�<�a�Ϙ?����t�^U $�h�J�<��eˊAN�<��g��Aqd��׈E�<�V`��!�v��5k�=�0<��&�@�<9��E��������J�j� �^B�<��I
P�����!H�a�b�y�<Y�l�W"�����	�Rg���F�UK�y!Z���r��"|��?�$��H� iu\�p��ٔ`�����OI�碔�MO��h<�e�l1`¨̛l�hĉ�"
�B��C	�(�'�"���'�S��wY����
I�L�'o&�T���M��:T	�A(xh�fmB1��O����Y�� ���6+VW�߫�LŊ �В8x��q+���'���u#�;5e?�y�+��� �Ml�����$[��R���{�W�	6p�4��-QS��E<�ԟ&���
��Q�BhӓV)
1ȴd�	n0�'�
0ʰ<���ԧ%j6<kI�nkͿm7���kM���҆�jZ�g�-�$阋y*�qO�e����f���0�dG "��L�0�J�Z�@jr�,3�v fA�ȨO�N�ʅQ�+.�� #�Pv�z�\e���ġ�)%Fv�nN�W�Ԑt�Ah�:�D~����4�Z������c��A���F�{�o� n�!
����n]
T�=Aa�R��'`��B��C䉓Z���p���	�{r�;~|�It����;6|�=sVCB�X����I'D����w�W�p4�ȕi�+Gdp�=ɰٵ�u���0Rt��ƒ�\9�C��M�V��-�B��	2���8Pc�$)��-���A�S�>���@I��]�C =
]�` �N��z�e�@"�~�pС��&Pj4�>�;^�(��d��Q�@�A �j��O)��	3�)��V���6&Xc��58�f�h��I�n��1ci�f��Y��b�����
Ub�هҗ!lm@0i:|O |���&D� ��X�e��%�v��l���׾�HW	&?!��ϣ1{��I�%?�$�rĸ<��!M�yfG�G��]z׃�9���J�?y0 υ��ğ
I�R����Oz��6oM��	�z�:d��Ő�TR��P@��!�.�ãS&�XK!�*�On)r�ݣk�h17��+*�0s��\�<���0ӊ��&���O���-��Ix���( w6�ۇ��%�yˊ:W��B%@W��P��mAi0��E|�B��(��)�"J�,�&�w.(�@�� Nkt�B��N(9 ����'�B�teȶ^��P"6��:'tx<��A	9N(��Z������L��(r�H�oTJ��C�3z���P�$��|�H1��_2��-&�a^bQ� �
�<AH3��<�䴔'��q���.�i��H�oPJ���8g�͢�
+�O<���F�t`� ��}����zB�Q�:�Z���,��.�(O���JU�� u�K,$t#���z�h�O
I�B�5�)�S�e��KǓ/~lt`�\#��[��@q���C׳o�lub�LT@��]Xl��*K
�Z�[���+_�h�,��ÅO�S�C��*l�� V���o��S1j8��N�_��U��S���U�QU���q��^�����G2��\a�I�S,6賲Z1h��q�v��q"ם�\��`�I��5P�@A$T�$qF.#"�ιȂ�["JE��%HA2'd�0 ጫl8�O���}e��vg֭rƾ�ڰHK�)��k[�A�7�F#�plZ��ʹ��">�;l���r�"ƹc��0Ɍ�h|�<�O�E�e."�)�S�.��v�A611b�C\մ����/�e+��p� !�QE��A�$Q"g?Tj��
�3cF9��-2���=مҟ�)1��Y �@�HC�&��̒��F�o���'��8�!+G�0_ ���� Qhj�{�'yk�d��lZ&r�)�b.̯8߮쑳��G�/����L�L�@f��̄�OKMg��c4��?v�r���#�E'��s��0���[�S�>�D�V�,��#�>��R�F��n����bNH�#�� kj�>�;"�8D���	8~K�!
 *۹
_�ݤO�AH$�)�SE� b0���V ̚��2)�HU�U�	 F�xi�	ЌYM�)�v�DM�YZ���??O�<�#$3N�2e��G����Z2d��{���?��aԦ�h첇�^*~�R���	90�D��O��Q�02���!O�vp�	A�Jh����ʁfǳI�$@Ӷ���m�`� 1�Oܓ&0f��Zw���z2�$(ZV�ӵ�>9�Q8XӔ ����+s�&�Q�V�s���1E�i$.�pW��O,>��|
��p����{_�$�g�[�Pp���89����m_28��>�;.��`3L�(^����ի�	Y��<%���U��]�qO�c�P����2mD����M�N}��%-oQ�,�B̟�a|p����ķ?L�Q�v�u%�a{�m��A	*� �9Z���{���R ���qf=1����̖-���%␅L'>��
'?��C�KN}��=a��۶Ss��2��YCug�}�M��M[ EO4p(����&�+(����G��I�h	H�#��pgp�dg��4�� p�-R���sW��V��Dx҉�M04��ԉɤW$�𒡟��� K,�Mx�HR,o��XF}�w,pIa�㈂D
��Ѓg��^=��ZL>я���P1�p����	j�`��%�\
����)N���rƜB����ww���p�#�z���&�I��qȁ�d��'삐��\X���t	(!ܔ	���&t/.����7~���h^] 3�O���E� 8�1O�	Ω>^����+0�2���X0�׉��'~�Q��?�s�C&R��R&���%(2�ȁ�č�&~�p�m�@�C�>y��if������X�
��F��ɴ��!�����ތE+ ��e\��!矯vQ��t�zli!M�I+hTJph�j�|�C���A�`�؄�V!�� 7��Q���G}V��j�']�����2?�
W?9"�I�rN�P���+�k�.!�p��'�$jgd�T�ק�OY\,�KO��LK�J�/'�>��O*p��ȅ�~��Ղ^�u�y�O&�!PsC!!���i�\T�`�e
b�ɩ hDH�P�?q���Y���e�ZDNS�>�� �W6�R"��d4�ۄ�SO��?�O�@b�ީ�*��爊'"u� �ґs"h��&�(:�Ys(B�L�,;���ֹ.�l��5*���Ma�t�LpD�|�x�o\�/z�u����_��-�`��B�BՈ� Z�V���T�	�Z�*�)P��-A�$i!@��I��$���<x�VFt�B�Bぼ��)d��Vx��j��Jy��`UBS&�t��H��,���8�J����kE>)�`�C��W�}Pf�@?|2��6K
�I��?�dj�tv���dn1��q�C�,�ʓ-|T��L=z����=e/ ���O�A��r��B�Xe!*�P���10�*��$���S��l����d��Zᅆ��I<�| ��I<"6`t�$ȮS�(��B��7r��!fV�<���8��D�6:r�̱e�I��f���/�dR�< L>��W��p�ß+��h��
�Hw�'O�P��tN�D���&�L4|A�%�g�`I��(��p�@��߽;��ٲj%~�C 8~,P����<�T�,�`!�a��0E�JL%?��9��M;��ɒY�� �v 5u9�����~����'jr�WGIP|8�1C4^.��{��8�Ȥ fD��Q�@E���J�@e�u��V�xB�-����P��ȥbL���d� �3}�#�6a�ĽzWI�mr,��tF��r��lbF̋7Tmӊ{������嘠� �&=R�	9@֐s�͉#a~ ��a�3A���lWܝ:���2*�V��1�@�uY��*ťG ���r��>1Q�[���dM�;˚�a��v��J?y�R��¡�?(�XxrTh�h��y�V�	�¡�h XypP`�'(���ޏv](�A	<��0�����y����1S`��I}ǌݙ��)�Ic���W�nb��͔�*t�Fn�'��H�b��Tꢅ�,e� `�P�T�C#~��6H+���u�Ȑ�T[�tR�MV�(Hz�NDGy�M	�e��\ɺ����ۈu��T"��ɻ�
�B��3�}�d�Y�b�d�	�P�mԼM3'�(�?˓B���/�RAk�R6jFH�R���"��,$c�n��ao�����	��}2f�ڹ]��[卪-p�D�7L2}�.�;���=K��a�ukE���O��Q-���X����3�)��ǔ��PG|Z ݙ�Γ1�fAQ�͟	9�GjΊ[�8�B�_�E�`�HńZ$r��ɯ@˴�Y������|��OdD�[u��0��0[�P��5(c�J��iXڅ�`�Q9s�Q@���-N|�?�3� ��`��#7˦E�C�D3W;�)�-�Q�I#w{ )���:Y���ݒ)� ���>��d)i�ޑB��ݛK]T���l�M�F��R�	4�޼�?E��![�'rV)�}�^��`�Ǧ`�T+u*G1!�1ۃ�
J�~m����^�No�����|+@$z����]xV�J�}��T#ηb�e�N�%#l���`���})�韢d�F�c�l���h�<�y�̀�E��A�1o��]����q��p>y��1P�\<1�m��Z�i;�Ƌ�m��x㏢?x8�u�|l�Q��X����IMFP�Dz�
�;a��g�ָX�"[%R��(O"�I��Z���c�ƘD"Y]�`��cS,",���Q�X�_Z�Q��F�>�6� ���
X��|�A�d�b=x�Ï�Q�.�al�\�ԹBB"ƣ�����B>6@���4��JaAD�P㬙�
=E�b��"O¹�`��u4�9{Łɲ�N�� �ͨOh�ZC+����-��愸(�g��q �͂�b
�>������G�p�{����|5���1�|l��S"~�!H�d�.4�@Y���VO�g#t��_�,򐀐y�I�5_�H(0�	�B�J!#�N�CռyF�� k�	,s���P+`�ǩs�Wp8"C����b �A�r,R�p�	�r��	Jd&`����B��ļJ��zG�(�Ĺ~�d���D܋��a�s�������?�����H�X�hL��E�=��1�К������ zh�t��9Y(�ը�[�X]G~�Kۇsvp��F�،m ����U۔T�FM::�|\Kc��-�(�=1töɸ'W���?%+�(�D%�+`�����N(��LQT$�'����j��H���X���y|qO�D�*cx�U'T/gP���'n� D@���G�[ad�\2���7��	����q�C�3&=�d����N�h�`<g�=a֫ZF�S�>�F�*��(���,S>��Bb(���&�2x��0�胉i���杢rH��ȯIȃ��Ӻ)��' -���陾J;�E���2L\�р!3Rz�詈�DI�J��@#��U<M�R0!��w�h�Yfc�� p��fB�3�P���D�#s P��ybZ>��o��OP8�!t���(����>̖��'h���UjW��,ɱ�*Ga2��L>�'��છ�		r�r�ɀ[�`�F�~�ɠV���'K.�X��(�W��'il��Ue�n�
!�M����V;����������S�OHڱ�N��(0J���!(R29����j=���^�.�&-�SԧyG���~�:�{!ۙQ
68�Ġ���A�,��d��҇F��~�h���_3A,�*�BʷN�8ݒr�B>!��3��� *i_:��pC�Ky��#�r	Qb��_xՙ��ìL�\t;"'ǱP%V���]��p�帟��������V�Q=\�D	���+q4JE "O�}��h��/P��sg�$1f-��"O޼��'eۼ�[�,Ƞ"	�Xq�"O�����"���@j�=s�\s"O�A�a��"�@PY(q�W�ˉz!��v�x�y��F>d%Ia7l�5[!�$P(��4��k�>�$��Q��/Z!� �Y��У�ȣ^F��H��S#6X!�ܽ_��,����'H4X�p��/`�!�$�~˔Y����,�"�j�a�!��*��X``�@KVx��
�[�!�Đ+c��L�v�C#g��(E�Z+vd!�$�:|xر0�#J���!���@�\!�L5�\�B�iA`\ S)P1|!!�_�g���b���;"�Qf���l�!�Ċ�k,]�W˂�X2Zp���UK!�Ā43Ȥ�9�H�@���c��B!�@�v�������!\�V�K��V1t*!�DN�L�
�+@4�*���U*!�d�z�*qxd���2q<����=
 !�d�Jp�mq��&8�hbr�]�\�!�� x,r9`5�;(|���m��g<!���,G��D�Q�M�a�<�Pת;%!�o AS��
�eC	K=L�!�d��@�F42��˨�Cə��!��K�ܔ� E�9:j<CV��&T~!�$P��A�GѶg;F�`�j>as!���vN��"Ð68�Q5��o]!��I`������H#P��p	ͷE!��T�L�x:��f�8�hw�!�� ��H4Ӽ�,%J̓0��zE"O68b��יQ�L��.,Hu�"O`���܇|����@	Vh�Z�BT"O�E���=t�|@�t��:qґA"O������i��A��.[�,IF"O�QY����y��1c��֎d?��)�"O��
����� �t,�s�"O�x���=rpQ��^��"i"O+j�*�3���4���3�"OR�{
�w����Z�%�N��D"O∊�($t�����^��)0�"Oj���;,��݊E����RR"O:쓀�P,v���E�7��,hr"Of$�Ue�"�2@�_h�H�U"Oz���O
k������.��P�"O�h��-�!L�¶�y�(��"O�@��`��%�� ��B=�؜��"OPh2��L�*@z����/$.d@��"O�hp!��&1at���? pU"O����Q
gB�k�͜���8��"O���N�Gx���5퍁$��DH"O�I�@�g�*r��	���T"ONI��>�̨i���,7��İg"OL�pˁ��@t�v��*f<)�"O�; ��#�ι����0'�Xѐ"O�a�Dƥ7�{�&܈n
���"O"�0��E�#��E����R���"O����,{����^�6D(���"OzH���Nf�4#��"O6с���<˜U�5AAU� �R"Ob ���
4���#�X��|QS"O��j�l�����DaM�*��jd"O0-�p��?�4��I�.ߐ�X�"O���m_�6�7�,f���0"O��H�)Df1TU��1(X�$R�"O!�4Eڙ9-��32(X���"O,h��ǃh��,Bg��r��w"O�I���w���P�oj�]@%"OҀ��"]K�I�q���d{�aQ�"Oh)��(_����c+�c�� �#"O�Aq��]z"e��
@8+��"�"OL�	���������F�/$�]ӓ"O��zv$�&T��baEL-c�P@�	k���)�*9`j�R�cq	I�E�:E@A��'v\�S�M�f�d��P�U%��ɱ�'�8�� 8e�")��*F.D[�թ�'>�Pj4�O%�pC?AҖ18	�'fВp�U.\��! Ϗ<>
8|��'�r��e��L���-ʘ!�R���'"<͠l�,tJ�k�f�%�'b<�S��?��mM�Pz�(Rr���z�2&�|�<���D~@\%bB,�/E��	P�c�<�e��3N��r�B.��%�"�U�<�6H�%��&i(X¡cP�L�<)*=x��%�Χ ִ� I�<5'��ayw�#"o����h�H�<��_�v��A�mc�쨃�@�<�t���!����h��`d�@eOHX�<YV�Eh�J�q��� ,�`����M��>��J�O�TLhtNI�m��ɘa�%T�����'@�+�lT�R̲�����;F��
�'�̀s��,juH���j@�'��q�	�'E�l1��{��J�I�4=�q	�'�(U�EV�>?��8�	�>������ ��fO����У�(��C0"O��%g���H����@9"O�aBhK�b	�lѳ�4�r���"O�q�F��M�,|��c�j�XL���V���	֑9��@qELҙZ��	�Y�!�MXV��P@h�@O�(�g	ؠyi!�䃻R�zL�W �)1 0PC(� \��hO�̩���jD:���	�h���P�"Op�bW��ҧaT�Rq,�"OnE�Խ_&A)f+� ��"O$h�o�Ze��Y��֒X�)"O6As� �`�4T#@��P@�P�6"O,�;��k�Mt�n>��H0"O�bfB�,(�v� ��T3��jf"O쥓A	Q/&�D\���Ƃb:�(�"OdU:v$�0� ��f��=���"O�@S�BU�������'L��xX"OB��p�?���fG�_�3�"O±��n�� �D��Mw�8 a"O^�X`$I�p���6⍀jn�ɩ""O݊��D��ِ�B2���b"O\!A1"�>6k�1�τ.`=�S3"O�A�I�e�̹,�+$ɢ"Oй��"�m,�Qdj:!�
`"O�q�A���s�b��u��3^�x=��"Oh�jd茼
h� w��9E��R�"O��BB�iX�ـbW�F�N�+"O<3��x	�0b�юᢅ"O�i6��!h�<"���6Z[��&"O�`A%�U&mY� 
����wK�"O���3�Q�t�DAzd�bH��"O
hC2c@�O˒Š�fW�q2A"O�]	��гj�(��˜&�y�"O����(�/Vl\"䤑�H����"O4,��c�$b�5p!d�d���S"O���ô7�Lsuȕ{�5��"O� 0�(�[�yH@�ٔQ�h��"O@h(S�X�]l-Jo��Y����"O�ԂTC�*iL����ߦA����d"O<��
J(���d�)�*訇"O,m���;q�<���A4j <��"O���B��",����Q�ڤSgd@�"OX�!�I]��,��0ɕ�gx�@yT"Oz�9��Q�s͔��(բ1x���"O2%x�BU)SB���焎|�,�T"O>��Bh��e+�����NÀ�e"O.$�A��5�s��6�,��b"OX9�t���c7�i�AJCp�с&"O���&�� 6�R!{G!�o \i�"O�) ��HB�XW/̰w�"$�"O��ծ�60�����F�?x�U��>��O��=�O˞ ��CW
]y&�Jd��=f����'����d��q���׏c�l�`�'X�I�^ �H�@Xˎ ��'�&��"��]ݴa����`�Bt�	�'.�@#1NG�!쑰H�^`�K	�'���#`�ܵH���:��T!o�@��R�'Ԏ!�3�"<ഌPŉ<��	�'��ɨ���+K�Lz�G 5=�d��'*�Ea���"J�`i�#�'8B���'����	Pt��Q�j)9%���'�,�c�H�jK��۠�D��Г�'\Vu�c��tZM"��	�u�"���'�~YBD�]�h��]���RH���� `eCӤ$8mL�+f���!u@�"O�<�Agط�lp���C����"O����&7��X�#EG$D�*��q"O�<��k�.|�dCS�u��5�"O�31�4��� �ڙ{��lH#"Ot��c ��B�P	A?�����'��I�cK�5�B&Y*!�>��G�Y��C䉋^� ��R��=�庠���{b�C�	�6�|��&@<Xw0x!4A^!I��B�I<b�Z�qc����!0��@����F�V)r��ӶB�4A9�I���	�ȓL<��ѵL\V����)H�H"�!��r\���h_�O�������N��ȓ?!r���!E������f�@(�ȓp���0��4��!����m�⡄ȓ�E�G�,}I*��!��݆�a �� OB�2H�$��@�<?D!�ȓM�l=�n�9��*��6T&�"O�l�r��&1#H(#f��q6v�b3"O����d�� Y�Dx2DN4 |Y�a"O(t{5/ְ;����vC�7Z�ؐf"O� �6.�T�n�2��	t3��@"O�����\�s#��Y���y���;�t�C�LLv�A3�'���y2 I�"��Z�G�o��R�S=�y2J"ld�}�aj�a1�d�AG҅�yBoS%�h��/�dv�����'cў�O�|(�t��#H���� �r�x���'I~���Lad��Q��
n8��'�x���CTQ�䝩����f��@��'��YSZ�K��܉Q�0[BХ�I�Ȅ��< �D:͈4yUmq��	�,B䉐qߴ9��T:h��̂3B�@�C�I�t���)W%?�ta��%j��C䉐!JnH%#�)o�@� �88F�C�	�$d��j2�]D�$��A��H�hB�	�t���g+�<
SAze�K�<G�B�I4��B�\�@�Œ7&�=NY�B�Ƀ�L�C�*߷&��"�-R��B�I'Q�d@b��W.*w� bEU #�C�I>��Ի,�!K�$i�,߶��C�	��uR�,�4`��1���B�	03WJ�v�Q8N���8C�ش'�B�I0o��P9�!�C� ��V(=��B�<E�P"�(�; s��҉��B䉽u���.� ��#�Q�B�Iz��ӁF������"B�uC�I	#��$�׵{�$��dn�
�B�ɴi���D'�1$��)��l+�B�	�>�>���a�G�Y3g�ۆ{6�B�	-rh[�7�K�o�ZL��d��"?�B䉗"�>�:b�p�2������u�HB�IeRj3K��d�
�a҈�c|tC�I(K[�9FK�1�H�0h�L`C�I5b�Ȅ!�`R s�2��b*�DC�	(�����/);>�m�w�R  ��B�{�`�����P��@�Ё�C�I6(`+e�Y�	Zڸ�rk��*L�B�ɦ9x􀈶��)C7�|k2��!LB�	�e�ah�%I�j=�4�2bU�N|C�I�_D�9�5ᄉ<;D��2c��h�C��7P�"�eC<@T�ţ�PS�bC�	�98��Gѝ��)a��M�$-DC䉖kFaЎS�!��E��z�C�)� ]GA��w�@u�V�X�6���xW"O��	��ϵ��)�H�&�6}q4"Oȥc�)W�:�l�E
B%�^�:�"O�pr�A��|��TB�f��t���"Onq0#*�> ����dd��}s�-�7"OHq[���O�Z豲��F���C4"Ojs� L8���o٦G
՛"O�X��_�Mr��	X�r#hi@"O�p35��6R����i�"O8@	��Yk���AG[�[˼}S"O�ؖX�N�L	e�H�8b�"O���tC��#�݊v� `h�L��"O�=s���#�D�
c�X���$z�"OL�&I8$��S1�Nk���"O2���|�
Y@�� +Z��6"O�B%��r4PcO� &�~(��"ObkV/�)[�ڝ���N#+P�""O���O��4��fIL�D>V0$"O��� BP�en����M ��H"O
��,�j^�=ӥd���vEP�"O�� �GG�c42T"����PV�u�T"O^��T�M=n��F1r�0�C%"OD������}�
9�רC괲6"O@1���C�>��]@'h	�<�b�"O��K��4L4�ᴦ��V���X�"O�m�PJY���\�T�I�`��'"OVE@3"�h_�5�"I�$�x�f"O�A`t�ӶV+��A��/��"OP@�t�S�IB�J0�~���ju"O��Z�j�.9Z�p`.�D�X�t"O���I�L�cp��64Q|��"O�e�CC �yC�ݑ���6	AJ�%"O����2`e�9j�1�Đ�"O��ꠍN�]����Kv&�}� "O��*e�BP0����А2@P, �"OqC6��,&$ t���*��!"O*�#-��4fѪ�Mش"lz�"OD��r��@0"a7;�Hx�"O�Ia���g��8�2aF��DI�v"O���o�6Yх��?d�5W"O��#�EǑІl�E��=c��h "O�9K��iN !!͚>����"O,����[�.4	afF�
�a�"O���ۦumb�z埫[���c"O�s�ĉF/z�"AW� 
I7"O���ۋ	=�	"!�6
��H"O��f휌=�e�Di�/����R"Ox�� "�\�
�"�hRt�Z""O������w*$�85�  ��� "O�훖��\*KaĒ�b����7"O[��F_�Z�l�q7��r�v�1�"OB Kq	�7B��|��BY�Yc�u"O*ܓq ӒIxQc̼,d�i�U"O��pхG=
%N)JQ�L�t���p2"OZ���J�E��L�_l0թ�"OF� ��,\5��A`��=a6�;0"O~���j����%Nb^4�+b"O2���E�6tJ ���N�6O�M�g"O���h����&-9���2"O�d�ӡ�
^�!p�GW�q�"O��0�^"y����k|��� "O�]H�"N�.��f\��B���"O2����R9���
�\�����"O`I�%�C1��0H��� Q$��Ȑ"O� <��R�w%R��p�Ï~�@@�"O<���]�^��P�D;n$S"O�	��"�!/8Q�L`�lC"O�i� O#�����c���
�X�"OL0;l��;�ISC��2FH��"O�1�!ٷA(�!�4��bF"O�t�a�E1�~]��
+y�ڨ!g"O60�ޏgY6���@_{،܂�"O�S3��&��|1Nڣ}�d�J�"O��ߜX�JLRQl
��'v�!�Y�U�0�ց����a6W)�!�$ChW��Ci�2z�YJsCܹ�!�dO��4` �,N�}�e�?#I!��:� 1:��ݶ/I`��s�J!N!�ٷc��	ь�d�p��T@.:!��I
>� �s$��87�N�A��7X!򤆻a}�����*�Ȧ욟U!�䖼��8��g����T(kI!��-�^�i���k������i�!��T}ЈS��<+�����$�!�9[�te R�3���Xs��f�!��C���P�@B
ld���'�!򄁟�����Rb$)�d+�#>�!�䗧X�0a��.8��|ɦ*M�M�!�D�T��<��R��P�c�H�>D�!�d��Ԉ�v�ăy�(����!�!�$�L�n���MǰPh��K��[�5�!�d��~D�SI�'w��� ��Zr!��
]i�e���:iw��M�S]!��=-.,�΁#PBJը��
�k6!�$A�F�F�A�148�=�1'ӡ
+!�P�}+���U�u+RI�F^9; !�dFtڀHí��"h�Q2cƋZ#!�$�8��Z?"\�p�^�B!�$O�pL�ӻz�L�A+��!��D{��ز#��	4��Ӏ_6�!��Fq���aQU���z������dL��~X��S(hw�R'�X5�y2��%n������֝`����aL2�y���عӒ�S�O�"���BS*�y��X���YC�E"O'
ySlX��yҩ�%)�aLL�,����/�yҡ	+!���qVY7@�a��%��y��C>c�j����Ƕ<��Y��y2o	��8X�ũL�7NH
coϠ�yRa��F�x�kI�]���r�X�y��:��]q�lXE��ѩ��W��y��$(P���Rj�+���� ��y �,8���ѕ��R���1�	��y"a�?�@0IC�B�l-�U*�yB�{��c'C�;��)ủ5�yCU�.�x���4���QIV��y",A>Ü�@aC��b6�)s�S�y2K����XE��F��=��ň%�y�-�=v��1I��δB���C"�ɱ�y�� �)7���` �3�� gJ(�y�d˧)
�;4���;���P�cΞ�yb�Þ�4؂��#$ �AX�'��yμ6�1�fJA'*5x,�QIB$�y���]p�k�bH7��*1���y��ȑN��٘��\��^��3(M��y�&D�M���٠Lș<���Ȑ�yr�ܫ���AHʹiĤ�B�y"�F,O��{s萤}��aR� �y
� j�qF�Z8�U��;$uZ�"Otu p��8#��4)Eԋ!��s"O�A�t���:4��K,*}h�"OZ����KǢ0��+�<@�"O��F�R�F5
P
���6]h�"O��!�@�/Um,2�.M#
�ʱ0V"O��I,&�(�d�PR�tUZ�"Ox�Ģ� `��� #I�	�h�iB"O�(�� �EYЕ�d+J7Qy����"O0]�GOI�N	P�F�Li $i�"O�1�i�1{ۜ��tI��;�m��"O�`-�	�=[���+.�6Y��"O���f�-�~�5#N��t"O��`B�A�L�B ��s�Ҝ�U"O؍����U!1��B�D��"O>*6���6j���Ť�	�81�"O�x���]�n�܄�`-�G����"O�Qp��"T��aX�S=V��̑&"OX��A���H\�9���#�Z��P"O<L��FX�>n�3��5jb�"O�m�WhaZ�4aS�|"�<�"O\iHQ�̗y���� �ֿT3p"OD�h��ˮX
�]Dn�2��5��"O���B�	3&t��H����{�\��"O���
Q6W�Q�Sj�(�Hۓ"O\�c�B���"#I����"O��#ঀq��A�&�83����"O���Ù8�x�p¥�����r"OJ�  eT�� ��pc��+ p���"Ojx�5�L)M�0b�P�`V�1"O� s�`�3;��i!��/N��5X"O.��4�ǞU�����\�
I �;�"O��ȰLS�/9Ȉ�E��@/z�"a"O �ѐ��RD\�2�U�MFp�"O�����#%K,�
v���h��A`�"Ox5���1;�xa	�jS1/�\s7"O0��̰#�!����Ѵ�R"O�ix�W���XECܢ-����"O�yr�'�
���&�R����D"OX�H5c�1\����؍M�buH5"O��(w�θinx��E�ȂI�B��"O5Kl� %]�Dڕ��>�}�"O*�R7쏔%�1��ϻiԨ3"O�a��G��5�`qVy�P"O�#���\7b�x�c��:�ҩh�"O~\����E���P���'����"OxX#W��#o������3��U�"OHg�A�PN�RgҴ>o��;�"O�<(AC��K�T��V,�6l"Q�f"O\u����-Iw�8�2��% ��Ax�"O���ã���%x�n&n��"O�$�tiV��(�R�K�S{P�(7"O�m2�W�]eL)��L��1�#�"O�i���
b\d�I�6	]�,�s"O\�I��Vs����N�Y�!��"O�	aS!W��)���́h��� "O�]�I�$Do�ݑ4F�R� p"Oh<���Ch&زKR�zM��	`"O�$iuG	 y����	�-&��*OڭQ�7G�P;��,}��� �'��-�"'��Ã��|�F��'O�T����=� Y 2���b����'���BB� @�zXia�ϲ[�����'(60A�iΆ��y�W�=[�h����� N��bK��:���L�i��4�A"OX�(���_��U�)K�Pt�̰�"O~��a���R'�ձ�Y67��E"O�A[0䓯8�y��&���r�"O<�r�N�1�>�५B<��D9�"O����_�^=.]#�jݩ|�0�C"OZ�����t��	�Wj��E"O��9����B�
�#��q��"O`�"&ɏtSbL@���J)f4Z�"O$ѩR��[Cyj�N�2z0ʆ"O��xw�ɳA�0����]����"Ofu�V��@�8�N�1�V4�"O:a�+øH�:ݨ���R����"O�1DŒa���xH_�#J���"O�4���ߥڰi��\%d>���"O0�i4抱I��0봆�bҌ��F"O��I�j��hf\�Ē Ϙ�2�"O�|��bӈH!XW���A��\�E"O�2�)R�j��q2���#��`�E"O�uaP��5*�"RJ��d0�"O��Kƣܵ�}�޸;T,��Q"O�a �8��L��oW>�!�C"O��Y�f��A�(�:O�~�>��"O�9j��ΑA�<��1��h9�`"O�tx�D�j��AK'��9p�,�k"OXU1��đ]0"`0b��'���"�"O��ӢŞ`�����[�hxq�"O�m��&B�'R ]�6[Ĝ@�"O�"�c=��
��f��k"O>�2qM�!7/��a6@F�\
l�C"O��MN�ڨ!f�:S�Ȕ�"O��3�ʄ�^��yR�b�']�����"Ozh�Q�/W�|��!�+i�l��""OX��S��;ET��3%&�VL��"O������K#b��	ͨ]��"O��2��șD�@�J�'��5�8��"OLɈ��U8!�\X!�ES8����"O�4�Ao�mjx���� 3#|>8�"O̼`�׮5wD³�ͰO{E��"O�:����o�:��c��i�K�"O`k�G]viJ)H&��T�vMI�"O=S���(P�0�"��+�|�B"O`� eաm��;��
6>�]�"O蝙B�
�����T�k�:��"OH�)��O%����	[v����"O�dI�*W�u�� �BHGX\Q)G"O�:B�V8>:n����X态��"OTaIQ"�b�ty�X)&�%�G"O�рC���R�P� E�,l��!"O\D�%(�Y*	�cC�vV��p"O��H�,��}�Ǣ^�M2	�`"O8-�Q�V,���P�_�<���T"O�e�f�Ɏu��EZ#Cz)x<�"O����I�G˨E��M-��"O2ӓ�I"�2�JP�%����"O�)ɣ�<Ў@��Ӥx����"OĹ���[�N��1���^=��Hx "O�88#i��B���g�r���kg"O ���/1�\� F]����q"O8-�ma�.-#����^pz'"O<Eit��)9�*�R5�� v����"O-��B�E-���!�9=W�dx%"O��2��sB"�*�`:vL4���"O�1C��X?+�2$��NM�h�PH V"O� .��Ą��GGĹ��m� ���"Or\)7���K%h���*	"�޵�!"Od��lY�{�~�B��՟t�B�;r"Oܹ��G� V�0�UȂ�Px1c�"Of�����	L�֌K��M)M��і"O�!* �L7 ,*�8	ȺѫAM6D����J	ՠ�ʔ�׵8ܑ�qb)D����Ly� !���dhby���%D�(K@
Z!*G����8e��T�=D��v閖
�0%]!Mi�t�D�'D�X���8[3��K�ah|� %%D��r�˕9}�z��d�T?HT�׊%D�lqf��c���+��D�L��k1D�ĲE([X�N �OȜP�P1�J$D�aFꃊ]�Б*v�E%?��Re�"D�hE��	[�z�¢x�ňӋ"D�<
 �K�|��|kw���(J�i!D��y�h$�Q*�`J��&�$D�Th��I�
�mj�H�t5�6�#D��b�N�D�r�jgW=BGX�;g/D�P��U�qN�Yq����ZD<�!u�(D�l*���Z��Ab�hP ��2�&D�4Q2l��q��M0GEm8�1�R�$D�@��#�0ф�Y�¸Kj����"&D�p�˅3�Vt� ʞ9J�A��?D���@P�Fj��QE�+P�&$�� >D��#�R:+2��i�真!�.�[�i<D�@���:9�|�e�[4]kJ�[ti<D������0H�;�H�2I����B(D�x�1�=Z3�4eb�F6��Pp))D���!�y��p5B07c�T`3C'D��i�+	<e��	��
T�Bk�@��?D�8C�-�=Z�����W�G�8]t�>D���V�#����勾_���">D��� (1 ��lq&k�(yԜ8$O(D���Q�#�Π�$f�5r~�{�3D��+�(1��
2�	�
Z�[�+0D���S�[F.�J&+r�T@q�.D��KЎY�
�d�W�aO��K'�!D���w&vn�	G�W	:���iWE?D��a��uzj��O��z:�ܓ2L<D�lC��B�n��d�f�1V`�ʃ <D��re �+Mf�����S�髴�%D��[ ���P 2�S#H|��ɱ�6D�3��]7.��Cp��Rs��yb�ׇB��]+���W� x�B)�-�y�� �� �#��-��N��y�lɢX�<iCF 4����M"�y���K���ؓOӨj��p����ybH͙n��;�#h&H���ǁ�ybhA�P��4Iɂ1�"��PD+�y�J�0n� 1sԤұ�lDc�M@��y��&#�ޥ5��%��p'�C��y����6�~�em�������&��y��	V�b]xv)��AqU ��yb�Է?l:8�&�v6�4�	�y�EU�"�~�xb*�S�*,� ���y����m���Jc6�y��D��y�����"3"�;�B8�l�/�y�ƑYt�����O~A�xs�D��y�AޏExV��P����`���ػ�y�FM�T�VE�tI�P"���yR���������wP�=�v-خ�yR%�T(DQ�"N4Em 8&mч�y
� ����!��J�H���R,����"O�]�P	�E���s�G a?հ"O���H�7HA���(/<��Y��"O|�)M4H���q�
�W�6YR"O�3!o�)K"��Z�[�Z��<0�"Or���4*������"O�����P.� @�l��[s"OdH�GbL�\+��tn��&_��"OF�s3�� #\���.^'xQLh�"O��B̑*:�e����>I&m[%"O�ȑ�`�������q�D"OZ� �VTYF�H�T����2"OD��W��3�n ���	=t9>�"Of����A�c� ��S���D�W"O�uk���r�C�>� Z!"O
��fn �=9�M'�-�\A�"O���c�VA�L)>xY�"Oa�g��~ȡX�BK�V�칸q"Oҽr&�/nߞ\"2!JQ�e�"Or}�S�2N�x��/B�x{�"O`�:pHY>
8��
5�ڌo�H��%"O��+'Z�i)QK�
�0�Ӆ"O�l�pl����ِ�/
��䱓�"O tA��Z0�$���B�B`��j'"O���� Ţ&ШC���jP��"Of��o���н�C��(|�	�"O"ѣ��1<����ʇVl����"O�D����x�i�n��S8�1:�"O������N�M���J��|�e"O��BK
�U�g�x�԰@"O���C�Zʘ��Qi�+1[�L��"O���G,>8����獭g82�"O�ɸS-�4N��sf�ʲ�v�� "OT�*b��ywE������"O���ꋿ?C�8f*I |ԁ��"OH�����5[/&���N�In�3�"O����gh�3�aڸrU`�Qe"O�AB���wS��z�ω�[<l���"O|�т̟#(�,
'��"�<�6"OаZ��O!�H�h�픋hbֹy�"OL|�J�hnt��-|INa��"O���'=R��y�Mπ1=,�z�"O(ESG�-��/~#���"Op�p��5<���5�O�jtkQ"O\�ӣ/M�|bR���� �"Oz�3J8I!i%	�s��|Ð"O ʄ喋b���(i���T���"O$��,T�z������la�r�"O�q�s�&7fp��b��I`v�"O���O�S!���]3RHTAB"O�5s���m��s�`¯1��w"O�`;�^�Ux�@��7k�4x&"O6(b�+6.�� �&�99�@`��"OF<90:�~I�#�1t\02"Oޔ� ��p�*�ȥ�� Y���"O�[@ڿ;K����� d�+#"O� �B��I�Y�gwO�h�"OD�s.̵l�"�0q'A97D��:�"O��� ��"�P%i��)��E�"O�b���o�6�xP��b�ؙ�"O�H+1�Ƙ�����ǯX���+�"Ob�I�%�,d�饥�J�j � "O�����o��)ф�)]���"O�L��Nh�I��RT�I��5�y
� ��:�ً)>*���H��"O�yQH%/h�Y�!aә�
�)�"OZA�p�� �t) ���1P6����"O�=����}�V8�.�="�)�a"Oh��c	!�J�3��1: !��"O�):�L�&������
����"O��N#���y�'U��z�"O���ꗬ'D<�s��8���d"O��
�͕,Ae\�b򨁩4�ś�"O6�i��8"8ؘs�T�x�(D��"O�a�<M٢RE'Hrp$`�"O�Sf��7I�	��&F�%GtP!�"OX��Ǣ8Ci| ��P-3�|!"OB�a� ��RK@`:�Κ�K2N��7"O�%h0-��,hb�lR���0"OR�K����b�(ٹv,êi���3"O����LH�*A��Ҙ��"O*9�wOY$#�A�A�ݫj��8G"O$�ٳ�)1��eEM�4�0�b"O
��nG�gr.���91^�(�"OX���G����ID���"O�Z�K:+�-�ah�'N���v"O�Ig����$�IK&M���*a"O �b׻˒��b�g�B��b�<�a
ڤX�D�����	`�N`s�iK^�<	�J؛\mp�نȈ@��e�<&��%/,�A!֭�#8|c@k�<��h��)H �P��2�h�<�cg���u9��%`��Xw�a�<��MI� Z���!�ǡ3.���FZ\�<1R�Ҿǜ��Fm�P��Q!�l�<�% (p˶P*�i/�q�p�Pm�<�R�@�O>~)��̆+3��b��^�<1��l8��s,M-����'@�<ѕ'�m_H0��+6=2��Ł�q�<a���j�l2hQ&mo�eA hMp�<YBmY��Iy�b�"W<	1�Ru�<Y�)��E%����3&]r���+�j�<��LB�̌AI�=�\ �K[l�<�c*���#1��>�)��e�<�g�*�a[VKS�Bh<�����`�<ٲ�`���(Aɜ	�DL`�<����	?��(�T4����@)t!��ʜ,��O� ��x(ӀV.�!�Ė-� �S�LZ�|�>Yyq $<�!�D֙;�����A�F��7J�s�!�68��`ԉ�:'����4��*�!�P,Z�"0D�ob���Ԃ�+${!�$/U~�`�0N��YV�q�̗({!�Ѻ}�$�.݄[��LS��{e!��A�=��X��!��4)�	_�W�!��܀E�����M�I,���h�:0�!��\�2@*��j ��g�k�!�D	:Y��DU)������!�؃!���&��aWR}#�R)�!�I�fw�]��fI!0芥"DmA�D�!�dٺά�Y����Kg"˵V!��Z3Kv%�b��}�
p�2KM� 9!�$
(;xB`�����0��="!�@�4�h��%��"rhac��"z�!�d��}w�ma���0n�	{�F��!�$-a�t�
&'�lZ\ 2(�!��D��ԍ��R!w������<7�!�D�<��Y d(ۛ�D�@����!�� ��gG��V鞸1��<*����"O�8��GG=�ʑ0wA��Y\�Y"OR�2o��v��a;#��.I�R�`"OH99'1��-��V9P�Nhh"O(��C��ziZ|r�����R"OF��C���T�xT+a*'�>1�"O>���B͘%�Z��Q�E	��hu"Oj���D.PW����؇W�~��G"O�D၏�&�� #��{���'"O�i��p��y#����7aV""Ob1q��Q��������~I�"OR	���_oCu�@� �.9�"OD���4,���4�����Y�yRϜ:O��X�A�i� xe��e�<)�U�r�����G�3ν)�]v�<�Ѥ@�+(���a�~�0���W�<����u@`,j�^9�8͇ȓL�P@�B�L�p!hB��+L�	���.�����X���5B�D���ȓd�A�DDoN��1�R�/����ȓ#f�(" ����q�/H�7��ȓ��R%)DW�,D��*�4��Ն��"�(O�`],�P'R�8�t��ȓ$�FA8��&22L���m�{�����Lۢ�Ҧ,^ZNx����&/��F�Z Z���N�m`#��W�2d��s�(}�g��+zCLh8��k2XQ�����&F�:X����fEuN0�ȓ+�̹c_6Sn$�����5de�U�ȓ= J��D�~����O�/y��ȓcTX0GǞb̤��e�04	P��ȓ'���Q��W�`u�&�<yՆ����0AR�07����ߴ
����ȓb�,�����0V���4F�d��\T�Da��|��T��٬N�I��N����J |2��J�D��\��o0�-��Eз �<�񲦉Q ���ȓ@%`-9r��6e��ѠL+ l͇�y,ā��"?��� I�/-2y��F�~�Q�J͔��`�h��Նȓ�������7D���!AV$��ȓXCRĈ	Y���p�҉f� 9�ȓ(��I�1E�`�@�J��W)��o.fQq�'�qH$�r��E�֙����y"���/I:�2�h�<Gp�ȓ��,�$C�b{b5� hX�@E썅�#��=��$X� D��"-�&I=>��ȓ/�� !�Ů7|ꀓ@D��~����t4%@� )M��%S�|=��
�&��ѠA���VO�2nي0���6ljHC�-q�14 ��H�Ʌ�P𶬩��˲G%�xa�N�g�!����p�D�Em8 ��ӕ@���ȓm.�9a�X�}�@e
�;^"���UL��VKK�\�n�c��es-��,��|	���ߘM��		%R%�ȓ{Vz4[�+ƭ_�>ى����uv��ȓ�.�p �
4
ZTX)�gP�ao��ȓq�֨��|�x�o���e��(�I`�,
�*�Ř�M��.e�!�ȓxNLIQ�(�m$�`����}���aY��B-Glh1� *�_�Nԇȓ.�N�3B�ݠ*�:�q�˚_������Я,9Zl@��Zy8��[�"O� ��u��-`2!A��y4NE�g"Ob@���<�<0�J�zE�9Z�"O��{���W�`�V��P(P+�"O�I�@E�1�9B$�`#�A�Q"O��˵�fk���'\�0j�I�"O~�)��߬X*�(X2�C�n�Z��"O��жn].��jW�X��t�P�"O��:n�O���[�>tFE�B"OJ���\��V<S �F�{f�l7"On�*V���{�lsA
�X=Av"Oh����Vߦk2爻|��I(p"Oh�#�7G~���%�4wr s"O��� ��*:�8]�&jy�䂁"OV��f��9�0�-gfnu��"O� �nN'B���svk�rg���d"Ox<�5�E	4{HarlA'k
�)B"OV��`���&���JE0U�pa@"O���#s��UI"���S��"OʐCU#)B<@
B��G�QK"OHU�2b[����� �(9�Q�A"OTP)s�S:[@ʈ�� -xH�"O�Hj���$����*�G�l�1"O�T���$"�`s�FY5��,��"OjEeh]����Е�̬�6"O ����
�4�hl�E��trv�Q�"O�l���&O��j*�.`mey�"O��Q.��{;��H�~���a"Or4"��ю_FT�u��?~sl��"OXX;��I�0�n`�4�\�i>��F"O85�F1��%ۜI��P�"OB@J�zb�녃EE *Y�"O�q����P�ޘ� mף;�B!��"O(���9V'R��ʜEj��p"O��T�1V���Z7_�n��"O@��[� ���2HQ-'� ��"Op5�p��9g;&���Ч�0;�"O���bhG�Ό�.�J�� "O(C�K��N�����x"�jU"O.�!4fK> �b6!E:%m����"O�9��3y�:8
�=Cp��3"O��	��Nn����-b$�Y�"O��zu)!8��uxѦm���A%"Opcd�T/aM�	����,{ �1 �"O��QC�KY����j���a$"O��e�S��H�"!�8�h�"O1�F�%�F������� "O���c�ݩT�X�4�ղCn�h��"O���v�$j���5Gߎth@T)V"O��C hF�=ΔXZU��:Ȥ��"O� �+�cv
ԛDd��l�N1�W"O��C�k��S����Ec�L��\��"O�Ԓ��V�e��$ ��<4��\��"O||3��7fJ#%��7�H��"O���%�Wg�)��CM�- ��u"O�d��ǉ�`�&1A�!']-H�W"O��!��!e�(���`��@� "O���A#%~;��#"A�g�8��"O�@GlG�IH��(vnS{�^�"OY����2c�ְ���w��3�"O�壤�V��Fa���?M��<0"O�h��\4��c `�;AnXi�"O��9�j���8K��L�>�ܓ�"OX�"X0�j�Y�흭_.J��s"OlE���
'
�I5l�S/��4"O� ���̆9>��jY�)���31"O L�#H�&��Q1)ǭr�#"O�!�"�41,�U;�g�?xdRr%"O����'(C�1�&=��z""O�U�s匤ݠH�Cf_g�x�2"O��x͍%.dı����ݼ$3$"O��q� ��)m`XZ��Oښ�4"O"���*��0��5*�.ĳ�"O�u�&@���(B?%�Լ�@"OD�Qk��f���V�
��q"O^l��%�-D5"Sf҆��A�S"OR]��2uDfe	bWB�h�"O\���쀚J=�XkŦJ\s4�
�"O¹Q�B�	"����<���U"O���K�ten�R���LF�x��"O��y7A^(
�<�R$�"ٚ��`"Oȼ�d.4>.4�JDD���P��q"O�`�LU	o"XJ��~���a�"OH)�!^�G6�äd�!'n��@"O���� �:x;f�wsΡ(3"Oθp���F��� � �vUV��"O�![��?�(mz�b��O@
иv"O��GCݎ(�I�A�(�q�"O<�t*8V��q�� �`(D1�"O��*��Q�u���!U��y�Ř"O��
���U-R4 ���:�n�)�"O��w��� ����×,D�\�g"O�ͳf�I,eA���+�*2��{a"O�}H�*� "��Yf��x?�tv"O�����=4��Y��!1Y��"O�l8C�ׅG����ԩq��Eb"ONM�m�l���j
�s>��*r"OJx�#�^�� ��b��$hA"O2Q��	R z�2Ș�ȗ�~��1��"OƑ�3,^ta��5G�-wl���W"OX!���Ҏ~.��X��ײ8�A�1"O͑'��T{.䂗_*t���`U"OFYЁɅ�0��۶@"�&T��"O���43Z$��#�V�vY��"O���T�B�_Fq��r}�i�"O�m��ܦ�*WP
^B���"O����B,=M�8���^&��"On�`�G�U"����sJ$Yu"O�!�)��U�+�2V����#�\�<�e�'9}�թ �]8bM&����Dc�<a�N�]Ht�����/r��i��@H�<��D��<��\!Հ�"�F�貀@�<y`�R:q�}
��>$'ڤ�.�x�<Y3�şjR8{�iӹcb`2v�<��.��_� t�a�rtB�a��t�<�3	Q�9j�pS�$E�->����n�<�C�ƅb���Q�Y�{����"A�R�<Y�,D6c���8�)L9Q��xs(�C�<�r�+2���CӇ��Je.$K�̉d�<A�'�]�vi���4b�p�3�v�<��3Ln�#��܅%���K��o�<Q�K� gm$�u(�&bJ����k�<9�+V U���`TM�<'�xe��ʓs�<IfP�m����f�;d�"�{Um�<Q�
�.U)ƉY�!5"�9�L�e�<c�ߎm����u�J�RTÑAX\�<�6��G� �p�W?:�nt��e�r�<9�K?V�����G:co�H�*Sp�<�c� >���t�1��MQk�<� �U+%OȬ}���Cb���kH�"Ov-�կM�[A)g$̥(�AB�"OF�z�!�|��p�;1/jm"�"O��[s��2*�V!t�`5k �f�<ٕ!5�M
��Vi6��UKb�<!�нZu�ax���k��#�!Fr�<�w$H{��;ć�K:x���H�<ied��0���ćY�|��f$EG�<�E�BDӸ	i�'� b�Idg�F�<��%C�HKL����׋'|��9��E�<!p
�;��QJ�ȇ
!���p��\�<9v�շ�ha�eɔ/t �O[n�<�����~a	�/���kFEB�<QR.�=�(�Z!+1��I ��T�<	մ"(&%���}�scOE{�<1R�'b$�d
лR�;åu�<�q%	��&�sJ�Mwl,��dH\�<��ύ�$Xr�Q��nɲS�AY�<aP
�$A+����1.4}2s�y�<���Y�n�|�����J�n��@bM�<I��7.gT5A��J�6���tmBL�<�(�Ҁj�B :�Ȃ��R�<�"O�1"|֥8����Deֱ���W�<9f$��f�DK�g�+l������W�<ɇ���ɡ3�ʱ�����CP�<���9t�j�h �
�ּ�VODO�<�7ˉ��r��'D�<~4Y`�B�K�<y5��k! ��ZXY���\ �RԄ�B2����[���zUbE�6m�8�ȓ^T�LI�o��v���e� GH���	�!��.��퀲�
�^��:o�]����S��L�@_��D�ȓK�(z��M&&i4t�!�Fq��?$h�ae?M��a8�	9&���q�6���ᔆmR�T��
�&�Ҝ�ȓ&��<@A�٘`�֍�b��s0u�ȓP�)YRE?5R@1�W�ߔ4zp��g,N=��K�b�M�s�S6z���2��e��J�J���cI���ȓ?S�Q&߁I��xR��2N$��r�V�kVO ��"���Jg���'�Ji��>4~Z��a��7��B�Ƀq�T8�dX�Xt~��Ҙ~
RC�I�y��X��
?Apy)��܏>��C�I̰W���~�8��b#��TJB�%vɒ��QaY�j�����mN�C��ئ<�h�dܠ��kV�C�	�H,f��,��&�Af�\�<B䉆s#��c�	Yx���3�� <�C��#� U�bY�> ������*Z�C�	%`�Чi��Xހi���0u�C�	��<�H@ں'ސ���A �w��C�	�|�%T��%�4�	�˩nh�C�FV�\���*:q�#�ܻ6��C�	.q�ғ��)N5 #��'c�jC�	;/�P�&E[��0ݩd*�'B<B�	�M����WG� ���G�8B�ɩW��ٲ�K `���!���J�C�I+4z��f -;�(UQ6�ިv[�C䉍	�������P.aj��26JC��H������'EB�Zg��?�4C�	�,��qS�aԡ/���U��r��B�I�:3
5�uO	Hn<�s��L�`C�	!Q*�ȣ���[�d��G�Q�C�)� ���$�; :�X4A�U�`��'"O@�Q��%d�)"�+�5��"Oz�c��?o���1n܋S�j���"Or4����'N ��7��Y &"ODC0�+B"i9�`���Bܰ "Oؽ��Y����P��z@#"O��5$RN�P��˳Wĺus%"ON}�����#bܔ8�ȐU�:�A�"O��c�ٺG�\���_.�8 �"O��s%�Qꑳ�!��B��"O��r�0�g`H�$��I��"O�Ya�B:v���ߟ6���"Oz�u�1��3(�:K��Q�"O�*�+��A�ԃ�`�Ա2`"O�!�!Bw��M됇�Z�,�p�"OH�`ᖎ-�4����	O��"v"O����M�"(M��	a@I"O�@{u�N�����.����YR%9D��(Ʃ,���I�,�; +�M� 9D����`�7�,�0f炮%$�}��7D��!�Đ S1Jp#s� �Q���R��7D�첑��uBM����=�Td;�` D�d�j�c�e��k 6Z� `��*,D�t�Rg�?�)�(�%O���c�%D�(z��ϾnX֥��MA�+r��i��8D���$T(}����E�1g����7D�\a� G�7O4�ࢅ<5�0y�4D�[�됧���D��
����F�/D������3ob�I�W�	&s���bs�)D�(�p�Y�v��p!>rK����H=D�`���Hr����GR�^��#?D���o7w�P���
�k�>@���=D�x9�c�7�d�۶N��.��Hy�`0D��� ��)�a�G��:.Լ�`�/D�Ԋ''�
���:F���@Ȱx��*D�x{���2nT�I��gɋI�εCU�)D��y����Tz<�a�Ų1U��p�:D��uM�*<���(e��xZ�c:D���EF�f�$�S
ƫI\�ԋ`7D��ɁawN�	���Z��pyG D�t*@��Z�pxk���T;��=D��X�mDL�����C�O�T����9D�@��#�z����'��� ��-,D�p+��ʲ+���bA[�V��k�,D��0R�X��0�fNZ��li!AB(D����oG=D��M��pmN���*%D�xّF�=DH��2��49zn$D�X�sd� Rz|�Ǯ>��yi� D��Y��Z"U�T�91�P n�IA0I=D��°���6�T��p���
���!�.D��ɗ��~�]�ǵO�`͓� !D��[sOޥ2Ɍ����W�$	A?D�P�_�:V
x����)ڸ!#w*D�H�'�EϺ��B*�yh���A'D������=��=��#�T#r|���#D���ubL+	�\l�Տ[��nh���6D��RAN�.A�t0䎙!G#�4	�3D�(Bǭ�N���	�"�Tjh80D��(4H�%q�ډ� ϕ�Vf(��,D�l��AV�}�4�2+�����Jw�)D�d�����~` �Љ3��=�F)D��E��`L0�#H��z���
)D���B"��lXx�e�M��*�J�B%D��PLL�_��{�}9�l�Qg#D�� ���4mZ�K�A v]>s?T`k�"O�pqg�B�:lD0��5�꤈�"Ot��V	�[{Xh���<ƶ�p�"OR5{����1B�]�vn�-��C"O��k�j�$W�JSm�2[%�]�f"O}Q����0Ҩ�TKֆ=��"O���5$u( ��&,|R5"O8=�s��oǸq� P����"O���$���� �@,�"D�>�� "O�{v��Pt�A��G�d���*O���c��*`b �e�ESm$�c�'Y^��v��&E�W�J�J@p)��'DL �Wg<\a�"H�w��P��'zZQA��

+�e@Z�@<j�'_F�yծ3b6���C�F���'f5����z� V�55f��`qF>D����Mˈ�]r#eP�V�t��=D���Ɣ�y_x�ېE�wP&}��=D�ԐgoƸQ���3A@Jq'D�QwE0[���V�>��Jp�(D�xk�֭S�2�2�Cգ
�L- C%D�X� ʟ:9�d�ǏQ� ـ��@$D����A�2MT���9m|�#'	%D�����C�:� ��Y6�f8T*#D���ҭ�wި�Z3I�,J ��!D��%"�:fB� _�>��s��>D�XkQ)\/*����AǘiҬ�(� <D��[፿}��#`��0RdI��H5D�����5[1�1�A�6�J1JB7D�����3F.>�+�,�-�t%;�4D����.R�cl5�G��6&Y����M'D�8�v/
�sn��p�gݯ<z� �m%D�8ّ�6!7�	7����E>D���d#�I��`� ؀DQ�����;D�,+�hׂd������as�$�I;D�tk�mˮV0�� Õ�b}�5�S�#D��SNg��x��В~ל�(5	=D��*"�A�!JdfE,;h	�R�:D����&�<qz����=G8��fE:D�� 0����݁�ɗ�v^A�r�3D�,b����91���D��m���%1D�L ��|�!E����8y��.D�(�iT3a3,E�晚7Ǝ���.D�<���#A������
�e(	,D��	�h�$G��L���J7s- ����(D���a,M�z��3���a:�|�!�'D���@ͼ8�����'��c?��@��#D�L���,����G�\�J/D�����X�P� A�FiD�yz�9T,D� �@`��d8@�%)3s쨝�Q%*D���w�.H��F � G�,4	��#D��ɣK�8���Iݞ)�$�Aw�-D�c�Aڼm���x&OF���*D����,T_*��%�Z�+Ȱ	�ad;D�t@7N��53	W7˸`�f:D��Z�N]k����iV�	�L���+D�(��H���0k��u�0d3��5�ɧu��z��zy���6�14���Qe�7�yrC@�WQ�@bӇ%�T��"�ק�y�A�^�R������jy!����Mۈ��s�T�2A�շ#I�d��L��F�1�"O�Ց�(I�vϠ�����eQ���"O5H�@0Zˆ����ѭx�l���"O�88A%.��\�cE9}H��T"O� :�5�ˍ����CU�%�~��"OД��B�"%td{ҩL3-��1+VOJ�DFh?��d�>L����
# J!�D�M���2%oC�h8�ꆃ��(!��X�6��c���T
-�"ڵ)�!�DSW?�$"�Dɟ4�����"Ja|b�|�m�4V��!�"��r� ����yb��,��]���, _�0	R�L9��<Y��IU��Pf@uB�z�CGL!�D�!��1+���/	�j��fbշp8!��RQ�1[���v�ڝ2ע�!O!��koލW��-l�����!9!�����v-�h(���.+� f"O�MCCBV+�D1R� Pn�@�d+\OD�
�8<l����'|3 9��'���@� �4VZ�P���U�_�`�YS+D���N&*��p��JT�+1\ A&�(��e}��?ţ���u���b��th�5���,D�V�Z ���fj\�� �V�V!���p�|�ф�]�8.B�Sϊ�Jr�	P��(��y��b_��I�p��\��z�"O���7@�s>ag�#�XH��"O^�+���q���
�:$�&��"Of�1��v:��0�	8#Ǿ4P�OB�=E���y��d�H�,�c�� ��y��C����镄G��x�H�����hO����H!�ԐyP�,���a6��1HI!�䒐 :��[HS��9bMcG!�$إD8b��6��}�ܹՋ���Py2�D�1�e�����+ܩ�ҦS��y��;eLf!8���͆�Õ�Y�M�-O~�O?7M��;�]�� F5h@Wj�5!��F�1�x1(C�
�C�Ȑ�ђ3+!��̢Uꌸ"�ț6U�r1�"!�p�!��.U��#��K�X���£6՛�
O�!0eT)d$q�f��w�t�87"O(T#w*��4�ܔ�����F�7"O69rj	S�R0�!�/�0���"O�A�a�Ux�Q��Q�|����'4�d��Hxf�bpB���i\���"�O�K%��bf@X�%;����A�'+1O����
�,Z@���#��Q�P"O�I���K/�q�Ƀv�T���Ot����(���{�� �$8��n��<�t�p�"O��f��-8���͚>���v�'����O	8 f�W��|�'�P��*�c� �!nQ>[��	�'2�h!��^��M̭*Ș����$6<OT�Rg웭?^"�sgP�
8��S��B}B[���|R�<$���+s%��[�v]�41!�D�8&�����$��*ĔP`	�6n����HO�x�?9Rf �Zᢃ�T�`&�95&s�<-������z�ڠ��y0�Q�=�!E(�S�qT.�����
{�Ibi�Y��C�I�id�� ��v�����D>��B�	�k���c���3mА��)�B�	I��JT0iJd�8���Z�B䉹mR�[Ō�K�dD�>.C�=cmZ�)�*%�ΐ��m �B��/@�&�+�Ahlq!e��E����hO�>=�!��Q�� ��Ηq�I�a*D��8�ݫ�$T���ڵ���&D�Dɠ��:
�ŋ���v���<��哼W�@�ƚ!c. H�$&� (�*B�	�7R�	r�=����D	F��C�)� ��;�O�[
���A�;��D��OL���	���#�`]"8a4�[/kԑ�PE��'Y2v`�P�Va���.�KuC�yA�5Z��s(�%	DXH,��y2��:8\����<��e�T��y��D1������%������yמz��kV�\�"�F=��W�y�,z#��B���6!����U�y�@[�F��V�'�4�rM��hO\��),4AY�J<<�M*��8+�!�	)\y���	�dpu�V�L��!�D	Y��zs	G&uTN��G��5�!���#�L� �EC&P6ڴ8�+yH!�Z]���*e�T����b�D&}R�D~���ie�p)Ke�\��Z�7�� �1�'��<آ���\�Ȍ$iǗ@��4I����|G{���=�P�$,G�; $H2��=Y�!�D�"L!���ҥ�8C.!)�Ƌ"���G��H����[��<�	D##v� a�"O�4IѨ\�`4�a�X}(A"O@vkPjc��ȥᄎ&��Q�'P��<5��'jQ�Jah���=d�B�	FZ��)�(0W�Ή��

o�,B��/n\>�c�^�CP�Y�!�L7'����%�IOs���ٟ'�͛U�I7?��O|�=�}J�
��r��}���T6FA���O�������{�&��O`�`�����Tj�������'����ۻ��t���D4,����b�'.!��=fyD����tvp}�"�V@!��P�|�Bq��!��Q{�u���k,��(ON"|�g�߄'uXRL��j+�h�T��G�<�eǐ�C���a���,r��2+�A�<a�EۧR,�P����d�C�LY�' $�=�'g���1��8����֨�*&?����-�PYc��� ��:#��E���H<��O�r�'ܬp�B�0Yꨘ��``����'�85 U�:*3=5�C5 �$Θ'V�{��%m�� 덦-���!���ē�hO��^����I=�@C�&V�~y� #"O\���o�@�ࡩ�+�v( y�"O��pG�5��1�J<72A�24�|��+	�8s��Уn�Z�PK"D�p�g��39:�@� n
9q@�7�?D����nuX��&�� ��=��+�O�ʰ�
�I�
x���,.�@�"OD�����@��$jw,C+\#\���"Oy���Y�� ��G����"O���0o. ��� i�2�t3�"OI t��j2���f�L�Uv�e�'�ў�gm�
U��4�V����b�>D���.X�t��:b�_6j���;���<��}�����8*)��1�nP;w� ���hOq�|��'섓S�F��"mɴRz=���.�ŞL�h��d��~@�բ���6��x��hO?m��Ѫ��Y����3�n���/D��� oR�/1�$#����5h&�3D��H���5�"�TʲR�"��q�&D�XvGʳ$��У@�K+g0����8D�4�&�Q�8�ei�-F�&j�����)D��A^�MF��C`C L�\,ұE)D�\�Ճ(}�xh!�ᆄEH<ȱ�!D�L�����B�cP(6(K�ZrO*D����hɔu��	���`V�U�
<D�0r@΅'W� R@�15��=U;D�� >����]	��)���8�@IS "OR�R��k,��A&�T��$!m$D�|2��Xv������k�B��)D��kc�^/ �`Q���C�*}�2A(D�|��N�7(�:�1WN�/M��y[1l%D���q��(Ud��9�HCX�v���$D���B�(z�nit-�LF��$D�0������x�*Gr�O#D��i�ʁ�D�$��@Cd*� &�#D�| 6�Z�ZFh}�k*s�e��4D��0󂋪*���`�� #�ޤrp�/D�0�G�J�C<bLX���O	� a�.D� ��Yt�����D�FGPH�Ł,D�d����
L ^���A�Z�8�5�)D� ��h�0��(�+Ә|4$�{2�5D�D�jK�)e�)p�џpr�
�!D�ȈVGK��b��]�A2�A�׆+D����7$�h��O*B(��k=D����ĿSf���)J�1�� ��o0D�<Jbe,/�(e�R*�`����(D������ELr��7
Y2BsƨkS<D���b�U�G_&�J�j��2J���D�8D�\2� ��}�Z���D��H\�d2D�<Jd��q+�MrEG��a�30D�����}T�%y�!_7f��e�,D�P��g5n#�];f�4�B !ա*D� �$�	$&�N� �XT\
�M+D����$	�{����
)9��Pdg��SA'��Y���S���Jh��a�(�\T�#bOB�!y����^�V(Ԅȓ�}`%��6�MB�nʋ3�܄ȓj��(Cc�����8j��R��X�"OtM�F".0�i��m�*P��"O^�H�gH���!H��*i�)��"O�C�^t�)sQ'Q�C�`�I"O���qf�n݆�$�K�=�,cw"O�}��l�z�

``�Bꊌ8�"OV��1Љ��Y!F���{W"O�x8⏀#��Ԍ�
=h�p��"O�D!��i�r�r7L��<	�x���'D��#P�?ba�]�񯗛p�:�`��%D���@i֚��g�<������%D�,X4+҃h�J`jG����6D��q�M��7K�m� V3sĀ)G�7D�DP�'�x0A�X��'���ie0C�	�`��Pi�i�"�$��U���B�	�G� ��ҩE�o�m�L����C�	���$*4�R<���Oͷ0�B�� J���*7�T�4���sfN�)�B�I�5��(��"Ϧ���k�tB�<=���lS�b�$� �R4fRB��+O\��w�Mc�X�9�ˎ8`�C�	$M��J�7J[.��%�!*�B�	�9���j�I%6�uB�0F�B䉥K�� Y�B1 F.��1 ȦB��.	��� ��l �4�c	IޒB�)T���'J��%y!��	N��C�ɭ\hlU�c��;)ƀk�o��'C�C�Iv|<:q� ���C�Uq�C�$��=�`a����y�1��$8��C�	�p)�h
CA��il��C���!*�,B�I�<�~����9Sx�0�wH�8��B�I�(u�E�"N��J{�����%�xB��,(.=8�b�g_HlHq�`�B�I��̹pd�3��27��/8zB�)� >���0I}�J��׺Qd����"O�GdA5 (T�EG D�L�# "O�H�a[����i�0Pj��"O�hg� �Ψ���J8dW���"O�ۓ%z�邊 m�UJ�"O~|�p瑤Fc,�*釣^|�ѥ"O��5f<�� `�)��4���;"Ov۷�1"Ȅ�����B����e"O�MZAG�o����?o��K�"Od0a�խV8�H��ҤKr�QX�"O�����7�8��se�!t��`"O�M��ň�K_ �8E#Ⱥw��@�"Oz]�U$΅ZQ<����m���5"O�Q,/;�Yj�	�VQ��"O�]s��:�r����S�_��]��"O���q# �V:�Å��/�F�92"O� �PC�9Uܥ)��mTlx�"O��tk��1�f�&A"EI2"O͡2GЫ<�yq��9~��myt"O�Y�+CM%�)Qь^2d<-ñ"O��2�K�M/�xx��XͶl;"O� ����W-�U*F�b��,�7"O�P�AoI$o�����o��y��ֽq�H`�w  �2�\�� ��y­ҟ(+�l����,F4T"�.���y"�� uF���IMh[XȣR�O3�y�6eE�y� ��l!Na"��J��yBi�6w��aG�:vV����
��y�꘎k����ҧ�m��pe�'�y������3J!1M���U�P:�y��#Z�8�k�� т�r�*��ybD�p�d�����6���Ѯ��yR���q�(��ۦ3l-�6�:�y�!�=:�bŻ�%�!
��RU�6�y��(&R��/Y�B�ݔ�y��؅,�pa�#��<�,9�-Ќ�yR��>yL:��ŵK_��"B!W�y򌋰Q<�QE�?隱"S�Z��y����'����P㑟>��qk���y�
��6�&<)�[�0� q���(O��=�Of��1`"�j�5yrn
f<�h��'Ϩ��t�*TVP�R g'���̊;�(O?���=�@Er2$��5Y:����O5
!��X��u'/
\h!p#�&h�l�,�D�5�g~�B�=��襉ϐ	n~�NR�ʐx"�V�F����V�\v�աQ,�2 %XŋD	��?A���PlxiDki�xh� �Mb8�H��E�/�}&�Xp&-�;)�θ�!f@��2T��F D�4%�ǧJ#�%���_�z����r����t)ķ���s�Oހ}9��s�Rex5�E�(  @�M:�j��"O���y^l�H�jӖ`���"���ᦽ���Xa�b��<Yo��3�"�pH�,bd��b�C61�H��ɨ+�>hc�� � Xa��`^�}@�%1U��`SK�<f�)��'͈y�TNUA����Ȍ9�h�;�}"#��$�a�WR���oQ�#2�\��SbX�=xfbĂZtZ�����l��I�%Q�~��ą;2<!)0΀';��E"%�_EB��s��R�O38)���e�+7 ���HY�"����Y�g� ��q�M�_�4e!�إ{��A�O���X��+҄�U���$��=�nU2�o�1,��0�tI�Y��y�/R�-��$���Z�5�(E�2�9Ӣ$9Lpɋ����0�\8S���,HƔ��I���CeR��N�D⑟]���OL�	bў^�����oN=\6�Ap.�C �ѭ��B%�R YB�`b��+n~�:�"O��Xv��W��P�w� U� ��Ϛf:d0u�H'x^p`8ňZ���PN~r�X��.J�dS�'Q>J2���O3�!�DA�? ��s�n�v�X�i"� Mr�LC�/Y?g�<� '���#(.)���6`���[��ӊ�(OP��(�\�J���Q}���Q�'�R�����+����Q��(s���3
2X����6���k 舻Uت9�~=���
8n��|�
\(6�BM!T#}T���
F���'����L�kfS�/�~�+"o�� X���OQ:i��d��6�����ޓ.�#�'V����(4<��i���hq���>$�P�*C�@������-R��'?!��!�&�yG�S>B��E���Z�8��x�N���x��P$&,�H���4��l_�[%�Ir�� e�p�{��R��	��b[�$"HV�I��0�v�-�2]�PF\�vW.��N?X)�y���:�d��bÞ@�ht���W&)ĵA�	�L��Pt�G�{�rq��<�O �+�W������g�I�8]�q�xrAυ(��m����x�>���C��P�R�&
1�i���l|I�&�Y�T"-� R!����J��s鉑i�΍��ȟS�}���+8��,�6H�Lc��9�@��Ik��	�0��8���l��a��(*[n$P�Oʤ�'�W.� ���aM�`Θ����z��oӛ\΄(�FM~B���gא-�2�<�v�C8H��2T+�`��dyf�qX��U(��B�R���g��@`G��	L�d�rn��R��2_����4�	-���6hG@)6��*[|P���#C10O��@Q3D�r@����*`��q��E�	�1kD�?�"��F��3�&� `/z�2W�"D����J�<R1�.¨^,*�C Zn�D���Q�W�6���a�!�4����$�� #�2�](a�	�0"˷s��x���\=K�tC�	�'��.[����W�١u�Z1@2@љl�^����ެx��='I��&��v鉠��QAw%��O�J-� ��=/����N�B=�`A �(����i�ʀ��֖�<)9�f��s�ͨf�=�neA�#��u�^)\J� >%F@�<A#��>!LT�P"��R 䝡�A��6��)�V!�W�_8_?`��"G��$J
P�""O4M��3}Bh��G�%�zk5+ӥKeD%���yH����V�Q>{;O���P���(:�Z���'�xQ��"O���P�5wwr v�]%��,�4/��\k7��c2�A��	ȣK��"�w��@P��<m��h���+?��[g0�	���'�xj�� �r���1%�mnj�۳��&�4M��,zE��llh����$�Th��
�@ݢ�`���#�E� �E'H����E���!�O�\�i"�t�3��(I�,� �b�[C('�����]�B���Ox�+��	DB]z�%�;����i��t�ȨJm�@J`W�"~n��Cศ�c�9""B�3ϭYZ�㞈�5�.�a�TMǘ8�b�sj�8	Ֆe���Q��y��$��~��ՉNE :X�����Gܓ �X�|�'� �Q�l+[���r��0?%���'H�X�V��6#�j�)�zU �d̄m2�q�sle� �ZB"*�����7�n���;]�	�O�����Y5~����s�Ȱ�"Ov%�G�X�+� A����$;1"O\0�-"�"�`���HJ�2�"O�T��ɖ+O��$R��M�_:���e"O�iдB��-�%KOT�|,8���"OFl�th*�8X94A�e?np��"O�,�G�V8~8.!���T�|�к�"O���GB����sC^������"O���2jT�(u�,�CX�g�\�07"O���QN�dU�!P�'���"Oָp'M�A��4i���q�<1�v"O����J�E-t��e�.\�1x"O>�9��^Q8�rË6t��Y��"O
pA5��t2�
DIY^t�ɕ"Oi��@V���	Yđ�T"O M�%.X�(:h�;�ѢjQ�L��"OPt��e[2��R�EM�?�| �T"O�p��I��P��-c `�%��"O$رRn(y	�˧E�^�V"OFxŏ]�m����֨erT��D"Ox�"���"���c�L"-T��hp"O�(	�ė;?GxxA7#�D�3c"O���[�ƅmNTkb�e!�d��Hcv�`q��L�<)a��کNW!�� V�0�ct�(��ɿ3���D"O:p)���8r�Q�«Ãk����t"O`d1҄	F�����2�R�"O��"Ʈ�0i�%��NT���`�"OԑrQ��.i�@���J�ܼ���"Oluȡ�_�B���84냹S�ʄ�f"Ox\�e��4,~�1�,%��bg"O���C�Q�"�
�nwr��"O�Z!�Pa�	�� )`�l�'"O�S�gZ<N(H��L�M��x�"O���,M���4��:JKl=y�"O��8�FF�S����/N"��KW"O�A��¸Y�����Oˑ\�&�A�"O��a3���\Hp�.�%)�\��"O �&FJ�d���(����4"OHɘ��\Ƃ �⬖�-� �q�"O4�w�]�t�'+�<1�j-��"O 
��68(rT� (iL�<)"O��%hW�x�|�sDd�+l>�!q�"O��sk�VBA��Ԉ~+p�q�"OkgLT�}k�" 
B�-��"O��W�ڑ �����&��3�"OZ=`��թ9F��#B�8GTұ""O�I�d"Ԯ'��)�&�-`کCB"OtibX(r�f�� ʉdƅ�7 !��Yd�{�&/<g�e��%6)!�d̊T���uT\���k#!���fl4�Q��р+a`4���+X !���kh��R��Ũx6�9�$��!��UmU����Rz�T"�7Z�!�D��p�XlǮU�s5,*6�T�E�!��H�p_�I�$�/]�l�ҥ�L��!�dQ..� �J`�\�|��N��i�!�d�+Q������5�\L�D����!��d�P���;�V�@����!�!�$TfV�h�&�ŖI@�b�*T#!��Xm�ɉD�ȵq��F�2�!�$\/N��ZЉ<�y�o�}�!��]�,�)��t�,�J��y�!�$�Q�X��KD�C�X5�2v�!�d�*���O�3 ��1V�KcX!�$_1!��I��F^Q�0�Ä7*_!��I�*Q�D�	Ig
�)���<	8!�$�b�H03�Ψ[���T�%p!�d��nA�旖:9xA����>�!�H/*����2(�3�1c��6-�!�ā/,;F<��"S�?�����;�!��=e�����" ��³�U�!�$�)J�$! ����O8l�!�D¶On"�
U�]!'Ժ��V2KT!�D�F��<����%ɴ+�	ZE!�\�02rL� H�2q���"��A<*N!�$՝M�V���*=q�����$X�!�;uu4	:P�X�� :�ԟd�!����X�qcGd� x���!򄚲6;8p;��D:;�)Y��#|�!��5'��EcTo��N�`��KH6�!���7��q�P��<�QS�H+a<!�dS'�ndsC��5 �â��%!�Ge
D[�甙I�<�hE��=C!�Z+}����%*F����ZBJ�,k>!�d��=�Px��Φf�����ם}!�$�V� !���v�$m�e���Na!�D�af-GB�3�X��v���Yn!�� j�����2�LY���UV�:T*OPa*s��[o6�����/L`�y
�'�@kΟ�
x�lHF#L�N�{	�'��[G�=�,Y�(�,Z�83�']�5�A �'9+%����
�'���s�̒ l4 5z�g��LӒlc	�'��H:@�Q(eВ(z%cд�p���'�T�U�X�OQR\�W�
�h�̉�'��x�(\+�p��P�� Y��p�'�4{�G��@�b���c�Q��u�	�'�ޡ�ECį:Ct�1��ܰS��|)�'�d��K��L����!�{��Ш�'�ڰ��Kˑo�I� V�{n��Z�'�̉�TNˢ
FR�£I<9����'.$ QON�m�D4�wIOg4e#�'�@��%�#��Ҥ$�)B6��	�'�v�*���u� (Ӆp�.:�'y�i�C��1����f�? ��'�&e(1 �{;��P�َ4v� z�'_$�B�e�6�窓�,
ps�'���f�D�S���mF%�	s�'�V���M�,��Y�l�8 $�i�'��Pr2���^���G� � k	�'�DJ��k�廁`�qi����'͒�P�+���������y� �
�'���S�J��&��
�q ͘�'Ѐ�iH�~�N����D����'5ƹ�2���W׌�#a��)c(�d�'��)#�I�\,bA��EOZ�ht�'h��Ѓ�F+C�Ԕ��kď@�^a*�'i4}�U���Wx���ᒼ<�2Y�
�'��$��#R(u�4C��Q�1��5��'S|�;�����l��?3��)9�'Ҵ�-T���e�9�n�Ⴁ�<�y�+��Yk 0�E��&;�����;�y�eؙ5���;QTE
���/F��yZiH��35k�k]��0o��NddC��:c8��𭇔��1���I�"C�I�21"(2�Y/iaxDp�#���C�	r�`���T;o�`�2��5{�B�	h��(�©ݡ#�DX
snR�H2B��7'���JA�H�v5���z�B�ɸ(U����%Q����l�*�JC�IZdN�Ɖǜ`�����S�VC�I�>L��]�W-����/Zq@C䉪ZrDdxtN[��C���V�jB�I%n�A�Lq̰}�0,H�#��B�	$��Q:ЬԬM���IT�Miv�H�?9M[�����-s�@��N�O�|����6T!񄜡	%h-�P�?'��R.�X� b��arꞭ7+����Ö�z�0 �1����p<�_^��E�H<ـ؜��1���W,H�Z���	N�<�R�VT�r��q@׮SJ0�2F�|��@�X��\j6���Ƽ]i��b�+�_���I��k�!�H0V8��H��1s��L
S��;q҆'�\2�MJ�t�q��'������VZ$i��YB��	�'�Xq���Z�{�,���%�e���N'<��i���'���ˋ;b�*%��%��H~ܴ9	�-�%�$̇���v|Z%ˎ}F|��V!E��q���@-C���o��K��t��P�OX�c'��:��O��|�eݚM�F��v �XpT�["O(�$cQ�G��� b�R$:�l�bA�ɤ8x�D@R��|��ԐtIvQ��)�3L��tl7��xDݒ,6���CS�;�,�Ѵ�ҜD�9��Ͱ?� y�6䓊<�>lr��ęo$D}�&�'0�xe�|,[i �r抓�Ql$�Sn��y⌎�0L8��@gʋx�I��aZ��y"h���i��$��b�*07�ϡ�y�+J��Q�˖��� f���y��C ��p��
|�^e[����yr陒w58�Pqc	5w�H@v�V)�y�ɖ:���vF_�lj�mq�C�%�y���q��	]3\�	�����y⤃�g����"F��I��}�fK���y�&�-iI��bsǊ�}Dh�l��y���3�|Ua�f��pW��Z�I+�y�����	����`�#�E��y�C���d���#!�񴣙��yBc#\i($Ä�,{��1�7���y��b���,���B�������yB�ȧ9��p` ��M
�#��y���a�l�"%Я�:�*�@��yB��51�x����
�������(�y�G�V)@)Ң�USX���=�y"돰pc0ƪ�R4�y1+��y�HT�	�Z�(���xL\���̄�y�+�@8�9XCaJ s�UhT���y$��(�"PI�v�X n ��yb�6w�4���m�gN��7F^��ybd�_���a.���{����y�/:}y{�%����X�a!�y򤝂r+��P�)�$���k�1�y�@��!��|07��+�����P�yHj-L�s2��&$��0�/��yBkO?HX�EI��a�%�͓�y¢_Z�T	�oΉb^�Un	��y�γQ�T9KtA?y�Ő!E��ybN��	�@ ��:)XZK ���y��^��\r`an�	]Հ�ȓ!RJH�aA�_e�0ѧo�R���n��� N �Xu;F�޶z%8��!�+�^�p���3l����ȓ�X=Q� ��,
%Qn^�B�*I��M���\��x���y����.�n�<)ro��"f8���T�zdv)�/�^�<���_�s�|H�q�ޟ%i�mgVS�<��/-01<�����d��;�eMO�<���,g=���4�I�u�ܓֈF�<	GD\�aS����8L�r��~�<�$O=5�p:A�ި(���:w�@@�<A�h��th6����T&;����Qi�<R���{R�*V��d�l�XB�d�<	�hS�4x8��T�|/x�0f�O�<��j7R	�x��#�Qu�H�J\�<���A�gP�ڕ,ҊS��\�<��*���dA���)��hp�I�`�<q 
�X�iF�ܬ2��T�CX]�<q��E�,e4<��g����G�]�<�S���z]�u�?w)�(V��B�<����

lK9qp�i{�BD	#��C��+-�r�cY�`Ȥ�x��,5��C�I#q؆��KA�DȢ0�G�\q�B�	8)`-23lǷ�(�3F@���B䉯oG�����r��١�mު9�C�;,���f�Ƭ>���I"�];LVC�	�-r�` �"v���'�2;B�ɩW=<\5�Q,涉�g�F$A�C� &(z����% ���z&�;G
|B�)� ����x4�BdLY�+R(��"O��0"��2l�Pj�<�E�"O�Y�@e�;���H�;�-(�"Oʽ�BJaJ@�h�ڋ,��=!�"O0u�d*O!h�,q�Q�	0��:�"O�H��%C7�e���'c҆)��"O�����$ =������oӒ�"O�ij�Aez��㏁-=xD�R"Oj5�T�n�@eq0�͞jA�[�"O>ar���wE�<1P�i>��p"O�1[v̟�aJ�#���A���C�"O��S��,Qܒي�� 5kD��3"OR�9uL�z�ԣ.�3�&��'"O�i�2�ˍ)�0őb�DQ�2�ʲ"O@��G�Q/^^ұ	���:���"O)���8%����S��r�V)8�"O�5��CX�mI(�@�%�%��ЙE"O�c�MX�!��y�� �(Ѹ(r�"O���ح�	B�ϒ'���2�"O����9^2 ;����&!�9�R"Oʔ�"��� bF�%�	�F��v"O*x���8�@�Ye���YQ8�8A"O�SnB*=�8�c0*�}�����"O���� v���W�A�=�j���"O��a
\4(�k�FV�b�$0�"O)i��ӫ@C`�[UD:O`>��"O��	Vb��M�
����ھ[S�l��"ON�:�JTm��#��(?��$��"O~���@7/�X �W��I��kb"O
�x���
9��"��9?�i�A"O��;"ᙣ]�J�9��n�b�QP"O�*�-�{y2ԂDO	@���r"O��[	E����Q�D�C�ɡ "Op9��HŘx3�-� zIn�;�"O�����N|m�i�d�L�20��"OЕQ%��/Lf���LK^�2�u6O`Ĳ�����X���B;Vi̩)��O��V催M�1O�("���k�X��]�V��B�����ڦ&	�&z3��X�7���h$Q����S6@�52��8 D��01ǎ,���x�^M�'��c>ik�`M�vnМC�Aެod�)"ri�>y[��<�{�'k�U:��� #X�)�N��z<PK�4J&��"~�dbբoZ�Ul��U���a���eўD��>w�Ȩ�U4��Y�KƦp��#<ь��?�:��<l�<z@ɕq��}0�N?񤒫�(O���I�Q��<wR%�&ɒ�U��3_�䰃�)ҧ[j0p�C����B�q�20
j�oZ�.~Q�"ZB�^�<�~��P!W��-9�@ �(O ��ӌe{b�ۅ'qМ���̏=�M�K�����?��󧖸�M�C�Q�
0[ƃ�Q���1#l�I��Q�b?u���52z�rD��#(XXz҅�>���7�S�OAtA�ː�+,,�ӥ�ĊV��#ٴh z�<E��˨w�-(C��![L��� ,��:�Q�l�çf���0�G��r]����0�n��>	����DV�E'��y�A�v���g��+��=��y�IX.`����գ�9T�e&Gރ��7ړ^<�O(h2���/*j�[�'��]_��t�'	�#=E�t$KR~䑲�T\�{�L]eX*Ey��"�'�����6�,���"���-���'y�xGyJ|�b.V�*�bp���3�J��6��I�	o8�D��kJ^:4S�Řq9�-��N���'8�)��n&�iO
1��4�zI9�%�Y��4b�ٱ�tu��^�<���4Z�d��jP�.j������Z�<q�曨�|4s�\*`�l�@ ��Z�<��_��e	�H��=K<0�bW�<� J@I���-ˎ� #JT�4�d06"O$0KҎ��(W�ѺQ�Σ8��Q;"OF)A�'�*W����*�C��u۶"O`�C%P��.E�7j�`~8x�"O�IRA�Kl������ !.����"O"��"�G3lj	��@͟]�2�I�"O X
j�<&Lt�A�p��dз"OY���<��p;S�˟$��t��"O�lZـ9-�q�W�Htm]�"O��Q�i� G~l �ϛ���h�"OƱ�Wc	�z�r={����Iu�A�"Ox�i(SFڭIU�lt��"O�3��K�\�A�Ư4j�9�"O��ؗ�(n���Xc�H\�@� "O�iB��lh��0���`N�E��"O"��g��7�d����r��ea�"O��"@�i�|�䭈*���i�"O C`"�8u����тl�,�&"Ofy�q�C~�ӡ�lg����"O��5%��A�Ұ3a�Pcn(�6"O��;犇,w�����x�#��-�y���Y�tآPZ#w�,�Y�h���y�ѵX�Չ���4YW Xy�*هȓad8�S�{�HrÞ�k,؇��RsG�?/SL0�5�cCppR�'�2 *�;OXء{�k����;�'�V���Ҩr-z�FE�"�H���'B8�s���.��`r���E�@��'H\`b�ȒC��%1&@'1
�0�'��Њ'�׆;�^�H%��)(� �'���#у[�@9�3���N���'����vEGRع
t������'��(%H�6�0��JW����'�؀Z�M)P�>{C��o�Y��'����>���LP!Vi�M!�'Nb5�o�Y�s� ��Pbp"Obݪ�ʋ)F���� y�aR�"OR�$�Aef�R���Lv(�R"Oh]0���vՌ*���z6�a"Oҵ(��ܾ#��i�([>v�pȠC"O����<$�y��M�US�1�5"O�X6G���t��0M N�T�"O�!���4VG��LFn�;R"O<�eEً\��\�'�%�y!F"O2�`F&!��X���>9�v�#�"OT|�V��T�l9R���0� "Of-�L��8d��b-�NnP�"O���2]u4 ���Xw�r�y�"O٪������3#[��u"Op�����Y�H_z`�z""O��R"��
�6ui؅QJ4ͪv"O�L�6�CP�b�
�l�X���"O���C�Y
�<�Q(@a�X�!0"O0�p!a�9T�|�!�&o)��"O�9��i̻;�i��9D �W"O�� d F�u�z�@ce݁Q����"Op�1�
ދj
�Ȃ!eB`���Q�"O1��&�	*)d�#��^τ��"Of��2��E�Lۇ�K��܋f"On�0j�$Crq˲юQ�mR"O����J��<c����JJW6�E"O��a"嗇� <�׊�$lД	e"OJyz˅��M�pKB�x�"O~U᥍�D��"Qk��!f���"O� �@[ƅ�rn���k��^�af"O]�f$��&���KãV�>�1�"O �A$`���ᶫ\|����"O�P�$��.*�l$iI�L�@�"O� B��O���F��U4�H�"O�D�C��\Rr�r�0�!�"O^ �C��1{G���Ӊ��<�18�"O�e�Ye�����W:(5Е�/T�1��;�L�j��NX���i��)D��	�XQp�Yd�f��|��&D�I��}�ҥ@bL_P�jD�0�%D����`��O0@x
��P�,X�r�(D�,�C�M�:��,��zY�9p��)D�d�� ��=�\�2ڰ7)��5D�`y��ȹ�8��d�V�\�ERSD7D��3F�Jrl3�wtN�*��6D�Ё@'r�n]�7eC�-o�*Q�4D�	ӥ��5�,x�g�S"(M�)�i>D���n��B��D�'��>��R$�&D��I��4C�d�kPQ�T�~�R��2D�$YD$�:\C�-�F
�豫*D��h�
�Y���	X?�
���
�'�쫁O�1{~�5�J� v�Tc
�'�<)r7�0G�Xt�E�Y�E���"
�'Q`Qs�d���< ��JR�=�:H�	�'3|�h�JYش��@��a��9�'��tcv�P�V[[��ޤ`6N�H�'q.��NI�W�4$[�ْ'+���'C���3T�ne�e�H�M���	�'PV�3�DβS=���Fn�C	�'�(���' ��
I�ƃ3T���'L�����4	�X��'� ���j�'���s��F�#W�Lq�̉%�P��	�'i��;�DM3��ل�'�Z��	�'� �S�I	kDt��)J',�(�K	�'Rhu6�V	��Dj��G)8@�L��'�R�����Z�¬�3�X�(��`	�'G�t`�K�8�Z,1���s�0X�'�T��G�0*<\�����'ºE�]�9{�M��Gh �
�'&��ᄥ���e`��� <@p�'J`,���m����"���'KrXL�<Yp�#%D����a՘�y"J�1h5���W�R�?0��֎��y�雅v��5	��f}�Q�e���y2Me݆�b��V�y�Q�� �y��z΀�@�­@RX��u�U��y��U�g��Y�S���3�� �#ݽ�yr�qH~�c ۱*���v'��y��
!A�y�s�&��ڒ�,�y�
��v���2�Ť~�ت��߶�yBM	���i�H�!,�Z割�[�ybi�n������EvL��E��y�����XW��
]����yR�ۢ�d��,��T�-G%���y�葆)	�q��"5�!Rv+���y�,g���[�O�m|���ȇ��y�F++}�Ax@�V�`f|����ߟ�y"�E"�T���_)p�\��A#���y�,Q��X�5a���y�g7�y	6lvFe�$�[=	�BzP ��y��лZ�HK0$�36X���N �y¤�!> p1	�n���,�Гa]�yR+=P�i��Jv���3���y
� ���a*�.Fr��a��0ih�!	1"O����*]�"��C�͇�+QbAB�"O>�:P����a�,�RJč�F"O�����Ďɜ��2��/w��P�b"O�!1Ŭ޲���g�pτ` 6"O��S�B��l�t�0q,�L�RM�C"O���(Cd�
m�&��$w<((�"OF�PrN��e��1���`g���c"O0p��Y�-��X��ꃈ}L@�:�"O ��"�#D��R
��GZ�i "OR���;.K�S�S&C���s"O�81c[9$ڼj��R!?��t7"O
�(UFFL��t�&��B|(�"OL����(A	fg˱s���q�"O� B�*�I�K�/�c�I�"O��c�"̔������^�U�$�f"OH<b�n���2x���?`�
5"O\�Pe�$ (��"gn	^Kd�0"O��{@���$��!J�I,���"O�=5�5O�Ti�@�:8>EJ%"OH�&F��
��������e�����"O:�෈�w���i �ʢ��m`�'���"a��p:ڼc2b�#s)ve{�';��S��^"Ӵ:�t�'��x�,��}Ǝ�±L�5f� �'�>\1��ڼb��с��}� �'�4)вi�:w5�m�WK�6n��HJ�'�V�"BX)���$�X�D-��':ܱX�"Y�*�pBWG��K��]y�'I��UA�}F�s��<O���
�'�b��&�A�rɠө�F~��
�'���ዄ ��r�N�?��q
�'/��s1�ɵk
,�Qb��b!)
�'F����H�tT�L�&i���T\k
�'��J�څ,ݾ���>dn(h��',�ؑs�#Tlȃ b;�p�'���a�ѓI�`xa5�?^j�`��'��ygd�& 7��؁+S<(�|�
�'(<�xDM%�|8q)�h{�Z�'��d��.yk^���G��^ް���'M��3��M7E��b܊ -<�(�'���x�b^�E��]�P�y@
�'��hB�	!�ؙ1D]�nM��'��!X�`���TU?U5b��'��1�A�Q:v$�(��Iœ:����'��	�3!��bat׿'�Fl�
�'���׭B��8�� �"K�Vm�
�'�V0"2�W�l�f�	�a�G"lDr
�'$E�P�.��lC�A�<qn�ʓnAf��K�B�l���.��ܱ�ȓI2(��!K�F��=��Å5�.Ն�k>\	���I�rJ|��ۥ|�Ru��cX��p��.6=N�b�U��ȓb9bl8$�ɹ;[L%c�݃p��Ѕȓ,�Q���@��3S�4�^�ȓ^!�l��!$�bHY�������'4õ�n���f�Īk`N9��D
^��u`�I����aT����M���ks��8]�T�Q,4"ɤ1�ȓ�����mP�v�ء0�jEՎh��J�X�C��2�Qh0+=�h���y]��#���&O�B��J
%N����V��Wi�"����m��b2M��;YR�R�m8Hʴ��3�:Ml̆�S�? �H`$
!��E�]x��cq"O$�&   ��   9  �  3  �  D+  b7  TC  lO  �[  �d  >o  �v  }  [�  ��  �  *�  m�  ��  ��  7�  y�  �  ��   �  n�  ��  ��  @�  ��  ��  !�  ��   B � � � %% m+ a/  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�?����~��璹W�䑰L|�� *�S�<�g�Q9 \��!+F!F����SřL�<!���d hxc�ϖ(��h�K��<Y&�7f�O���R'&�����X�{s<e��650B�	�S�QA���1 �\ ���-E�O��>YM>�&��8�P�S#%W�{x�Yz�<��N܀�1�j��r�Q��bN`�G{��Ox�I%������U��$@M�0�OH�����n�@>]�t��"�08pa��1 ����9D��pH��d}�t�C�&>��k@"�Ą^�'�1O��;�f�}�ZC�"n�h���B؟��	�z����h[.�h�6Z�]����O��(��|Bd�	�ܕs�m�0.xx��� \"��O�#~�`ʻh�&�öO�={�N9VnEv�<��H�-�ʉ��^b�8#d��u�<��L�0~6�k%��sT��%�y��d2��[4�Q�s� 8\Ȣ,�fo�(`���T ��> N,:4'�ц4��}����A"7�T5F���]��^�N���
�m�>i�c��|�n���Ϧ��Y�<���!z'`H�bj$h�`%}R�'���2���H��``��]�z{$���� ��i���{���%�5x���"O�T)u޳Q�ʝs�O>p������'[�'�^�I&�0*&�ӗ˹C�"	;	�'Ih}q�&ԃ�D��✽CU����d���O���q���RE�ȉ��	T!U H0r��';��Kѫ�|ˬ���3S<� ���V<��'�����O��:cΑ�f�yB�j�\�*��x�
�O�c�b?��Q�16R�ː	�/ZA��Sa�v�����|&�&
��8S��1�n�d(���'��zQm�*-��c� ~�lp�ի�y��'��X�`��- �:W��$2���'�E��'x>�w�&���p`@�kv$sK:�O�7'?q��5k����  B���s�Q1w�jY��H�)#ɧ����CB����
��~�̵Zc!F��hO������E#��
 cۊ;��q:��['x��	�U��	�q��E)eeE���cP�ɗ?�@�'�Q��'��H����dŨa����lO�0?q+O���į@$���cJ[�K�́ʡ"OXYQ�*�"1 RqU	��p� x����Z>Ғ��2k�yyR,�$ �q�
7D��C��G}1.\�lz��ђ�E�O:�=E��ܤ�A�y���a�܂S��B�ɞ-��X��z�(2f��7nn���Ķ<�Ot�"��K��Y�$�L����"O�@���S�F�� ��E=!���"O����	>�������)HK*$� "O���]�@� �
P��
p����I'���'e^�S�`�ƮC�C�Ɍ�4��G�2�Ĭ��G�_>�C�	�@��IҍB���d����-C���=�
ç_���8���=1.9��L�7p�-�ȓ�����L��I�Q���A�U�ȓ<��JQ�ϝK�4������*�ȓdشP���Q-�A#��>'��E��_�(���E���`��7z.����I����*r=ĬkW�@f�6�$[ PC䉑/�H��p�� X9)GNp�Ң=	W�S���|;�l_	B�XրL�.�B�ɲ�� 	��̞`�D���4X)�C䉅<�(�y5��P2��g�G�x�C䉸Us�y�(�}X-�X��B�I#o;+���G+ʅ��͏*zXe(�'v±�c�����g��R6&�C
�'-2�I��kr�ss�W���1�'N&����^�e�:4К
�'r�9�6IF�/.�8�"(V�bɈ�	
�'��1r@\8�b䌕S"�$9�'F�`ʳ5^���aŒL�,�0�'���Z!�M�|�d�r6�)I��c�'Ĩ,ȃ�֌D7��dj�:�(�'����Q.]��񡅈�mԬ<`
�'�"I�GI� 9�UZ5�,x���ʓ6�z��R,G�4�*,�<#���ȓ!���q!��^��V�_�e6����F�����*���Č 5�*4��V�x�$�
fl�$���Bm���J��M�Näd.� H�1+��H�ȓ5�F��ȯjK
,�BJ�
��|H��fh�8��ıRa�> ���ȓIg��)�	[8 g�X�GĚ��ȓ��up@�7�)�3,и.�~���k��0p#NK@�h�fӳ��ȓp��E��b��~�B��Ц��zJ ��ȓ�0��h�dB9���ݬ�δ��S�? ��+$���%�d�5Q�>́b"Oh�ŕ%�n�z��)B�^i8"O���tJ�9I��҃�."�֜�"Oq���3z��`j�	�����g"O�,��bӞ<-�!��m\c�����"O�ٹ��ԝL7�E  cT�Tw~��"Ox����E;J���a�CaX� "OBYd-Kw�TX3��+rb�"OfT�wiA}���9�I��4�s�"O���d oB\聢;`�hu�"O�|{&l�$x�L	1A��x��"�*O�\��垄w{�őQ�K�O�8p{	�'��ظ��ۿc&�*��p��A�'�FT��M�J�$ 6�˪[K�
�'�`B�HY8\=.ܪk�Ms^�@�'�Bd���cZŤB�u�a��'���Е�	�|�|")Ѐ{"	C�'��u۴�يbG����]AȪ0a
�'f�8�T�B:E�$2!'�5��qI
�'R�9 �D�Y� xCj֘&����'��84��JX���ң$c��;�'�M�C���Q�a���x���'}B�J��%7 Y��_V�I�'PE;��P�\Z�x3KR6|#
;�'� mB5�<ęISN�mp ! 	�'|��[��ȨM��(Kbb�d����'�
� �/(9$ [p`Q�BM�y��3*�b���A_�uNnٰTo ��ye8=�@A��r�Ή�w#] �yҭցq�B8ŏ��l�:�Jң��y��ӕY�"=�u�+ti� A3�	��y�Q<9h���M]�s��ex�<�yr/�=i��<!S���c	�� ����y�dK0S�t�ȱI��~$��E�<�y�o��>��(�|�\���۔�y��:ӑ/ �eo��� �B��y�g $�)X���^�2�JF��y2E��!�p��ӝU��)��cΑ�y�A�<n;�"ƾ{�4������yB�(cĈ�B�cn���5@C��y�n&*{�8��Q�l�"l[5jG��y��ǣay�\���>i�����g��y"R	%nxI��bT��KFh
2�yҬ_5�ꐹvOK�V��sEn���y��^� �|l�ւ\-G�|(#����yB匍0-�P�
@"��ԋi�y"k�>M,9kᦋ����S��4�y�b� s`i�$F"����l���y��^/�H�f�Z,zp�@+ـ�yr�Q6O�j1�W�+fF���΀��yR@���ޔbӄ��M.
�
����yB��?c֌�[�MC�N-��Zejֆ�yǛ���,��k��T��(�Q�y�N��X�l�R�";�9��B���y�J���,I��U�^I���&ꁩ�yB��R���
��-^�0���
)�yd��5|E[���X�(���QV!�D4n{���bI�L48 �	�!�$A�s�ԁ"H�g��`�\��!��ِc�z����8�ҨbB�X�w�!�ڎ[���X�>�R ['�R�V�!�
)c��Њ�E�H6��%ˇ&�!�;G�\m���-!0��N�!�dI:�,�Q���i���C���+�!�� .yq��Ͼ/��(;��]�iY�Lp�"O<�7L�#}­qEoɳD%��i"O>P�a	���Pǧ�Dd���"O��(��� <�h�'憂<�ޑ�"OL؊&��D�k��ܭ[��(�r�'�r\�d�	쟌��ԟ���ܟ��	<%���e��P�~à�D�	�����۟����4�	��X�	ܟt���0���6X|�Ge��erQi��
&{�l9�	�|��۟t�I�$�	՟�������GT�]�6:S�~-k�j&<����	ҟ��	��t�	̟4����t�������:R0-�$�
���՛u ϋ�8��	ݟT��㟨�	�������Iɟ���p�]֎1<زA�o�17T���I�p�Iܟ�����4��ȟ�����I�M�L�zroI�g8�m8e�#Vn	�	쟠���h�	˟��IݟD��П���;h�`�Fǜ�H�� ���&���П����@�I��$��۟��I�� �I/q�T�P����f���P��+`�I����	럸�I埔�Iğ�I���ɾA5N��-�yX>u��D�����ퟌ��ן|�	����ß ���4��~��R6CF�E����(+�u��ԟ����������� ��ß��5>��y�,�4H�t0�)�P7 �������	��I���I؟���ԟ��	,�8�j�;OY\<��A�$S�=�IܟH�	����	���Iԟ�ܴ�?q��Yil��G!�-I6����O\52���Zyr�'��)�3?��i�QBd ��<�2W�Ѽsb�-�6L�4��d���p�i>牀�Ma�S�L+0�Ղ�/���A���p7���'N�Y2������
T�����*E���S�lB2���g��5J;�or��2�y2�'w�Im�O�I��h��BT>+/�<JcG�������'��lz���q��\W:�C��P)H_X�����,�Ms��i��D�>�|¡ު"��̓F�"Իh�U�IP��
$y���͓.�6���O�F�@���4��$�
"� ��▃9p�A�(�� `�<AO>��i�Р�y2�څ�T��&@ <8޴�m	�#��O� �'��6M������$
�39tez��͈a b�߀Xj�	=��)X�� �db>�	0CX�d@�	�+6���gU�n-\)�CjT��0�'$�	Ɵ"~�RN4����G�O�ҽ�ť�od��0�������DCæ��?ͧG��k���+�Ļd�r�d]͓V�v�a��$���Pz����2��'r�^$��e3~hZ��C�X�����-�tD{�O��y�=.`�'T>���G\��f� J��^�'4�>�i��C�)����wg�0ht��/�J}r+nӆ�m��<II|���?�t&
z��@Wƹ ���pI֗_��hB0EX} ׍K��$F��
y¤�O$@�'�*5�vK���ِDX85�@�r�b[�d�'��'mT7M	 ��$/�9z��M�p�X� '�Z�x�L��IK�i>�I��M���il���v�2��1�d�j�|k�TB��I-D�ZE�^�W�*��0џb�I�*.����)ۼ���
`T�]	� �0��mϓ�?	.O��S�O2�q�'��@W�I��B^] �yRb�伂���s�4��T=��I�AS�'�@z'��O,���'�ɋ�M�Ӳi��e]/G��)@�'^^<�5���1���K�`Hl���Yd��Sb
� �(��`���x����Qy��'�pt[�fDqG�t�\�a~0�'l�'96-M�1O�'���jb�c��`�� -����'y:�q���nӰ��g���?q�RT9��h���!X���s&�.�>��4e(h�����;k���:L>��n[�K��灇�6�6���_2�?���?���?�|�)OeoZ�
p�8J�
O�ݐ�M�5���,?)�i��OvH�'͸6M�&#.��q�J��1P�`�D�Ĭm�#�M���	-L�'�X��B*�8�hY0\�x
�պ?�̸٧f
�;Q�	X�Fl���'��'���'-��'A�34r�e��K	�6�D��G�_�J�J��ڴ����?������<Yf��yw�X8X�̔k�aX�rs�m��-�7m�˦ ����ɉ5j|Ȩ�e5OcB�/~���s�4U���?O���.�*��X�Q�>�d�<����?	�N�g���(�䕿%�r�G��2�?y��?Y���d��Qy�l^Zy��'�I�%Ό4-<��#�FǕ,���dS}"B`��Mlښ�?i�O��cȌ�[D͐nU�JH� R��x���W�i�Q��X�*� 2�_�[0�O�U]`���#Ua��Yv/����Iʟ��	Ο�F���'�<MCA��(S�@�d�5(yJ�ˇ�'�7m]�%�����M���w���@U��*X��A�+^,/	 ��'�(7M�즥��4l�:=�#|~RI^����x��Tc�)�`�՚3>�Yʔ&��􌡧�|�V�l�I�����֟l�	ʟ�����"�r1@R�ԧ=�JpQ3�yy��o�^�ɇ�� ��A���i�AG=W�,K�C�Er���U��+ܴH�&)�O�"}���E}�(����V�X���b�a
4'<��r��	���	�����K(J'��O��q�@��I^2e
4H�f�<����?���?A��|j/O��n~�R牧Jh !�E����	��N;:�"�.�M��B��>с�i�z6��a₤@�\Nf� ���c��l���0W�p���d-?9w#4D������L^k� �:�CI�F,��X!,BG[���03O����O��d�OV���O~�?�&#�0a��Apk.Dq��jV�d���ٟ(�ݴW̼��'Ԗ6�1��G�$Y�EMP�5JpQ��T�I
r�	U}��k�αmz>ѱD,S�k$�ND���n��L�vY6���%`�b������k��hOf�D�<���N�'"I?Ea|Ċ2CA$"?��͓��8	�v`8��'E�C�Xq���-X|y�j[�Bz���I2�M�w�i��$>����ʒ̖Y��� �MU�u��	b��|Ƙ�uKZ�*��I�?ѐ���
�&�`)q��;��:1���+�l�SlCVy2�'c�)�3?a3�i@@<����-M[�<��ǍM*D["��ߦ1�	\�i>�	��Mca�!/h�9��)3�"!��k��a����'S���F]$�y��'aР	��`�C�OTq�ŉI5BP\�;P�1`2��x���O�ʓ�h����)P�	cŘ@�߲�$yc� �Ѧ�jB�,�I�?&?������3�TaA�� ��-A��t�'B� Z"�& h�j�|}�O��$�'�R��U��yr��.lJ���G�}��m{A����yb�T�Cj,T����ў���\{1��,z�$s�$�<B�B5�w�Ȗ'��'��7-�3�1O$�֥�.�A��9:,��� �	*���Gæ]�۴�y�Z��{���d�T��J#�8���{�KVHE�h�(�	���Ӻ;YwV�,)@��l�����}�p�aI;5GV�0@oF�\w�d�O����OR�$4ڧ�?�D�ˆ�H1Y�����=`���?y��i��\�AR���ڴ���y�Y*��4f�$���aP)��y��f�}n�&�Mぢ��(�0�ϓ�?Q�N֔7��ḁ���/���k� 
1��Ĩ Ľ"���I>�(Oj���O����O ���O��X�m��p�tQ�p�p�����<q$�iE첞'��'���y�\�G��I!�E��t�4� �K�PsF�K�voz�D��Ih�S�?���YH%�EJ\'��,J��ȶr��!��H�*Y�tՔ'��i��OG9E�h��Ŕ|�_��ai�f`�RBfE0(G $���N��0�I���IП��@yb�l��͠�7O�a�6.
=QĵAV���w�*lr�5O��ny��.��I��M�"�i¶6�W4<�.�w@�'l�>4Q���z!BA�����{_�	4e��4�$X$�H%?��^c?h���T�m�1R�iȴn�n�@�'�B�'�b�' ��'��������"<�x����u9��3�Or���O��l�B�ɗ'ɺ6�(��	<�� %�O}���ܭ�T��IN}�dw��Lo��?a�T��99����ɟP0mL=��x���H�$V�L��d@����&[o�h%���'[�')�'٨��j����Q��]�s\D!��'�R[����4GU�͓�?)����)�(v�Bx���

�����	��	����˦eX�4]�����=z�I���Yh*���o�`�qB�/��D$'�<�'$��Lbs���������˔5t����m0B�r��?����?9�Ş���ঁ�ǎ�� i��	^3K(r�"�-�y��I�'{�7m5�I1����E�qK���RM���Z*lrm�#�K��M��i�xU�@��������k�ꕷ\�b˓�"d�Vg%$@�ѣb�o7T=���d�O�$�O���OZ�d�|���ŧ�@ર�֣�F�bs@"���cԞ�y��'`����'҈6=�咣!I&��ECp�ޘ.{��9Ԁ��%`�4w�V�b>��5捰3���I b��D�֣�q�^0P?)J�I�k}�X�J ��&�P�'���'7>a�S���mT@���ߦ3������'�2�'Z�|�ٴA*����?	��$_n��e�S� ��GEҝnU`�rȨ>�#�i��6�_՟�'�ԭ���P���٘���j���'�"�?f�\H�0,����?!�M��X��ɓ���*�)�+N$z4!�8R�4P�I�������	\��y��RhSܤ�����V�f@q� XYRkӔ
�<!w�ig�O�D8[�J��f�ۤk�FU�A�@�(r�L��ٸߴw�&H7#z��R�'҉¼��S ��I�"A�F�J�x��B�O�d�KT�|RS���I����	ß�I����#�} <�Hb��Ij�;��y��oӀ@*���٦��	ǟ�̧��I��dؕ�%N}��h�'�`es��ˀ���yK�4`�J~J�'��EJ�42o� ��P됑`b�Y���,Z�&�����F����0�Y�\$�O��u����� sJ�XĘ�CwB8����?��?9��|-O�m�#;B����??J��6��kj��E 1$�I!�M��c�>Q��i��6��ߦ�h3nŜ0���Įd���ܓu8��3�s�����0~i3gJ�3��%�'���m�9���Q������rv!sC%t����Ny�\�"~�� �4��%�僂���,��d������<��Aߦ�$��pt�ףzRg�A�s�)tQ�<��O�o �M��1̌<�0���<A��n�Zk*]?s�H����(�T×Y�rA�c���hO�<��O\PY�T�L��X2A��|(�Q���f�����'��/d@v50W�]�>x��	3y��E��	��M�i�d?����YD�ӻ���'��HMnш@��k�hH�νY
�I�?��0
��x��%��رɈ�`"���v��4
�Oy��'��)�3?Iаi��d"�mʀ�|LH4��E�0@��7���ݦ�Iq�i>�I��M���w�Xy��J��!��(¯W?Qp���'P�Gks����@�� �+Qx\�&"$?� �<����L�漹E^���:��d�O�ʓ�h��lx�bX'n�ඃ�
4�g�O˦��@-�	R��]Λ�wR`����',��Pl��/�\� )v��}nZ�<ɪO���<�dV+~w,\�4O�TehϢ0�PXaКA��Z&3O�,
N
���=��<�'�?����楈�nF>8_R(��A��?q��?y���DGʦ�R�^۟t��ݟ���W�z�����؆5R��a��O� }�I��M#`�i���>�L�'}�ӄ B/#�,��&N��<���I��C�΄a���H.O^�	�!ZF�"3D�$��)"�!�B�n���b�K)����O���O���(ڧ�?��N��9 �YƄ�� 15�gL�?)b�iK��y7P��{ݴ���y'G���2����$�z5!�����y� q�d�o�0�M�n@�=:2���?ǫ��P� �~~J�ZTJ�b�(�a!2��h�L>�)O,��O���O����O؉��"+����i��
�r���L�<��ic�9�S����b�'ibvj��>:��e���P
�bR���ߴH�&j�O@�����)�E׿; �RPn�0Y�<�bC�0�H��4F�<�NQ�F��կǘ����Dڊ��X3.�f�q��_�j�����OD�$�Ox�4��ʓ]�ƨ���y�*�3:%��#�1|���R��yriyӊ⟤@�O� o�3�M�%�i.Np��`��a;NAH��ў*�t���	Ȉb�؜'�I�)f���hР��aC�	�?�(Yc*,i�e�N�n��(���	%�����'7��'�"�'i�'���B�]�"�Ж��0q2�1Ox���O��o�@-8�u���'�	7J%0��2`E=��;�h��7 �����$��P۴�:`
G�x�u��?G�L�4(�I�W4w�v,U���P��9�g��7��E�L>�/O,���O����Ol��'V+5Lb��l	�����O8���<�3�i�V����'�r�'@�Sm�h�Se�5XtZ���83Ҟ�5����Mk�i�V�D>��㟤��b�YsR��F/��7��Q$��8M)(��CV�=��ʓ�b�DEZc��I>yU@�$Yx<hAB!�Nj�$�?���?���?�|�)O6�lڜU���n<SQ�p��Ɛ�m[%l ~y�b{��P¬O6<o��΀��S���U+��M�+���;�4u���Y?��!��'�2�N?���J@�_+6o�	�)˸I���ԊA����$�ʘk:��	Dy��'D��'7��'�bR>ɘ�j0:v\hf�Z7Fh�Ӣ���M�&���?���?�����9O��lz�!떎�<��]�&��"6%^]`����M�!�iU��$�>�'����gϦ�C�j��<���+�rq�/K�Ȓ��<y��I�j>��I�������O�dE(T��-z2����͛@
 �(�����Ot���O�ʓm��&�H��yb�'a"&S�Or�XAS�T�Plv��5/�7d�O�(�'266�\�������d	;G��t)�lF#k���jD&	�$�OL4���:}r^e�<���[� )l �(J���;iV���Z*hd��7�&�"�'��'
����<
�$2>���q��z���0�+����S�4`9X��'1�6�?�i�E�u�.}(�؆��Bd�A$z��ݴ(��6dӖU#F�c`��Oz���'�.Ժ�C&&$k��I1Q0l�����n�f�On��?a���?A���?i��#�`ه��)=��f	&XIZ)�'ND6m�3F��O���.�9Opt��)]8M�xi�,��](t��g}�Ga���oZ;�?�L|�����Qk	�b�A �S�@�]qU��=K���W��DR)���B���<`HB�O�ʓ@�֔�Eڮ٨q��޻D���A���?	���?��|R*O�nڪQ���	�|_��Pu	�� �q�N���~�ɧ�M�B�>�q�i��6�����S�QYHSdI n�zi+G��-v�6���j�t�	�r$����R	��'��D�o�QS�#��`�!BI�$�&�4�r�l�I���	Ɵ0��ΟL� �֎oU���@��
S���Y�M��?���?�4�i˺e(4P��:�4��t�N�Y�	�hO"�����n��Y��'��I?�M3��i������)��D��'�R�ӛ�T$k��G3�Ӏ�0zy8�sȖ:p�B��|RU�d������ܟ������"ԴTA�(�AVv���ٟ��	Fy�xӈ@Qb�O<���O��쟦����'�"بT"��P'=d�����O��mڤ�M�T�'t�Ol�T�Z0�E!7n3>L�ћ�J�%���S��!aR���Ӊ6��K��DS�	#f�j8d�7*�&�s�½mV]�	ӟ������)�Sly�K�DĢ��Y�5��|�B���xajQ�Kg�˓,O�6�'��'��%՛���7 LLM�q��6K�L+"Ŝ�L��7���ŉ��O�>�:����9�mL�R�*4�c�Nyb*�i��m�ǭD�+��%����y�Y����蟬�	�D�I��4�OY���`�2�6�S�)������v�jɃ�3O��d�O����$���~�������XMt�§Ǎ!-)���4=v�&D�O���|��'���N\�PXR0�I�*�v�۰e��G���^"r�v:y��D����!N>�)O����O����a�F͒1�AO�.6����+�Oj���O��D�<	��i$���'R�'z8�K�'�N4��T�:�`�%��PK}oo�X�mZ��?y�O�d���M�F���RbVCYN`JQ<O���
�x��� �<�Vʓ�*��S��Rt���cô%3%/Y�^C`��GӎCj�S���?����?Q��h����� z��t
sg�^B˶'�>&�x�D�ꦭ��d�Hy� h������<��Q�	I�t��#�	 �牺�Mcf�i��7-�r���f<O��d[6|>��`���;�� �}�$NUo�zA�A�ԡzDL�hAl6�Ĵ<����?a���?����?q!��=���񆇈)\��`����D�Ӧ�ᒉ�sy"�'��4���lY"�x�p�gP6e�J�؇�H5Qu�_�&$x���Ib�S�?�S�56p#Gl8���( �.��G�<pa�(�'P �@v���z����|RY����G�m���Q�,�R�<; I���d��ɟL�����ryrFr�l��)�O M��C��8�k�OH�a��4�&>ORlF��E����M��i��7� �Y�N� �@�0��`��8؀���	Q�$�OL=���߇�B�� �<��'uk�4XTL	hT���p�t��q�D�OD����Ӎp��-V�4iYBij�'Yv]�b���ߴ �4(�'m"7�5��H/(`��V!
� �"-�Tm�6V,���X}Ey�lo�ޟ0QNBA���֟��X ��P��3ָ����V���e ��
.EE{�O!���pqU-ׅ%Y��x��ӠS�Jղ�h�X$��46�$��<����y�ȌF��d�GC�;2`f�(��Mq~��>)�i�7-s��%>��d�L�R�ޟ�x%j�L
+�r	iAϻ��Q���<?A��K%E���9��Oan�
��\<�J5S5dK�CR��,OZ�d�<�|�'��6퓿^1Q�ۊU̘�1���X~^�������ٴ�����'o�7��0KМ����*'Ɣ�#O�g`o�������v`��Iǟ�s'��/QD|1I#&?� d���d	6�|�X�c���T��?i-O��}�@��+-N<��!���3� ���I���'�-mz��$�װO<x�(�]"x=ҹ�`oϞ�M�i2�D�>�'���m`��
����<Q���D���q�-mƮP+r��<�I�$�d9�� 5�䓥�4����HU6p
d��%H��,G�-D���O��O�ʓ5����Ҽ��'"�!g��Kg�����e�e��9%���|��>Y �i�d7���'.~Ѯ��OIdшW���f�!{�'��D?W��̺v�_�D�	�?]��U}�n��Ɉ$�H�I�� �Ē���Iϟ`��ߟ���Y�O$2�5��I�X,x	��� ajj�[��gÛV�ԷGA�I�Ms��w�틀⍬Tf�۠��Eh��s�'�6m���5��4u�ޙB�o_�<��z��Q�d�����D���������+
���gKɋ�����O��D�O����O$����3��X���T� ���Ï"O�˓Ic��Ԝ|�	ӟ����C��~��d:e�^p<a�f�S,y���M�F�iѮ�/����0�IB����Q^�m�9 �a�p�6L��]>OM4˓R��g��u�v4�O>	/O|c`��_����`����2$�O&���O>���O�i�<Y�i�p��'�L̘b!�%� 1�'
��9��Ҟ'��6�3�����D���H�4o'�f�1xę�b�.I*�`�*�kp��{A�G��y�'��J���5tP�pT�x��8�5f杲������.>�,�2H��y�'*��'��'����ƽbW�آsl��p�I�䃊$zn���O���1�NMyR-rӪ�O����DR��<��0�̅N��xE�@�'��6m�ܦ���#��Rga}�p���[�d�	V�y�)zg�<l�tȳ�o� ʐM��H�z��Oy��'�B�'yR�ʓ5�A)6�<Q�P����׺C���'t��M�u���<����?a�'�����00-��ϖu��S�m\~�·>Q�i�l7� Ɵ�&>Q�� C��ea0eW*�kw��n`��3�*��wt:�P��Igy��O�Zy(ӂՆ&��'X��ĕb2�����)eo�)�A�'���'���O��	��M��Y�~�M�Ѝ @@G$L�%?*�'��6m=����d�ݦm���%r�FŚ�B-9a`��MC�i�<�bҥ��y��'9b|����)mR�
5S�$�ba�j+6��C"b�Z����g�H�'���'��'�"�'b�ӤB{�@� ˳b�}�Ǐ�x�Z��ݴ'��T��?����2)����.���0b(V>?p�Er�C�e�2�{ڴ8���O���|��'��V$��(Ⱥ͓^󶬻쑯H$Jy�#��.N2̓5���c�)>���*O>	+O��$�O�=)a&A�h��Gj@:_Nd(*3��O:���O��D�<Ie�iL�\JUT���Iq-0���MV4�� ��b#R-�?�tX�0��4S��f�O��� Ǝ#D"�	r��!KD���?9C$��d���@.��d럪�anOQ����:-<�2f��q^���Cϛ�����O���O0��)ڧ�?�@ʌ���K�B��.��gEލ�? �iI\z�OJ�oZB�ӼS�$��"��@�F�b�u �D[�<i�it:6m�ŦIG�ތ&Ѱ�	֟���5�Z1H�-PMJ��pU�@�p)�_߂9'�L�'���'��'r�'Oz|��瘍 �)R�$Q"d5�P�P�ߴnbڵΓ�?a����<!�*R?]t�����r�~�@��Z#]����V�H��Ƅ�Mӡ���O/�D�Ov\,[3�N�qaJ�q"F�m�~=��DE�m�Ɇ}J�
���f�$�̖'eF:��P��I�5쐛y]Z��'���'���dY��ݴX���̓1Xʘ�	88{\�2QC�[��l�қ��DVd}b�o���o���MӰ*�#sz���G�!T���ӆM�T��'��<���}HP�Q�n�=p|2�
,O��	C�[�h�;�,��2�d=තW�<���?a��?���?A����B�#V��C��(IxMi��E�	��'��Gq����A�<Qb�i}�'I��X�U�V� �p�@�|M.	����O\�g&��k~�����E�F	ba;O��Νy�� 6�S��,$��ˑNY;��tm0�jW�-�$�<a��?A���?�E iOj��7�P7EN`��a�η�?�����dئEqv�q������O�J��f���7�������o��Qk�On�'�~7�ۦ}����ħ��7�B#D�2�S3쇣m�"h�4I�ϦU�6-RQ���6Z�$���9v�]	�Úv�A|X���(V�Rjty�ĬY^I�Iɟ��	����)�dy�v�t9��S)g�+�(E"�r}�G�G���&�M��R"�>�c�i���
�?4��Hp�aEJ�^03sNs��m�#Y�v�H��y�p�	%"�j�Ёǂ�)(�'^��'0�UAs�F8����'p��(�	ş��Iԟ0����"
�u��H&p��ph��%�6�I?���O������<Ɂ��y�E;��@�NI�	>v9�r��0#F7-���K����4���	����X��a�D�����u� �p���$��A:�G�~:�)ZS�W-uL��O�˓�?1��{�)`-�+�N]�C�@D����?���?y.O�o�wĴ1�����	�=VP��j�\�~)z�#X�%����?��P�P��4`ݛ���O�x`L�`�_pVd1wN&{�.Lϓ�?g��#��<�L�"�����~�Cw˖�����ٽ'�¨+TD.R�����ϼ^|���O|���Ot�0ڧ�?���J���t*�7��(�p�O�?���ifN)I�V���ش���yG	O5tLak���5��k��yR�kӢ<l���M���.:J��?q�P� pz!;��'y�8��I&1L>��֬�Ye���L>�.O0���O\��O����One1��U&	8Sp)�G�j@�@�<���i!~��u�'�B�' ��yrm��Q�#m׬;�y���
~iP�	ߛDl���Ij��?�:p�6d�t �c<xPSb%Z	""TM�oV'N�b��'������e�4���|�R�\*�>E�r��R�X�ALpp�������˟��	��myҭvӀ|�ԫ�O��pj1Du�٘wJ�*O���!'4O�n�{��9���:�MK��iz�7M4e�����ةJD�ґ�d�Ve)G^4��O�] @�}������<��' k��=L�&8�&��z9:�۰AG
"/�D�O��$�O���O��Şr�	���N�omX(��kWdʂ�9��?���"���A�;��I�MJ>�V���,�JRh �A�cڛm$Z�@ ڴFR�F�O�h�KgG���y2�'�J`jтdvP�@ؔ<�k�ǁ\��	���)[k�'��ڟ��	Οx�	yU���0Q2�&�!&Dבf�^�����4�'s�7�<����O��d�|ZG�
2��X*�
U��5A[)��ɶ��E���j޴>�����OQyq���7B�p�˘��:���9���Ц{��	�?�(�H̚Q ���<�R�K�^f��T��n� �N˟������Iϟb>��'�6K��za���1&��U{���Nl�ű�T��4��'��\8��jަy �tJS���mX(ȭ.0�t7-Ц���B]#���@�Ѩ�	Ũ
*4�-O��M�3첸J0�ُV����w2Of��?Y���?!���?����	G�&��A(��91�=;��&<m�*{d������N�s�$������!\�eRt.0r��.�1�6�b�&���G}�On�D�O�5ʱ%]��y��#M�4 ���T�@�"���y�,A�.�����80�'��I̟���]��I`��8W(hy����5(BM��˟��Iҟl�'~6혫9��D�O>�ďM��I��mI$\��	+�a����T�O6ml��M��'!�I2YyΌk%@H�'hFAy`ό��d�$OP��Ug�%���M~
r#�#`�A�3ʵ�0�%�R�0��::B����?���?)��h��N��h��1�9JtY�ǘ�JTL�$���AB��&?��i��O�.� ,�4�G���I9�9��W�K�$	�q�۴�§#- `��O�5���I�~cN@�NL16�@a��P8��r��w�6�O���?y��?A���?��k*� ���
[j���+�(l��D:,OB�m_�\i���� �	�?E��y�	5?r% �� ��0c�!ۡ*��6c���f�2`�	C�S�?1�Sm��D��įtK�}�S�LF��Z'J��T�'Lⷤ�T�$!��|�T��s놡x��G��
�A�g�x��䟈��џ��rybed����Њ�O�� *��}p�[!��oU$�£9O�oZN��d��I �M�¼i~7��|� �+���I�B$��c�*m��m�l�B��D�O�Юː5�,��<)��R)k,�Z�¡��&-P>���\�h���O@�d�On���O`��4�@�z�V�¾?4͋�ĥ �H���П��ɰ�M��R*��Ϧ'�Щ�+�d�N����*~ZV��c$��?I�O�`nږ�M+�',�| ��ϑ�<!�$����vh�5�v���#��#�KN�B��S�����O.���O��d��bmA Էo�. �&j�	�p��O�˓h���k�2�'�S>[u� ?��QW֝�.�RF4?��Z��qݴ ϛ&��OP��	$
T�B�P]���t�
�N�̡�G�H"0!P��<��'iй�$T���A՞\��
Y7@x�'��M��lQ���?1���?!�S�'��������W�UW�&$R!���z�`@�[�~FD-�'��6�&�����$M榍b�F04�M�7��/m>,�P���M��i��<Hp�K����_����)X_Y�}-Odx!���$�����&F X�`�9O���?����?Y��?����)S�g3�af����T�S#��b�Z�lڡ�����Ig�s������c�DY�bo����PX��3FbN+�V�d��%�I{}���[�H[L̩��� 
؂�P)Y�	��e_=@�L���3Ot�����>!�̓v�+�Ĥ<����?T�ׅ3`1
%.*ej!�� �?���?����$�զ��t�������v��>��闚D}е)B��_��i����M��is���>)P�W����i��m�q!A��x~*Һs?��F�]}�O�v9r�F�]��_�0tnI��i1 ����X��'�"�'���ҟ���À ��L��߃g��zhUܟ̸۴u���k(O�Un�M�Ӽ�J֍E�8T	���	k�XWN�<Y"�i�P6��ڦ=*R���Q���I�Ps(GPp�9u�ƶo��0mŌ7�ʱ�p C�>,~�&���'���'q��'R�'{���U��&�X���O�V�!j�S� �ܴ+�t����?�����<�q,���� X@*

�qb��J�B���2�M�ַi�R��0�'@��!K��I�cH``��
k�� &	2}ԥj-Oԍ�񅇂m��y��8�ħ<�W�(g"p�CC���0da�
D��?����?����?�'����z5���+�-�S��$A3#�8?j�������#ߴ��'@N���c{��m� ��1h�ǊWx��@lH Q�P����g����ß�EK�N
)X�GPy��On�֘;>rijq����\4�Ӯ�Ac���柔���,�	韀�	U�' q�*S��س��¿Qf��Γ�?���r��6������즉'��YD��<c��S����S&�?٫O�m���MK��X�h `���<!��*�h��"��;Ά��%��aM���anJ�Dc����l�9������O��$�O^�H�H��'����*4I+%-���O6�>�����<9���'CT>���k݁$�!�䒋n'�A�U�/?�w]�@�޴7�V �O�c?����s
y�凚���((�B��Fl��$܏]�і��4.�L9z�a��|� �4��'���2	�d�2ϣk)b�'���'����R���4b@�Mñ/�/^Z�Y�m�n�9#�7��d��i�?�]��(�4Z�x��ƈ��d����͎+#`M��i�7���iƮ`c3���ką3N���lGOyb� �[=���%I^�Vd{���y�S�p��ПH��ǟp���Oj�@1a�n�JX��F��D���Fl9����Z��Y.��w��TA
G�s�nD��!=}����mb���m�#�?y�O�)��`����VBThs3:O���CA7[K�"$al6�3S8Olt�g!�MRnY��F,��<��?D��2n@�7ɍ'���6�X��?!��?y���֦��Tcd�P�I󟜰����M�F$ٞ'��P:�	H���ɖ�M�2�ib��İ>��M�0]�Q ��N�Gk��H��<���I�l��������h-O^�逗*C ����O���UNB	 ���i��8`0�"��O����O>��O2�}��=,��N�*4G��c��3*�����wۛ�ȩ���XӦ��?ͻX?4�	G��_B6���ĺX�*UϓP��Vkaӊ�oZ�7����e���	ugl���խJ��dɒ<"c�Z�f��U��p�IBy2�'T2�'��'�R �tUd�tO*0=�p�jа!@��0�Mkp��h~��'��艨�.�;y�:̣�e�x�0�S�LIX}�Ew���oZ��?K|�����$	�.|����U�V2Oʤ9 �_�"Q�x���Gry��/J���%JT2��'��	�wX��s�Ԁ9�}х�D�$C�l��� �	۟��i>=�'X7M JT�DP�l]��`��rh�x��"��+?� 妩�?�u]� �ݴb���c���S,���%I���$9tQgD7��)�5O���yR��Pj˓��'�@.v��E��������E&��ȓJ���F�JX�T0�7E�.^έ��	J���3g�K� �����7|4r����U}����Γ:L梬c��R� �p��N�<�d�c$��=h"��PQ�6ty�ؼ5+�R�Mι()hX!��ʔ	v����*S��L+��L'М9!��`�%k��gyp��hƇJX�ڥ�R�W���$��i��Q@��$�M���?�� �@�C3�x��'!��Opͺ��H�P���#,�
UG�iR2�'f��X�K��'���'�2�'V��6H��aX`�#I�7� �g�����+ߐ)%��I۟`'�֘:c夨��j�dhr��v�f�>�l��0�S۟@�I����۟��I�<�I�.��r��˦a�֜ؕ!ǀ*8�*J����'�2�|"�'���ә��A�R�R�,rd�b��&$�`��'M�'v��'���'S��ū �"�ӧ@�4�R�"mV,U��K+C�\On�$-�$�Ol�$A2���đ&E�yqGO@�r0%Jd�Q+~�� lZ���`g�8��'����i�4p�㜪M��c
E� �^�
�'������b�j�H{���%�n?A��ص��\�sM�-+�jI�s)D&pi�k1΢3�L��(�/"�*|��
j�|�z�Q0@�Vl�1�Ӱ
�P��eLʴ-�����ʩ"�����VҌ;��\*t���J��ئ&��աC�߻pVpj�d�4��P��`��0����"�N;^<��R�C�$r�!����>����럼��ܟ�1C�PW8�r"��3n�vi��ИS �k��W0r���u�ۼ��.�\c>������K)]3pAɑ-P6_�ZD����	�`$�6ᚍ���b���NjQ?��I&T�ހ��p&p�z�'ӫ��xZ���Or�n�������O���<
��̉ ��m^92h��i�C�	�Y�v�[b		�y⁮L$X��"<q��I���$ue�U`Řo�d�c��;qv��O����T{0�D�ON���OX��;�?9����eM/E)δ(EF�h�AFUs���D��n�yB �Y��ۺ.G�b�� ��� �ݵds�H�$�6ٳ� ?74իvg�Fd�8�7��&kQ�	�./̌S�y�)]�R�\���Q�`�d���!��>�B
k�ʑm�?˓�?q-O:�y�-S�{(*�	�/V=XP�BO6��τWdt�S�(>T�j��Y�^+�Gz��O3B\�؂s���M�鞥kdۑ�X�7� dY�ß	�?i���?���B0����?ɘO���₞ N��AÕg�+�j袂G�6_2hP���h9p/�u8�0Ѓ� �Y|�1��ƵD{��d
dt�ܒR%!��b����`�1աt�'ע����g���d�m�@P�!��	(hdh �=�d7�9�	7�H��DonU�#C�)f:���z~!�ĔZ��)��ά��DQ$MG5y� i}"S�S3���M���?�(��՚�C���;��
�Dd
��c�F?L���Ol��Rq� ��P	8��5:�L�q�1�p'�,Q�� �Pl楛�&��YJ��S�ɞ	�BtS� Ǒb*1��A�6Y�i�@IF�{g
}���ջR���Ë�$R�tp��	��l��On���O�ʧY��C��>6��Ut�Ǔ]�*a��������{LN��g@�h�T ���^C�	E���T�6�F�#!�)`�d��w�.PPtD�R'�dЛ,:Lmǟ��	G���H"O��'U��9K����c�'G�(Ґ옘}�D���D"7�{w��"�D!p���{�t�p����wB>Q�����s��X2]Y&��a��\���	U��"	R0�Ł�� ��Ͽ�
A�O�heåCn[v1��AɣN�$��(��n���$2�i9��
Dl��H��c�d0�`���	ß�D{��B!m����RK�$4�$J�Y�1O���ɦQ��4�����'"��4S��ݐ܊g�_8>��Y���?�RJ޿yV4����?Q��?yw����$�Ob1P��&ш���Lʌ5q�k\@>�yыQ�M�*}�V*v�2��� ��a���d�?���d�i�F�i���p�Yzb� @����k��I1dӟL�+׋�-k#t�T��>��!�r���h���:�B�xBIr?�l�ޟ��IT�ߟ��IPy2���`��L�g�2�i�D��xR�'� =P�X7"R��׆ 2�����-��|������zEn xh�a�ۜ��P#���8��X�Iߟ���ȟ�@��Ɵ����|2�d�V��I�P�>�k�K�	{P}�-D�0@P���Q�'ʂ8"�'2 �0��9{��jTB\	(  	�p$X8�	�`f�lv@�I�^�"8rbP���Ey��'��O��-7�&苢b�*b7nAc� �,IC�IL�$�`��U�l2��A*�@F�牵Yv��<���/`���O����|��#ڤO!va�Q���^�l�)A�6M�n]���?��D��rG풶yH�a�B-ٱY�lHТvӰa˧ȉ^�^i�v(�_�X����(Op#�/d�)�e�U�_�~����,��6m�(> L�Q`�YP>��5h��[
�\���A�I�Z
(��Ŧ}N|���%|�%�EƔ Op�����`��5�����?E��']�m{G���3Om�����I�f���O��=ͧs��CfӨ�dM�|hҀ���5�6(5+�	�h��tx�H�t`L�<��,#DG�-^��x�b>D��!�[=���{�Y��@i�7D��1��BK��f�j�
��?�!��fq*��&hX$8��dY��[";)!�L8jX�/���|��1���!�dU�$-�/[)s���Y�(a�!��Z�����ΐJ\��g�:pqPC��u*��pA\%>1+���-�JC�I.o�M��:�F�{�Ԍo�(C�ɿ$l8�!č���=ˣdR�`QC�bvl )E�>gv�a���P)3zC�� p`�����]�'�"V�.B�	�"��"S��,b��Pր�<�NC�I�Xl4I:%J_=0�L��Q&F�QqC�I� 1���I5yD��1�<F�C�	 |��rE �&~M`%����~��B�ɻ��@c�G��Lqx"��t%`C�I=_K��6��1��;rՆ  B�ɥBj�Y�aɶl�����
Td�C��<Xi�f,OS&}3�Ҧ&��B�	�&s��
'�!r%4�iuO;�B�I
_0�5�G��9�����@W
B�Y2��r��>W��	�%	,i��C��1q�:�2Q�Y�f��XV$[��C��%zCvA0-�< �r�BP���B�)� np��オxs�QC����k��I8�"O�!��(��yR�9\)�ȱ "O����
Uy ���I�<8%�a3"O^)P�� �\����v��A���"Oh�{G��!I.� ���9jd"OF=�Tŏ�o�&��f�&�,8��"O�1 ���X8ʶE�c5<�rV"OT5�Bg��1ӨD:w�ĐJ$����"O���tۢ��0|oαHR"OF!*�i��c8\#HʪV^Zl�"O6M�Ō��&�t����܍�F"O�{���N|�1��P�/��x˥"O�)y@��8B9��R�挼
	�q�B"O�,���%9GŢG�Ǹ^	L4r1EؒI�nQ�w,@:Dz��I��g�&��c jV;��	��2s�
Yc��F"f�!TB@�0�~(��i���Ɛ
X��m[�U�<i
�.}�,�Z*�O���  )[#��y��F�<���6�=Od�`�	G;r����� 7� IH���|�)`�VƝ��fPdܓNc�PhO>1�LK!�c�rE %k��=�"̓��� %���xc0l��6�19"���Fɾ�O�4���C�ܸ ����l���UK��Ol���E6�u�� w�H�"B��V�;�Rp��&�$� c)��a}�h�W �o�R�Bv)�,��S�> X}�Y1W�2c��8Fa�<a��0��ϊ53Up(1����p<����u;�L@���r��gp��O.c��<�R��	'�������0�Ow����3��\c�J�"$|�rw�'���Hv�/h5���5�͝/yn}۔�N����8HR[~�5�����Ol�3��<ͧS$���`ؾl�u/V>C�B��
��eP�1g(�L��'K �g�@j���c @�`X\ pM>���DMP�C�E�I��O�\�`9,O�D
1�p�!\w2DLR�S�E��H$�0H�bɪ:)���B�A9���@L�D������X1������>�pS�uP��$!�K��c0FF4Kg0d�U8�AɴlNư<�T��D��A�u�ɰ�aB ��OJ�G��`��K�813�$N�2#  ��h�.��x��L�x�ʍ���%:\)4�B�@����<`���!�ȃ-|���N����D�vdx��gN�d����H�$%\�	�CQ�o0z�bt�l≂_`�r���%\Ȁ����q�rc�P�����8	���2ĉcZ�BF�:�:I����?9��|�h��-c@�&����A�+��`���ӗ��Ûi�Ԑ����<|>|���������5Wn80�
ÙQ
 [��;~͞Yq��a:w(Z!$��xZc��!a��^1E���$O �V�[��䭟ЦOV��'E������-���s���#���R�N����ƍ�{d��x&C!pu���w�I <%��go�)rF���V�O��]��|z��δd�AIE�R1<q���U�����%���x(t//�8T��y*p'�)U:��DL"nqO萩�蝟��\2rI�tFT0�a�O����O�1��/k��Uc��_�&�.;��|�'��=���`fʉ/U5
�pՋF�6�2����Z*&&��PQ�0�	�l���~�G?-^ �p5K�u�.AyE	�.}Ԥ����/3t�P#��0���������`�`��"~����|"� v�d�<9H?��Ou�,[#OY	^w�Y�!�u:MhV�'�x܋�nͧ$d�l�0�I|K�U��ǘ�F=���h�:��pJ�#��4��uj���R��A�O{6R�uB�
S�>#BTX��J(- ��Q����:�j��I<-;x����F�\�TY��Zm�������ˁ���d�V�(�� C�:g�<Q�'�"����;w�Ѩ"�@0K�	+r��{�ǜ(�y�vj֨K�� �Ɋ�'�̸�
����'n�Y��O.���jQ�3M��h%P�pX����Ve�<2��L�f�����a����0@��7�T<gF�g�'��O��'��tA^�4�d�S '��) �9��9u�鑡G��pv��"�F*A�� �P!���Qv&ǘ	��:��O
��O����5n�D)Υh�Ǔ'�\�Q�/�%u+LXk�D��9;<$���҆�m�vz��z��Ĺ�f5��&x�d8�*��fղq�*�9.�����Mk�+����'f��enZ�eͪdN>� b�+͖$�d|b�����J�����dY��`��s���~b�R�o<�����K�T�Ԝ3Ʈ��(D����M���3F���Ƅ��c�
!:$�hX���Q�@���q����K< �$ɵ�	E�$AЧ����'T9,����O���x#_���䲄Nӫ�zI���Df�y��>�(�sv͒�/�\���_Jc�\�`�[$x�q��/,���ND9Gz���קܑ�ē2����_�c�.��'땥Y�ڈ�>�2a�:Nȉ�b�_��KHܓy�I��T�I��sFF7c|2�&�l�� ��&�����Ϗ|M�hkqNǶ���j�(8���ʋ�:�	�0N��*W����1��J�HK|��옉2�h-��g�\��%��i�� $p� �J	=_�5!o׺|k����dU��(O�O���A��r�(UC3�̘i�4����'d�P��nL�qShP5	0v(l�"B�^S��Y�ӫ:jv��|�ӻ*��J��Y��	�7�T�#읍�H���Qi|>5 �G.��`)=�O��x�)��iQ@D�a0H)�g!/�`������?�ǎ�?*?�8�GG�:=��qD��'�|P��ȁZ�V�%?�ٴ舸u�2�ۑk[�G�Dj�`?D�$9!j�;����Ee���@��>@�Ͽ�2)�>}���]u�:p�a�ǋp,�%�VdL4�!�\-!P����Ƨ�]��_�zH@�'�4� �Ǐb5��OnQ���X�<�f�)7ڕ<z�	��'�~ݡDM�?4haZ���e�R�[&,(�B��et0���[�7��\��*rN�d���Dkwў����sF}B����hY�52Z?��U q��
e�]�5B�`wA'D�H�� mR|�(��(j�L��r��O> �"�W��p�����l��I���银v$L���a�>S����f�1�nB䉬N�(8JE�Ӡ's$�0� � ���� ����>x6O�AC	t�|FyR�ĥ�5(�/��u A萻��>!E���.�L]�t�B����v��\:~�i�=g(�4��?-\��ĐD�|�Ƣ�%#���q� �3�ў�0��
_'���g�f�-B(�n���b�v�
�%����yr�[�N�6�[� �����!���y�`Ø�R�Y4��[X��'5Y,9��@�� A�	�1I� �ȓ/nr�D�@��HA`��|�|��.�~?��N"K�l��� ��.^�7�R�pG@�YJ�Ibȓ�p?�O�8u����(�:`8d��ё?J�y �?}�1�'E%`�e�A�Y����>|���$�n# �$�R���'T�8\ç`��xp��{�	�.;�X��wB``u"֥s_� �Qf��[P��'g�QC ��������I�6d�D���.p���"Od�j%�V����MH�N�]s��W�	���dK!!������3'.PE+W�>X!�$<u)�� R`��$���V(@�d�!�$���jr%�Y���r�Q�!�$,B���qq���U܄��b��v7!��e��i�d/��9�`@Aʤf!�2l?��7j8[p�r�*!��$mz��S���v<j: Õ!��a^|3a�L�Z9\|��Z�!��ҤO��·�p��y�CGY!�D߄w'v{��6R��C%��!���` ��svÐ�ݎY�fѱT;!�䖯X_T ���ݥbt���)ZW!�_�C���Ӆɚ�du�fC�1[�!�D��9��9��!\��٫�â`�!����A K)ˌD��̔�o�!��f���s��&
���!߭X�!�dKEK<,�q���E)�����4v�!�D}TXAq��^��,�m�dW!�dҢr����"��l�\19�i�*U!��U��Ha���^��0'p?!��+"�T��,H�n�DS��@�-*!�dR+Vn�[�ˁ?��$�&!�dET�@J�@S�`�n�;ѣ�$8�!�X<e(<�g�ؤz�$qB�K1q�!�$�:�����dF����"���f�!�d[�O��8n�
���v�X�!�$K7_۸�.��$� Ś/Q6��"O�9k�"��y��1�R�	d��st"O�x+E�H�|����({��5#"O�m%�۞o?d���`��x|��'"OL���� WZr���@�-We4e��"O���b�_�j6
��Yq�S
6!�D[�X�h ��+�)?��$�E��b-!��  -x��S�],��PJ:E��"O�IKr��6�T"��H�Pp�a�"O(����ǂ(�@��1I4(�X�"O	�E ��EC�Hxf��,�\%h�"O�	Цo 0��8��M���A��"O�(#�b[1��y��-��z�>���"O.���β2�̬��fA�ft�`9�"O��P�˞j$��,��UT�jW"O6A��AM�{>T��JM�rB��#"O6�X&��2�=�`�� K��b1"O��y�윊%��}���2&� ���"O�9��Ӂ2O �	4i��y�"O�	(RF��f|�@j@����ې"O�A�@�Z�f8�r�G���
�!�d�X=��R�C� BO�[��՞�!���,�ys��Z�$2���GO�pP!�$D���3A�l��9f��%5!�_�_#V�I!��.&yB׌Y)!���9+ PJ4�O~��ؚu,ͥ>�!�D��NV����y��0@ᇑf�!�D�]/����۞�<IkS�!�Ǝ���(qi�#�.� ��L�t�!�$�!_D�	���P��qfi�5*!�$�f`h�F�� �(c�!��,jnNQ+�A�mmh$�˘S_!�d� V�P3�ơ}�I��*��!��!� ���kD�{�,̶*�!�d2X�*U�4@P�@�����z�!��U`n`��I G1�M���˵p�!�L!bR��a��9y�`��$B.�!�D@�tr��Q�͜�Y!���W�=�!��I�-E��Q��&��S��!�d�QTJ���`�l�آ�AY�!�D�S�T���c��i�yr�	"%!�$%rv���7^�p��P�-~!�D��A5���Ì
-k�^���G� !�D�8�F-1C*��j�����!�O<>��xwJ��;���3��=%!�C�Y+Ƽ����Lפ�Xs&��y!��`��A���˿5'T��r�C27!�$��q_��ؿ@���' τEL!�.��g�}��`O�hP!�䅚V�*5��l�&8"���mT�@C��D�,IOV���*��I]v��riD�ybo��"X�I�ᄥtB�TM��y�dO���{��S�s'� � iH<�y�'BҞ� �B�. W����N�ya�4�Ԡ� ͞/`,]kF����y�#�F�� G*D�v�\31�*�y���$��c�X�.�	R�Z(�y�mVw��!Έ�K��8Zqm��yb�W�u��H��Om잸�0�ǋ�y�J YX����-ڄ<L�ɚ���3�y��y�b5�kI�6�:CF�ң�y�˛,V�^Z�!.e��p6�y�@�m7�0�c��q�����y��I�`��Hp�J�4��e�ūÉ�yr'����5��� eq�BI��yB'��Op������P�O��y�"�2u4k&���%/Be��CZ�yR%��a�ځ!�E/��Az�/�/�y�����ȫa
H�&:��QfO��yR�ĹR�:��c͙H�(��n
��yb��52���q,���rf߂�y
� H
�ٚa��O�-h!�5��"OA�A�	�p�z���4|\#G"O����.\�x:��@�\���ڲ"O>�J��ɘ�"T�%�0S��\B2"O2��D�Dȉ��I�.���J%"O�l�u�Z�L"rL���9Y�t��"O���!�53��Is��#�8X3"O2��4BD�q�B�ZP�ՄX�:\�W"Or�#�Z(�NL���,F�0��"O.��#��*}|<�Hd��8Z:m4"O� c����Y��Y�p�_�t@�Ҕ"O`�k�&�=J1c�-��x1�aR�"O���d� ��T�-c�8I��'D�ȠW�»2?���O���2�c�+$D�@���M��!1r��A�!��`%D��:� �&V�D#�b�.�$�2�(7D� Y`C2�	7b\+i���y�7D�Lz�#�+Q�!�C��1�����()D��i� �6���(R�H�@�)D��C��/���U�N�
1ZL34D���%J"�������Q�0D���m�0Ŭ,`��e�>9���0D�L1W;"6�rP�",�nĺ��,D��˰�:9'l��ƥCfzQ0�(D����(�,sP��iW��*	=X`B�4�IK���S�:%�8vO�6R"�\��f��o4�C�I�1K4�%� �5&��:q�.�C�>,�X����4">ؓ�EK(t�C�	&~G1�FT9�*��`-I�&ޚC�	��$9�#�^/V��⧙�U�C�	�u�$1S ������\�̺C�IU�J�q���lUEC��7L�C�I�
���:PI�6e��8 fUj����0|(� ss�Šml*	2]����'6���κ32h��'��C���3�N=�y��u����B�e-��
 ���ykޅ=\) ��
X�@����6�y"�\D��L�K�O��Sg'�3�yBJZR�YT*��N	>���@
��=�yR�N6�8�q�ڷv
ZYs��H��ybÖ�mL����c�"Ȃ\�Ȁ+�y�*I�YV��5�7iohE`����y2��-��x(�^Z}���ẼCHB�I#fR����8�� �6Z>B�	�J8z)�sj҆ut��z�I9qLC��'6 L��n_3[��y�oS��B�	�c�f�	'��_P��2��P�C�	�sA�]i|0DX�JX�:��L:�'�hlQ��^x��<���!�،!�'�����U�
������z�z�'ָt2�f�W�FD�я�*vj�'J��Vmv�H6-�2 ��q,O�EDz���2}��	@p�̛X׸�1C��h�!��/C'Uy&�)h���J*'!�$T�F?f��ev�����Q�!�dT�"���+� ���g����!�$�+b�����¿�p�J��!��ݯq��UZQ)L�}$�l�è�4�!�DV�WX��2���-h�(�J9 !�$�U���;�ċ�J�c�eP9�!���>y�� �<x�X�u�B)�!�RXD,����r�J�	B+\�!�$÷_�MY$h@�#n����ŷ3�!�DO�����v�	A�8�萢D�!�� R	 V��t�*3Oߛ:t�82@"O���G^He��'K�lV|��"O��3��J��`�g청�W"Ol1�Jȳ����f)�l�N%��"Oܘ��R�wE��׈��U��!�u"O*�%�8vr�X9�B�Ͱ��"O�|JC�V���a`�̣ b�]k3"O�	R�Kf|h��Fާ|Kp4��"O~�;�-"e���q�d\�x��y�&"O\)J�"Hh�3�"��CC��p�	n�O�,��M&$A�	�D�!7L}*
�'��T�t�ȶ{i��0@B�6d��'	��2	�=��\�c�4�.�@�'A�Ъ@@�"4/��K�l6�A��}2�'�8��O&n���A��1��'^l�pQʔ�`+ά���߳��8R�'��e�gɅr��1��R�6.��'�^�#Uo��E~�I��g�"W���K�'3�	�ᯃ�jp,��!x�+�'qQ��!�D� L�@�⨘�'E���v#7D�biY��6�$�
�'�T��� ���D£�G	yVD�
�'�P,�,R9C�6�cvb�hk:
�'�:�Ѥ�H>�`�+�o��r����'�{�CJ=3%
�F�hx�C�'��9ٔ�&w�&���ɼd�D��'�r���
�|P�!�S%�a�'�L�i�o�7I�&���[�{�P4�'d�ܨ�V����ɷ�كn0��'>���G�-4�b}8T��	e�t���'��Q(Ŝ����K��F���I�'f�h�Qi_�7�>�Y�C*F���	�'�]�DJ	rp��YEMՃ?'&�b�'��t����b���I��7�`��'X4D� B�-EZ�J+d�X�'�f9��5k�"�r�� ���	�'Ȋ@8%˒�-/�+�f�6����'}xX䎆'Fh��GA�Vp�R�'4�Q'�����"%�D͸�
�'�v��B�xh�Dc�'6+��Z�'�t���j�P XB䒤۴pS�'��`���S<�X[��W�F"|��'k\�(�.��$a3f I*fY�<��'j��AO%����u�U�^�ʰ��'<V�0֠֐G� �pu��+[�8u��'&�yT�^%:��<X�'��P�n�
�'�N��եT��܋ekM<8Æ��
�'p�-��@i�3JC�*d`���<ȉ���`9�)7!<��Ņȓ'	���1$�=l]��2�G�~�&x�ȓ94��a�GʼѸP×����ȓB$���g�׉^���:�K�t�����O�~�׭_9~��ʵ
Ł*^�q��4~dłv�P1A�1B�kG=����j�ԁ4�B�#�-JW9H��ȓh��:$�8;*0��ɴ"n��$R�H2`j�=δ`�Q��2yjx�ȓ�d�W������3l�jaԅʓa���DB���@q�*�|��B�	9Ұ@�i�%-Ī� D�t��B�	7M1�9��2_l`zF�H�\B�I/%;@)�qY��,�pQ5n&B�	'�|��7�?=���0� |�\B�ɬ1�>䁤lQ��*�
3}G�C�)� �Y�gWI�	��� �qyZ� �"O�|����$�Lڶ�V)�4��"O,�C�i��@���k����H�"���"O0��L�i�`��s-R��-"O�21Y+ƕ�b�F�`�.�U"O���QH�<�������I$@�"O���&�;%���ӄG�?7��r@"O��D��?&�)�dH;Sn��G"O@��Am �@�N�ၔ��"O:u��H\�9�j�$�����"OZ�KWg_�W����ǽ2۴
P"O��a%c5���I׋�%%6>P�p"O"��6L u�F�r ]4!���"OH�H' K+q�N\���|4�"O���v�-��P�� XԞH��"OPHd�ҮH���Cf*��x�|p�"O��'G�vउ3P)�Z�R!"O�P۴�J*6�Hx����wH�0Qr"Ox `)=?J�,���5\9�@"OԴѷ� 1v�y1oJ$��&"O�ύR߀�*�ɨ,Bd�2"O*QQ�ޜ$�	PW�Џ@�8x�!"O�)��N�A���c�b �`���"On8*1�%���V�d%��"O�l�E)�4���+c�O�4�@"O�,�d���	�,0�.R-���'"OX�s���2]��Qr���N8�s�"O>��̔�s�:�kg�0-~3d"Oe���и(�����7'��9P"O�Z�
ºK����%I%�9!"O��R�#�+�x���%u��h�g"O|3p�[�}���{�@��L�1�c"O�B���c�� R�G!U��y�"O���0LQ�Aǎ�s�XH��I��"O�qxBcZ�[D��!L
2^�	ғ"O�)P�-�-�\8���0Z|���"OX5�7�>ev���b-Y�%G��r�"On��&���a~��c�KG>
5���"O�,9���/^��2ʊ�]�d�z�"Oh|
֥O.Oj%���®r�V��"O��T��]��e
䍙@R:�I"O�$�4�R��˴�<�T"O9��8���w�S�`ϦMb0"O�,��m�R~D����&!�b��"O����+�9�xى�ϑ�ri�"O�����|�"|Y!�B1H��T�"O�-�@���;�`$�/{�r��"O��˗CX���\1�Ap0�.D��vi��a�̩sN�Gu�����.D����с^+vx��kY 4�H1q �*D��;A�N=�=�	��^�V�{�*D���E���hZ6.��W��5H��<D�����v���`E+ts��$D�@sa$��{��xT�I�l���
�f#D�� ���C�>�؄�Xc�)��'D��T_:��6���έ2$D�T�o��(j=Cf���r���T`<D�$Td۫�X0�C�j���ц?D�D+������\�lBUn�]��M0D���U�eS&�TI �Q�ƹ(�H/D�Re�}�� ���J�?�1�#�+D�,cG��(MNR@9�b<�� ;P�&D�P�L+He�U Q�	�
a�""D��xU��	V���L>E����ǆ?D�� ʴӄ��+=���G� 2����"O 4�TFI�^+ި�g�]�U�0�n2D����Z�0'�u��#Br6����d?D�̩�Ю,L$�0��JW��K��>D�#���f���Aǜo�h���!D��jW/�;X�.�z�+����+D�<���R1]F1 �m�e�J���6D�|*Ì[����t_�!�T�3D�(R�؈O-J��([�u����1D��x����y*�)S�N#�-�Ԋ-D��K&��� gܼ��C	�@�8��I?D� y7 ��Ĩ0�Ƭg��tZ"�>D�hz�I
�'(�ɀVň` 6���;D�|�����F�L�+# ĿG*����'D�h�T��U�"m�0b��/>��	8D����g[.$4<z��%r�t+�(7D�4)����f@�*d�2S�=��B5D����/�1od@#b���,ܥ[��4D�xF�P�m�f�bŏ<zg�A���3D�l��#ŬN5 
eM�'-�%(�F'D��Q3���@����KٺţG�(D�D;D���.ys�K�8�L��T�'D�(�Rh\#Ъɨ �҅%Aj�@2%D��3�薠� yh��VqV�{ �$D��R��
{��@g�źb�b��!D�x�[�%�䑚GoV�m�@�x�� D���e��O�(hX��� �j�[0<D����I�~���a�"L�|(B�;D��SC�H�o�$q�V@�
X���i��9D�d�$�S0q:\���ǫ��!�}�i�g��g����$�:~U!�V�I8Բ�oA�!��i���/8!�D�s��8v%��*#��h���!�D�2/���s��%�J��4'ĵ�!�\�FC�ѢFG4�2Ui��R>�!�d
PMD�J��ŉ�&�Z���!�D&i
�R��� �� �A�k�!�dWg�@��b�}td��̀�s�!�³2ܰ��,,�̸&�Z�Y�!򄙅j|T��ŢՏ|�\ȩV�I�~!���(���8?���tI�S�!�DCye�����Ɨz ��P�E@�-�!�	F��Is5�+tF!8A��-�!�$��~��c��� D�8�'	�T�!�$�+x�����C%a�	��	��!�d
X�D�x�.Z� ����g��:"�!�$+X�n(��,Z�u��p�e�G��!��/-zb�
E�]�G���0FB
!�$��r�ځ35�B�=�h%@�"��C"!��0F  tr��ar
�*P���>m!��ٺLz�4��̪=><�`!��wa!�d�0':Lx�ш8A��`����u�!�U���<�#�+coH�+O�A!�dH�D��i[$HS�x[*�K��Z>)9!�$�<i�+#'X�GC�iу��)!�$	�Y�������.;��x#C� f!�d?ծl"��Y�w�Hp�K�E"!�d�
���+��_(�)�1�P�50!� g�L@�䒘}/�}z��O�g!���> �^���#:�j�Q�ʄ�X�!�5HA�RӡX*r�>�f�W;�!���1�$�
�H
�L�d�*6M�3�!��&�P�+1�I�C��i����!�ϏZ���$M#*�� ��O3!�� <����u*"%k#��~�P@RU"O���L�*[3HYȆ�mr���#"O���Y"j$�q#�A#8[���"OZ䑱�=�DC�)C�2NnuQ"O�a��K�3_Brv(�	A=��!"O��c-^*/~�����!Q�r��@"O  ��l	�{�ʹH��ڰ$�����"O���BOY	� �{��ʸ8\� 0"O
�J0R�μ���d��R"O a�����R��	��a0"O�àfC�H0�Ղ��şO��{�"O*HS�/ld�sf�V8}&`��"O�Y`#��7ms���$�
:>�)xc"O�H5�&*��۶g�i��q��"O@�R%�2~�vac�C�5�f|��"O@���FT??<
iBU㖔3�L���"OP��1`�g�<X����v��	+"O�ͨ��� k~���b��5"O�[��cK��1�m�
x��"O����#K(��c�D�U"�"ODi�A_#_ό<EB*i�Z�y�"Oj91���%R��uyt` 7s�l�g"O�q����<@< ��L��J�r�p�"OT �g�˜4���!+¼|塀��"O�u��S�e
L�ǩZP�F�p�"Otj� 5q���P+7(��"On��AjQ�'�R]��ى_��-�"O��)�	¸9,�!�!}���ac"O�Y�B%ۻ0J���55�Q�S"O@٨�eD��(�@&^.����C"Oz-�!k0^ɨ-�P��'��@��"O��[�Așqa�BС�	1���P"O�
�AJ"c<0CT(=�Jd�E"Od� Z�zfHũ0A��0=F-"O��Z� ��Z(� �Q6m<c�*O$��"ƆtF�Y�v�ߟy�4�
�'3����Q6H8��fܷ�T�
�'PZ"`�/3�y'&>5ގ��'A.�kC������WD̷ ��(�'¾1��� �y�l0�	Hx),��'�\}���I�|P鐍��uԲ9��'4h	r��5U����@��6�N!��';ޠA��J����"��^�jD�	�'�@�d�A&%͖�ҫ�;m��m	�'���� s>�����_HL(C�'T��{���F��0P��X��,�
�'Gd0w @�n���n����L"�'�����]�R@y"*ĨzI�8��'r�}���ԫ��S!F�%c$n�x�'���RVlL����Y��<]�FP��'��f�R�걙ր�(P1�`�'
�05��,�Ę����0�	�'�F=	��B9a�S1lП�$��'�`�G&��Z����䙠nqb���'H��)��Ao���z �3�F��	�'9�}+Gg�WAz���*�7�J���'�0�0� �6�2u�* h�'����ͪ=���Y�ʈ0���a�'.�,I�Ș�p��Q�S�D w@�
�'�Ԝ��"MY�����fPJ�x�X�'Y���w*͞n2832�оpL�q�'�l(�Í�c ��rmS�l�@9�'%4�a�B��tH$��c������'˒`A���=Y�	�AP>�`iH��� �LHf�F�F��h*�φ�vr��G"ON X� T�H�NT��l�rz��5"O~���*�'7' ��e��=	w���"Oj Ƞb�4S
���c!�!c�F=�"O��X�D�A��(Ұ�G�$b��"OT� ��5/-�q�Z"�ř"O��h7h&�$x���*q�"�cB"O@8�teM�C���Q��>[L���"O���գ	LX]����,��"O ���`�>J�rl���A�_(���"O�m�f�[�ҺUjelΡ[�=p�"O���d^M��Q�W�Us��R�"O:1 !�m���fS�W��d"O���ܫ�^�9�>g E�C"O�(��d�/6\�P��5^��"O�}��灢3"dTy�%T����"O�A��Ȣ4�n����E21��+�"O�㴥�	z��Z�gې<��ˆ"O����؇H�X��
~P*xa"O��BDӔ]`��J�"I�)l�:P"O��J�G�1b1�pq&��U�HK�"O��з���[�ι����:�"U�F"Od�p��P��y�ǟƞ�@�"O�0���
kdXZ���"�`��"O�ժS��k��+S��=�Zt�"O�@J֢A����$F_�r�$�8�"Of|�B���bI���K�h���#%"O�aY0dD�DĬ��ʅ�vV
LBU"O~���D�2- �
���fP���"Od4A����)��_1:T���"Ox��1��T:|�34��'M��b�"O0��֢*�j�(2m,E4�$�@"OpD0PF��e�X�`�j�)�p"O�|p�Ȕ�74��Ӎ_��|AV"O�I��(اo�|e��GP�ν��"Od$���P]�!�5�*E��<ڷ"O���`�H"H������N��K�"OX`ש/#
�-ZHچ �����"O�X;0$N��`��0͙<U����"Otś k�\;�8J$c�~u��"O�L:/��w�թUa�p6��"O@�2F�Z	����"YĻE"O�I�6�ݹ�B-с�ABy""O�ܘ���'�"|�p�%J�BE!�"O�dKBD�;,��@`	�d{
}�"O,����YqTD�3Oļ<_����"OԼ�"* ,��#���b�� �"O6̀ǭJ}�!�R$\5pH5Q�"O`�Xj�=r��F�e�da�c���y�Ǟ�/)K���� ې-���bH�ȓu\}8Q�>�ZH�'ͻͼɄ�J,��)�2}=(�1,��?}���ȓ	C�L��!@XJ��ؖ!^#=����ȓ(|�IQ��NK��T�A��)��\����SB��QŬb��$>�~��ȓ&ú�r�EʬQj��p�9I^���%;j��`[�IO��wAV�}
6�ȓD�=i��ú.� J�X4�m��/��isa� %���K����ު,:g�]0IC�X*�o���ȓ��M`1�A�
�� j�)�+����ȓ3�L�b�@ЊE'�y�C��~ؔĆ�Q�:����,?t��g֘s���2�,�@bm��h�^�s�ٗrl��S�?  u���ʪwڸu�Qa �0-��y!"O��*@��D<-I�.��d�Yb"O�bV	L�?%�a�RN�)PI��"O�؇�$�������|�v�à"O�qa�I۔�Q®'dvdIsD"OX�8ǇրU|�ucF�A-o�aIW"OTpq��%d���`3��~i�x G"O��q����v�|���	!�D%�"O��k`NN&S�z���� ��1	B"O�� �6��q��J���ab"O�)�TiО$��E ��Zzp`"O�p����7ތ���A��~Mv�X�"Oh`a� �1I���v�R)-l}��"On�S�G׆x�,lS`���`d��c"O歸W���)h'A�<fX <�b"O޵	A�ƯR�,��e�#O�i��"O�����%����e �8��"O�� �M� :B��Tc�WI��"O&�FʈY�0��g̷/Ȼu"O,J�b�$q�l��&KNP �a"O�	8CcP�qqd$Ғ�
sdԻ�"O�GU�X`���^"8��<��"O
]1�O�
(�V��d)�(H���"O��qC��^4�	�ʑ�.d�5"O�M�7������H��@��̱a"O��A�ӴE}D�
�ŝ4��ct"O|q��ܒa�r$yD���IR�"O\]B�"̴/� Mʥ�Τpm�|�U"O����F�}0��$��]Ѫ�"OV�;hP`�p�c�\`�+�"O���#�V8�q�e[�i��"O�	����M d�f��,hEh|�"OV�{N5�.)����	- HI"O�����D�V܀UƎ"z�B"Ohd��7RMĭ��ɸt�p��"OL�
�)�)�ڵB`��q����3"O	㲠�JQMۇ@Z'�@�d"O^�ԍS=Wf��T@��< ����"O ��K�y������<���"O`�b'��'�ҴX2do,|"O�$�3,]4��I��9C��R�"O����ہH���ꆭR.�%
U"O�)�!E�T��T�'��t��"O2 *�l�.�4��J�?pIA�"O��ek�L��d�h�k�~�
�"O�A"@��Q��=�ƈ� ��Ir"O�H����+0�`�5�J�P�6�:r"O���4�J�6��E�
w��h�1"O�MP�dn�����({�" �!"OQtIJ�/��@��_�Ʉ��"O�Q��Ϸ^�D0�l[��)�"O�ɳR!��~�V�r��<N��"O�i���
{��p0G|���;"O��)cn�(},Q�b�6g,���"O�$�bN3��� (Ҥpq����"OĠ#�N�p~h�	5��L���P�"O���� ���M�����p"O|�Q�Ԁ~:� �= ���"$"Oj�"		B h0d��D���"O^=򶈈z�E�P���Q;4�0�"O$��c�(.����Ӥ@>�Q0�"OftZt!�0���&�>a5޸K�"O�"�E�m�$#�
i+(��"O `x�4c�t �g��O
4��"O� �MRcתG4�hB�"֟}��͡7"OҔ�&
�a�X���JBP�1"O�٫�N-�+�[<?.(���"O��I��^<4-���˳\8i�"O�|��D��Yځ)�H���(h"O I�� F%=q�Ac���/ָ�˄"Ozi��̕�f�zm9�V,^��y�e"O��ca�0�И`"�3�}kE"O���q�(}Z8�)��ԘE��S�"O��tjJ�w��@*��q���"O
P��=`0��d��G���(�"O
�P�^�(�a��Ʌ^�L���"O�a�t�%5�p�Bw��X8�ܩ�"Ot�c�/��~p��E!(x5i�"O���IP�`4R�P<`��r"O@-P���i�N{��R~�9�"O@Ԓi�@��1	4�[�&I�3"OJ%yr��*��U�V%�
wg�͑D"O�I�%�0]�VH�4gT9��"O�3�µA��A7/ȅ
VxX�P"O�8�RJ��`P�y��@�2i.�K�"O^h���K��($k�h��p4"OlPKB�ɭFu�@��<P}���g"O<03���T����q��<LG^p`"O8����pd�I�G�0;?L,k"O�<���K�e�q���v���"O�Zپ+况)�$��xոii�"O,=���6g~r�H�]���*�"O�y��7I8"�Ȅ(�|��"O�$���%i}�l���R� �
�z�"O��C���#E�=��ɞ>ѱ�"O��y1��Gm^'#Љ�����"O����C�+�8���Y<:�ܐ"OV5�4C����#�`�f�4 H&"O�8A������T8G ׎,�V��S"OЭ�,B.6X
�x�dǓ7@��"OdK��?I#8�a[���jP"O���js��H0�@��ڄx�"O��r���J�m�1���Rh1"O�9�/��E@�� �!@?
x٠"O$Pj�eن"�D�t0��1"O��H&h��H ��v PČ�c�"O$��D�]�tJP�s'��|��$&"OV��c�'��4�Tɑ;D��� �"O�`��B�9��%���C��@`�f"O8��ήW{�E��
�$Y�D"OlE2�[�E�<�P��Ҟc�L�*�"O��Р?Ĝ�Sb�(m��@b�"O�tp���D�R�r�"�A�z!���Z�R���$�f;B�֨<v!�D�Le��H��w���cPdV��!�D��#o�}��j�:K�Z�e�	�!�� �N�p#f��s�P��Â�0(!�d[�HmJ�S�hڂ@Z���ىz>!��[w��4*��^.a}�mB�+�$S/!��6��+��kk�����%9�!�DѬf(�A��V����[�{!�#M���{ͭl�����7j!�ʦ\�h����D�B�?Yk�uq�"O��C/�%<z�Z���[ZLA"�"OIp�k�p����E"<Ry��"O��2�+xH(�c�C�~��C�"Ob顴�(6�M�4�K<o_Lr�"O&S��F9�D��4���{$ni�"O� R�AF�5~%n�D�%�(��"OTUС�ɡ)��s��j����1"OJ9�w+����(q��5rd̊�"O�]�K��d��T�&#Ĕb�0Za"O���m!s��pvt r�
�=G!�sD�\Q�� G2@�T��i+!��N!}&��b���^ ��`�J@!��]� E���"𑑢�?�!�d^�7Q���ëQt3ht(5; 8!�àd�樲dh�?�: �čS�aF!��N�u�o�i��X�-��-!�ă�	.��w�]���PZ�Ƅ�:�!�d֝x5F	+���"g��g���>�!�]�h����d4K�><��@M!�Ǣx����"b���C�p�!�drk.��ň�1 �`@p� ���!�DE�;�����^h�0 ��F*k�!�C(R� P גV����Ï�;!�\�`hd{Æ����4�n�/9�!�$C�Mshx3g̛�Tߨ��ªR�G�!�Ĕ�.xx���I�g8X�(g�I,j!��-Gy���(�^� ���p�!��+��P�P��.�Aŧ�:f�!���tÔ�0`�K�
 ��@�W�!�D��F ZRhA�̼�&�+�!�d��z���F���� ���x�!�ė����@��ӥG(�p�Iѵ�!�DC5d���%��>P��#�.#s!��[$0���� *�����P�fa!���QX8�����*1�I+���D�!��	,c=��3�S :U��"��C�!�$�5M���d�)6�����AB9�!���F�v��g��8�u
�8�!��:p@9k�����	<!�$>toب�!o�;�y��A!�B�+��Y��$׼�bG�!�T�n.���a��{�F��%^9*a!� �U�`7[��3'K�K�!�ÑT5V��3�A,
��U 7i^��!򤍄a��xEg�(���'�{�!�$�=M�d�+W�X lӎ̳eG�cˡ��<�Υ�7`  ,@JP�S-_�y"+�h���RU�?$R\��G��y��L�f���@�!���� [�F$�y��ͪ��pj�����ʋ�y"�0q�VO���;�./���'�4 ����%(�H1#G��/^�m3�'(�UѰ%ٽB��) ��L�YDT��'\����^#(���V��O@�٢�'X��굉�>&;Zey��?�I�'�d���S:0���d*O:w����'�~�K��_:d� ���hG¥��'	"a��6r�غ�g®,����'�D���('q���F�)rn@R�'����+�0^�������0r�XP�'�0Y���Љo���h�6+
�P
�'�b���U-�Xs�'�;9�hC	�'����ӻay��3& 1!*L��'׾\�j�/:1��ɦ鏭0��L��'����CEż2[*	��T$)̨��'�6�J)[LЛr)�qx<x�'��:4*ۆD���R�$�bRHpX�'�� ���5=S
 ���!l�$9�'X�u 4�ڜO�����e�6�Е���� \�!Pg��hTb����'XSV��"O��:FB�4�]���ߥ A,�qf"O�<��m*�D��L֊��*�"OЬhF#K�~��	�홚Y��9J"O@�� ˜�K�!�F�7V�d��"O�5��F����-�r�Y0N�Dy%"O&-���P��n|��D�=R��X�1"Ot��v��^��CJ���"O ;���el���,�?lsbu�"O2��PMH.��$y��ԉ�����"O��K۲6\�Sb��x@�"OJ@�pTe�Y�*�8w�
�9A"O�40G&U�*������)Ryx��`"O 4R�r���pn�`�@@q�[����ɶ',��SGLP(�1R3�K!��B�ɿU��H� ثB�y���?8��B�I!���+�
gB���p��B�	�a�T@9�25| ��hWM��B�I��a�r&�d��Ubf�+,�.B䉝cO�	���
VѢM
�)SK�B��-F����ۊS�H�XW�$C�I�\�|��egT�6=65���$(��B�I*}��!*�;��0�(�U�C�	�Rx���eZ,`��٦V��C�	x�l�:�L�9�썲�ȏP��B�	>}ń��% \5p�z�����y�B�	�-٬E�X�x�r+�D	�(��>D�hPE��� :�L!<.�Dj��<D��3b��	8pX��D�Bx�)�6h.D�4��cD1	�d�٢/�*9���i�b8D� ��)"��5�#Ê�z�T}[�C4�Iv����ď4&W��#���1a��*q�1D���MSjz��f�Q�|i@��-D��z�CGU����B�
$`kq�8D�$"�GO�t��7 �w�HI1��6D�8��'\;EP�ĠJ<HPn��$'D�XI��F�8Wzi���z[r�&�2�Oz�	�eیD
��K��B��R�)i���O���0<��LO7j2���:;-n�a�m�<��iסGR�89�mR�D�d�R�M�j�<���R�t&�؁��E�p;:a橝o�<��	I�N���Ѫ"c�Ȑ�g�^֟��IR��hOD �� �\=i�S/�����RO)D���T�G�9)�0� ��g1
�;G�%D��DF�vG�i�.J�VQ�k!H)ړ�0|"�i���Kv����r��M�<	�#@.�Xܙ�o��0ҩ�I�<����(��!0��YZ� ���Io�<�ݰt����R�Q�q��+T�cy��'k��x�G;;�`���Ɣm*�ܣ�'$��bf�ظ����I>1���'�(��U��ck����7C�I(�'�"a��� �&����LG *�C�	�=I��`%j/��:uEC���C�	��D��8r�C��Y78B��:b�L�Co�-P�M�Fb �]�&��hOQ>Ap�%�4������W�9����!�!D��;ae�:��p��AT�:�b!D�$@r^4)�6h���.֎����<D��0����s`>!�G
6֌5r��:D�,۶�C]_���F����>D��
BiB%{�򁨷���d�KS�2D���@@\}��aR3ī}-RR@2��?���Q����d+��L�\!A�,L~!�� �)�2���S���т�[(AZ�0��"O���sE=A� ��МfNj�#��|��)xO҄8����~�r���"16�C�	�(C&p06��/�TЅ���Z�C�I��a��K�V��[˞C䉯l�h�Za�*��,�MUi�˓�?Q���Ġ<q��ā�>>�"�B�M��tL�Q�H
��'���i>!����>~�|Y�$�ے!�!���q�<�$FJ�b�����Z�$U2m�m���<$��F�TgI6a	�m�%��@g
ź�yb�Y�|#h] f����p�6!ۏ�yR+Ľ�h�[G� �� �l\��y�/@+OF�I�mֺU
99U�3��<)N>E�D!��w��P�dETA�IQ�Ģ�ybʠQ�2��SƘ�Tz�Lz�b���O0��'vU��� "��Fz��Ҁ�Y���@y2�b�/�� bV�84r�I�dֽL��H�ȓ&P؁�C�"vԦ1�B��U�X�����Iҵ��K��HE.@��ȓCo6!��kQ�0Zf1
q$E�WS�A�I[yR�|�������� ˂����Då\YΕ�6D�Hz���]rR��%&ݲ	✵��<�
��$J�jI	^��)kw��+)O�؆ȓ���r����m���^����ȓb&�����,��J���Bԇȓ}�X��!�jk� ����?�0��ȓ���	t�Ҷ�J��W� ^�-�	T��������ɟC�䨶��f���Ï<D��ɗ׫&"c��{dp�o<����<�O��k�H��.y��Ȏ+vu����x��2T��2P"�1"N
�P�j �y⤈!l�P�j4�Q|�
�'D%�y�%�hOZ0E���X��Q��"�PyBO޶p��˳e4oP���J`�<Y�Z2 �l�̙�\����!WX��hO�Wp.0���Ą?d����ˌk���Ɠ5��U�U�A+����� +i.,�'d���gͽH��� H?a����'�u��L�V20 ��3V�J���'�ڠjVÑ� ^� :�(�"=�xT3�ŁQ������()����'�#�!�Ğ�i��uW\hら˗qў���ӲK�P�kW�F�q��d��)a���=i����d�<)�O�,(JĤ?V���p��d��}B����$)�O�U���"lE�%����qB"OT���}���`��&�U��"O^�q��
6y��t@G�(n,��"O��G�D�y�����?C\�Q�"O����@�#DE.�����D5�S�),?�pyJwR�1.v��rn�]!�P%;�Xm3� �2(V��7���.!�d�7�6̳#,E+�fh� �z���ȓ)�rPd;����H�@�2d��#(y�#HKd�Lͪg@В��!D�@���ĊJ���E�	I��y$��O�=E����1V��)5KȠi�Lac�
�j!�$F�g�l�C1��7�4���;z��	O�'��	�<�!��$0AR�@�xE1$����'/a|r��	p�x '�C7�R�03JV�y�`�kݮM��O�zY�L*�hي�y���tj�p�!�V�j�~l	��	<�yrL�O9PAzn�0S,���O���䓂hO�,?��ͅ	VB"��(���2f�]�<��C�L����j�
8x���W�<�  "pdqHXQB%d�T�'�1O6](b�!5�C��<ސY�"O$X������d��w��&�v�@'"O���CF��%VʴU.�}ʾ�"O�U�C㗾Z^@��1.�7Ӛ%��"O���(�"�ޡ4b���|��"O�Q�	�$�B а��X6pIj�IVybU�8ϧ]xꉓ�Dԭ6��˔�@���%�4D{��DՆ\N�s�k�:�t!֗k�!�d�,�|�@4L�cG���7x�!�$B�b�H�!G��a5�Q��	*R�!��0�j�� C�������	Zy��D%�Ӝ/��a���$%q��z�DG�T�؅鉾%���Cu�n\Ա�2��_l�B�I�o��#ҏ�^����GZh��$�Ot�x�
� e�m{���?	�Ԇ�Y�#�ҽ�����/W�����*�-`��D�b������ �ˎ�ȓg��t(�gF���p+T�
u,���6��-����r֔� ��X�u�ȓi]��pTN�";Ѻ�y�c�#Jlh=�ȓ~J,j�K%��Q���k����������%9�Qɶ��J����ȓ(��87�d��$b��1"O���S�xV��:7 ��|p@�"OB,;r@߂#�"a#�
�>^�r"O\�*���}�x�aw.�<7ΐ�c"O�ѡcMހI�t�և߳.���G"O�+��Ͻ	Y�i�TF$y.}2�"O��y�%��A�j�q�dĜc|�Z�"O8-�jE��dx8u��\x�(��"O:H⠃Ƥ%ߜ�����a�"OR�T�38T��p�!P�?Y�a�"O�}�� ���T��XK��H�"O����ğ�+��ܠ�֚I��q�"O�	Z���6C���hb���Y\� "O��TE\4@\���F��&F5�"O�l1�θh`���=>�!2*O���X*�������d�)�'�N�߸5���4,�������hO?ـǍ����&�Q�Bm,�؆j�y�<��@ʲ�,� ��̆m�*���Q�<���ەmb��V	E�F�����T�<�gf��c{���$�-�A��mKV�<�P�3zK�LHh,�)�Щ�N�<�4ˋ�_��"�W�=�	��	L�<�NO'1)��Hue�>}��� 7N�H�<ɔ԰7��]g�
<!���#�O�<��ʀ�u��C��"�jcb&�L�<q��ːyX^�`痻@6^���F�<�f@�83��Ik�:��e[ĈL�<� G_5}��(XCdSD��9�f�HL�<�&��nT��v��35���2�OG�<)�H�V��%S�I�^�<�nHL�<qq��47���J��}Q���A�<Qc��b`�!�M����Zt!Rt�<q���$stH`ҁ� &��4�V��I��V���O9��`s��8�u0'�WW��l8�'� �S���e�)�N�#M����'/<ɕ��~i�I �IG�x���'6h��pB��IvJр��i>X٣�'Rݨ)�,o� �G&��ew��{�'��)ؔAE�Ybǋ�#o�lX��'ۊ�1�R;n2us�dM�<��1 /O��=E�� P����	5'L ��K�e�Y�"O,�آ֕�(�+��z��x�"O�M�gѾ:��EXAi��B�9{"O��jEK�����ڏE����"O6���F��Xr��P(�I���p�"OƐSD�_�Wը�mr|()z""Oƕ �G�% Sh����_?0Kl8���'.ўb>a�'����p���6�{�f�J�ę+�'B��čۜ@)`aY�Ӏ;�
�q	�'#�Qa�E�2G}^4S���46�x(��'`h�3nN @���k��_&��P��'Ъ�pK�[5��GD��l�
�'f����0���W��*�]��'_x��*En]p4�w˔�L/���D=O��y��+<�j�̀:v�D�"Ob]�f�� ��5pg�F0-w�+�"O2� �R�a�9���yk��D"O��Z��X r�&a���8`Q��K�"O~��B��=���&ƒ�$=H�
�"ON�ম�r�H�>S!���"Oxe�6 V�!E�|���E+	~U�"O�����óT:9�g�ġY�P��g"Or$*bGЙnz]��h b���B"Oh�jr�� Mw��: a�#?ӐM�F"OD���МX���k�	��9ú͐!"OX`�m��o���ҴiHC�`e�W"O���N>@"r���`�"�@�"O�Ҳ쏈A�ڤ+�@�(J��0�c"O*�i�D�A��`܆A2"O���R[���o7|��"'"O<�*��əB��TX ��3IEdc�"OP��v�\+~+d�Z��B)z^�ty�"OT���jѷ?��a�
L��`"O�$J����ˊ��2�K�5�I�"O�m�a�R!T���ҠmE>cvl`"O`Lzf�V�aE.�u,Q��,l��"Or�{��Pz#�$�!��g��"O��XD���V�^���>gcl���"O,��l�<ô��+�<p�"���"O�S���[�� " c��[�"O:�JэM�d�/QHu�j�"O^E���E�$���U��.U��"O���g�T���@�AG�5%d�z�"O�JDB��q�КQ���/�Ɲ��"O�x������{%��B�� "O�M�VoKy�V`�J����3"O�A��P���|a�^�9ɠeS%"OvX;����D)'Ы1e~��s"O��8�=pN͋`葥f�
���"O���W�@m�̺�gؑwX`��"O�� ¼:̼AaR�N�m@�͊V"O,����f�	�����U"Of]��C�8��*�)٘R]@�Cq"O:��R-�Q�@]��	A$BPa�"O<���I�,#�d|�v�)q;&�B"O&�jg��*Ss ��v�H?L-�)��"O"8�C�$J�MZc���8�D�r�"Om��OW�qjYQ�j�D�8�G"O U�5�	(A�!X�ʶ�0Ԉ�"O��Xs��������֮a��P0"O���VD�`��Y��P  E�%��"O� Y�\M[T �'�:�ً�"O�Q`�͕-V:��3�C�I�|B�"Oj���cQ�t�PE�֭�<V��P%"O� �1ӓk���7>�vq("O|���;���HQ˄�x���r"O>�:,Ȓ�ޠ��DR\�r�Xg"Of�׀o�� �E )Z���"O@�zu� �.>NT8�k 	,X���"OT�!FQ�u�y�2% 9n&�1�"O����[1�:!�AW����q"O�
�2H&@�`���t�Đ	"O���f%]ؒJ L�^�zh!�"O�`Є���#�H�ŉ	?��谠"O�UȒ�8��i�'=q���Q�"Oha���>$x��w���y���d"O ӆ��7}z^e����# #8�c "O=�d(�?r���t%��0%B0J%"O� '�@q4����#Q�.$���"O&e+�/�p|� ��u#<I�3"O
����R�P �ʕ��%gRY�3"OH���s������8]l�l��"O����#�`��t���d6��rU"O.���e��3jW�G5"�"O�I�G�) t�0�/8�L��"O䀹uA�1�t-��cU���"O
\� dJl������	�r$�B"O��ؠ��/g�,�/�@V2F"O������]	��zV�]G��"O� %l�!M� e�7m�>��)�G"O�k�t7^�p!
�oH�)"OD�F_�c?n4J�(�'1��D#""O`P�TM�U3����G`HF�"O`5�D��,m��}`��'*��T"O�z�&ѯ�R8�S��?>Ջ�"O��GϜ	p"D�3`ʖLZD\�`"O2]����,&�� 8�nA5�!�"O���nE��%�t.ۂ�N�Y"O�i�Gj�5U�БS]v�����"O����F�U�b,\P�L "O�-�5G�/��j�*��0^� "Od�sk�@�~@b�	�v�H��b"O ��(G<W���E���fT""OP��g�N�?]T�;��_�	��q��"O(�2���+N� Y���m��	
�"O��׏���\X�d�&6'�}ڗ"On���k�"2���U�L �Dq"O���FIX�]Æ|!�eϡ̨�5"O$���җV4�ecW����*G"O���� �?*l���D��-7����"O>�8�f�����U�0>@�Pt"O�� ����a�0µ�_=[S����"O�l�N��ɶ&�F0��"O\��� '4����D��^A���V"O4�#�,���ã�6'"���4"Ot�*vj��@�䖳(Ҵ��"OJq�		;Xđ�QM�)L��`g"O�9�3�E%^��z##O�w��I�e"O�I�i�KRI��Z�j��"O�2��J5�����fOy��`@�"O�uk(�#�K4D��"OHA ��yt�����!�}a"O��St�?��%���E�&�"Ol�K��
.4��`d�W����6"O����"ڠ���(��'u��ز�"O�d.]*�� �Ls{��!�"O^	���Z�*D�	'�*��MX"O\�l�L&x����/AI�3"O� V��C�X�~�w�s,a�c"O���CJ�:Xh��Aɮ}(`�"O����� T^��Ơ�H�!�"O�ͩ2�	�{�h|�f��j���"O��X7	Q�MGp�[ Z5Xc^���"O���X�pbP<�f��ey4��"O�8ʥ�N[��]��E���"O��q�怙r�&���o��#{2�� "O��@1�Klz��@���-�z8*�"O�0�T�ՂS,8�0�2�BP��"O�P�S6F��)*V(Y��z0h"O���1�٩5��|')d�#�"O����*D�n(w�_�~��1"O"��4��A2as&)>�4��"O4⦬PRy�Q���?�X�"�"O(��̰.�<R�T�?�8���"O��C(Eb�Q&ĠQZ�0�"O@��*��LdrP�bE�|O���@"O�@���Wbq��U%̄2l.�ط"Op��F)�0���Mh��"O���n@�O���d��LKT��"OF*�Ë�� �#�5"���"Oz@��ㅱ1�Z8��0W,T�q"O�A�p����0Y���#ثq!��9c���+�78�b�{�\�E�!�DD�@�lKDC��:rX�*��M�!�Om��tH6�M*���g]�!��-���(�d�%T�j��&-�0s�!򤜙P�V�Е  L���"�+ߦ}�!����lQF���~���ہ o!��@�L�R�b�e�q  �j!�Ӝbl�-�sE9È+�nҬ ^!��4�i1�ƃ6����v�٢IT!��x}�v��������/VE!�B�3��̚&/x��u1���a�!��'��TB ��C����ͯcW!���G�4$�n��^���C߲p!���pDI'�R;{�&̚T%TdF!�D\�%h��VΎ2"���T� !���!1��d�b��x�J)"�IF1�!�H�~��I���X�_b�!�D]�@�a�U�ЩS��,~�!�.Y��Ja��gi��"��!�D��/qj���-P��`"[�e!!��'E\L���)T( J�M�3�Q�7!���j�\"�H�4�hB$�D6�!�$�(22&�9tOZ1NQ0�j��$:�!��>�ڍ���G�&����р7B!�D�~X�թ]�t�����i5!��#���B&1%��)!��r*!�䍚
��r��o�Hȃ�Bo!�$�� �,ty��?�>� B��^�!���C����K��r�4��t�҃5�!�X$3�
5hX;A�`�[fė([�!��V�v)h�j`����ƹ���K�.u!��	m�
8��Q%:��S�/��K�!�������4�p��Ɂ �́|�!��I:M��<S ��++����2n�!��M���q�d�JScҼ|�!�ݴO�FU[A��&S�,�9��<b�!���I��p���ǧg��Z��Ը�!��I�.��gh��"��yc�kI�!�Ĉ$]�,ڒǕJz�����=I!�DG1&����A�N={тTI��Ub!�� �f�g�:�B��ыhr��r'"Oj�rd�VJu�q��j�]�DR4"O��;C��p�J��*�Dn��Pb"O ��L�t�f���ǒ0Vk�Z4"O$��(J7>P�9DHA�,b�9Z�"Ox�Q���x��È�)b��v"O������)!T(�yև�\l��"O��F�TS���fٞ$U�a32"O�p�$2�<�sQ&?eO��Ks"O��%ĉ�M��%OW0�H
�"Or!���0+m��/M<y"d��"O�,���Ǹ3x �9��P+	@`A"O� r��X�@\SC@�q��y0g"O��p%5��WN[�^���zV"OHq��K�m��Ua�M�9��;C"OFX�@��(�;�bS�G�(��"O��Xޔ=�r�4�E�~0t��Q
<D�ġ$���u��dE�0�f<y �<D�`�`Ȧc�r�xխD�O�b�I2�-D����L1�l)�D,R�R�{�",D�tj2�×l�*0B�l��"�6P��+D����E� ��D�D�R\�h�	(D�(k�k��.X�6�P�x�d���%D�����J��DE@F͏��L��m'D������g��*T�	s�F�{S(D�T��(ʼM^f�S�*�)s<�:U�$D�8aA�!ը����9�zu�`G5D����ɟG�J�У~��x��=D�|��eO!b�D໲�7'�.��Ӂ7D���e�O "S
{/�%(6���0�'D�\��/��t�-
	 iH���b�$D��P�
݀YG��c��v�X��>D��Q��L� Q����j	Ƅ�e#'D� @ f;3S��+r�S�g��:g� D��b�lY�^�`*ץ�4Z�
*�*D��
���J��,t숲
L7�y�R�\	,*��+PUd�Q	���y�#.
�	�/IҸ��L_;�y��7p���p�L�)I�������yB.D<*u�,�����R��[����yR��s�d]��wF.(w���yAƜ;lR�5e�)��*�!ȕ�yR�S�Ys�QkgE+��=C����yR��>:^�� �M�wո��ǏE��yB��&L���z���"բ�r�O��y"��+}D�8�� �zY@�勸�y2-R�����Ԁ)�A�5M@:�yRf�i�Y�@B�:Ծ�%%]5�y"�ږz2�Q1�|�I4��y��H���!P�߶<��Uw��2�yb�:�n����E�.3�pWE�>�y�h��H�����n	�'��(�k��y�DJ�b��C�A[r厸�&˟�y�	�7H���g�56�� W*��y"������`��=(�q����'�yr����u����	�P0f����yI�ba�9��� �XDµ*E��yr��)�t�t/�
K*^��bm���ym��L&B�(uF�B̮�2��y"(K�2o�̢e���@V�h���9�y����)稨��N82�f(#b�:�yb��%"dv�𥃌�6��gٵ�y��'M8�[ѭ�(*v�0�ՙ��'}ў�O"�1��Ӕ�2d����~���HǓ�HO� .e��M�H�X�����)�D�7"O6� ��A�$�.T��F�v��"O�`��2J<@�vI�*ז|��"O��0�.��Wm*d�ƧIj��E"O�E�D	=0�ru
��ʋ{����s"O�d�f��&���cED�L��0"O��	T��<�dճF�Ow����2"ONy��B9Z��
�`
�2��S�"O���Bg��-�Ƥу��4J'�4H!"ONUj��� G:x:�܇u����"O 	!K���5�G���w�i�"O-���J���<Rw���+�r홒"O*샤�K��"rc��t�	v"O��[�e�Wlh9��y���*�"O��B��5�L��7���K�����"O0��ƬĊ3��Yە�*D�`�Y"O��ؑc:6��(`vC�</b���"O����F���I���MS�Xc"O��z��2Ač���.fܼ�"O�1��H1	P4W��B;�R`"O�\�V�Ȣ#�I�ׇ�>^6�D�v"O�T�Q"]9�Bx�&ˢ22x��"O�x��Fe���s�4�,�"On9(6��'&���@�y�9��"O��jg�]c����@�x;�@��"O�x�X9ﶤJu��14F�ñ"OP�$8c������=!�"O��3�����*'��V�B�KU"O�h{w'¿,,lYr���c�"OĔ��T�1j,��K�6�fa��"O@1��#_,�\���J�r�H�"O���2EO�7'V�H�4).Ա2"O�X!r��	`���DX,���"O��{�$S�Fq� �3���9�"O�Ժ �&�Y��ϝ�-�x���"O� ��B_QeP��5��Ȼ"Of9�3�P�)��=�l�4��� "O�|���^�;�~$��*�� � Ű�"O����թ1@��X�ɯZsd,�"Ov4�C�D�8�Q��V�:I\�["O&�p�j*-���v.�9٤���"O��0��Q���iI�зB�J�Ye"Oɺ��<G�4=�@�@�I(�"O^���jǰG�d�K�����"O��rIB��X���`n(�'"O���ه,�"C�H�$ �H�S"O�}���ߟ�NA��gˋ;����'���N����hWHN�jyb����ju!���"sE�Ѭ�o:n��nI�gg!�ʩ3^�0�J!	/�
W�:E!�R�n�|p�$�C-I뱭Y,!�dV�f���E�ԩ��KvM�'R{!�D�>\pp��)�'V�ܻ֍N�$]!�$�=���a	�,H�uX�,Ѕy�!��דZL��5�B>FH��Q�n�!�ݿ{O6u�e'��d/,,ISY��!�$��F$�P�Wp!�ظ��θx�!��ID��	ud@�*&r��b�=0[!�d�g������yn*� vQ�#V!�d�?B�Tᢢ��0qP:��b�ȆK�!򤛉e�������3|g St�Y%!�d[!T����g�Q�{2��d���԰*�����-^Iv�ؽ�y�Y'?� ���ýI ��/K�y
� 2�Jf��c�0�VM��l���"O
	1�i\��|�yu
6U��(3�"OpHа�=
K,��CԔ\�F8�"O�1���k�zh0�Ok��a�'C��2��H�� �J���tJ��~E!��1s�y� !�9B��U���0<�!�@'a2<��tF[-�d�+BXws!�FmZy��,@�hi� �ĝ>W!���&sy�yЖE�4x��\ᔧ���!��;I,U���}�s�!�Dۀ}�>ecp$׿U{��I�ʐ��!��$h�z�%�Hx��&�K^�!�Ð_��[�)�#Cɦ�H��t�!�IT������X�8�i��L�!��>rp�
� j���
�+�`*C䉕ъ�AG��b����'�17wC�I4J=�-Rw��6S�D��C��_�B�I1h�[F)�5En~�3s���"O|��'��ft��&�H���j!"O�]����W��jO��&�>���"O�Сs�i�
Lٕ�Vu܄RU"O�Q���-EV���\65_����"OB�B�ɶ�ֱ W `Bl�q7"O��`��?th`�����$t@s�"O�3�`�.7R�`�a	�YgN�)�"OP�3fΙ�:z��(�	oX�p"OF$
a�>h��2"�S�e�|B�"O�dc��ʹ3mbw��<)D����"O��$�UB� [�lMC���"O���� ����;�K�3RF����"O����c��/,�aȥ���q����-�@�S�#��/J���%�,A m�ȓ��z���.�d�HQY���,�ȓLil��a��
���Ҋo�졆�S�8@�6ÁY4,`f���A������æT�%Nܣ1J�h�h�ȓUH�1B�B��$�� �+�
�ȓg&�K���	&��GN��t]���ȓ.�Y� �#��YzQ�U완�}���M�s�R�h'��)\�H�ȓ^�%��+�.Ne�Hi���<q�����)S.�/%��\��gY�>z�B�ɦ,�bp��k��1�FX�c� ��C䉲(��K򤋼w�����d�B�"P����(��h��M2�C��_Gnu�P �X� n�kh~C�<P��qX>����VCDC�ɕ}2�b��g�A���|�C�ɗS�<Ax��^�4���ۚB䉔��سwk��N�p"/ʐdpB�	�V�b} ��B.J��͂�I�9/xB��%)�䄐Aƛ�BV P�g�D���C��#��`�BX�)��<yǇ��ՈC�	�O�H�M��p��(|XnC䉰֥��ÅE���	���B�I���x� �.�8���M�C�	b�"$r&�
��B�Z�� YE�C�I�X�]���sh���lه|7�C䉨cp��� cb�m�EF¨%��C��:Q�PT�a�
"��cRN��B1�C��<nEޕ���y�m�W.G|��C�	%J�����>>x�����C�	-8�vR�-�;2����	L!lzzC�I%�����öc��P��-��0�C�)� D���F�)�&A���!"�=�a"O�<mûr�Uц��3G |i��"O�@d[�7�CEʹ'�U(3O������s_�����?�8��	~�^�j��Ќ,�r�"�n��vVB䉿
���h�HF;J�T�Y��]G%�C�	�M����C0R�8�3ŅW�vB�R`�rp��~~~@��L�$l�RB�	�b:�!�)Ė�(�S" ��|B�	��%`��ʅ,��pP���U�C�	?0�������:��ԚEfM�^�B�I	.�>-ȔB�.
���A��J:b�B䉐3����bٕG&� Р�=U�B�4S��kc�_!(����g�è�B��C��`/�irz�3�GT�kLpB�I��p0!K  <tX��C��|��B�	)VHh�"r%��,BV#Γ/$ C�	�c'0)@E˖Bj6�K�I�vBC�	�^�$���̀Y�Y1��;m�$B�	z?u��/ϓl��<+�%>
B�I���0��go�\Y#ͅ�A$�B�	�zT�#�M�O�؈���aNB�IH�j��@]� 6��*M��B�	�[E��A�oF��C��ƈ�vC�I�F|��C7)#5�F@8� B�jC�I3��Db��V�5������8*oZC��T	$)P��)$^Ұ
���	�tC�	8Y�mr�aֹv����ШQ?�C�WP�t��B��=�>$���O��C�	�
�0���ǆ�p�pѢ��y"�C�	+%��{��2QA����)>�LC�I�J��Xt���xۂlc�C�Q2B��< 7�U	Ra���Xi�*!��B�	�Lj�s0ӸmN����M�(�HB�ɭ
�!aS�ɡl�R�z�*oOB䉾Pv<�!�HEH�.�0��C�	�n�l���*�")���R`�X�e��C�	�Z�!� ��߾�:�AM�1��C�ɕP�!C�I&{y� P�Ȩ+Q0B�	+
YP�G�H���A��%W�C�	�"w�mR� v����Y86��C�ɞ*�����X����Pi
�	��C�ɶ;pNm�B�u�F9�F/'Q�C�	�t��P��X�P���D���C�	�L�:S�M���#���TB�	�R�0ܛ��. r�0B�eX�7��B�IU�L����XE�q%��+��B�I=bt>�*t�z���J4;[��B�	�C�H�)s�
�k��pQԣ��E2D���&냾p�ʄ�CeȕD�P��G$D��0�6+�p�0Ħ-� � �'D� ���)�fT˱��V���Cp�&D����銫uX��;$�Ԍ,;����>D��q��]0f#�(`<B�a�9D� [��V�>�d܊�a^g�\�ao3D�0�7g@2K8�P2�eH�eb�T�a.D�X	r'��Y��H[��ǿ#�`�{�.D��ѳ�ըa��@���N4�r�k/D� �D.��_ߦ����ܽ�@��'�/D� �#V([`��J0�X8Z c��&D���F؛]\{"�� ~6��Ӊ(T�����J+BD�a̘&B�Pܪ�"Or͐�DA�v��Q7��:�&a�v"O�q[&U/~疈����JX��)"O|!y&gJ8��P�~�Z�yU"O� ���6M��In�H{@ϊ��LX"O�H (	�4 �A�8�$��"O�x��*�+'�:�ҳC�!n�r�
�"O\��� S�G���aU!�����d"O��V-]�O��}In�X�$�0"O��`B>%s�Ic�5w��Y"O�dK�l�1vV��7Z	�h)�"ODE����[y2�ᱮ�'K�¤� "OV�hb� K���(wL���;"OL#���X���+J��0t��R���֪��\S���|�'�	:,�By�M��������Z�5)��dݬ|���Qq`ݖJ�丰���:_�d�jV�N��a1�J���E{�O'nɺ��&	�(��Y3a{"���2,�U�H̲5��O*�+qjs�S/r<|��aĨh�z���V
���h������Q��,&�J���K�(v�\k�'K�D�F�J��/����R�K�{�>���%��>i��-��A�hI�js�&?Q
�DE*�a���!���%g�ФXd���G�)8���"�bDZ�MDD.��<Q.O��Z𪆞X�ֈ+�i�#��K��'j���t�̐v}�=y��V�T�b�i��9�>�R4�ׇ{��X׊��t�^��|��i>%	�F_�]z$ӈ" oh]��=���"!l`Mä˝k�i�@��2��0"��V5��iJ�:ATm#ską�T(!�ߘ
��d5�S�O��x �%���;Hߢb��͐E��q�q��O�g��5fmߌZ���>������ˏQ�V�#��S�>���w"�fH<�CG �x��y�G�X�.��M~8��靆HyD���ʃ���0���z��a���d�9>�r�%�E�h�ۤˑ�QSay���5��ɰ7I�!
��D)Co�?a}h�!�]9]�Н��g5i~��SVg֞�֙�%�'�h��f���,�:6�T�|�T�H<�U(l��要�/Z��<�7��#\�h���/Z������r`�����؞�x�'�&�yb��%/��-���61��p7(O��y�"*ݡ`�\K�hϚS�����O5ڝaS
��~���x�a�!=��f�*+ލ�LG��C�>n�KcR�=+�g��ni��?%;`Xy%N�0q^�H�̗�<k�s�C&ʓ�@��C*���J�Ka���ɋ�^0v'O����Y�N#��5%�I��\x��Z�7Z�с,TT����LE8����	�0I~X8�B1����B�'�dZ�`5z��#�	R|��ȌM�yv�>?Y��S�8���k�b��
ZL��֤�
n- C�I %:��n٫2:�CDg�Bߢ)A��=I튅Z� �?A0|9�mZ�!'�Ov `��z��z�E�J)�e��B���"2$�d	B�$F,ȓ"��QT�#����K%E �#��8WY�K0�[�5�h{d�@�'s@M�*7w��0 ��۰	��U*�o�|=I �5e�˔�+oݢ�*` �<�Y�F� I�2l�(�ԛ�HQ%�p>p�� _�������3��h��oGt��=6d����o�lz�AP���;�.�KFo�����"�Fa�dC�&1^|� ��3,�(E��e;�D8�/Ź3��L0�L�Jn cƣJ7�F�k�I���ҷ�F�d9������DF�cq�� CNQ��f�c�Bh�2�WmH<�  %�z�a��� ����R��h��I�Q,�U0-�Qo	.�^�VJ�%�v�Y��ė(uj��Đ1��Q.X2Av�y�P5��!�X0E~l)���Ⱦp"�d������X�WT��;G�K7C����I % ,�a���(s,����DЮ|�J�O������/~�Fjr қe����yH �¯�� ��G6o� Z�,��m�p��"Oڙ����cD�j��ܻ+�0pY�!��~�r� 6dQ�u�©�R�C���?e��cޝr"n�3L��@z���7p���>D���$�&=��@�Ǟܲ���PJTaR����,L��)����d5�DE*��Ӭ�12��JᤗICR��ɰU+���`��`��@H��pa�㒖lÎQ�Ќ�8��AI=*m����{�}���>]�t%�V�_|���@�@��(��aY|��Z��4�D(?ƶ��Ad�0Fx������y�IO*{b��eX�I��Ѧ-��u�����1X���D��m���9O�r&K�n��A0+\!�ry2�"O���#F���F���V��h�f\�0x'�ƏY����`�w8�л�PKO>D
�g4
D�eh3D�lb*DD�j�Q�D.��Y{R�2D���!���>ژh�E���]at�>D�@E�ڥ@/����˲<w����=D��BV�\�Fhɳ�G!`��K:D�� D��w�L
�ܚ� �',� ��"O�`t%�0.Z�A�"B�U��Ŋ�"OPe����4��qO :���:"O���o҅Zc&��SNF�j�z���"O`���!_����cֿ��L��"O�Lw��	C�LB��^&'���"O��)�镗X=����=:��0��"O��,d�t�j�Ι�S�B�(�"OV�C�4	$x	�-�I��EHA"OE��7ʊ	�]4��W"O�i*�ʏc~���r��Hd"O���
<L�$�Ie�����""O0��� |��2��\1��5Aq"O�A"Qn5�������UY��E"O��(�D�	��M�)�1
P<p	 "O0<)B"Z4"Fby9���?[$y
�"O|ICs.�*Q��⤢��W�W�p�<�􄁋)�����m[�N)��Pr�<�v L*����G��A@%GU�<A������Sv�E4E��Ed�[�<� �M�?ʮD�@���Ŭ�P~!�N,U��j�S1�8�k��@O[!��۞# � )���1�TУ��@�[!�$�3Q^ Jb��"-� �!��
�ON!��%m��K�_��Nu�T솯F,!�$ $,�Qr�e �1i�K	!�d�&��܂�d�6D&Ԡ�Vɉ	M�!�䐃[?��
��������F[�!�M�q�ͻ2��:��k�̐�!���eU~8ɷ�F���%�g$�ná�$�(4Yz�;���6b�@œ�aR�yr��1|N�#�a�-�"`"0��!�y�,��gD\��铴>���e��yҢI��jM�f�Z�7_��`����y�k1;�`0sO=_�T���c���yb�ߙpc�	��!��M�:]�'�ڂ�yC�>��q T
�0I+�t��C��y"��6��ڷ�l`��-�y�[�xR��f������6���y�f\�p��0Z0+E�^ATu0&�H2�yb"�._�ډ�4% Q�X0q�����y�Ĝ(f�[��_�O~6|���R��y�JY��T�*�@�����n�:�y�ޕ��E�(2����ө�y�^6n�m�D���x�@Q6�.�y���4I8�
VN� AmNy{C����yR��,+��2�	A:<���B�B��yG\�,�!��\9��=�A"_0�y$�e2U{�΃*?��lC�.�&�y⊚i5�aR�Z�*�`=*�`���yR�ByV|������NJ��y#�8T��;r�^Rth`����y�M�<[�m�[(e\�̂�K��y�f��Pb0�X�.I1�9lN��y҇�d����O��U���Q$�y��U6"���ڝ(\*�AC��yH�*'T4q��-]����$�y"F��d1Mٽ ��V)V��yR�@\d�0'Y�`�|�æ� �yb�+�b-�V��?6u@1���_��y�!_-#�~�*eI ,�l,�� _��yB��6�l��c't�~�	��X��y�ң!�*���8i0�E�cgA�yBn�d�*�!c @�X�a��Ǌ��y
� D��G�(��Ŭ��PC�U��"O�Sc'�;��% �,�yD�4p�"O�I��B��#��C��]� ��Z�"O TZ�� axx�֤Ѭ%6��"O�I�gE�P��h�$�(	n�X�"OT8	���pI@���V�5@� ڦ"O�!�3��)��,J4�	�nB��p�"O�a굂ėX��Sa`�`JZԺ�"Op���'ۗ!j�����_�<|qT"O<���A�&q
v�A4/�0A8���u"O��j"'��`p��h�8'�١�"O!�X= ���''�l�����"On@���!��0a�hV1�a�d"OhH���ǹy|:�rť�E�"�Q"OJ��� 73꺱���OĚ(e"Oƥ;��;[2�k�k޵
ת�iS"O ARV�9@LBa)�	}�y�"O�0Å8��a (�;p��u"OҹH�f��m-0X��h�
C���K�"OV`p���Qk�LТ�J8�vq�"OL���"�=M5�S��&oIM�<��i��,���?� 
�(�!�a`��(+ٚ�5!��v!�$S/s{�� �i����ˌY!�$@=m��2A&�/��ae��0Z!��ڏ�����vg�}#�,1H!�D�Qg$��SJL�ȡ��}�!�$Ȼ�l$��0{>�� dǈ�	!�dҎ5v4K��աaC�d�'��A�!���4���Qp�4�ި�u��4=�!�3)�HݢeNY�F��#!&Ý�!�d��, r�ӭ;�$ � O��!�$�)}�,A%��2`r���/�0�!��U��S�fW�h��ʡ΄�1�!��"�X�Κ�7l���X��)�"O�� ��B��>U�Y)O
�I:!�CCHY�d�R.=1�pr��Ȁv*!�d�$A4r �-
<"lx�Ѥ��!�䒀
1�T8���B���A�0>�!��?7w�  �%�%Yu�	u�M�!�D��}Da���9o�͋��׆P!��޴	m�%��=C�C�C�(&/!��4v�ёg�jgX�!�Ø` !�ʗ4�U�R�B!��z��7�!�I�R���{���/H,���C�ʥ�!��3��@p7� 0w,U�FkQo5!�$�7�سǅ܉��`�
�Ir!����z�|m@6_+��KfH �OQ!�d�PP(� c' ��9+�(�H!�Č�7)~x҇��0�(C���!�!��F0[�~��ud�n�n�:� �"h�!���
B,��{j�*M����J�8+�!�4P+䔪�k� ��r��вG�!��/;l\���' ٠�Y'%M]�!� l_��)�+��W�	q���!��L�rt5B����#���`u(؈is!��'N�S�D�q���	V'�+c!�$нZ$.Щ���*uА� ŶZ�!�5Hts�Rp��r�,�!�$�;pp�T��" [B��p�F�!m!�w������
,��TE�48}!�$ի{�r� �L)����1fl!��5#jv��d��B��+���I!�K	o�
� x��ȃ6bս�!�� �P�)c!-��a�2��c"O�,b��N�^�k`Ȼ=.0��Q"O���F�3r.�#�/Յ@*�\�R"O�
4��:yl��rs���W"O���b�?W���$��d� �"Ox�Bc.��f%"�!�D�i�h���"O�1�0�$f_t��(�7z ��"O�50!��|Ǝ�9����08�r"O��@�!�E�(��FY�s��9+�"O���
���^PPk�*��i�A"Oƨ;!��z)��(�K��ӆ��"O�dO�H
F|j�m��e|��T"OH���Jd��ʒ/M
�"O�XH��^iY��&k6��R"OLeQ��S�sƶ�2b�#'�X�"O��͙�A	����F�V|j���"O�8��A~�6iȢ%ߩ&W�ȲU"O�m��?3��c&$��Yv���"O��4���
�МV�Ի[7R��S"O��B� ��|(#��J};�"ONTr�@S,�`��n�SV�@"O���6��.k��R���H�Q"O����X#c0�ဗ�!�A�"O6M��lΫ�-�0R�������y�L�(��T��8���`ք�y����X9��1c��D�L��y����2�N�cVLЉ��Խ�yĖ�nwv q
J-`�����L�y���2pp���>	5b,�SFW��y���A�)�A�a P�3����y�-�05sp"�f�x_�t�T�y���w9�i�V�Ju*����\�y�j�0G�H�P���S�6��R��	�y2�A�P�L	��W=��c��"�y�b�� ݰQBB�\��l���y�*��7�
Q��D� �Y�����yr�A2I�>u@ k�|�HA��Յ�y� ܛ{W\��w�}^��T�׹�yA�7��ձ7d�:\R��SFػ�y�e�6�jB�* ��}a4���y2`SC�A ��~nU���+�y��с�ԙ�D$w�(��,I'�y��Ұ.Zx��ǏS�n�JMHp�&�yN�`v���Bb7FH�7'�6�y2l,2���Fć�f�F���.ߑ�y2nB�8��]�edE'�]��]��yb	�<I0�ؓ�"�x��*ԫ�y2��MMЭ ��q� zf�F��y��_t؂}kweɛG�Xx	B�Ŷ�yB��	/ȥd`L�>�t���m��y��M�t!�c˙� �2AӰ�\�yb�Q*�8�i�'%��p��@L
�yΈ^�h�f
��Y)�hÍ�y��L�*��@A  �B��W�E�y����:��,cV���q��V���y�� �ѧ��<#�11�I�y�K׵F���s�`)=��Q�E��yRJX�� ��܁Z΀yqA'���y�&X�?8��c�5$r͠�2�yB���g�<�ӗ�+$��xA?�yR�A����p�7 9n���	J��y��O�V�M�P�S�l�Z�%����y��rZ@�5�
�ddH;�O�;�y"]��)
VA\�l��M'�y
� ,	�HԺf<�+2��<BFኂ"Op�F�-m
ă�酣^��5Zg"O�̨�B�U�6MF��c����"O���FCE:��1��,�%XJ�"O�xA���x�-Q���	_6b�ط"OL���"���� ʁ�4�9�"O���d��<���9�JL�F����c"O�X� j�=��|�cF�k���aQ"O@��wkݪ
?��P���Y��qI"O�X1����LP��B�r�"O�A�m�hl�򍓗b�B` �"OXk�aU�k�e��+)�Z��"O��i��L%V/�T� ��A�̘1"OJyS��g�����H�+�ؐ�"O<@����%�Y�L{�c5�E5�yBb�1/�������	R/j�C�y�Z���yc��;L]��Y�	�)�yBɞ�m�6)�%Q*F�=�#��yBAD)4H�遢�13D�D��y�OׄnZ��h��(�Q����y"g�Y�������$��m`&���y�E��S�Ҥb�@�&���1E�U%�y"0rZ���Ӣ�=	IZP�d��yr�B7#������x/��I���y�FD� `f&M�Eښ��q�
��y2�)l������8:�� A��,�yRn��=�P�[�L>�A0�?�y���sc��"�A��7��0�V��/�y��8?��E���C1�f��2���y'H*f�<��AZ�����%	�y���xp��&G�>U� ���\3�yr��y�v�j���eB4��H	�yr%�0VX2�GA":��u��/�y2�Xw�j��@F�tR��8�BI�y�%��S��T��i-tb�(�T,��y��A�4ߚXBH�iƢ,�TΏ�yB��+5$*� C��t�P ��#��y2�	�}���	���l��x#�Q�ybK�F]���L2rS@��2�W	�y� DB$v��)Ek�Z�P���y��86Z0p��m��Xt"8�y�)�̱�͖�b��Lc�b��y�m��]�u�-\	 ��U�+�y�拮Xx|ؓ'=D��5�UJK��y��J����#��9���q&�0�y��FH
�iU(16j�8rŀ�y�u��<��%ҕ8p^ `�³�yNڷ�d�â�=���*@��yoK! ��� *�>�mb�D%�y�ޚ'ݲY�� 1����"т�y�A�B��b�K�#h,��3�y��+n�iR�j Mf��g`ݹ�y"ȕpJb��Q��FW�D�V���y��B�c��G�<%v XåP�y2�ך�k��D�3p�9����y�kQ�Z���� ��#����y¤͇K��D�$��#�|�x���y��?�򱃴$&���ą�9�yb횑�1[DJG�����d̜�y���I:�!�qF���rыS���y�I�K ,�d���EJ<���
�ym"
��i`ңHO����$Ȃ �yRG-5u*�F�Ԯ9Y������yrcI�lR�u����7��%�����y
� "dг�%]ʜ��&_�>jL�"O�a��#�D�L�`��*C�x�"O�X���ǛJdΐⷈ��p4  )'"On$!�Fĸ0���Ň�+�m�"O�A0�ݐpb�g@=�DU"OD��3#G�J�`b&��D�nɂ0"ON�{#�?;H}o4R�`R�"O(x��@{��``_&�A"O@}S$D�(�t�#-�l�t�#"O����C6S�z��M�Lz|�"�"O��aևJ�u=r��K�X��c�4O�#'�V�Z��%�QG��&�ɉZ;@�R�� or4�2  �	��#?�b�2~g};���Hl�	�M�J&iBj�qdfL}��Q)n̓L|��A���$��!�L�t�9>�Byc���$��s|@��?���و�T��uH�>�B��Ԉu?�ʝ,���h���3�B�0<�r��'R=(5�@Ѓ��C/�	�?E���*Bn����b$+�m���A"W�<�4@��O%���r�ү��P�a�S�.L<5�{� �&��O�Ox���S䘛j* ��"0�t��M���e�C�S��Hl��" �g�Vq�M��
����<�����(
L�8�ǥu�<�*�*ߏ(����p��J�S�O^���s�>n�9��V^�r��;�	�A��'�'=mP�Ѱ-L�gTN�j�(B��	��&���� qV��Var�*l:�	k��3Z]���ܺ&�.��eR#*z�r�0���I���(��$)�o�<? 0J�Z�L��W�'��(��#��S��OQ?��F ('}��`kFi�F��l�8`�z�'�@�)�<�'/�v92+��j�h��U
�n���J7�	0<Q>��O�(2�Ç-=���c#W�d���� "O�p���� e����ҩ�<x`"Ol���牅?W֠��ҷh�@�s"O�=C��Af�i�&��*N6�B�"O�e0�#P0u�Aã��&��a"O�]��6�V�A�'�H�1"Oph��AOΙ���#k>н�"O>��\J\�
��RݚQ"O�I2�b�:s������3 dʜ�"O�ܓ4�-u��W�@7R�4�"O��g
�j~N�eT,8���h�"O~011��SV��ٕ���+�D��$"O��z gðV��;�Jۮ8�ŘG"O����gVⰰ(C�Z&3^� "OΠI%l� @��N>.d��"Ot�a��%�ژ�1�U�K��M�E"Oa��J�F�:�*U�#����"OLH"�S-
��q�Rk�-&�t�"O�xڶǃ&µK�N7H�Zh+d"O���ֆBBԔѐ/Z�1. �ʀ"O�#�d�xSR��3] ɛ�"OV$�F�&k+����>Uu����"OL,�a�DS�@LH��к,o��`S"Ohe9֢� y��c`��=Zk@�g"O:��e��2O���F&�+:S��+�"Op�BP�=��2��)jB4�J�"Oذ��"Hz�������y�.$�,1�$�60f�1�ԙ�y�l���X�[�"�%�e�0/^�y��.k�r���Lد���a���7�yE��e{�B
!�p��J�yb�C�t�j�P1�l��V�)�y���d!��S`�Y�^����%�yB�Ɉ')ʁ@��W4Z��%`��y�땆1���iEǇ�#EZ4&^)�y����Xn^ KCM�Hz�	�Ø��y�A�0l� ��U�:��9�o1�y
� T�@��(J�ƌ�&[Z`Vd�"O��Q�^s^z�@1L�E�����"On���4�v�x�	�6m*W"Oh�{r�2S� #<��� �"OZ�p�oM3a�<���ؽ����C"Ob�d��% 朚��|+���["O�P�&4o�4�DF$�܀"O6ls(� �>4�G����L�"O�psB�6et�l�vÁ6�(-�"Op�d�ٛ�h�E�%{��$��"O�`�l��X �yP%2�����"O��Ӕ+^$NO"8�g
ЃH��:C"O`�y�,U�j8��B٪9�"Ui�"O��clĭe�b�����&�ި��"O�A)����_U�l�bU�Pp}y"O60Q��,�H%C�ii���"OH�S�F���a��⚶bZ���b"O��#U���7�T=����0SF�P"O���Rm,|TH�`˕
d�i�"O���Aѽg��LS
I�.O�y�u"Oz9�3�IB��@2�IޢkC20Z�"Od����'q��!�)T�T<���t"O(�umU�{#�!��胸L�Dm�"OޡK&�UWf�D��Ǝ�gz(��"O��GdY�r�ܽɴ%V*&Rz	83"O�]�B�^� t����MK�|��q`�"Oe�ŉ[%M�٦l�=�RH!C"O`�@g�P�*������C)����"O�! �
'����b+͒l)f�5"O�������T���"65����"O.��em�/s'ԭ۶hܵʞ��"O���́�8&lD����]�� c "O6ī�<Ipt)G.ۚA�vC"O~�c"������p��P��"O��-'�.�g�t� ��"OR1G@���a��f ,c��$�"OPa��^N�k¯�=� �V"O��q�D��2/�v�Ty�"O�̩6��t.0�����2?�|@��"OJd��N]�f́a͋�~��)�"O�2D��MX��.¬f�Ɣ*T"OJ���eN�g}pb�ƈ*�<X"O�=U�Y�?LV�R��H?6���[�"OMb�8Aq���/\�E
�"OxEC��,G\�qbB��,��"O�����ϻH�mKA��$#�J��W"O��	p��\�<}�$X�U����~�<Y�c�[��\�ބ&�D�"N3�y��ۘ��uzt%����#c'���yr	���U��CZ��&O��y≔�EOбi%�<�ذid)��yB�Ԭ1��p�F�39�D��GW�y��҅u{(qk2fS�,gVyz�L��y�0!`LZ"1��,J�˕+2���(
�'����]'K��TB��S@��'Pʽ�խ :�t�s��S4����'�=ӢW�"z:�q�BܣD�����'��msTΕ�6IZ�Q!�
�6G���'	R�[RƋ��ع#��A�4)����'W,���V	wI��h���+>J5�	�'�~�*d�H�q�<����w� %�	�'
��'�8�J#I]�l�� *	�'Ht%A�لQ6���� �](EQ�'g�����Ƃe�\hɇE4V��I��� ,0s�%�	c�2Hg`�;;��\�A"Ov{�n!.�2!3�/,��uY�"O���6�N�0L��5��pi\1���'ўtK7���� Ǝw��I��>D�X�����i	FI{'C�����?D���0���@��JշN�2��2a?D��(��3/�V ��cS�Z�����;D���#N��-ynA���уn�%ː,D�0Q�N6%�ڼɀ�T*b�Nl"�L,D��@2�;$V�gmS�]`>d�L)D��i0 X���[5D��7>�I�$4D�������J1)2��)-���J2D�0	��ؠ'nU2'����0�c.D�����3=��y�H�Ht��7e*D���	�=M������	8� Ѧ#)D� ��CV:t)B����=?�ސ�F&D��s��K��
���$̴�w�%D�h�@ˊ�Xm!F�+7vZ��0D��A�+�V ��-�*>6�c��.D�Tc �"%1�Xk&j�CV��B�?D��å�з(�F���!��J��s ,"D���g�Q!&^���dҧ<v�ӄ�!D�H���_܎�ٲNw����S�?D�\k���l>��8 ��2`H���>D��a�ԣMݚ9��	��4'y�'!D�,�Lǣw�x���Z��d!�d+D�P↋�K�L �4$Y�U"xݻ�)+D�<j���{n���,֬+Pms	4D�xC���^�,��f<��;��,D�X&W�<�ViV($�����>D��Ӧ�qbh찐�S�𳤭=D�����::N�qҧ"�#[� ;qD<D����֕F�A�SkC�D<�,U�:D�����Z�T�܉(�	0�"!�G,D�`p�i��]un��%ޛ3T�sR�(D��� ���m�nmq
Q&2zT@��2D�P;���d��\�AR�O@�S�(>D����HC�@��%S���/<L>�9�A8D�����5X��m���_ X ��tj7D���
�3�*%���ؤX��%�@4D�(���2Lp��q��!W�U	wc&D�P!Ge��v��:GQ�F�����%D��� 
Hh
T�F�Z>�$xa)D�<
f��
[*11�I��;� a�tn9D�0i��J=>�e����1:��8��7D��[��:{��0���KRu��(D��Q� g�ND���̋9�rZ4D�����J�.�LQL 6�<��D1D�(
@��N��Фb=��H��9D�4��/?4���۵�H�0B�T���%D��)G��(q��4Cq���Nr�,��l1D���G����M�d�J+xdQ�0D���S,̾30��0S�* �1��2D��4g�^޵��mE�9���9��2D�t31�Ҕ$���8@�F�:�Y���0D��HgJ�'Rk�E�b� U;�e��#D�ؠ�M�G&u�"B@'�r�#K"D�̛�N]�W�:�� Y�c�r@��"D�pjF+ j��Ht���?$L`Rh?D��:�A�=K��KA��"1���h*D���3dI�R�9��ܺ_�T���e=D���5��)���MM�#4`�u�6D���&%J��]��(�&4q@�8D��;G�"8j��h�R�l�l7D�� <��
3S� ��D\�aNu�0"OJT n�/#Ȋ�"u��(��`1r"OHy��M�	A �I�%�j0kR"Ozء3��W��B���^]��"O�P6,E�W�0A���<�ތ+�"O��ғ@P�9�ҕJf%�)A���P�"O��u�^5����dǱO�n���"O�=@UM^�qY�
�c� f� "t"OƁ�TJ�q�4�����S���`"O���a՚[ а(�(R:)�F���"ODݣu�I�t8��t'��o�MH"O&���֢f̀�bF'��uL�24"OE;�ȀJڰ����51p��$"O��a�jA��‣�\<p|L���"O�͈���f����-]vj%"O�Ua�N�!% �`bK��WB,��q"O(�rg�[ ЁX@͇�4 e �"O�a���"�p1�flY6[#ܑw"O�Q��J<u'�!�Vf]++�
�"O�0��ƟZƍA�o�N�Ԩ"O��FH��q�
�����T��8@"Oh݃��/uB; ,S#->�,��"OD��獎�sP��`׭�y f�b�"O�YR�k\�V���I�b��d�@�Iq"O^���5:�dq�Mk<�j�"Od��c��5qB�@��hS�*��d�"OP�i�E
N�z�8A.�4m�r���"O>5)���9B<�58҂ݭ��,r�"ONL(',�0T �0�O�)zF�z "Ox@d(˳cV�p(�"��J���6"O���0#ۂ����s�?�`12 "OF,Q���L�����B�@�L$ۢ"O^5�q��0y�j	!5b�4S���Q"On����G�1/N�(�f��S.��"O��2�B�Q]L��uf'H$Hai�"O�iCS��@{�'�$�
�I"O��#�\�i�x��O� b��<�"O
�ZP,]�>fe��m|w�@w"O���K׹*�� �5���%�$��"Op���֧%Y\�3�݃v�Z���"O� �'   ��"H�8`6"O�����׍t��1����4]_�a
�*O��V�Ι�����%$jb$9
�'��BQ(�2��')��&��J
�q�\��Dԫ��I!Wd�?h��)�tE�@o�MF{"	�hS?���^�r̀�p��E{�`�6���-�ĦOހk1e�^���=a����ӻO��]`Bmò)����'�2��i��&�4(��a�i>]�T��b�.e"1 D	G�d���5JDB"���B�xoV��?E�T�k}��	6Cـ�[a��V1B��Z_���h���`�T���0|�w�ƣF�
��G@K�ײ}HQᒽ}vn8bd�~b�,݇��+��I7	C3,<��Q���"G�Y�⠟t�2@9��S9�h bd;�s����u7�Ƈ4.��S�jV����F�ڷ9�jx@��E�f4i�h��m�y�ç0�bhDZ� j��*]�XaЁ,�DЩ�.!F�,�z���U>���1#�����I�Lwzdb��	�x��;��
L����d��h���&D�ZlHů�:x���fc?8lJč�T�8|����n7�U������ 2|V��� y���A�R��*�G��MR�`8L�Qj=���{0 A8CF�(ጙ
�ܺQ��=�Mw(�( �9CA�[6�����7A����7*��[e�<�>x��N�t��i�������g��(��@s f?
���'���+��B�= D :��%\#���8��B��03~n��q�V���А�+M�B�I C��X ��7+��d#A%
Q�B��o��[�ćaL,J��F�R5�B�	>E����B�<h���bB���C�	%/��m������dhv��0x�xC�I�|�k:z����F.J�WJ.B�ɂ-^�&cٍB��壆�@��C�ɑg��U��(M
X��	b��ؘC��8>	��BKU�L����	t6VC�Qyly��Bױ*�dboM�%YTC�	&I�Z��ۛ��L9⢋� �C�	) �����kF)$!�w�
8�B��k�V!����<�@+e�]4j7�C���J9�7�	�`���A��B�I�ur����;{�^�k$h\> "�B�I{(=Y�B�I׌u�Eښ'�fC䉃k�>L��FJ$8
Lբ��X�K�VC�	�����'��{�.��1	�P�2C䉚/�~�-� �Ѷ�ϗ%�L=�Ri/D�pA�J���6fA�,�&��G.D�¦�Y�N�h|� �̴��l���/D��R5�T�Z���jP��np8v�-D��(ƥ�4��|�B�ͦ$4(��c7D��Y��֚�4,X�\���&6D�,��a�-���&�TE���K��.D��R&��])�c�.Z��� �(D�P�B�R;:�y��I]O߼#&D�D�K�j�,!��-�3\Rp,�8D��h$�)V8Ft#J�d2���Pj*D���-�^��سNO�)Z�]9g(D�X2蚃kF�8h�`��M��b,D������ܘ���'i� ��C0D�8�c��A��U �
�&�l�R� -D�h��Ǌb8\�K��A�83RE>D��ҶfI6&ds�����غ%E>D�D����Q�B��t%	�u䢄�C�=D�d���7"v�x��:9p�$0D����c6�=E�I���h/D�<1u/��@��Tj��ɄW���HW�.D�$��K��j��FfHFA�J-D����P�W'�,ʥjZ/>dʔ *D�0x���>Xp��+�8�&��&D���6�Ë4�v	��M
�?UR�hc�.D�� = �bė`���A��ѓf�Rqٷ"OZA�ugԾ7���+���*7~�Z�"O��J��Q=dd@ "��8r�8��"O�Xc�,�Q��P�$鏹6`�i�"OjI1�E�m������&���"O�a�ӡE�'J�гf���hK�"O�h6K�4d�h����if���"O� �p��@Dޭ3�O���T;�"OlLbcN��G�pe����)O���z"O�	�'!J�J�]���
G��%;�"O�h'�5�xA31@]���m g"Oޅ�F�ѝ6T��
T�؝=�*Q2�"O��v��S F/�4��1�C"Oִ�"�t�B|{EOC�(�<E)"O&��q�XH!0����2|�
U8�"O����μc�X����.�)�C"O*���Q�_0A��M�"%Ϻ!9�"O4۷o�14��r@<R�~$ #"Ov z�Ń#HBB0���J���"O��&L�?Ƃ�����8�ʝ�A"O2�(E�{�dY��V��0��F"O�
"'�M(`c'F5�,M�"O�|r
<_y�����M�S���*D^�D{���\f�������jd
���+�R�!���,��pW�M�jS
��;�!��
t��$���s�V99!gg�!�-Q@�;��`9P�5fm!��/o&�K��)\�0��1� Ve!�$۱W��$�Q�Q�f���Yd!��)G$Y$���"�p���+._!��_h��TjˋZ.�J�oԈj]!�䗪 f�h��ͯz����B.]@!�$��Cܡ�Jր]�X�a'�8!�$�I�U�g�ܼck����Ԑb1!�$��\9��@nZ�]Y�ϙ"z!��	�HH�	Aw��;uF�X�u���}�!�N4,��`��c'�� (�'Y�!���~�a� � �y�p!�$�7 � �I���j�؁��%@Q�!��ͼ���M7 �	P�X�!�S�m��*sR@��HQ7�E3r�!�]�k�4ԓ&��!�@�A�bT�[>!�����2�X��ԩY���#X!�W'A˂���efA��U*H�!��;0v����M���q���xw!�d�jޔ0A�+z~�[&[)x8!�D×h���!�_buY��6!���0@��J�Ej�Yv�%~Q!�Q'WĜ��_F��kr�*K!�ĔY0�U[���/'g��*O!��&sc����\�,�t��&��'d!�U �Cg�C��;S`B
)`!��9�`Ŋ��Q&�B�;�oI�!���@���kӓY�f��p��9=�!���j�Db��w:���CO�l!�W��\<B�d�p�r��NR!�a)��05mX�V��X�� S��!�dA_����AH�P�Uk�@�Y�!�$��C�:��	7{z�11ņ��!�$��ҤpB��T�I��ĕ�Q�!�p�^��a�um�k�C1AR!�/I^ ���Cs�1S���	)!�$� o�|h��z�F][�BǦ/!�$G"25���g͸0�.`PR�X�Gj!�� 򝳶(T�u��ci�*n��E"O�c�$�&��4꧈I2D��Xf"O�i9ba`��Ex�gX7� �b"O�`��x�L0u!L�cİ���"O��âD�/z�ĥ�s��.H�(`!#"O�4 ��]�6�ԕ����eR�I �"O0�r'�ҭh�X�l��j=���%"O~���S1C^��
��ҿ�|��P"O��Yp�K���a���"O<mA&(,LJ�mt
�6���:"Or��O+n`��Ո��X�|��"O��{��Z�)��bƋ9"�8$h�"O�䑕F�g��a�1� ��1�"O�q�5eV�T'�t�� ���ɵ"O�9��ʥc��l�e�4�84"O�ܠ�ـ?��TbE+	���h"O�=0�_7��q�e������"O��͕#J���a�K	a&�PP"O�	���8I1�PH'�1@!�d�(��$Ek+"�(�-�8�!�dY0;���u�^	�i�$f�L�!�$�^�H�(U�XN�|U�C����!���1��g� U9����s�!�� L~$h�ę�4�Nk�(V��!�d��!֐�C��0�l�i�Ѿ!���:)�4�X�-O8C�0��QT�!�D��"����%Lx���U	W�FC䉜z��\���������S�U�C�I5w{PM�eS�u0�W� 7TB�Iu���P�+U2i�׽D�6B�Iզ�I���{��Ѓ�(�@C�� <�xc���2���SW<C䉬`�8"!�х v	�JxR�a�'Xq$ǆ$A��%ӵ`�M��5q�'�ԭi3��;_6���E�%JR,��'�
m��a�<PC��e�Z <Lʼ�
�'<���$92��!�"�8/b~)[�'���JAɮ^��y���;*�څ��'����A�˦�c�ON&���'�0DK��x� �Iҍ�I����'+�E��M�6I�1 ���9	�t��'�J]���O�_��@h�h�1Y 8�'��`��!=���G`П
��Q��'װ-�� ̲8�VI��Hn�0��'�f�"&��7a�f�AG�<a�Qr	�'	� �O��kq$r$F�GE�M��' �I�dԢ-�`#G��$��'����e�=`5"�6c@N�ŉ�'<C��9��v@@(	� Ph�'Ԓ�)��M672�����8����'�<���m��h-�e��F����'�r��P�ϒ_X��5
�
�s�'��)sf��s'DT�G%ד3~�4��'��h@"��0��c���"t�ȱ�'�T��`۾SL��a������'.ļ�G�0ⱻ�dŰ~^��S�'G:!��bD=L٬|@l$q���z�'���S)�!��,K%�!\�<,b�'�<�x�f!Aɷ*1b�@%���yHH�µJ���6%e�0JD���y����k�7e�j �s Լ�y�IJ!e�>��3��-XgFi���y"��Dm���Z�Q���ӵ�y"�T�c6H����(H�X2�
�y
� ��B��w�4R�(�$�d��"OԜ �*�>@[���)t $ �"O0�!d-��O,J��iA�,��a("O���a�vt����0f�p�Q"O�=h���[gVQ����L�21�4"O��x��۱Ef )��͐(#ƀIu"O���U����Kwl��K��,��"O@�K�n��Q)�L��+��c�|��"OF��Bd̞m3ЭЕkJ��85�'"O��[ta�t�̸`��B`�W"Oh�#�I�1J�<���,�l��"O����3N�pc���(m>$å"O�d��'���#n��X#C@�z!�d�-���
����J�w�!򤝺��ě��¯:r��I�oܢr_!򄉔c� ��J�O��q�5o��&!�4;X��%bϡ lDp���H�J�!�dQ1R�n�2NP�[Xൌ�D�!�dR+��q $�H�����W�T�!�Ds,��@�Բ9��)qQ��W���L�7U�xġ �B�\�8v�M��y�D�	�̈W/�;0�<X�eR��y��4a��4��i8$�n�Zq��yN-B��D`���9��"���yr�#��e]0~�Mi��(�y�I�K6�뷈�.M ��p�Ĳ�yB 
��x�Uǐ ���B�OQ�y2���/��A���ϋu������!�yR�0|�ޕc��O'@b��{'=�y��˰8KE�F5�ة�gù4� ��ȓ:�J!N'��dQ��Wƞ؆ȓn�1т
ȟP� !��PZ]�ȓx�l����]��h:�ْc��i��'��h���$j:j<:$l�ivT�ȓ��� @�?�     +  �"  �-  ?8  %C  �N  �Z  af  tn  �t  �}  U�  ��  D�  ��  �  <�  |�  й  *�  n�  ��  ��  2�  u�  ��  ��  9�  ��  ��   c � o >  & D, �2 �8 r? �F �N U D[ �a �h �n Bu �} 1�  `� u�	����Zv)A�'ld\�0�Kz+
�D�/j�2T���#Ĵ���+�?YV̒'�?��]O+��yk��P)�T�pH(�����8��)L/	����'�� m�E�e���S7X����1"���r��=�ʝ�A;E��8��/ xS�'S��pH N؜3��<���:`��:�f�ǰ����(4lc��˻Wn�1���X3_�����i��A���,D�r0o��a��9�I����	ݟ���/|�^Adpv$����\Ӑ<��>�e��h޽�Ms���?Y�� �F�����	�1IR��t��-��聂0K�����O<���O����O���Rk�N�}�,u�BLҔ7�Rh�#��pɠ����xL Г7ͥ>YN��7m%�,�F�SB5sO���B�|���a"�+���~��&���!j�)[��� T�瓏.Y��X�O� A�Ձ�*^`�$�O���O��$�O��d�O�˧�y7+��6���Ŭ�j���♂�?�s�i��7M��QQ�4�?���iF�	Dx��|1�@B p��x1*Fyn*u(�&�=rH eHUJ�F}��bӔ(�p��OVip!
�yoTq �fɽrI��sYw(��!Օo�d��a�ϧ-�N��
vh���KV�I���&)��-bӮ��?��SԺ���%&k|	J��<�c��>* il�&>f�HR�Ł'����K���c�ʗ$c@�q�4tV�Gc�d���E�A�PU�1c�H�� �EQ4��С���o��MC��i"�����d׈�[�g��g�r����۽L�C�,Q$
�ه�ő\	���$O1t��@2�pӠ�lZ��MS7fL�C�29Qh�= ,8���mE�/�6;Oq�⟾ ��-P�<tH��ؙQ��.�<0�o��F�%�;���'S�&��H&, Q���|�����'�O|�D�O@���Ŧi�	��D���є<�A�<@v4�oD�X�ɺn~N��	��	�7�F�!ط64���O�0�MS� M�D�♁e��t�U��@�/Qi��O�'�(OH��͆
ȠX�����k�6-���6cT#��)[d"ē0��mZ!���<Q᫋}y���<�d�&��
a$�-'l�!�,�ܟd�I�D&���	럴�'|�"�"��9��#kʜ�A'N�^��'�|Kq��cr�'�t�s��)��|ҵ�ӐI���7e�K����a��O"�I$Њ��i���	t�mC"��O�����һjά\3�
�O��N˂M~���e\	]$����4��O�F�Q�-�'*��$�D_b� �@��`���؄�@Ӈ��R�E��`��$�� ��G�
]�­����2{���{�ΔE�d0�*E�7��$( (��E莘��|��'�B�'X?E��*�� ~��d�0-:�y`0�;����r��b>�i�-`4�!��ʧc���[ᬎহ��ɟ��Ɇ.�=(E��˟<��͟,��ڼ�qk�}Xx��O���!s�y��'S��au�'`������I@����~�hQ�!�|�,���b|�0�I�I�69�1�1O�)��/X�>S�5q4��pXBB�V �'�]H��ϟ�'���A�捁t�|MS4�P+�㘝8r�)�5�\��i]o7���_;&��{.OB�l���M3J>ͧ��.O�,"�/�l��=}a����(�"w��T�'��' �	[�4��
A�cH�(d���h(02�1~)1�G؂f��!�m*<O���Ȕk���nˆ\V�({r� 3|J����QZ�|�6�/�@�����D%CD aX�hu+E(�����Opnځ�HO:�ب�/�	V�]��h��V1h�ӟ��IƟ$���Y��yx��W����AӦY	B��Od�m��M�.OJ`@���ۦy��ܟ�����)T�	6��?.Ve)�kӟx��9Rg2��	՟���;B"ߔ/l��(�̇�;�z9�r`R����a���V���r��CF�x� �1�E$0L� 3�J9<�ĕQ��*ۮ|ZrퟸTZ-���P�!.�Q�!+~��!.0�$���H�4�?Ydeχ	0��f�A�E8����ۘ��y���	e���>������$X����m<���U�2<O&���<�4�i1�����
 �N�#Q�_*u�T@��gz�h����I�j2�,b�i]Iy�O�T6-�HX��Kb:`�s�+D�W��b�d�O|�$T�PɈ܊@ �4%X����RV�=J���Ô�,B �*�a�F
��HU�9K�	-y���؂l�Ds�C̿i�L�תO/ϊ�����?mE�P�h/r�H&�)>�|1:RD3?q�Lݟ�{�4��O�1�⁒�AP���1��ݧ$������|��'��'���'��I'#P ��^y����% ��q��ҟ�m�����4�?9�ϒ1P�|��k�0w� Ճ�Q>g����'
��'���E�μe���'���'���]x����PCH�u�*(�d�S$w6���,�84J6۔_�T��B¢|�!�$>F��L"�����Z�X�
ub�Ĺk0Db�+�v�,�v�)ư���V�J��҉DC@9��+����o��]����'�B�'��$bĨop�I��[���֝|��)�E�@9��D����	 e�ʓ���nӶ�O��)�0˓׬����N�.Z�m� ��7��݊��.|����'��'��IT��6�D���S=q̠�l�V���u���:�rtFB�J�T	&�"<O�!c' ޕ�!�R	j�|�pK�7��Fֻ	��0EO�1���"��!:C��&��.L����aꝠ
N�ы��OH�n�'�HO#<U睤=mVA��6L�����̟&���	ȟXF{"�L�?�h���@.��Q#� ̨&�"v��ė��%"�4��O�;X�o���@�T$ A
]<�Ȱ�c��N�(Q�	Fy��'sR;��43$ ^u��/|��7!� ʔ1�kV��r��aS���'z��AnՎ3�,����]�w ��F�wC���#H��L5r�;	�a����<w�x�40�'���P��ɶ&���M� �b��I>y��4�ɱw܌	0@+�k�F@`�	� ��	�M�3\yL���ae BR~TY� @�Wh��V�P�c�G�Mc���?1(��� j�O��ˡLF�䬱B'�B�m�J�Z�o�O���X;H��VK֒f+zٛTE ,e"�Jfh,����O�j\���˘n+�q�W��=c ���O�l�È�AG�D�P��xT�0�!�M��~Z��<t"�H
1��=(h�a�j4}2B�9�?�&�i�.6��O<#|¡Ʉ=�ŰR��*)�({2��ǟ\�'��^��ߘ'���"%E�Q+�}���&<̺��Ó�Mr�i�{���H�&xDrBD�|nha��v��nZ̟p�'��	%�O0��'��^����H
aG��6bʱ#�ni8�cЈn0-��n��
���m�(��	Mw�Ae��	�I�ip䌘�� nj!Z�`�W:���UA
rD�I����v�'H%*��'͖	[��[/po>!��{E�3䌄�m�.O\p���'��$�?�O�$�Y� ۰$R㯖�oG�<�C�O���<)���Ow�ɩ< �����Ge4�I�L(��ᛦk���]�}�O���_>����S� �d�XRN���@[l��L�֬���������?=��ȟ�ͧO�T,P��I1�<{@�K&f�f��\�!�8�0�B��A��*z�l�F(�
YoQ���6@�;{�F`�@L�q}he�W��(ؤ��������xDA��{�,��˄;M�Q���dM� @r��B��I>�x��3�O}X��Jh���x!�Q�.�F�R�,T�
�����j5LOj�$�rf��ep\����m��ɹP�8�$���'�d�%A������� �6�_U1|�ɥmӔ~:r��4��R�'�
����'�"�'�Aa���k&0���,ާE zeX4gS-i�\�ۅ���NJ���1�	V�m���H��(O���C�^>v � �ܐ4V���M���ꝈSgO�4'±�&"��l�9����(O<%���'��7�[����	"s�)V�#9/����T!-8E�'s2���#�\P�����n�Tڃ�N)�8��d���	�#T�8����>�r9��c���M�+O=B�ϙ䦍�	ϟ�O�je1&�'0����>^(�1�&ٯ6�̐kQ�'��cT�}�EkB �5@�X�jP�dN(��W���Sk%� ���P�}#Rя^�n�^|��b�%�D]��KH]|x�k�%$[+6�O��@�4J�:)aL���,A��@s�OȔ��'j67m�l�O��i���iP��C�c�t��'M�@S1�Oe��X��kO,R�H����*�Na�fIl�nc>�@.�:s�pJ P!mrD1���������X�	; K:�s'�蟬�	�����Ѽ;�㌺G� IB4��2A'�j@��*I<�,��M;
	�IdH�x��T�i�,�'���*uGY
L�e!H2\��\zюR3`�b�i�j�(��ݗO1��6�[!��$߾=����J�9>�F(:�lEB�ԓOH8:��'�1�1O~�P�T�D��r���dv�J�"OНJ�jT-�@��C�ip1���'�2�;��|*K>��ʜ�G}�`3'�H�7z��!QON�g(8mh� @��?���?���H|��O��$n>��w��T�@ȊwU�_/XA�u.�>Y�"�1�	�h�U���\o� P����D*~+��`��g<����B�1r��f�q>� �"A^�N�����J�ir�ma��D�F8n��2�F3#Z��#Kׄ&S"}K`�'J����	7aj��䠗��h�ȑ���2!��[�O)��7�Gkyr@�V�)?�'��7�4���2~��OR��wJ$�G�^�a�yZ�g�<R��'�����'r"3��at�l��ЁH'b��ؤ��M�!9G��	�5������t�?9��Ҧedf@ ��ȥ}
 ���l��pB0/��U��@iu���SHD����� ���'&��&$�
�۰���bǈ4|�h�Is�|��'�az�CVkĤP�D�J��N� ��?�S�'�$8�Q��!>�@)qҠ =)�����@�W��l���8��A��a���RÕʂ=2��Ǉ2�SD�i���'-��\&%/8��Tj 4�N�3�D�~ʟ�|x�bI6{�X�œ�Z&��W��h���<)��h0S+N�8��� eo_Y��kOD��g��1Q`��ᰄJD��'������?�����Oj���D��Y�&��wrf��
 D������h������-Q�dRC�:��/�>���'^���*��0H�bަ�����4�	�$H(��b/��H�I�������'��$e֭���]�NJ�P9 �3X��(�`Y�+69Pդ�7 �\'?�y6�ƌo2��7% 	�w�	�`� ��%\
�Qf�-N T�
Q!�/u�t�@�4�654����ORU���I b1�3�م���DFu�@5�'�(\���"ϟ�'�+bK-~,H�e�"�E;P�Mfx�,�b��#!]�˲��\²�I���ɦM8ߴ���|:�����_]��� ��4gLQ��C�q_�+Î�?=|�d�OT���O�����?	���tJW���p1*A֐�2j�'s�v9�Ӌ�� �R�ȣ���Ƅ�{d�;�}KĔ� N�jp���o�pmiR��5Ꞩ�$�I�!�����ڍ6Ͱ�;0(D�JNk������=b�(ݓ2���q�x��hI��'�����R+= Hr���4-�:��mh�!��'G����Iׯ+fH����p��'��77���(lC:i�O�R@5Z8���.�6�� �R���'�Ny+`�'��=�9@����X�r��B����E˃z�
Ń���:!jLx���<oh�E~R�)z�
�Q3eFd�e9%A�O������a��9b�1� #���a��Gy"j�9�?������M<!�D�D� �+֣
�(D�'�a|�nX�`|t�%&
�7�4��A��6��?�!�'�@�j�0���W���<Q���$R;4~l��@�	H�TɈ8!��Z�t@��E���O��"�'��EJ�'�*['I�4r��k��W�drn� &0��IS��?us���P%�T� b�L�U�b)?)DǊ�Kg؀�s匏XB�)���Xu�|�dF$�d�(VDzS�� H�����I���D΁A'�s��F��2�d��l����#'��6�Ba��"O0��fZ�g��$��-
)=�Yq���%�h�b`3�ű\b�T�ƫJ*'�ʴf���d�O@�$P71��İ��O@���O"��~�E�Ǆ�T��BJ����ݣ��ӭk�fgN¦����ܿ{�B��|���"O����0$�t(�bL"W$�ӫ!y�ʑB#lK�*KƔsr%N�:�2zwI�)��'F��i(��3�I��J�f!�0�\�j��Tʂ�M3dX�(H3L�O�� &�8`U��6�2E���U=P���Y�<�3��x�)�(S ���p�̒`yRI'��|���d�>����ۈ7�P����Jq��a�X�sE����O��d�O���;�?�����t J�\
5�Y-f�*M��i&o |
�Gݚ>cZQ5oM���(D��Dere8RA�d
�G��(97 S4�qb�'M�x�V�>~��p�݋Pՙ� �;�?�Էi��6-'��)��O�����Z/d@&���zs��ӓ��'��1[s���h0
ӃL�x��AK>�ľi�RP��ٲ��$�M���?��ήV���F����x�<�I����͟P���|r^}�I#��\�� }*��g�Z@��k�]08,�#M�]��0�a�Mɔࠎ��\T8��ҋ�y����䅏w�6x����p�V�P׮G
]�吇�<_�x�z��dG�G�r�䇾�V�I�'��>�xujs`�;2�!��Mk�Ju��ʪ0�� ����6����O���]f�@U��l�d1�xI�|���t?�6��O��Ŀ|�eo�?ar.�4�1�M�]D�ݣ@m��?A��:�FfU��<����@T?�O�S�%$0��#��bW`��b.��{��h�pl�P$o���Sb(�'Gو"5*�?/��0PS+�%8DZy�'Yd���?s�f�1�'�2TƼZn��F틕t���ѓě�y�� r��c��n;p�hSf�,�O��_���)U�Ny"��ԩB�^#���A�M���?1�}k��R��?)���?Q��g)�j��ٚ����ge*�`�Bؔ�H���Qt?9����j�|�<!�U��d��Y[��K�+�75�R���ģ��Qh_�c>c�4�! ֯ ����h�
�qE͜�e�-O�L5�'���O�Ob�q鈪�>	2�+ӛ&~�-{�F!D���sOC$($��+s�\�0Ҳ�V-TO}�"�/ěv�'������ �6��C@
|�9"4�M�U%�Y����(��矤�Xw�2�'j�����Hf�Y's�Tz2�Q�hLH4��W�
�;j�:�p=)4 X;)Y���3s�x��E(_�_�đ���=N\*�zj+\O�i��-m�Eڱ@�6{�x��@CſV2RH~��%l�n��q	񟖘�rL#�%k�囡��G�f���2�ɋ<�(���B�a�$(�a�?+%X�O�ml���'���4��~���X$ $��Jk��pG�]g:����?���
�?����j�=��0ƪ^m�m�'��z��8�v%�sJ��3Vꔅ�I�+�!x�-asD9�!�O�@P�h�� �j�����X��	#d�'�2!��3웦�<	3�.u�5��$R��h�"�U�I۟��	�,��M�%́cJr�Zv��Q*�c��F{*�����!��0����� 5��D_a���$�<�nk�&�'^�_>yq`J���顇[5Y��mh��P%*7�T1p�[����� ��ɣS 9pE�SaU��M[(��ʧZ�����t'�ų4��o��`�O�L���Be 4����O�� C�
I�x�1�H2m�-z��� s��=	p� Y7��,9A�O0mZ��M���� ���	���ޕwCReKa�|"�'q�'�� �P��3s�Ҡ1�C�B���(�z0��x�<�O�u�#:2�� �N�J���G 1��$�O`��ӜDh�(ã�O6��O�����Ǘ<5. Ba�����Va���y�'���C��8k�ϸ'�*D� .,�� L�ڱ��L�(>����v�Typ�� %S1�1O� �`Yub�	$.RL�B��RX��m�rx�'��x�����ɟ�''� O�,��6m�:9z��Q�q�4�w��iBv]@@���bԦ,c3ɶ<!"�i.6�*�4���i�<���8B�����z�ir�`U4%<m`w�X+�?a��?�� x�n�O��t>Q��&�<v#`��?���I#���x�� �
)$�$X�W蜈�
I';.Q�4ˠ��/:��`4�� y:T�)��!˖�c��VQ�9��I ��pa��48la�?���$"!�\��#$y��6	T^�������E{�)iYM�gNT������5�<B䉽)$J� �W3޴�1���?SjT�OJ(n�˟�'�n�WC�~��u����EK�;�V4��Ή ��!����?��	��?����ԠF5y�B�+���:�j����i�0�	c��iq:l��)CSV0)t�΃0H�Q��Dվd���O!g6��`�b�B�����q�n��c��U�(�'
}�k�@�c��]�IꟌ�'w,�6�E	񄡰4C�#J�}iO>��w'�E�?�r$�R��dq�ȅ�I��?�@���q$!��'�b?��Ku��֟(�'N`8h�.}Ӵ��O��'oĲ)S�a?fġ���L�쑖-���d�����I""$����N�/��L:r��!��%"�@�)Xp�O���'�U�2�!Qb�S���OZ����I F�.7�W�L$�XCU�;�0�$�Tg�tBI8p �Q���Z3h`����2�'՚��I�M�D�S�|Z�	W)�H�[��ց:���!biXE�<��I��\�V8�NB)DKx��	y�'팢}:7��cA�@th\��ib�l��M���?)��4e왠Ȝ,�?���?����y�A-^��bg΋f; �H�튫2XZ�KcBU�XiA��bڔ�S��䇟�X�J8��BD�̳��X&Y�K�nA�4��]G��%\D��f�v�k'�P�L��c>�$& {��ē�t�,��N�0sFC�S�7�Cay����?!�'���|B��4y�څra�H�L2�<�L�Q+!�A�
��K�0T,���#g��(O�Dz�O-�V��[��/�QQ�$�
��!�7 ;���Z!�[՟X�	۟@����u��'�0�b�~9	��ڦq��"dL�;��ayc� '��u���W�'�	��V���Ey�ŗ �s�U�
������Sf� �R���`��s�Ĉp�
ŋ6�F�0Gy��3b_����֨(H�����u8��q8�b�F�Iv<E�-�>Wۄ�2�"���y���	$�t�R��7E��@r�`ߕ��:���|�Η.{z�ꧥ?���0
.�0T�8��Q��&\��?!�Q�	��?i�Ok�q�旙��A��W�� N��w�H�S�jӂ8� �3��=��I��h�b�'�N��,�
g�0��C[��`�شBK�B����E3�钲ѦDh�H��EQ�',\��w���<��G�*
bA2���.E��ɓ@��S���`IǥM �D탨qc4��f;�OHl�	�d�F� �u|.$c$QTCH�Į<���FR�&�'a�X>�f�	ꟸ���sSHI�cN̼V8ZUb��D���	 �L�g%Y�*X#C�֦ACQ?Q�Oa�)����Hi��)\D0z�OH1�Q-٣6�dj¦>>���T��Y�i��h"V4<�&m���G-R��	�ix@�$Ʀ��M|*���*�O ع�D�q-��h@Ė�5A6xKN>����0=���R`'z��@m	�TB�����s�'�b�>	��4�̗���3�-A�9'�apƈ��YR�F�'�B�'��d�6k�)	��'��'��n��7�tz`HݮbTqA`KZ�S�j��a�ɺ�
%�u��=�|;��)?���3� h����%`G |�El]���ؐ��=>.�e��e�% �i*��O*X�4h�Y~.���f�!5�r������O��D�O��<�&l�g��l�&)�I�t`�F�N�<�2D&x�v�� �R�Vv��F�HyR<��|�����8��@IULR�V+xX�C�A���wZ�c�>���Ox���O�E���?Q�����S�]��-Y�mْ 92�1��J�TT��N�"��}p��^+&N�C��ɯtV��`�:P (h��B;S�| fA�7/�04�M�q���s�\�'ؼ�2��>5D�����6��T��.��?��?	�R�ӝlٸzu��)}l�@儆{��C�I+5�|��j�)>\fԩ�(N羓O�)nޟ�'κ�Q�l�~��;8�!��/���-�B�<D���?�Rb@,�?A����G�I�D�q+�s���14����@�GမC��D�"`��E7��-u�9b��Ժ=2c�ӂjw��:n   
�A��M�@�V 0�ӌ��O�$��'-����o�-2{����e� 8�xY���&���Ov��2#U�4C�H�
r�0D�ʖF��k�O8lQ�eS<�x��Ɏ�c�Q��'�	�F�"UR�4�?������:�b��J5�&�)T�#>Y���45Z�d�O@\@�:A�R�B��F8�*J�T�?q�t*�4��ģ�О���r�H(?u�׺q��[�5�e�ᜇ��O��(�둘��!�S���i'��h�O��C��'R�Ɵ�� T4��lM�|��r &�cǢ��"O��B�NX�B��@�ݥL�B�2�	��h����De�,+5ڙo�+M�(��}Ӽ���O���Q�L������O���O:��{ޑ��Ț6��h6-ܳ"<A��9�fu(�K�R����&b�c>!&�D;�$��H��`��Y0'h�b�cS!Q'xD��n�b9��A@̬A[vc>&�@ʂDPb�PR�K�bӜ�ه�`�I`Ӑ��:�3�I�2Ӣ�a��ˆ(қA��C�!;L9���)Y�|�B5cZ<�˓X����O�I�1HR�+#�.+l`�H3F�v�]� "ܳ;-*���˟\���#[w�2�'��iJG��`0eN�4ym�-�ѣ�%j>|	Z�k�`�Dؚ P�p=Ɂ�U+uҾyBf�?Rƞ��P���)S�+���Mj�
5\O����&F�UA�d�0{~�9�a�%$��|�p�m_�Px����7��B�t�s�g�?o�"�he�';�O<4���+d�1�v���tȜ �|��z�����<���A8Z����?�@g�ӳ_�Z%���#S� ݨ�o=OA[��	��J����2{�l�JL#zk|���?n���r�@C{���#Ah��~����H2O<��f�'�1Ot"��L(y��)R%0�J��"O��ܷX���H0ElR�v�'���d��]XIh����>v`he��-n��'�F��e�'U���O��'�����:HF]��AX~К�j$��?���NZU��k%&"0 �M�=/��� rx�\0Z`� ����	-Wjf|1Bh6J���ŉW�O]�����/%j��]�Eیq!�OD�2�'�b���<���|�V��J�������X�<�$���!�����I�F�vL�Ō]T�'!��}V�ј&����	Y���˦��ȟp��`�hy���!q22�O�R�',�ɘ�T���K�6�K��c �,	�J̙+��h���l_�DC�I�g̓g�r���MG *�S�e�pP KE-^M�����7�ub��i�g�ٜ������~m�<:T�ie����e~�2�?����hOH5�5N˚��Q��1pc8e���1D�ܠ�m�>a��(s R}t���<YT�)-O`�!��>8��q�X���	��yӦ ���O��ҧ�C��v�L��4AEh*�ǿs�'�m[B�9A�5<H 	��Ģ�?q���?A��?٢�u�X�"�$�� �D��>�Р���x�̨��+�<�`��p-ގ"�@Gy2�)L�(��-@� Ҹ0`"k�����*TbʜdѬ� b���9`/�"LxtDy��G�?�@�ioғ�����C�Rl�h��|�J��R���	���p�U�6*$��p�Z�/��$�xy��@�;�z�`UJ��l>�ɻ�KD����N�4��$őnF$�Ħ|j�G�?����檀S��L�~����B\m��1��Ԡ�΃��My5H�z�~Tb��D�>0������e[�	s֨�Z���1��X=�y����S��Q�&���)�TU���ǃ^>��EN�V�'R[��yOT�J_�Q�A���0(H��$�DQ�	��M3V���R�'	�nP�`
��`�Zf�M�.`��2!�#�_�E���VO��KAD{�n3�{r�3��մ+Qʭ�r,J�F�80�ֈA�?��^T5��O������?i��N��.�Oh�&�ږ(�bYarÛ�*��`�
*V`Հ�	[�&C�!��k6b�'#��
��:}B�W(o�
i���BӀ$H�!фR~�]�e��;|�(�Q-�#xRΟ��)p�����I�x���%%�$L���R��7<��J���Iӟ�F{�:O�){��'������-.2M��"O�h5F3{���
�F&�I���'�:#=�'�?�)O��X�.�!8���Ƣ��b��VVb�b�8���O ���к��?y�OX����K �Ʊ���rip�)�h�x���ۣl�
p�1A����r�"?�ע��R�<����e���h���<E���b��\��|:�IKb.�#L�	��<��O����!(��Q��%��	$��O��=����X���:Ђ��8O�)���;h�!��Ƭ0Z��D�ԕ`�����˼]~�Ɇ�M[���K�U���Bk��$i>%�B���^�Ɛ;���^S\ͻ�B�O`���Ot���O�d�.K�[�:�[�h:@Q�����������JZ~`�PƖ>R$�{c)K�}EQ�$��}z����b�&3;�dz3��J$�c�V�.2�M �sͤ�"��C�Q�Q�X���O���3���a�Tː3I;*)�ve�@ʓ�0?ɥ��){M�Y���'lĬ�N�fx��
+O�L�C��^7Č 
�:)�!Q�^�p`���\Cq�V�L�O�	�S�O�B��PJ�E	.�:p:�p�_7a����j��X��a߸(B<�Z+	j,:� V	˵q1�p����)	��#ֈH�tH�y$7O�$�#r�D4��s����2},4R��t��\@@��Qn�5C���QQk���yrdD<�?���������� ���D���"�"��&~�K#"OZ=����8��PI�Ҡ�r�	"�ȟxu�c'�`2�9�[`"(�����F�v���Ox�U՜���O����O�I�O!�sg֐r-��"�Ǹ}���6�N:
��(�� '@�����|"�6.�PaTi>}��0l��*��=,�6ẰL7_!���˽)Zb�+�M�=<��P�Ο~|�V=��IN�@$K`�_�0͢�.�" ���������G{�?O�!r���S�����q��-	�"O��w��o#�m�G($soQ�V�'��#=�'�?�,O�D�������KB��0<��0��= >� ;2[+��D�O��D��x���O���JMj�J�,��}���=����Bk�"�q�s�K�eУ��ծ���I�8XͰp	��1F���Z�
��r$X}������'rr�������6�?n���ǉu��	�Ȼ?,���� `��?���O�l�L^2A0�ass/�4X��d��"O:p8��^�FM��A�^��P�P����4�?�.O�U�!�Mצ��	���'	��f��q�J�w�)j�$�	?Wr���	��I�*aa��l��|B�%��Q�8���$̃g�h��m�z�'�f�R��I�I�0��=�4��N^�|��4��O����h�yF��蓛Y
�`+�[[�<a������P�D�|�huoZUx�0�*O����k�d *�(��R����џ��ISyV>��O��
��Tz��G�>�jͪ�O�П�'��S�'d*���%� =�(���C1d��?�ش�ēh�d����F�2An��'� a�`����٦}�	��MϓW\`�	������͓1@ҀQ6��V��؉�o�s�aP�N!�M���Q�����y"
�������7џV�]�[N�!�p�˾i@ �p!��mģe�'B���?�$`�%�I��(�S��xyt��"�%P��7*D�& � ���?Y��}�L�P���2�������/?�ش|p�]Yw쉅3��b�
�$:Z�dtb�'��Q��Š~���?!���?��,_Jq��F<M�,u*�% 7N����'�?��`X���XR�����ܴN��y����ҹ�$C
M6�B�"�,O���A�O�LP�'�	\��$hݽ���P��E�4����5�
	CH�8���@��^�<iQ�������u��'��D�!���is�j�(f�Y�6� l�S$ȓ;7���B��dw���b�4�sC�OP��Y0��Sğ��I�8g��N��2 ���=r��4g��e"�'8�̰4�i�6m�V��HΟp�����?Ur��Y�'����U+�T�A��V٦-� 4�MS�P�ț�'�M���O�韜�,H�P�s�#K�B��h�q@�X�<٥��1	pP�W8Wv��E�증���x�������ߟ`���X��˟����<qR<g����L�-o 6��O����O��$�<���?Q��?�ֆH� ܞt�5��@��zf��x��V�'��'���'��'���6kJ�mPW뛀7�Ő�)K��6�'���'�r)�~r-�f�'7���F̈�~0E,��3�̱�O����<������2� ʐU��!��ЈO}\�3%�3��O����OR���O�ʓ����>%����)Y�>>�%s`�
��$�O��d�<����5�T��u� ���gq����׊�y�ϘxI�Y�!��/3��l+�Ε��y��O讍�qO�~~pU����l�<�#F�u��!��Ȇ{S,Y�0�w�<Iw/˶e8�: ��?)���"e%q�<��@�-�P���	D8cK�=��,�o�'��'#b�'2�ϻd�  �EтO�Ѝ����Ab7��O^��OB�D�O����O��D�O��$2L"�`#F�1N&��v�q� =m��P�������՟\��ן(���������|J���-u0��S~�rU3ڴ�?����?���?���?I���?��{I�9��5{�rD	�qڄ���i(��'"�'2r�'82�'���')�Y����Od�eK�� 
�"�(c�@���O��d�OD���O��$�O���O��F杼Wyؔ����w�(��6���u��؟��I۟��I����	�������nFfp��T*p�5�� W��M���?q���?I��?9��?I��?y�o��m�Y�]���ٕ$��m��T��ǟ���֟��I�P��˟�ɏB������*P?��b��%�4E޴�?y��?����?����?a��?���09����".����*�_<: �i���''��'��'k��'��'76����Y�Ar���d*�A�$�pӶ���O����O����O,�D�O��$�O`utH��Q� ��m�* ��8�Ԧ��	��@�I͟p�I��0�I˟8�I���mf�d�C��G!��`g��	m�`~��'��Is�O>I�dX,\�Z��t+-Z}�\R��i��I��yR�IW����w�T���JQ50�$ ��B/Mu��x���M�'��)�)�H��a���O�$�)��sBM,���zS�'��`��0#����i>̓"�$̋���<S�4�+JG ���|y��|¬oӆ�"��d>� .�a�@E9p��[S�L[ژ��3��ry��'
�?O�˓+$p�jf ��n2݈���_mL��'��U��R�34ry��O��Q2`�j��t�|Y���7t��u�s�5^�@l�2I�<y/OB�d&�g?�g�V<z:(�lK��Xl@�`�ǟ8��4]�d�'�6�9�i>=+�C�6��'+ʎyn� ��0O���fӂ�$S+2Vڜ����h���ގ'� Ѱ�=�BKÖ� D�Q3 W4��C�I��Ԗ'1�&hYc��z�c�7MI$�4Q�d��4[��`�<1���×'?�n�j�N�7_z�����{�tʓ�?�ڴ�y�铞R����$+Q:md*���A�F��<�1A.N�n�9���"��1^�d�@��$��l��8��,I�$ ,�r\����D�<)(O��Ovo�f�n���*�L��"��v��6-Ą<���ɦ��?�g?!��M��'��I��_$��\@��L.�~E�nL%-��̓t/�䊐�Ś��
�����S�����J�3�e��l�o]��{� ݝ�?1���Ľ<E�tU���E�x����<����F. 9�������<��m
/U����K� VY���VG�<A-OZ7�X��	���0��e��q�֝a��%��.�
#J�D�v{�ȱ%.�5�n�	r"�1Ae�'j�i>�'��\2e(LX�1���$z�⒬_�`m��|r/vӺ�ۂ�9���&p!��Dܶ%�#�|y"��<���M��'��O���n+4��̐�j���fGT�ߠ���H�)^� X�'�
� ^wްQ�n!k�O�a��OP��t���5]׫��5��	ǟ\�'������̦���/�^7j�h��0Uu��<mF�f.���4��$�O�hbq�μx7��.&��(�r�7�MC��C��L�����<���D~��ҳ�̰_H��'���KWꜘ(�0v�U�3n�Cu�'���'�B�'�2�'_�'w�ӻ`:�8��8M�h)B��C> )ލnZ?��\�P���,�	�?q�����O��̭^�Lm ���-dC�QQ$+�ch�6m�A�޴ ϛF�'��$�O��$`ӛa6��'��X�Ά�n`�t�f�J+L�Z]k��'�l(��*�
G��|�t��`�Y<.��7A�+n�Z$G�7i  �Iny"�|r�v�<qK�$a*r(����Q���
a�'k&�'�dey��'A��5O,�v�s�9:�)r��ː3hb��I��(�ӀP�6����1?���`�Qͣ�y��:jz�MywN� ����V��?����?������<!����;?��2�'jQ�A�!8��4@,���?�����|�'�% Sg�\���8s��b�bC�f�Ӧ�m�|���p��v�`�	�6R��$�(����
$�SU ֨C�@8��b�'��R���|��S<C��lT�i
�a��\y��s�L�$�(�ӿR��M���S5"n>�H�ϯh�4)O��y�T��H��?-�	�ul�M{��=Μ1m��y�����jѯ$}��H����+��]M� ����ޞ��C�����ab文O����<1,O��Op�l�!*�I�[a�	@ D؞9W��JD���W�\����?�g?	���Mۙ'�D����Z	J�H!�#�A5��� 
דTZ�m��?���!�H����\I~r�O����"1�$uZs�B*J)�y�pH�%0��'�ay��)���!֐A����3�_��hT�A�|�"vӶ�8���t�ڴ��'���u��b�Nذ��n�:9��'���æ�ߴ�?)�
)�N Γ�?��I {^@x5GߧS:vT�	�+f���3r E�Pw�}2M>9���?�'�?1���?	'��9��ݢ7盻x��TYϐ��?�����^��0�h���I��`�O1�A�!�V]��=�W+�(]t�� ��?A,O4m��M[�'���Q>��%{(uP ���T�+6���$]Z�S�MW-�8�ɠ�Bb}�������Ll�c�t
��.�Ta�N/�I��<9���$6���<��4#ۺ��0Q�@u��Q��<�@�����k~#f���$>�4��D�On���*[6%)1�٘T��V�fӮ��B�16�4S8O��D
==|z��2(;�I^88�D�_�_�lL:���)��'�H��Qy��S
X}�y��^=�@8�'+>d�|�mZ�4�zc��~��5�M�w�����B� �X�[���lgܰ���'-�V5O~��?Q��ן�B�ĭ2n$�?V:^�``j�D�y&/��`�4�IvȄ� 鎙e���E{�O�D�u�ҽʐ�eY�BDI.ע�����d*��\�esh?扶/�H��@=�Hl��cT�P��IA�Ɋ���O.6�q���'Ph)�/�!CM���ᗦv�@��?��.��݋�c~��Oa`�U�G��#(�R�F��{�~h�(��
I�IAy��'H�>�ɠ&�RBJ�Vլ=���
:���R����:?�v�i��O���4Cz-��H���X�0�N#���Ҧ��ݴ�?Iס��l���?%���r�`ݹ@�`�#U�ā�ԧ�R�$hA�<�����O8���O����O���E��0�JҮ8DN�$s)��V��vi�&X"��?��O�����?!c	DU�Hd"��QM�R}�sh���	��M��ia�$2����b�i r�豱��/_3R�����Ttъ�,˓HDb�c�@jxlT�O>�+O���&�Hb���G3+6x����<���?1��?Y(O�n��/[*�C�? X����ş9^����E�fǴ���'�T7M+��#��dWͦ�XsC�˦9`#�<g1��aG�v�����j�<8lDaCy���I��8Dz�I�=eI茔'�����$}�]]I�	�6%�Y�6��!�'qR�'��'��S��Ol���s �#TҊ�#�O[�2P�1��!F9<���'��c��|>OF�$���m%��ڂれ��4��j03�ƈ���P�?Y�O�@m���M���a�J�H]�
���؂)ǿ:w��H�Ë�D����(Q&z2İ����6��$���'0r�'�r�'s<d��D;��ä�(	��%�O��.�bT��R�4e���'��8�/�+Ӵ�U��_��a�ş<���'�F�țF�kӄe�IH��?!jMc@�=Ӕg�( ydlYE̍�6�2�d�NKz%�'�����Gg0��%�䓡{j��Q*�=P��IQ�$B,D��	� �'��������i	�._���yaD���D�����f˂ {��b���4���O8����ԏ"�fa���I%��	`�c���L�܆���2O��D�wB����[���I2	�p���LY�܊��T��b4�	ꟴ����Iៈ�Iɟ��IQ��DҮ"�vTr��Y�xi�G_%,��g��y�'9B���[>��tЙ�� ��탔O�@M�4jś��c��In�����?!���ʔ�tf���I[�h���t��:z�t��6�W؟��Ϭ_q�wK�p�Ilyr�'5L�b�v��Aؔ^��rD��I�'��'��ɣ�M,��?����?ɕN�r�����W����O��?!/O���b}B�p�d���՟(�O����J)`٢"�����Y��?�J&Aɐ@��j����dz>�P��*r�T�yL��䝫's���K�(q����O@�$�Oj�S�O�Ā(Z��i����<�v�� ��r�wӖԁӗ�x�4��'��$�|H1�E	��{��0EeY�;��Mr�h8n�%�M��G
�5�PM�'���B�i�/�XijaK *p?쐧1��Ԩ��'N��'��������,����h�ɝ%$��d���r�ހ����/�d�'XR7Ky���O���-�i�O�(��g�2h�&�1@��}+ ̨S�YR}2ki�ΔmZ�?YJ|����ҁL�e�`J�k��v���k�;��(5F����$ү��	;�&� &�=I���$�@!�+�,u�N1ZW���?�(O�˓��j�������~B���yz8�C���kN�uz!���?��i��O��O��dv�,�I,��,�nL7n�
d"��
9:$��DM^��O�9!�cY-��<H������ٿ��EY�j�rs �	���27����py�[��~z�զ"t쐢D�	d�8�j�' m�	�M�D�@~�
b�2b�����6yV�*F�B�D��v�O���M+a�i�M�<>`S�'RI��\�
��Q�+q�	ua �N����2f� uU9��i>Y�'b�P�P[B�� ��bl��f�#Y]��|�d|��Z4��.�
�m��t:+�>bk0)E�Kxy2i�<!��M��'�O��4�F�{� \�eQ�ɔ�فLޱ�nt���Y���KUn~R�Ox�r��_&`�|�OF�A�K3Mf����˅X� �A"O��R��F9DԤ��4,���}*��\�R� �h��|��ՒÀ�6G���iŭ��Hm���D3F��)X��U�D�2h(�%�w�d��Ȟ�K�d��T���d5����O)r��W�X�x��"H9`Ճ!���F�D���#:�\0��P6>,����&Y$A� �XD֥*�d�4|p T��V/bX�7!�.���RDE_�P`{E��+�����?q3F�	+&�!bv���<����?1���۴[D��b�I$~20����8
��!���'���'�П0�Or_����Ǝ1)>Z��-N����!m��?9���?���/\�0P�9��aH���?aF���ꘘa�]3h��ٻ�̾
�B��H�C8	��?1��?ͧ�?������'S`H�B@�-B���>6:i��'���'�B�'w�I����g���q�.t�7(-2�q��N|վ���V|�\�4>O�I:�b�~���Ǉ�^�$�O&ט3I�2\����M�|Z�k̾6��8�� &������?a���4����O&7�Z7Y6��uL�z>��!O�j)��Izyr�'=��I�Oh7mN�#~�1��I��
Ϥ�P��
F)�p�(C8A��sFO��v���՟�Q�@$D<Z�f��`m���ܥ#�D��,�40��4h��?�*O��d�O����O`��?�ݴ?����ƩJAo�(p��F4L�����'�RR�H����@��5A�b@Z���� ��6�5g����+�=
��!Bp�M�5�q�	؟X�/<� ��S�q����ٟ��	�?un��8D$3׮B!@;� �2�G�ʹ��?	����O�˧�?1�O�Y�$�P/Q�b  �I�
<MڣN��u_��Gx�g�'�<Q�!�=9I��i�L��b1��'ؼՀ��z8ZY�C/l�X1�ۍY�Z9���98
����̖�8e/�w$`!9C!��>HH=` �އM�p�!SA��}��H �?KMX��a�Za(x����:Ɛ!X.Ҁu��G��I@8	��)g��@�_JX}1s�L�@�U���=w��Ag"X�,l�CC�c-�����ldL�G�iTr�'B�O��'M�6�.;'aֵmM�0SP�|2�'LR��#O��'0�U>]�Q��NaęS�`�-mC��A5�K�,�����Db���M�-���D��D��'�Є�&]$|�@ȃ!.@���b��?9��j�(#��?����Ozd��G� 4b Ջ�GC#2f�$���'�đ9�jp�~���O|���� &���I*C<�:Ĉ'h}"� ��N ����I�1����Ο���w�'�?	�C(|xɂdO�[��m�� �1$�a��ib�'��5PO.���O�)� ����c�L\� �)'�Ȱ���'���'(C�G��~��$ƶw���A�ZS���ǆJ3s�1���5.)�Љ`$�{cp�Z&f'�<3"�I�Y����O��$�O��/s`Y�	2Z%H�B�[�n��	/Z�d�O��$�O�d)���O�x��L����I0@��h�+ç�O���O���O��jB3O����O>�$e>�1GgI/=� �㎁2wЕ�g�O��{�6!����?a����9O�9L��=��$��#4�Q �E&G���Oh��OH�O��D�O���O�y�f�I���Q0)�|:ژx��Ox� �<A���?����?I��j٠��Z Z�J���3r����TJN)�$`���Mk�����'�2�'��'���,?���@�'�t��O9�d8#�@K��h�q)ID؞<	B	[�}��a���T�Qv�����8$���f�U���xW�_�TC(�+�H��W�pe��Y�}�օ)��8����P��e���X�H{XPk3J��C� qC��'t4|�PÓ�Gr��k�Iח!p�q����!��EO�\������3\d� ��Z@�u�R5X(�:r��
kC�4y���Zq\�Rcn��9�(X��$�O��$�O���ʺ���?��-Y<��fĞ	SX1�1k�X�6��I�Ar$�b�.Ү�6�iL�6�+gQ���� F�o�<�Y�'ŃӺ�Y$$C��pAԩIU��p�
�O�lڌ��<�an^Ϧ	��d��X,L}�陾TN��R�`���?�#�i�2Z����ٟ�����,fpd8(aH�,s�L����NI�"B�ɑ:(��ӡ�,w/\\����e���'�7�ЦE�'�2��F/z�6���O6-�	z�l�Gn_�sfTQr�11S����;%��e�	֟����\�T�.Zz��P����9A��(�7Q"�ه��(���za�?J5��Z��/�Q�d7�<{Y�hQ���.0���+7El����a��Y�A�W:�(Oz��1�'in7��ݦ���Ӻ���9�� c�&��)��z�Tv?	�����h�T�85J�+h�v����8s�ސ�s�'��	������#�S���xG咧v���-OjԳ�d]զ���Ɵh�OI@̛d�'=�V�S�ژ�SR��
m��D#���%����۬� 6�X�;A4��q�$�?�Or�OȾQ;�l�1z���o]�.�d�O�4�m��Nˊ� #EU�T�N�~��Bż�񫃍�\��]šFA}�_�?�'�|��)�$<����"��BK�9�
��!��X�O#��b� W
��8@I?�Q�����^�Z�2]2�@�G,XNĘw�����韘���$�J_ߟh��ǟ��Iw��nđ�u� �+QtX���T�DMֈ���ќ<`S�W6]�ҹ{ז~r��B�V���'�H��Q��V��á�MA,-*�*Z7�@a�C�������*��'^]��xn�"BlL��wsLY:�&��|���HĦe��,J�ڬ���YU���D�O\6MT�	��lk'�H�3�>L��%��Q]��3�O"�ҦL?4�	!BJ�R;�ᨅ[�\n�MH>Q���:,O
x����~���Q�,��P�&4J��$���T.�O����OP����k���?y�O޶({4�[?\{<١�lDe�.59��yc� �&a�ɞ� ��x� D9���k�'F�p�ug�
G@���'�u��ɑ5w�(X0�$D B��U��S�����o#.�b��˃�zӔYs�Q|h�m�eNI��$�2sI�ǟ�'�����?���L����1����j"��=g��C�	�u~�4p �1}��!S�B 3�v�'-�6m�O^ʓY�p�ۀ�i��'ɛ�l�"Ͳ�N�t����OB�˦���5y�|�D�O��d�)����f��N�.T�U�`�֝�*��rM�B���R&X5;*"?t�?R����)R�"�t�O�r	Bv�H�8xp��b�_�8�b��P�K�bet�z�m�ǟ��;|K��ڥ@W��ԃ�B���Ȝ���?����)K# �d�c�l��m�)�g�˘)��~���;� 	�a��
q��Fg`�j�����һ{V�
�O|��|2s�\��?Q�4 ��sd۟�Ud�HUfVU*���\A�@�
I��l16!Y%Q��X۴�"H��)�
��'Z*�����"�`$�3�f���'}�PT�8sR�z�C�5f�xq��B�JY�y��'z�#�.|J���/7]^���$"�l}Bb�?����?���H�����o���b��N�2P�(}��'�a{r��y�m�������gbŌ��O�,Dz»��T1�g̈́tP`��L�\��E(�՟�	��RE΅O��d�	�\����E8���q+۽�іgI�(��H�Fn�,��s(E�~v��K�$V��O�0����Wy�oJ�*�챹3�XM������L���T�d�����9^�z��K|Z�O� G�˓	��Qsd��#&�2�3�nB�6�,|� D|���dѦz��dτ��gy��'��f���$Q�)R���-���'ǂ�y2�q\dۄ��:��S�k�� ~��Y�'����'z�ɩe��9��iв}{0@��4�(Avc�)��͟4�I՟@�]w���'-��^�d����-�bDjWc >ъ���F���0��@�K�fg�Cp
��I���򄇂�0xb��S�s1`[_�̱ՄT
���1�Ǘ*�Mٱ�Q��r43��2!LF7��1�T�AcŞ��d�@Ҕ]�U�'����T��iC�Ppa �'NV�z�'�v"��Ao���`Mv��O�R޴��]�0aٴ�iDB�'p�� ���V���B���/�}��	���j7L�����ϟ��F�v��4s�)�17u����I�,.OP1fJ��\@���6$3�@r-.Tɨ�<Y���~`�A���/4\B�J_7ָ�#��dc�dZU���~NY1#
91�hQ0���S���'t�O��u�ɊqB
�U���'�^�0���O�i��O�>���D�C6���A�!�npa�E;�O&���r�%��1r�6`��Hu:�`+�S�T�����M���?1/����r��O6�P�z�Ve���W�p����H�{�
E�	�y��p%	Ú;�d ����/�MK(�v��EP�N%;.���-N!Z����\�$�"�YJ��T��CŃ-e�c?͡��X)��Q��I8�| "d�>ه����I��M���H�"<y���#:�5I�*�%��9"�>���=)��^x69	�"\�=�q�M�R�ў�I޴��V��� [��Aڱ �#D�lS��AO�j%��ן���zqjl[t������əO����a܎�4���N�|)2�Y��'ڪIsۓl��@2�E�V��j�J��&��{#9lO����Q�d������6��x2'�;�?�˓X�0�9�"G�5��¤g�$7Ph����Х
�'(@r}��"�X���*'��"|��hC8m�\��M�v4��
5��A^\Y�a���?��?��pl��OT�D|>e�������+�,Q��<9'$�:MQ����^� u�#��i�2�@*^�J�uN
!�z�ySa�����l��aQ˂p q��$ʓ,�Ho��Q?,$`4lA�%��a�q�%k�1�
OFHygk:T�$`%n�U\��"O&���aͅP����Rmѝ#"�=�B�>B�DD�hi��nߟ0�	ަ��D
] __�����(u�r��Pm��?�b���?��?�4�P;�?��yZw��#4�ӃN�J�s���B�ܰ ���׺_��>�WaC���`V�_�<EΜr�;�	*��IڸO�^�K�	!N)֐��{�l��'�h�Ů�X�����g��)�����U�������{2/ʘ���DX�L��4;�5o��aɧ�O=���䇐C���U'�4Qz�U��4��'{��s��E�7���/�N�H�>�P��>qa�׵r hP�9O�8��EJ��h�Z�Y��L%v�`�I��@�ȓ}͸�е��.'��[����%6�Ԇ�x� �3���"e{wa*6�4Q�ȓ5�L5�2�ѕR�@�qf�@�%�F���Dފ��0g�/lsT(q2���{N��ȓ�N�2a�ͽk� ۡ�'2¬�ȓ}c�p1�W�Qs�]HŃ��*�D���]<8�r���F�Qj�d�+4���Z��\+�a;0v�!��Y���E����FܽJ�$�a�m�<4���ȓt;�'�5mjL����4M��ȓk��j�)�/[րYr��[i�5��'��]��-
�/H��HoS�o�l܆ȓ=DpC�AۺH%
����{'\�ȓ^����X
=�� j�i�����*���Y �T
�Pm��]��["��⏍)},���ӛ_@&�ȓai�`q1���#P�Q�t�0}��u�>����E�l�a��G��L��q�ȓDZuq���'�|t��K�&J�ц�,Qh�����r��r!|�	�ȓ	���Ʌ�!]�ԃ��^2������3/�,��k%ȉ�}��9��&]򃅝=	 x��\�P�U��(������	X0�u��ML�g��͇�f^�|���X?��-T��ȇ�1I4UXh�wTୃ���vZ��ȓ1� -sl^= Cؑ�E�L)�}�ȓ2�Ac`���!)�њ����8F�������v�@s�`u�>K�0��ȓt��i�׉ӻ/~z�J��4!k4���Q&��yw�ȯ<bJ��f%݊K�A�ȓme.�у"�
+8��������S�? Ω�bG��sƵ��ψ*,(Sc"OV���Cr���D�Jr��S"O���M�l�t,`!)Z,P�z"O"����� Y~20+��ϵc�(���"O� �AG6DUˆ6�A��"O �U[9�EPG$�,��Mӆ"O�|�`�	z��a��7#B�q�a"O�3�E6��Y��-5�U��"O���5�H�*�@���(��q	�"O���p��- � �ID.Ar: ��	r�jQD���&,�.Icd�4Y����'٨���J^�mg��q��؀�'�Pp�hEL�S�O:�LHC�_(�]��@':{�l�	�'���N����I�?6�}�I�!3D͓}haz��0/���z�T�
_�����#�p?�h�d˴<z��\xT�`m�X^��� D� ���U5"��1H�3��Г�<�(ȊU%�2�'L��}@V�F�,X-3E0���ȓz��$�ΐ~ZHxRa��?\R��r��ȃ"�)�'8\�T�P�w��Z4.�1c&�%�ȓ/,\3�NC�h|%���B8�(%� R6�E����1aB�gu���䗯5�D���,(D�4Y�L:@ׄ���o�S���(#D� +u㔆#�)���:9�����>D��x�fR�������"z�l �E�:D�Ȃ��ؚR^M�#�A� �@��k*D�@ˤJ0c�v���
^	)��8���&D�x�B�@2Ė�: �C�UN��q^B䉌�P��GA(-��1��,6�nB�u;�D*4܂%,��,g�TB�ɻ !�)��7�p�;�ɀLϘB��#���gL޿hɸ��1&�1�C��F���ŋ2-�t5J��%"�B�I+�m{т		$�F�N��n�|B�ɖg#XL��b�Xa�(z#O��fC�ɼT���ֆ\�8�,�R#d��>B�I2$��X��X�	#��PDB�I,�Yʂ˽ T���tֹ��B�	�p�6�J O�~!�̂�k_�oL!���k�V)Xr���[�EzR�@%+!� �VҐ�@Č	)5�<d�7��)O!!��!N��2�$Ҧ]fR �t���7*!��1r�%��NhR�.��D/!��e{���3tSJ��G�3'�!��ϳz5�j#�S�y%\l�`��=IN!��X�?d~4`�X�R�ܜ���N�|�!�Y�:���� E�o���a�-f!�DU�6����fɱ/�Fd1��
+v�!�dX8�q���=[����b�!��(�@鲥"�h)���3z�!�dH�f�8��q%R�����ʫK�!�d՞;|d�Fj���H�87�R��!�$A59#ܠ3�ǎ� l�5Z�K^!�d�!qD�m�,A���!0'�[C!�DJ'�T�ّ�/��UjѦ�v�!�@
NwFl�㏅ vSb\�t!��&�T�G瞾`Y2�tD�&j�!�����pP�pBD�R��R�!�$N�:���6`զKC�1���3S�!�d�0�����T�מp���ۊ!�DArKpa���,1�`�'�$�!�d�t9�j��R+/���3w�
��!�d�3�@p+6�5�8�&�WZ�!򄎹t��˱FC�V�"(�L�!�� �lz��P��ȧ�7TQF�jA"O���O�G<�a�E�k`����"O��ra 4䀸J� ��;] �H�"O�������z��p*Rχ�e�N���"Oh�/"�jdq᠈��"��'�M)T���ܱV�܂y�P�$Dܲj����e�9D�P�e
�FO1`*�1VcBوA�#0�}�T��=���|Z�J0P�~�!�&���\1��,T�<� �!]|��,H�3�8�)�j� 
4� �G�@Ɇ�3�'�"}�'��ԫ%�,rT���D��f�X
�'��9�ʌN8���*����X�șR�����#Y+C�����(,O��P��ǯ,��)2�)�$#D���'���'v�p冫d�^yY��N3O��W�M��yd��W(<�% ٫�p�P� �N�ƹ��A�w�O���ഁM6Z��
�����|�l#� 9z`I�&�-(� �e�<��NV�MX�
��D�c��'"�N`��eff��;�:7yvm�J�O����o�а�qN�i����O��C�$̥#|�8�Lܩ-#P��J�D�G�F'�ֹ*��� !�PY��	�S<�LsD���	����!Ԡn�~���1+|�eªD��*�jG=inb�e��g��|[a�P"N����fF�gY��׽ZRv�2�;��	���I��v"h�;�#C�^�����+KvI�@KWB�;c;8�'f���Uo�B-f�
`�Ř����o�"� ��P2 ༼�Q��P$��I�	T�[���)R���0�O\!� @�kG�E2����T �)��|a� �s(<��BY�)�H@k6+�}1���IX=���6c����  c���X�Uq�"�q�'�
���(ԙ`��� S'����Pe�izs��YTH�30�͢G-�t��4,D��ઊ�_�Zt�e�D���y��T:��>��΅"c�ZU$���'�th��l�d��V0B �@n	<_8ā8�,�/���)������' �H�vJ��O�d(��en�ȓ4�a[biڨr�c��?+x�0��5#����� �6Z$���aƌ7���|�'��y(��y��/�?a�ؕi6hH�Px∍�!e��3�.`~�POc� `�F�%��b@V��ƼQVj@�#`��{�L �?b���Fj�����nF� �ȇ�I�M:|��
Q��l0��ONv��d�Q�[�r�ʐ�H#J����o�����kס �p>��j�#~Ԑ�C�Κ-n�̐���v≝4X�ĩQe\�i�LY �0e��9�̜V�u�'SI�pJ���P�>�Jp(��
G$t��k�j��"�B�Ԡ�vI���-���G!� Id	̨m��=��NѲj�1���a���s02*c��SN��
-9�Ojh<IV"*/V~��p���VPA@fŬF.����
-���`�6n@�:tB�-Sr"=�# T�f�Ԍ��'^��f]������	G
�[���*�3�ę�4u��Fz-�,b'ͽW@�yG�а>S�@� Eά3&e�_��m�H�_���P�5��A���`U�]ʥ@���Ϡ ��q��%ć`��U���'M!򄘄,4R��S�( ���P�E����%�*��O��>��u�SP�$ۮG�1ke׹C��������M!�DG|!��E��@�d��*�r��
�Y@�y`��C�"���ϨO��3�/�e��-GvE{⃍U��|�I4v^a��O�~����+�&ka�����>4�� �m8N�a�dP�)�V`���A����&煒�hO�(	�J��� "��	�T�MA�� VpXɨ����T�!�àa��ի�A�{.�Q&l��+�����⟢}*��	O�x���֛B ���_�<���-v�4⁨����SN�T�<)'I+m�![�%�<B�h�Q�V�<a!��¨� 7JـNMj)�U�P�<I�i�&��o�lh���
R�I^���Oo�t�ѼЫ��.(0SB�*�yr��.bXh�'Dŏ@p���;��'��z��u�\ؚ���wZ01q�E��xG9(���a�,T�	+�G���C�I4=WX!�n� g;j��6탷;zC��,=�
\���I4tE�+U [+�B䉞l��x�C	Y��%�ӷ#�B����1��J�g�|�+μ_o�B�)� |�Ӧ�X�%.ũ�FZ4U{���$"O���ڌ�� 3��Ҥa}"�b@"O�PP�0vI<ݒ�)�8D�ܴ+�"Ote���� �ĹQ"����໕"Ol�A�'� |���Ȓ�d�rmp'"Oʽ��/�=R��GX69�be��"Oy��=�lp�E�&R�Z�Jq"Oh����1f��I��ۚ��0��"O�)�tnG�7�t�"��0u��#d"O�@�s���;R`�I�!2~���"O�j�-}Ơy�ơ ���!�"O��{Ӈ��f�xbK��[�`���"O�� ��߁��%i4
�vB�B�"O�Ó���$�T%�é�|>��"O�`�G�
'�:�HuGE�W^�p*O�ɠD�Cy���U&����'#�1a��<M
Zɨ�*���|j�'>RA�w�_�;l<X��gH+;�V�C�'oڠ�ġ�8w���!�Nl^��I�'Y��9�B��k��؀7��l�Tp�'�&8���-;�~�hp�^���>D��Z���:&��A��ß/'Ƚ�2:D�,J��S�[�<K0�t	���3M:D��2-T�Od1P�!C�����;D�� �aW�1�QrE��R�� $7D�Ě���4o������o�Jt�e�;D�l+pfҧtʈzԎg�����I*D�,��$L3��ӠcG8�̸`2�)D���KIZV8e, �;t˥7o!�d��*����5r�� #Vk�^:!��R�%��Й1�4�f�� ���Py2dGI���fK�LtM�Wٙ�y��!P�t,��*O�M�N1��Y��yR����p�:W��]+B+���y�C�-tQ�ۦB�8F��h������I�v��թBc�Q�`�u��d�J����#�8�x@[�A&�t9aנ<D��H-[P�
��/172�(�  D����H&k4�(P}%�YW��y�j�}����elϦhH�90fk��y�ON'o����h9KS
�yr�e�A�i��XNX��%�T8�y�dʝ}��!aEA�ED��4`��yb/15��U�񌖚@��T��Kч�yr�=?hz)�s�ؿ3����2��)�y�NխG���f�M�+�֑j����yrB¹9?�J� -Z��|�A��yj�`w\s���Q�H�1#���y�ݕ BDH�΋F��Xa�C�(�y��Y9sE��c��..�(p���yM�'�Թ�u���&�Ĝ��R��y"�A�.X1РNY"x�C�yR�uQ��f��v����B��y�d�Q1����˴���zF�S��yb �`U8i���824�Cg���y���lx���
,/d�z���y���U���vH�8pu���Ĉ��y�O�*a��A�R!Q�z����֫�yBIؾ8t���W�o=��S��y�.I��ݱ�!U3e�����@�8�y2a"�����Q�LJ��6���yb�׮�(�B02<҂b�!Q
ZM��f�R��s��� J����挆ȓz�rс��	7���1a��P�ȓ�≘�J�+^�5Bg������S�? l�I��E
NxF�&YZ�ks*Od� ��}�ܸQ%A��-��С�'�f��u�Q��c��I�R��]�'ui����)7l�����@��'r8� ���}��i���R����l�j$��F -}.LH����y����)I�Tar4��"X�JV!�]N�1J����<͎��-F���>��%V�W�"�ّ�̦�l�A�EP��<�����'��QFD�T�6|c��l�=�J>��ꄑ*ִ�D)!�%!���I�'Y^�2V͊ `��!!́d��Q1�'l��q�g�)��!��^�
tP��X<w����|\bG���<��c�/.2�!@�Z�~C�8��J�<��*C<B��t�3�lp���k��'�p���,�?�)p���,��]�PO�uG��	����i >1ٳ�L�1���3����YF����}��nG<� 9!�Ù784X9DJ�$k�a~"j���z����Ƃ[HT���
L��a(`㊃��'K0�u�Q!G��@��ܐ?Pa J>)�� ��wݷe$�-	�����K�NtX�����ҟ�/~qO$I�ϟ�Q����ݢX�3�|������zN���%�z�@-�s�9<O��03mٞ����b�_���x�qOK�-�)B�P�l�)6�M8o��֝���O
��T��*>�B��2(�*n�Q�� <OB��
Ј4	�̋�-�h���� � �J�;�(ؐ�V�<	�x��5u��Ƞ�bA�*��8Ќ��%E`b��F{�OF��uE��c>�рF��^�8`yvΑe
�4H�{�@�E�%�ZG����	ۓ��v��	0ǕfH�+q���QDxb�d��x	p/�<��#E�ԕs��N�<��)�3H����T����q1��k�9���O+�������<��bC"�HL��
"�"e��$�>�?!v�Ԥ@(�a#V"B�,�2���jSl�'攍��G�_q^�r�旐� 1P`�'��DX())2�dL>�ك7� P�u�c��Qsv8�&�8�D}O7}��1o����cW:-:��;��Y2PJxiXF([g��~���<�s\>-!ش~fp�A7��c>U��ˌ*g����JAܓs���b��Y%P9��ʬ@�fU'�$���^wҕ�wʔ%�X� @b�~ҧ���?I���^��)��ɦ�fA �y����Ebѐ��3m.cE`���
��U,-Y�*�:����y��ܣ\�@��`T�lԲ]s�C3O��D�;�F�B%�G�>5��̃��OVq��n		v��"��N���c%<O�Ia��HpMX"W���O��j��E#���ӌ� 2�Q���� �&�\5p����yh��Z�P��܀0JR�'�LY��D����O�˧x�V�"�Y2~4z���" �d�뢢�����=Q�J׬5������W� �� KNw�I�No�	"o�� ʹ`s�!7[�7�=}B�'�7�X�wҎ���E�&��;в͓"S�b�wH�a���_��+6-�<���s�X�x�����t��8X#�X��QqN�����c�ZV=H'�"6n����P�Z��y���[�S ��0��9J��䫟�x��|?Y����o�P$ir@\K�T�{��Ĺ��h��Ur�'�Ĵ��FU�w�N�Y��Vx�]	��U�g�~�
�D/
C���<	��T>QO|U��ʷ/B�kf%��Ph`�B�`+�	t�| y�F�=�*Z7#��n��O�Y�Gȃ�|�v��*����XT�$�O��=<���eG�,2	���Q�U��\���i�
��Y*&�BG�۪;�xP�a�\�v/�y��j�4�����8����sm�
<���P�c�1^����W����@,e�v���?x+�Rc��:R�,|S�� z�=��#Ax�|�?�c\9&�ã
g�������Ϧ�)&ϔ"��OxU@�4_�R���Ow�ѹc��/ov�e��GZ7�
� #�	3�1O�d�����{n �ֆO�Q��q2�EYA�8�Va1� <�X�� �v�J�p@���lJ��'m�
� �T"j�F�
�k:�dk��Ӂ`���B!���-D�1�I�v�>�\�ş?9�cG2g�@1�3m�&�R&�|�� q"�{SV�e��@�D>ʓh�t3��:x�un�<-��-̓q�
0Ie���g�ц�΢(^uE|�E�G�D�$�4q<�E�	���hO���@9A�І+@L� �Ѓ*z�
��S�l��	, < <�֨׍P��n�J(�-�E�پ[*"LA(�5~�qO��F}��
���T@Uo�Stis7A;T�@1��.��'������:��ᚦC��I�ؠ�*O��kȼm<�M{$��?~�F��`͹?������)d����(T�̠;�oe�� !��;a�M�q�
�C�͍.P�n�(���16NХ�����4��S�$P�X��SG,ǞaJ��c�(���?��@5Dr���	2�&@g�'�j�Cǎ�51�;�S�z���SN>9�C�֠�Q��&�'&&���HƏ����*QQˌ�ȓG��<p[?��<�K*>�"�x�ޓAw��VD ��L�,�sՖ[F��`�A?C�ր�	-4��� F$���5`�-�W��<22*,�dT�j�phR��BX�ܐ树7��PPg��Pbtm�o$<O�RTo���tl�O6��̃P��q�ɑ���"O� `ȦGz����O[�Фȣ�|��_/Хʧ	_I�O�(�g�\zmBS�/5kV��'����Fh��.N���͒��:�'��,&�'��t�C��>�E�W'$"��Ȣl����@-Cbh<��+�>b����^�QQ��]�;<2�!2"O�	1���ԍo�T�P%țE�4��^�t�ϓj��- ����"']�|�^�	@>��c�
,m��P#�&D���c�<p ıZc'H8%�4*�#�$Xe��5(���ȟT]����X��8�"��Re\d�v�'GR�V���\Ψ�Ë�:y|�k��/չQC	�g����V�D9}J~b�d 4���:�-
���tk� %Y.$�+Awܓl��鉑��9}HhPr�G�C)'���#T�epN����"�x��'��`��މ^X|}C`�F#o�"�ΓU�8�$Ջu���&�	m�|X!��>�R�Zi�:)����
�c���
�0�5KV��l��?��a	�I�$��!��9#1�F|B�O�S>��'nؔJݚ|ҀKݷ+$�C�=�@3č��.����HЩ]�8ف�D\(�>��E�X�ء�c�yʖ%H�|xꄅ�[t,�p+,�O�A��C�l�P��l�'M{�	y�N��3��8��D^�Y�p��"��&k<h�'Fػ4��'|��b�/S�������!��-����ߟ��@�a�F�]�r�8&��%���P9R����?
��j�]�!�F�9Y���d�P�a(�����*���fAs@���%A�pW�;��2,̞�4�s��4L
�RPl=5��Q���{k.�8���@�'J
����iT�$�O)*�&��.8[$̀�*B+ꘊ{ �Y�"��#EHE}�����tD�Ph,�8C�+�.cR���OK��x����J���	�90�`\4c �"](*��@�S��魨+�b�q����5<��z�U���s"}=�'`f�"��[s�:�	�����n�I�ORt9[?-_>���ܬ��u�g�'�����O��䞾#��z��Ӯ:�RH8��Z�f���9��W�:�_$��u�I�F�n�8�!*�Q�iL���jY ��`mZ�?��|C$�BZ,�h�;l�"#>vǁb��*'A\��ݠ4%�2��On8qBhȄt��b?��П5:��U�81\�h��^; �[��3�������Fq>�ݒ(>�	C���|���I�x�"��Zר���~��	N ��E�u��e͌9�7B�	�@+�Ht�qO�Z ��1�)ib��Ox�J��|b�$U�i�"DhJboL��yR=O4�ᢅ���FTJb �dղh�&L>n��	IdcT��y2 <d$��v耼NJ҈��E"�б�GN�.�$���qO�tP�'�X���!>��R�"S8L�N����*�v��;u�26�͉>�`�FM�]��u`���0r���F�Cb�J�(��� 7����OHU!b/-�&�֝|��ja�ى%<�<���=�bS�O��V֜�>YƋ�#Z�Z��7"f����L�v|��8y�>�����`+���}�D�B��>%?����0Q���s�&˴I�H�X��ӀQ���f�&�ɈHv�l1EK�3v٦L�C�՚&�OXd� ̈́2�2Qx楃QyD��Ք>���C/�r�9���l�d��TNFj<u�&&��3x�I�C�2�"�H+BrYJ�nԚ��; 'Þ`��  tmF�G|2$��PGdd9��7�.!��S'*0� `Ҷ��q��k0t�k��&l9� �{�'$���c�R�i��`�(�{���E�4�Y�6�L:��		}?�#��Z*=Ht�W�ل����"��ЇL7�8u�E_�0�]���L�A�
t9��*}h�ɐ,�Ԡ��F���ɴA��'y��ъ�I����k#�J'l6 P�&C-p��=Q���V�b42FO;A՚9c�	�B�+�P[�oQE�J8���Ii���*㤞��0�c��EV�Y��r�����ɵe$�L��%R�@���L��E��]YB�ٔ	�"D	�&ON��E}��ԅ䞩�`,	*$\�gi�	^�@�	y����H�%>���$�!$���d$"�7�ր�E�& p�酮ԇz���z���
P�h"}�!�I5v����%��ZZUQdOq�'=`82 A0��Tϻ[���:��H6>R䉣aM�d"���E�	�����������c<J5���KN������:�x���D���V��V���\p�,͵��'�p�;gǨq$Lʇ+i��[����<1�����:���0��B�}��nϛE����Q~\Y`�P �P�ؖ��`Ü��ѵE&���-�8��2%xI�ɣ6��t�	~ i"版`)8�	8	׸��#�2����Ã?�6">�D��w: @��J̡F��\��L#Y��O0$xSH7�)�t��H)�9���#M�`��e�='���JQz�'�j<Ѐ���\��;,]ܭ��ӛK"�'�W�ԀR�ܸ�����V[77k*�����914HT`�D�z�tL�F�$Y� ��L!ViW�Έ�E��x��'КE���X	FTx�7ǥvGh���J�s<)ŀ�~b�����w��� ���0$�Z�ڨ	�%R9:{�<��IâP�Ѣ��`�"����CX�l��E�&!�z��Ҋ�66b�t�)�O�h�m-�ha'nX~Bm����*6��@&�4q]���3��&>�C�I��\�B�	08B ZK��`�B�	�%����/d�hlP����e�B�I�#Z��j���=�
�3f
V6�B�I�Kd�
�k@�aa���@	�m��B䉩o���7�	H=��������B�	=f��ء����>�"��c==ɶB�ɽ@���H��Jq��0)�J�Rt�B�I�E��Y�&	,BǨXr����l]�B�3;�d.H�P��. ����"O�D9Jo��PE8%`ā@"O���P
�6��B���>G"�`�0"O>�SǬeޔ���͗8u}l�"O�%�À�:;�����՗t]	�"O6iS�t�,x�%��zb"O�A�G���f'.�y�%y�(��"O e�˙�M��:��ԀK�'�|�U'�h�v=�E����'G��#��ut�ݑ�&ג�N!��'	��
AM�i:�0��{^4��'�|pz�N*s	H����V�E���'���X�/�$�:UH%�U�؂Z�'�h�A��G��ya�����p��'I`��J�Y�����$�3հ!P�'��ŪQ8�p�"�&{�|x�
�')�x��(�?<�)�b�D  y�`
�'��d@T����*�#]C p�;�'�.�Ze+��R"$��B�;t6ps�'�d2fH�%.6�٠#��@\(��'$@��$��>��ъ��8��u��'�@��S��LPB02t�=��'8�I�f˨/� �x jD$#6h�`�'!�EH!��! QД�ޡ#�m�'����,"Ya���c�%-D��'p@%f��M��@�
�Q�'/���MҺ
F���s�H<d�rI�'ӊ ӱ	]�Y-^�b��8Յ�y�Ï�7
���MեN|�R  �=�y�"M�i� 9+B�����'A���y�자vD��f�*T?�����Ĺ�y�$	�>1�PX���;X���ȓ�+�y2�8oIj�1�)<���i�˲�y���7�8�)�[3ʹZ!JJ�y↎3lj�(y'�\A���� I�)�y�9䜤�Bf� -X����'�y��ȰTp$�k�!�z0���y \�yM�p
� �0�S�h�<�1�\w�� �!숎u�vL�ʈL�<�B� )�i$$��`'d���RC�<�ԉاn�V�zCA�L&dU2p�OC�<ys�q������Z�����u�<�#��F��:e�ԇ�N����F�<A�E�;zWLr�!ˋ*-�9��G�<�G ߃PX���KfV X�7�~�<Q8�RJ�$1�b��o�-��x
�'�%r�.�"mr��+ �\�&�Ԓ	�'4�����ޏ%���$L��*�Uy�'s�EJ (V�
���Ч��K3l3�'�Б� �995t����E���"	�'���ٳ$U-m��C��ތCɊ��	�'�Xp���jw�͊�f
<�	�'yX�zV��;���u��0\P"Q!��� �����zlL�������+S"O�9�Q���MIe��1��|��"O�,!A/Q��ir���<���Xa"O�y�$^��|�ӖT�.b�2�"O֍����1�xt�
6@a
`9s"O�u*�C\����s�䃌K- !3"O2�hWcE1�B�a��z�y�"O�X�R@ʜ;��<Za�S�	] Y(�"O�AB�O�cQ8P�VXDx�٧"O����h�� jBGY�Ma"O:1�&⌐57
(�@	̓W�"�3�"O����N�5|8���Q�8w�޵"�"Op���A`弉�(�+f��hB"O�Y1���{�:���G�.+���h�"O��;C/Y$R,�r��)4�NK�"O\�yD$H�pzQ��Fi a"O��ZEd�����׆bJ�X+�"O(U"!�B6d-@c23z4�"O�!a���ةk�A"n��"O�bǘ��L�P��E�d�˲"O����dMFm��+fAҹ+�4D�c"OY�q��#S|�H����C�8�Z5"OT�qB�U�E��0ar`�"O$,����3���4N�b.E�"Of��T���h�F��.I❉"O����
$`/��Q�*B~*ps�"OȤ�Ħ��Sf�����F�
l�Jr"O���ć�;=��1FF#tMT�r�"O�u��	))���+1%��f��M��"Or%RVꄑ.��-ڗ�@Z�"O�YB���-���O�J����"O�Z� �$�d�j2E��k�| �u"Ot*���:D|��G�ܫP�δ��"Ot�s�ZY��� #�ކP���@"O|	�N�.T��1�>a��""O��ְ5N� ��/'��@$"O��'�F� ]�H��/5X4"O�}�׮��CqR<x�x�z��"O�Y ����L;^@�B��f��lX�"O.й�lBL%�UQU�F<y�]�"Ov���T5,0�8���_@�NԹ"O����%X<Tp����A|]¦"Ot���F5����t��m*l-P"O�qY��˷>L �O�R����"O�	R@�Y)k��tА�д\	�yI�"O��i"��'ìPx��ϼd�`"OD��F�pK 혳B���g"O�`A��;�v  TlX�Yq���P"O��dC�)�晘�aEC[���""O�8��I��>d
� ���Y��!���N�r=X�捠_������ЀM�!��M8h�P�ӥC�+i�������#j!���B�y��b�0\��9���?M!��]�JxD|q���R�
Ti�^8�'0h��D!x|�a�W:f J�@
�'�)Q�H�yfp�3�]Y��	�'p�	hq�Y	#X��2�B�`)��'����Iޚ\ ڀ�@�m�z
�'=.x`c�[;&�-�qnA�k#>lP	�'��#��
�� �t��u��'cL�`�ǮU�lX�":q�'�>BRF��*�Lm���)+��J�'��Hȗ�[�(|��ۛ҆��'�V@O�5�Vݰ ��;!z��r��� ���� �	�$�1�aJ�R���P"O2�b�!U�L�J���84��� �"O(�x�,�]���&l��${��	0"O�=�N���TѢ�k��_s�j�"O�!�ӪR]�K�'/j�y�h[�y�"�*M�8ు�.�Ȑ��M��y� L�%�&͑!��n�ՊR���yB�ܡȬ��7���	��c@��y�%Ӄ}�����צv@X�Iƣ�y"� 9~j4\2Ƀ�}ɴLZd���y��XEDH҆BT7@R�D�c���y���w+l0aQ���K� i$Ŕ.�yR�#��[4�@�+�P0���y�b�=Zn�`�AHջ&�8�GN�<�y�@�~�b	����q��x�6��yң�)�^I�5���9YxQ).���yn�:P������+������ya�-�BDB�)K*K�Бg���y2�ў5z�\�
����	4�V��y����i���3���B@�Y�� ��y�Gͤa�H����(%�Ћ�̘��yR��1hp���N���$k��[%�y2� X�윪��bA6��杅�yr�R�(0pgM�_ƞ���$���y-=KZ��u�G*D���z�C��yB�A�r�+�HK&��	0@"��y�X�t��x
�aY,>r�`�*�y����kC༐s�Tbtݒ��@��y`_�&�x@����\gd����y�
�]1*X`T��?�r�J���yR�LbT�{���$@����l֌�y�l�.��oQ	�PTb����yB)�ET�=���#�0E*��N��y"�� p���a���$�}�7ā=�y2�(��)�B�å~�p|�UcE<�yb�Hn1����w�)B2�5�y⥒�nNx�aT�( �`��!�W0�y�M.������{��������yB�J>z��ʰ?y]���`��y�Q�0ӄ��E) #t8��*`Gè�yB$��*��S  HҔ��cQ>�yj_)��)�E���!3$A>�yhB�܄y��٢N�s4A���O�"~�W��"ri��g����d��C�<�èZ-Z�����JT8N�n����BAy��)ʧ	{8��n�:8�<+�&
�(x��cP��Pk�%���d�M
E�����~>����6��*â�f���ȓ:Tڥ����,R��,S[�0e��g� �"7�G�� pfMB���1MJdY� G01��=���X$����R��	����@2D�3���=G����ȓX@=x���Ln�PK�-��F�4����V��`%dT8���չw���ȓU�< ��$9�qGB3B�e�ȓ]���v�N�o�����+�_.�h�ȓA4���C��4m��,j��)Jj���C膥�4ƒ)iĮ�ѥ`�f�؆ȓQ�� �.��(����A���8T���V�L�J!�ݜ�N��%$U;T Nȅȓh��1� ��|�b��f(�P\D�ȓL���AE �#_���rb��/��(��M�.���,$���8�I�(����ȓf�kR�T�N@TN����M��S�? >|h�ka���%-�%hd�w"O X��BĔH���W������d"O��b/�%�v�� �t�N$i�"O@��V����]jiU�
m�C�"O�H�fo�U�x;�F��O�8�G"O�|ҀE�EiH��k�>K�Hx`�"O��.��I��ȃ��mx�"ON]�q���;>��Z�X)�"Or�S�Ή m&�y	�M�Ti��q"O��#O	9�g�XbO�u�&"Oΰc�I��,ha�k�ED����"O����T&#���D*�!G*�h�&"O��!J�7n�����4=J���"O� Y��Gy��( ̀�P��Mr�"O@u�v�6c쮥�a��E�$hj�"Oٲ������@���ac�!��"O8,� X�i��f�_Q�9r�"OB�2Ɍ�(	��B�X]���"OX�P`�S����R��wOv�a7"O
i��o�2#K.C7�!*�Kq"OH�ɗ˒%]P&�e
�g�P�ɑ"O����NE�űb(5�h���"OH���G�}���d��p�T�W"O!����`a3�f[�#֐}IT"OQ/Nbd�1�	*���P�"O���tBH�K<dq�'ɢ��P9�"Ov0SS�[`O�8�K�"O���Ud�;k��4b!��]�P��"O(���6�����ĩ'��E�"O�q)ӯ`.�D�L��z�p�1�"O��l(YGX��J�6R�4���"O��۵��p���%���Y�"Ot�(�$�	Q8Hb��l�M"�"OFiB��%"�4�0-�B$>�91"Ob����
Ns��.y�zL�Ň��yb�ھ1l�YlN�^���Yb���!�D���p���x ��j!L#�!�dE%E��	w�5_�Zڧ O�<�!�dG�Xtƍ���220S�ȑb-!�X�!��}�Yu�V�@l��H�*���|��G�M
k�XA�Rk����=W
lh�+OF�GB�je�����ԅu��^.ӭ��A�ل�B��X�`CE�u(��(`��=D.Մȓcd�)��,u��}��D�;$*0���tLǃ\���4��#RLkF]��7T����P(.?@]B'.��@�ȓ���K6�6|�&}��O�.؅�����
�N���[��T�nC��	����	�L�P\���roB�ɱK��AX&� $
���ƨV0A�
B� A���#N�h2�-�gDҐ�B䉢'P]@WKJ48�Y��Оs54B�I"#n�J5'ވ Q֩˕�,.�lC�	[n�`�U���Fԉh���6MۜB�I�!yؽR��L�"�f�5��-��B��+��h���Q9h���I'hW?p��C��1(��	P*�d^�S\!��Z3"O氺s�
86��,²�_,d�"�"OVE2�� tJ�8�@9C���+�"O�;Ѭ�Q�0Ĳ�� Q���V"O�IA��� �� ��E�"��Q	"O���-�/L�t�rbG��Ht��۠"O����g7_�J���c6�(��"O� pD{�d֝c�X0����73�U�T"O��F� -��K*h����"O0L�T�]�*A�a�&ʑ��"OHyɰc��_�N��#	�DѠpp�"O<��J �S�D�pÇ�>;�xh�"O҄b%��m��x�g�qƶ���"O�İ�.�>`@�`
F�.D]}Ѷ"O�����n� '�M�7f�T�1"O�L:4�>��-s��8���[�"O��z�Č�cBjP`:��M!�"OT�͋96��@��U�L��P"O:�J�K�B� �V�ݡ1k���"O��P�ǒM,i�ND*od܋�"O��s	��m{�� 5͇�u��|�"Obɒ��Q)|�ѻ�fY�<U@�[E"O�5�,A�U��Qs�eЫcM:�A"O�EX�nE��2�����K��!�D�)jx4��A�ŬK$ k"JAL!�d��V�C�,�=0:����V/!�D�6m} 񁑉Ɖ:T(17A��!��.Z���c�)ˣ.���)9P!��P$}F&��I��~�\i��O];!�$ɮ�(B��7x�hPrk]<.��xӐY�'�ߖMx�@�s���]�L��C"O2V���ns���)[2�=	"O>�	T3{�@ۇ*Չ(���"O�S28DaP� ��!L�y��"O��%�)'BI�&i�M�,��v"OHl	�O�}��@"�H]<}��'�!��Y,�m�@H�����h_!�䆧'���RRCǂSy\8:���do!�!.Q�=��E�;d�3��8KH!�dÚ5��i�Ej\R�5�pMj�!�R2�2e�*�����#�V�|$!�,�j�!�K�4F� x�`L@	!���1pe���5aZG斩ce!��F��,�5��z( �{��(eT!򄘀)񶡸��	�&��s l@!�)�(�4%H�c
6h؀�T��O��	]�O��a�d��5H�F����B� �'"�%1��6*qPIK�Y�W�4���OH��DT)0��E�!��P��C��Pyb�G�p���Ս"�tᑔjU�y�dA'A\ 	;`	�KZ� ��bK��y�mF<K�Ÿ�FȢDSM�����yR։M���;%h�ТkS��y��
<xM �Bɉ>���"'N��y2)@6+ Fͫ�G�<J.�k�Ɋ��yr���8��� /,QR�D�u�V#�y�/�;>��xq$ďPFY����'�y�mK�(��X�@��!�8��$E@�yBH_��X���>o>\Ѵ�ȶ�yB.K'E�EӢ�	p��	����*�y�k��/�r4:R��d{��g�����)�O�f@��7�:��Ы����"O���SD����H �^�D����"O<��ƙ[&��3��7^��c"O�p���(z��G\���"O�q
V ܙ"T 8��/1�P��"Oj�ѡ�6H�r�PВ3�� *U"OnM!A��:�OD/�2c"O|�SEE�{��]���ܳ7���ۑ"O�X��#_Y�f(2�
jp��'J!�K�Z-5�c��u��I9<!�� �l0 M ��KR�@&�0���"O&�aM7& �Veԗ)y|��"Of4!� O�#�q�%��0~� �� "ONL�w��};�����ˡ z�x+"O� s�<#��<��J�8Ch�"Or���� �!2�H6kw����"O0�ÁCI}������s��'"O�LᤧUc(���F����x"O$Ћv�ɎI�4�"�^CS�̙�"OԢr�W�|��'*A+;�Zm1"ON��+ŋt� �v��!YjR�(�"Op�#6E20ڲ��oɱWF,���IJ>�mк^A�m�pO��;�A��y®��nf�S��j�n	ó��1�y��|� ���F��Vb(� ��y�Ń�n|�i��GЕQ�t0�w�(�y�& 4QXk��<��L��Ę>�y�,����Q�ӎJ4�v�
���4�y�V�%�|M�V��10���#5��y��.\n0����&B90�M��y��C.oN����НR2 �"�b�,�yb���{UJ8��ϵ^��q�aҐx2�ަq<�(:oU+ ��0	�8��C� l{p���"�()��:�N�
��D{J~:�fU�=��p�n�N���16�R\�<� LI*�t]��N_/�i�B�U�<a"Ұ@*Ly�A�B۠u���Q�<�0 C6:2�È�'��c�!�E�<��(>6�΋+_ �6�v�<тAx���#��#�ɊL�<!���,�`�� "`e��GF�<�g���h�y:�gK��� ���W�<I�]qh!��a�n��bd�M��&�@�����D��!�'Z�&U2���n#D���cܱ�8\�oE�M?�=��� D��:3��4N�z��#�V�)����;D����kB��t��C��`����6�6D�<QQ� k�T� 'G
�d��R�b5D���qc$J)�CsCM�Hp,4�ĭ0D�b�n�HN�"�,�g���ʰ�+D�xZ2
�j�P���m[�:�����,5D�����ҠL�����׻t�=3��2D�(��L�O�f�Ѧ��h��a1D�$�6�56(ȹ�feV�>��v0D����ʦkO����剉v2�:�O1D�$P�@�h���qtc�9&���$1D�4Ham���y'��)s���p�#?I���'�
lR�#ɛ{X�H�0O;�4B�I�G�h�T�X14��0"B�G:C�ɌcL0q�(��Ҙ2D���G��B䉚(���(G!O�q�n��7���6����}�5O��ɘ^] ��Խ$�z��!
I}ȈB��-X�F��Q�_���󬉁o��C�	�8Dqt�L����(���W�`C�J=Td���:��X�W�W�8C�	�8}�-��#*?�ܐ��O�5�C䉶�@�8U ~�p��3�-[D"ORаŌ�9F�����k�ov��2"O�Dj£Td�.]������U�d"OD�&k�{�H�eòF�NP�T"O�u����_�X�B��]y���R"O,�P݉ZE�̉�%[��bQ"O
��ӏ�>&J��qwg�Ϯ�*OP	c1�]�٫BO��m����
��� ��pQe� z�=�D"�Ovp��"O�ݒ��I�P|���M��<)��"O|ؘ!
_�>�b�J�!�9n(�hb"O
�� �K�7��ɺ��\�4��<x "O�@q��ٕ-��h�@+����C"O��J4�\!W�t����|��p"OB{��D�WI�̛րP���"O���g�4x�|����4&����"O�]9�d��#`����Zm�Jћ�"O*܁���u�xTP��/@�P�"O�a�CK0`�(8�Hٝ.ţ�"O�[筙&dB���
	�i2"O��"╲i���eȲ\�2���"O������|H��d�!4�R�c"O"����
g�e�EV�	�̣u"O(�Z0�
�f��5��B�`�v���"O�${ՋѺ2��5���̴CӸ���"OЀ� ):9rt`
�B���s�"Oܐ`��J%U� � J�u��B""O��3��X�h��(Xb�ʛV�]�"O:�h�`	(%�A��`��@��<"O�4�T鑟A~j�toT�z��R�"O*�c��~Д����j4�˱"O�� �,H=\c�8�`Ӥ	c �pW"OL�sq%5��p*���� K�"O�Ljd�H�4 ��b���2�$���"O��쎪"��yQ�L(d��哕"O�QPeΠ`����;�����"O�|�uk�=_��"fEˢY��Ȋ�"O�0���i�<�2���6Eu��e"O9�G'ٿZ�5#G$ؚ+�ʩ�2"O��"$A�;{^$SӠ�i����"O,��F��J�\�q��sy��2d"Ov])��[s� �i��4&`,��"O�t0�!K�I�J�C5��RG:Z�"O4�cF�'ScrE��c�I�e�"O�X���CQ�.	���:FBp���"O0��e ]o�����4����"O�0V�R�Ah�X�V �[,��+�"O��Q�3PL���T#jtT�b"OՋ��S��r\IaK'x�:� s"O���c��C��"�aA�I�Ti�"O^�A@��;�V�"�O@Y�.�{5"O<X��nW�0�<�T.�u���F"O���D����1ۅ^3�:��"OP8p�عx�TH��t�M�"OPqI���,o�x��4��<Z��c"O�lXu�}�
���
eF�Z�"OZ�UrI�]���Q�&_@�Г"O*|Ȅ{�t�K%�mS�,�d"O~H���ȫ%Ja�L��&<��a "O䨚�(�"]7�Y���V0G5�]��"O��[��b 䪰�Ǳ<�Е9�"Op�� Y��KA����S"O��S�m�8�f��6�'�bJ�"O�X�@á��!��M�_Q��R#"O��*2�]�	:p;��~3��qR"O@�P�E�9g�Tm������{�"ONE��D��~{�_�>w�*R"OZ��v�Վ  �YR!�dgl�H�"O^��â�6z��1����4�b��"Of͛B/��l���(A�E�I���"O�0���K3n:�9R��A��v"O���^�4��Z���k7��r"O� F A���K���⚃NȤM)0"O�(�����y��� �^��r"O��c��^�k�H40����Ӓ�#�"O��X�%AC�8CU��#Y�(
2"OX���n�1"��-����29�i:"O�I��$}<)�*G n��"O����E_lҜ�:�)�6���"O��I�,O�g���Ȏy�麧"O�a@�͚4�^�a*]"nAW"O��;Q&Tk`��krC�'L���"OT%�ӈ$���)�&�kT��k"O�����I��6Gb\�b�"O4�s"T	���ב5K\8��"O&�z%�',���[�a׫Фl �"O�����Ԕ�� @���E"O|���BԐB��a+!�O9����"OR�ѡh��Ţ�! ߾K���RR"O*����� A:�E���Ռ�y"	Sj�=��mϰ]>Z jd�H3�y��ĭ�Ƚ��.Y�W:�0$*X*�y�ͧnp���M^e�@)�%��y����TW�݆J�&^#�C�I�0�x]3�ɇ4Pt���W?d��C�5CDT�+F3JJ���k�C�ɵ�ҬANN�j�1�͇��B�I:9�|�Z��/N���ѧD��B��P�V!����B ����
PC�	g��y�[$,�h�j�N̊F�FC䉗h�B�*��uDf,)��DZ� C��'.�-���@�~��°G�JC�	���8��-�� A��3��!*C�ɝX����&Ղ�DȒuݐa���d���#bC�81��w`��WV!�DF3$%b%BT"HG"�PU���]�!�Η��#�OS�B�}��.�U�!���H�pH���Zp�#w@�M�!��xtT���Q'G)$��㌝"v�!�D�*��	�"J�>'��p�T�t�!�ܼ$Z��䇚�7V|!`E-,�!�Z=X�x0���;a5�8�N��q!�d��g�^I�R�M����'�s�!�U9m��p��E {����#!���(kR4xg�D#�����&��B�!��E�p��ZDk
�6�H����	"o�!��N�T��$��
s�U�E��0t!�MR �,�uIgC��s���5 J!�d�	��`�X<
Q���IB!�DCI��M+�ߖn�&�61!��l��@ׯ�;ԊA���%"!�$X�oӘ�W�V	`��a��&�!�D�&�~M)����!�<�h���7V3!���`*ԵJRIȔ�Ը�R��.�!��E�h��hp ���Z����o�(�!�t�<�!  �RBl�/&�!�d"v<�0�ȐQ=��JЍ���!�$F�7shKg$�8B"p����S�!���$lG ��Ȅ�^���h��=S�!򤋿y ֨�Wl��h�$����V$$!�Ε]��u���[�`U�)y(!���`i�@,���%　��W$!�d�D!2�9s�$CՎ�C M�!��J�u��Ez7H�?��њ@ҏY�!���.��` t�I.a�Ri�o��W�!�DZ�w��	X�C�6G��iA����!�� `��dV�a��4Z@D��My
ٰe"O��1�-!ar�cA�Q�:��"O�h����`'H8ӵ_�V��t��"O��G�@,bT��&J��Ʃ3"O`�h	;��(F'F��F\2�"OFdPqO�`�H�A��+q�H�"O��qc���}�
Pa N�x`j��"O�q���R�f�l��ř�\M>@C�"Ox�x��L*m���� 9,P]�"O�eH@�'_��*a#pX�"O��r�#���l�Wcɋ>��@v"OL]��X3��7脽n,���"O��'@9�x N��)|1J�"O���E�{�tRǝ��I��"O�����9��9�6F�0]2VQ�@"O؉Fn�n�9�W�[�Q*�1$"ORB	<d
��@�ђ*mt|�S"O"5����+d��⠜�q^ D:""O���a[��x�$�ZIL���"O�e+��!v��5 g���!#�@)�"OP�ʆ��8-�ʝ���Zo0I0A"O���,´sC@O�f�"O��5
�^�$�U�́5��$��"O�b,ˎo�p���n�$#�"O����iԽiMΘb�ĴZ��<�f"O6ed+[=y;�xB$R)g$��(�"O���@
(tcFL�~���"O� �s*�N��D��k��,��P��"O������7Těb�J�K�`�A"O4y`��Q�Yܪ�� �o.�9c�"OJ0	�P&��hѰ.�*B`��"O�ؑ�ғXd���$} �	�s"OH�K3��QΜ�A��1 \��'"O(���H�/������!�9!"O����œ+�P��!��Z��X'"O�p�VB�HAt0��COI��*O� �`e�<j��Y����`�'?z���e!az\�0A� G�*�'�¨Ype�QxRH�'
�6*�)�'v�(&)��QS���Wj]���`H�'�`�2&ɴdPn #7`
�N>LR�'$�%��ʜ�8/�S�k]�~�P�'	|����/d)�V��|�5)
�'a��WF���kE@$c���	�'}��H�C��1D�Zb��l��'���V(V4Zќ�x��P\$���'���9�a
8'�
H�gdE��H=c�'K(y����^�:���Eݢ��'$~(�g�+���Q�9B�8Ě�'�5��9�e�G�$0ڵ��'Eޭ�e��[�� �a@ֻsȈ`�'�l�y���)����ө�1c�^)��'�2`3�C
��L�x&`׼MY����'V<(�Y�A[�d":�aR�'�:(hƍĻH��)�T�2���'�X}ҷ Ԡ.�\�����1&�2�'�Ɓ�C@�w5Ԋ�(�r�d��'�\@{�,�P͌M( #�&ᖝc�'@0�ڵ�X�W(.��gE�P����'t�q��Ƙ��p!׀�*A),�Y�'R	�Q#�3��IWK��b�
�'�>)iD�X@��V(�shLt�	�'G$*�ٛWb+��N敛a �d�<1D��{źыક!A���g�^�<� �HC�(\:V_�)՗L��%a�"O�M*	ל�RE��KL]"E��"O���@y�0Țg.ڏ_8l%�"O��sV�W�|3�V���� "O�
�ܫ:Y�F��z�q˝z�<�b��"1�mٲ-Y�KTl� �y�<!�
�1E}�IJ'�!nt`�f�q�<�1��y��aՃ �D2dXŁv�<�q��Z�x�)?�h�!`�Zo�<!DGM�e[�0�Y�(���8c�NE�<�vE�F� �ťhQLXHV�I�<a���z�����áFF0���H�<	�ذ�Nt[`o:3����N@�<1gi�8]\��ٱ��J��m���D�<�E��"^��xPj��M�ud��<q��<��A�c���c��9:����<��W#|��$z��7�A�ARG�<��9<$#�Ì�-"�e�B�~�<��+I�,��l�KP3��u�[{�<1��#��K�1Q�|����w�<� f�,[�ج��dĮ+����7��H�<�dJ߃�D�C3�H�)��<z .�@�<�P�>U���e/�_�hZ��H�<qt*Q-�����]�F]i7����y"�2R:=h�i��2��	;`��y�^�⡋��ߌ(g�4�gM�0�yrHS� � ,�'�`��	�yB�V,dR0�"f�#��Z�Fغ�yBD�L1��RM��M,<�v����y�az$��
ٿG� �k�/���y"'�-?O�L��睠pH���6��/�y2����Q9qO��T�������	�yR�R	3�.�u�tN�%x8Rx�'Z��!��ݮ?���G�7D�-��'-1P�܀Lˀ��TɃ�w��'�Pu�D��/�d�C�+A(wy��'��8)6��7 �X��3%�o����'���S �';:3-�'x\~���'�����-�7~ɸ8C�GvLnT)�'�pY#��_�WK����늄:�B���'r���]�f�$A�e.��̲�'"T�#.ʇ_�b��W��>+��y	�']04X�܂@�f����ՍVk2Ԡ�'�8���G �2�<�A� �P��p{�'{����"׵Z�{��O/S@z��'���R�
5���cd�ۊYs-)�'j4u(挊�^�,���L��ea�'ߊ�!��	��F��4y0�	�',�bm�Yp���`�Q�t��1"
�'x��V�\�FK������.i=B4
�'��Isi<V�B��섬d��!��'_���7 ��
���T��`6f���'-<�׮�3+	�Tu`N�Jt�+�'���Y�)Y��yzTL�Ji��i	�'fLl��N�:Sp�xhġ@"/Q����'��!�A͇,7yV)�c�R�.հ�P�'��x�1���h3��MK��� ��|�<!��+)L��:PlPe�ŋa��q�<y��J�>���d�	c�TՓ$�\m�<1B`
Bņ�q�.Z�l�)*�(#T�X)u-C?/V8�%Õ�;�P�f�3D�$���N�K�Fš�!��nZ$�+��-D��+�K)uV��d�$x�&T��[�1ƴ�*� ���~��"O� ��Pƍە6�th�,�+d~M��"O2��V%5:���cN�Ta��� "On�K�jT�"�l�H�lͱt�d�`"Op٣�ˇ�/¡�%��/w]B\K�"OB�'�]�{D��8���NV<��"O8�rQj�1.O����X�\z�"O,���"H�shbDZ'��4����"OP8!�D$f�f)��&ߥ�Bu��"O�M�.K89����C�H0b!�""O�hchU�^8�ucb R�B�"O�xB�G�n��cM*�"O���T�U�X!��g��e(����"O���`� ���r%��qj�y2 [mVN�0��;gruc��ی�yB*��d�>]2�&H�G6e� �yr��� �^A�W�<����X��y(�4�,�%BW�,g�t ׈D��y�O�{���3�I�S�&̓ƅ���yR�[0�ĨX�DD�.Y����y�L�*����F<4�b%��!V��y�͗�s�T�21؃{��6Ȍ��y"�ķ{ϪP0��Wz��	���	:�y�Άz8��D�S#[�[E��y�# �*���Ŧ�)Q��ԁ$c��yRN�3-��<y��:� x��yRjR6@营�CkZ�H�.���y�CQ��k� Ĥ�D|�¡�	�y�@Y'^��2L�,[l�� 2���y�mF�L�RA�U��Z�xb� �y�&��pk�YcFI0��@J)�y��3c�Lp�C�&��p�WgK�y��&����+(h�
�SG��	�y���/H���/Ȅ�붂R��y����o~�����1H2���@��yiZ�����"R0�hI1d�/�yҪQ�)Mf��v���,��2�%��yBiE���@�����R��Y5�y��=�](#���j6� �y�f��v�ԡ+Ud��)Q4�"&ǀ��yB/V#E����@�ZX�s��^�y����S�-������S0BfB䉚r{�#g��+��}{��ԉsc|C䉢Q� �ƬS=q������02�XC䉴����ھq�U� �B�:�L� �/s�@��T��o�2B�	-8�H2�e�B�~�h��$�C䉳7X|�1b�y�r�B�*�T�C�IRC*)06d�3Pd���ll�B�I�J���aŏ>+�\��&���rB�I8�b0�ĊW1]+|ŋ�)W<)z�B䉻XUBl��0m�p��LR�=~B䉴:��!6�rgJ=frnB䉸a���u��'&���5≹#ZjB�I�^P\����d��$؃���D2B䉹Y3ʠ�3E	?ƀ�'�=uR�C䉝a;��c�*�b����I� *Z\C�	���۰	_�=���J��@|bC䉪N��0�f�~�t ��ߣx��B�	��iq�ݛaL@����u<pB䉀Vnĵ����I�R����D��B�	�T؉��.���2������d:�B�#�dxa	1p�̹2ě9H�B�I 9\�$Q�N�C&���B�	=:k�	��н6'�}2���/"��B�)� ���qcҡU��Qh��/%�,L��"O�;�-䚄ـL ����*"O6�jp��v}�@3�L<D�"Oژ+�/e���@`oH S����2"O���'%ʉ4�IX��N ��e�A"O�mj�ĝ� �'C�*l�FE�7"O��B1�R�Lz����Og��a5"O�y�R�N9A��*cᔬu 2x@�"O�-�� �8��i���S�:��p(�"O���!�W��a:q�ö�n��"O���$�wz��D�܅q3�`�3"O8��6K�m���
5'D�<`�!d"O�%Z!`Q�o�*��[�뾠�#"O��EʩW@�[�Cb����"OB�c�  U&bhm�h���"O�;a�V:Fd�P��!�)x�"O4�S2M�����$�QA"O�|��`_�+��� �|�V���"O�����)m�8�B�R��ԥ��"OR�B0��v��RT�Ɋqp�|q7"O����ʲB�`�`UH�oe���w"O& �#���U L<j�j�)	GѲC"OŰ�jV�{�>������A���`"O�c��ilȢĀ��� 8c"O�Ѹ!O
,�z�C`�)x�P�x�"ON ���۳���*��H2g2n�cw"O�#q-����L;u'�݊�C�x�<�!�Jf��6�V3i���4"Fr�<�ы���DRBJ�=:p9 �h�x�<�4�ߌjpf�0��F�|Θ�e`Jl�<�"�f};Ubö�4�ː��f�<��ai��9�J\�]��Ö�x�<!�� E��V��_�xuSS��}�<�F�E�v���I*U�ČhBCW_�<AvA��!g���,�Jx�yQ�Lc�<a2'�"
�`pe�a�
�� Xc�<��B��B�X8
�¹��͐GX��ȓT#,����%�Pe��)]���Թ��@����L* M�9F���Q�*�9�b^����˅MLq��Y�ȓW.T"�N2a�� t녥1ҾY��l��I�"#�,�@�䇤Z*��ȓ��@1�.�7B�Dp�G�X�;�@��ì��Th
g��ȓ��G�,WZB�	�z��I����Y<���׭��0FB�ɾe��`��GM�K^b�֨gf�B�$>a¬H%���9-��eL�k��B�OTȹ�fh��� �0Tu�B�ɒ{�n����ϠQ����b�t��C�	�@2��z�l°x�ʱ��C1o�C�	4]� PXTNM�JͺhC*?�C�I�n��Q$�	�e:m�v���C䉪&3D����{ld��Ç��X��B�I�Ğ� $�ğ2Vqz�Kn��B�ɲ�x �W ɞI `��ēg$�B��T�`Ua`m�.]�}C3��;&�>C��'h�BwS(9v�A�b��BJB�I��r�����9-�i��I�R�hC�IpS��Jʴ\������81FC�	-`|��'����E���euTB�	�{��= �o:Ll���L��BB�7ja�"��ӆL�j͢&�TjhC䉗]�2ۄE�J�r8�`� �C�	4N6��灈1�@�ѧ�f�C�)� �]	P%�$(i��t�$�̸Hg"O�m�g��LE��	^��,�&"O��rhʿ���`aǩ�R���"OV�(���>hTX% އ3���%"O���"�K ��Pe��Y)���"O�H;uk�*�H,���!'��c�"O�\�����#>~�R0,�<M�`�a�"Oj��Վ��Vi!%"�6)���I�"O��
ei^���z�`̑U|�g"O�u+U	V�Q��U���G�bH��"O XA���)�49X'G"b;��9B"O* za	��p�ةb�+�	~^��"O��� ov�a�aJ@ ���"Oj�B���{X�nC�w_�`��"O6��:�J1x4/Q�hJ�['"OL�IէT6��=P�N	5�����"O@L��LބAP�H�NN:�9s�"O@��J_�n��q;�͜���Qs"O
�	��	�]$8�`Tk���X���"O|ȧ!ߥ	�))sl��j�(�"O:]c�S��5ck�f����"O"����T��GI)R��Y�e"Oȕ���.]D8����pB��Q"O*)	�ǟC�P����8*�$"O����gS#��Q�EB̲~��T"O�t~Q�VΕF	<�cB�[�j<!��E�4U��+#�Q?W��!�@/��&!�ϭGn�� ��%k��T�w��q !�$�Cj���MS Rp����MM.&!�� {9$�ч�Ǝ�0���!�=sKp�k�D:s���aȿ?�!�ǁE,Ќ��ַ`�yxQ�V�-�!�䛭MU�ѹÆ�Rh �`@��g�!��Iti���c%�~ ����R+�PyR�^�k������	D^���i�6�y��ǗL]�}��H�WS��@�ϟ��y��/y��:�K�H0�fcȝ�yrhC�r�y�DHD�\�A��6�y���)�FI���G<�T��E���yϙ�k��ۓ�P�4�������y�Ŕ�2ڬr\��9c�P"d���'��!�%!��FH4E�Rdŭ�y2�'#��*���*x��bM�	sNI��'F])�c��\j�Z��2*����'�%Ч��1�r���Dx�'�B,qF���tn���q�p0�'��ڔ"�7w�VxZ@��94����'�f�6��tC)�d!O0`��xS�'�.�A��@\}�������'\� � !�z:HE�AŇ��
Y��' `���D�0�Vy�"BGj�	�'�0�c�31̔A���c�� J�'��d8��ݠ%	
*�aP�'�@����a�J-�!�[�X�� ��'Nˇ��oÆu3�䊚^���"�'�&�`��$YTh��K�Uj���
�'�$1��BY� R�1�$ �w�j9)
�'..�����	5��S��S�a'�B�'�B�⯁�e7���3���^�0*�'/R�0U��4�pZ�M����Z�'T�q�-�8s�D�1�֫R��@a�'px�{d�-����O�����'t�;�fIW�J4�$'�%6
�E3�'��%���˂-dQ4��?5g�8���� ��������- �FA#FÐ�i'"O��A�7Swڅ�c�F��@S"O.l
 HmJ�S��A�<����0"Ov�8�憹tԀ�%�,o�Ty"O���U��Nev�)�N�1r�\�"OZh��a�\y|倲���1E��"Ot�� �,d 0�R�3A�^��G"O��5��L<�H�e��a�,�c"O��Y�e�tKF�k ��@? $��"OepglM��u�k0a#��p�"Ox�$!0b[н�g �t����F"O������9Y���3��.ז9��"O|��ǆ)$�@I��#
�l�)r�"O�iS�-L��sb�^ʚС"O4��Y�rpLh	� �?ɘ���"O���UY+^JeK��a�,9C"Od�q5�	XXl��ʉo�`�4"O�x	Q�ߘZ��u(�'��4��\�"O�4��E)!�E���7~���H"O~9A2��-p<N�q���[mxK`"O�EP#O�	���#2�%Ydp�$"OD{�� )LeR'�[�B��A�3"O��9R����8�sl&6v�b�"O����Ӊ228<��KE>[c��:�"OF���$^�.����%K>�#�"O^=����g,(�'�x��h�"O�JD�
v�ti1 N,l��h�F"O�U��n��i����1�p@�"O�AJ�q�b��g�����#"O$@�@�6+iDi��Η+�z]�G"Ohx`1�H7>�BL3�H.P��E
A"O� �
�S.��k��QJ��]��"O����o�+e�	"�KɑT��@t"O8�J�� �~�8z�DD-|SvH�1"O,1 �ٓ��5(W2���"O^4�t͔�/
e�Ŭ XFƩq"OP�a�'6�hu����;C��0�"O�83��@crUs��$lڢyI�"O� �惕5��hC��U����D"ON`���	:�j�cb���-��R"OJ��O97{媷�C8n̎�3�"O����OW)oݱ��T�v"OL�{��^��F�{�,_�cP�+q"OVQȀʒ�)Ru�2��I|�zB"O�e���J�b�K'Ϛ�^Ң|��"O��F��(E��ˀ.G%��q)�"O�4�'�F�Pٖa����)�� !"O��Xu�&+кݩ3�[�P�`"O�mi��@�M��xb���Y���ӓ*On	:���8T'���@�3C�ڍ��'Ĳ��n�3�p(x���N:����'*�pA�h/G�2y���Q�D,�x�':���#�$(����b��hmV�1�'��	��į=�a�э�Wx6dA�'��d����m	f�`��Q���'.���g��t2��­@V���P�'j>��U^!�J�s�Ɓ?�h�r�'7�e�3��%gnup�dX0
�L�'z�A$�]&D0�Mҹ|��h�'Y���O�)g�zE�6��GZ0�s�'Waٶ�G�Ѐ�h�Yt�D��'`=�t) &$3|Dц���g�~�0�'ۮ���f^�z
�xv� �dp����'Q��R�%�  W&D^�M���� ��{�.I(l���c�Π7���e"OB�E�
�=?t��͛>J�x<@p"O����&/�&�8�+��E�����"O���℄=R�=����4���q7"Oޑ1p6��� [�#vQ�"O��Q`g�Q�8�����Hx�$"O���,�F,bi� yE����"On�cw�͘;xH���!ȥ�Dap"O�hp��`Q6���o�^�B�"O����i4uۢ���o؃I���&"O��� *ju�q#O ��r�($"O���g΀"g��� T�n�z=�w"O��J��L�*R*��W �A�X�"�"O�0�:M����gO<���"�"O@��F�u�������+��	WO����[!��9!��$<�Ek�XE!�ѱOKp�bEȢhi�6\�'!���Rtr�G>��"@�\�Ew!�d֥@9�<�6̏�%F2�X���7 !�ԋ+SZ���*d#bp��L�!��Z9EW hի�5�%Zpk�}!�D��ASRXH2�p�pMs�(M�uQ!��O�jp��1��Y�*��ah�Z@�	U�'��O��ȁꓗ=����-ǵb��C�y�	�0tXZ�tÄ�<<�Ө��yRT�}#�)P��w<)hA�̪�y�@��Jr�����}������9�y��Ɯb'��[s�6*�n�AP��yb!�K<���BY���T�E�y�iLQ��a�̛�Y*$���	� �y2!0Zŀ�xS�^(N6 ����&�yB�ND*�[f�A+ ���k�yri�M
DH�&��5]ve����yr��g��H��7er5 R
��yR��t�5{��=�`�9�&�y��I"$)���ɚ�6fx�!���y��ζ\v�&��8����FA��y��R�?DJ��	+�عӤ�L��y����2��!��l��)��5���Y)�y��S�NR�x-��%�>�
����yR*�
pC��C�X�*(Y;F�֐�y2F�(��%��0K���y�A�.lڐ�g��+�XU×o\��yb�lb.4�ōL�3����\O�Igy��'�T��R���T́B�W1 Uy�'a��!�e�T�<��m1R��	�'����Gb�R�<4B.ŉrz���	�'.�X�cT;t�X�'�|�*(����[��^P�Xv��8��լ�y2oé7��qg**;�uP�ǟ �yBJ�(H�.qd#K�2H�1�C��y⁾*�8����Z�P�*���)�yrj7_���	�j�Z�0<�D��y2�(Tuq���$V�P9�"З�y�aZ�8�8!�2�J-��4���y�Gߕ8�2�Z��%K5�]�&U��y�BTK��9�,Y�O<I�p!���y2�܇dAl0�Tg��~g�ԡ�ۍj7�	Lx�|�t�!�`§]0&���Y�!򄌗"2��xh����qe�<B�!���66�Xe�6�̿D-���UH!D�!�Hu��i��˅Y���&��:�!���(L��k�O:3�W�!�d]<a��qse��r��cܥV�!�� \�����J�*"_��xK�"Ou�a`T	�` ��恭&{��`"O&yrv�F+)�݃�Bnw X(6"O�Y��#,����-��A��"O���fF�7����B�A_�yJ�"O	2���>Y�����jQ�-:�"O�ep�)��W֐����Um�4�"O�I���՘dO�.JT�q�T�	jx�Lz�eפ)Q.��2 |�kVn'D���iX�:_�x�v�;9�4���%D�D� �Z�D1Pe@�mۺ�+b�#D�`�mѱ��
�d����24b!D���(�m�h�cp�K���$`D�<D��{V�]l� ��I�]�f4Ҧn6D�x��Jʐ:+����F�g`Z�Kg�3?��n�����<,��xs.Z�4�����Q+@;��M8]���;R�ϽN�}�ȓ%�`S6�T:	�=��LU�>.M�ȓR# !V�
&D̡3�B���y��e�ꍐ3����N����3M
L�ȓ(�pXS	7+в�2�ѱKf�<�ȓe~>Yq O@�P�b�@%5"r��NC�}+�-D6��"��� Y�H��K��{u�̹p���x� ��Tp��ȓ!�t4�g�CD���g�T�j[(��ȓ@���AW�K��ׂD� ^p ��d'")�&�c��dIF��h�!�(D�i��H*�1��h��qU����*"D��1��$
�1�B�}�2??Ɉ�ᓒF�у�k�	���Q�۸	V*C�	�O�5�����Xi��Wi�. 
C�I:
s��fcX+#~�iס_X
�B�ɂzf`�X3BG�7u���reS�7��B�	0L�|�0(˵L��P�d(60dB��?Cϊ��B@�A*ܓ���l�B�Ik���E�ء'(��ĉ��YצC䉣c��CƓz腃�c�/{y(C�I1��A@�`��)A�P�P�*B�I��$cD�N0�т%��N��C䉂e|,��F��uXĂ���`.�C�ɦBl��K��S�:�8�3���>}�nC�	�yƒi�P.��V��Qa'F3)bC�	
W
\C�!7c\B�'�5v�B䉑�H�f��,�<
qOߍ	vPB�I>C��e�k��a=�$���±,�B��V����ɲD�b`��Ճ��C�I)V���d�Z��qAd�Z�C�X��@���_+�b��K�E^�C�ɾcx챳L�*?�(\�r��e=�C�"!U ܻU�Y�UUF��&Ň��(B�I�Y�(�%B�m5f��E�df�C�ɿyv��)@�ݙ^(�R�I@�+͢C�	�<�q[cm�{L�0sC@�MC�C䉔i�f���öPR.M@u��&dxC�I7r����q	R_F,3�흣,-"C�ɳi�l��1�jLk��1 ]C䉀j�������4z& �� [�rZ�B�I7Pn���gR�`"��!���C�I=Mۖ�Y ��ҹ`�MĊZ�*B�	}
���?*��B� 4r�B�6;^HK�$�u[\+RI@�!ɚC�I�9�.����Q�������޹YC*B�I�jwҩ@VnOL����<,B�ɌJJF �V�3�\p[�`�0?�C�)� "1ӌO�*6L5��ܳ{Ȋ\�A"Ovy�t	�j��R
>��)�'"Of��3@��x�b�;|y@��"O�۵�P�9�nѡ$�Ώ:o�v"O����l��;�PH{���<v��`�F"O�B��t-��@��]6&)�e�0D����	7����7d���Awh)D��Z"� U!��ǥ[{l���B�4D�\)���0Q$cI�v�����B2D�$�oѝx�\�[�BJ<Ed$�rh,D�Pd�Ʒ,h=�6̆�t�4���M?D��
Q3���!��':�SqL*D��KBh��-c�L�Pl�\z�T�&'D���4.�=� ���J��u꤆?D��6�w�f%�cF�-�	`#�>D� ��GN/XC6��!*҆n=ZP��8D�x���@�@ϊ@`ty*D�P���«NH����φ.M�^L�u$(D��1���{���6�3/�.�R�%D�8���ݙR#|HKҡ��	�D,��%D�qU%E�T�����8�@�&"D����b���Rg&��� D�,	��D>G�TUq��
F �5���=D��u���3xNA���w��Ѱs@0D���.V�/�Ő1�� t�IC#-D�����K�o��s�`U.�TY�8D�X���=và�Xc�UMY�a�5	7D��AOߊ(F.���	Պ��A�K(D�@��lU4� �a�0y��$�3D�<1� �,8o�t��D��%y��;D�\�5��1)����&/��d�$"$D����5ZPM��` �Q�� � � D��R��Z�)��?	�`y�2D�����+k��q�J�8 hDb0�-D��uΆ+ͪ�����K7j���n'D��3��@c"jPQN��J&x`��$D����e��CB���1n�q��� �e"D��j�S�%�(��34b��f*"D�(��R�ss�[��\�T�HX4n!D�x��VD�P��Wg�*Љ@�4D���S��̨��F(8bF�?D�8�w º͠�����U7^ 8Ua:D�X����O�ԍ��
�C�7D��H���$�b����]�U1pg#D�L��e���\���犇q���o3D���$m��22�m��(���`��0D����I�?�@e���+
hla��4D��Z%�fx�ς� �P`�1D�h�b�I�T�Nlx�,�Ct}���3D�c�H�?�P�V_�>9S`�2D�`z�n�v!��x��:�j�(`�/D��0dÞQ��8�a�{�=sF!D�h!$�ڥZ���ԩ(�kd�>D��Hv���$�d���[��=D��kc� y<bT����@�ư�3�;D��ۗ�Ry�t���"r^�Q��9D���GלG��ɤM�H�򭃣�7D�DKbi��R������L �䈒I5D�|�w@�؂7A�r�
�2D�
ՎU�#���}�.�5(!�2&�n���M�.mAR�X�!λj�!�d���8���p4B��b�8ti!�dĤZ�-�4%�ZȖy�p�\^[!��H2)c�iHl���P��0S!�� t4�v�@���x@�ꇮps(��0"Ot1C��ߜ{��ܫ���J]���"O���7O��.���pj��DY�"O�<+SE;&KZ �P� �D���"O�u@�,L~�1)u��,:�i�`"Op�˖ �P,�s��"O���e�$�t�XUj�5d�|P�"OPp�6��0{&���� r�����"O�E��F'������Y"O�=�7jݸ-�*5�S���'Q
�"O��;��'k�8�Ä�Z�D1��`"O��`g$'�y�#��� �Q�"O��Pd��~F���GG|d��Z�"Oh-�%����d)#F &3]h��"Of��� 9i.<�Я�8Xԭ �"O��q��7�B`OaH�K�"OV����D�{ ��P/�(<���"Ov��,E�� ��M�E0�-k�"O, ���9U\y���?R��$"O���V�� b]�']M   �"O�1��Ǩ0�J�Z2偿8B�2"OZ]��f4G�P#�4i� �"O> s�� t�`�`!���X�as"O�� ��͕i�L���4{W�m��"O����Ài�"�ӣ�W�V����"O�TЧ$�8=(��0e,MO�U+`"O 麢��>����N?Cd8D��"O��'� �4�*�!э��ER<H�"Oz��5a����[�]4X�X�"O�����ς��\3 ƃ�Kxx�3"O�	�3"�/-���1Ŕ�Ol	��"O���$�K�~�iX2�W)~԰��"O��)�J%W�>�	փ^�w����e"Ox��,u��,�Т�bnxP��"O�����X!K$��#`��._�LZ�"OP0"l^�%|#F͸Pb4e��"O~���,�"� ű�g�o��x�"O�h�bl���1�q��I���u"OJ!��İZ�y���>�hx�t"ORlH���
22# D6zi��03"Op��ᄓ$4�{5�׍;2఩'"O<�8�'K�>� Њa��#C�dy�"O��#D*	%����C���6��qK�"O�堧��!b��� ���N�"�"O"a('�,<T���$J��@9B"O�T�g���D|"�'ƭAt�E�g"OPr�'������c��.Xl	��"O$y�̜*K��R�\�q`�i�"O �FĘ��T�ab�+��xba"O��s�.�����	!T"OHݢt�Ee�@�k�'�  ���$"O���u�#���K��3����"O�\��ʉ5DX�9��M�YB"O="�(��t#DH�,=2��D"O�UI�-��tk�xP��<�a8�"O��/U�"t�AweE�^�l
�"O�r �[�9�R�O|�d"OX!��O�J��k�b�k:�)�"O��!dD�l:�M��BX�HY�@�"O䙠ւ�G���t�H�,���"O�i�gܜvk��*��A�ڇ"O��&�Q�!�v� �P/6v��&"Ol��'�9uZ�óg��]�>HX�"O��H�
2HQ��$�<~G���"O� څu��"��w��=�e�t"Ov��sbźS��\cb��]��d1G"OV�3�G�T�+qa]2yB(� �"OTRC�N�;+���׀�*c1��H�"OB�f�[35���s۬v-B"O`E�T���K���!�;(�� �%"O��KRKL$�0�{���?GH�"O��&G�* 6n<)!�(@9f"Ovy���(wR5��#%��<C!�+y����t�t@���!b�!��s�`=A�N�su� ���^5�!��Ĉ6�T�RTIP8Ԁ��LO#!��߯k�8��	�]`@ZԌJ: !�F�V76ybС�|�T<��,�p!��Z�D��X۶f��0��$�%���!�$ J��W�b�tP1O�)�!�D��^Rb��;sG���HE!��_��xX;2�X  ���I +dG!�Q/j�*�7OT5�JI&	4!��Ԓ'����"�B����1�5 $!����� �
�h��E��1xv!�D@$t3D�zQ�v�ܾ-8�`@"O�E2-�jnh���6v}� s"O8XR���xޒ,P7�_�l���"Ob+��	7�.�e���f�\�
6"O� ��76:]@d��*Nn%PT"O�mcuc�B�8ȱq'�WV�x��"O�e2D��E%z0B���`?����"O�mB�dȧ*��œS��n���s�"O�qsa�V���Ё$
�m�܃"O>ԓg��~�v 3�U�\2���"O�0C�.Ҽph��)Jd!!�"ODt�%ܝ��f�;Y$v�07��W�<�f�D<7aʥY`ǃ�P ݒ&�CR�<aqL��j�4�mƱO�N$�D�PE�<�cG�:ߨ\��w,�)ь�C�<	5ꘒV���*��%�
���|�<��A�sZ����1x�8�1�A{�<�.��3^��4��'>!���Em^n�<ABkB�2�Hj�g�'-c4�sF�<q�#Αr�y��'~�� .�z�<!��C&Ҵ%0& ?Ble��s�<�$�ݷO��h��l�.V^kCD�K�<Qḡ�P�W̓5���W�JO�<��*��P���G�z1�<J��M�<ق�PeP���5�s���C��^�<Q��Ւ`Y��h���pA��1 r�<针
0Yz.ł��_N��Ă!!�j�<I��آ� �����Bl�"��n�<A! �>{�{�o�@X�!4aa�<2�S�}�b j��R�zO��2�F#D���Vo��zZbXhҀ��x�$� D�����'x��vnM�|��Zu� D�H�Iӿc҉H �0SL.����?D�� "k�|;�q����;F�+c�>D��b�I�)[���-D;�&�b��=D�L���@�c�A��#E�:D�x��f�c�.|c�M\(��ؑ5"7D���6�E"��up&L�0���"�E5D����9�H�1ɝ�r��$��J?D��#�L�X�ٱi��5p~�
�	<D��i�&��y�	��U�R���c �:D���Oڪ`  I��X+�N-D�,� �P>D_.�;b�S�y��A�,D�� �-�cѶL��T���]�"t��"O���`A�c*�0W�V���"O�myw��4D���qjćA 1!"O��'�#F�S���S�@a"Oި"bʇ�_2!)�~���{T"O�y���Ιe���r5�O�媥QA"O����Jr���K����z��9��"O�(��I�..o����+w�:]�'"O�٢�
�>j�WgH�hv~R�"O�5YU����$G�,\TTAf"Odi@�/OCv�pǈғy$�5"O�$�3L�/�����,\h| ��"O`��e�_�r�X��2G5_r$��"OR�[�J�7��a�6b�@��S�"Oh10T�F�h�� �bG3eUl��Q"O��S�����c���x_�jU"O� ��Ǫlp��m��{N���"O�����R�ke���F�O)rZ�1�"O�u�c�?K���`�b@$��"O�05�P����Ʒ&[ $�4"O �&l�&4H��I	�j���E"O�Ms���2s
�Be�܊��A!"O0���ō;*���Bu�@�92�AXr"Ozi#b�4*��k� �k#^��a"OH�.
 B=��5 �>G�Q�6"O��{gI�'Z���Q
� |�5"OF�S%��/w��y�3ÜD�"O@�UC
�3U
��-�Z�H�"O�I��@�0�0�k�LWB}�Y�"O*��nA1<����((Bw@�`�"O@ԀfWn�����S�a"O��{GE�|B�CO�A9���"O�����7Tݺ��%��05`���"O��1,ʢ�M1�	��(h��"O
tyrZ"o��	��I�w�Tp�`"O�X[������Er�VD��'$��K���M$& �F*�3me��*��?�ļ<�J~�'x�d$k���s��_�)V�E4j�Q�ȡ��	Y�h�����2C�B���Z�8HԽ��'}����MA���9"�"f��n P#q���cSXb��;��ď�M��O:e���+�P�+dώ�ȴ!#"Op�����-*�l�i�hQ�Q��	Q���6�����f@�6�!!*�o��R;O�E��y�������n�.yi�"O�1%��A�hC�R�/�
 y��3�Ӻ�wR�1���!��8��Qp��@�-ړ�0<ɒk5nh�6/2��hF�S�'{铡�I쟀!$��\Tli*Eg��*� 9G�*D�� `�I fG�P��I�,zf��7"�	�M�O@c�D{ª��rq��gY�;�.���(P�O\�=�O9V=t�;v
I��7�L ¡O4!�E`\#��S�� �z>q���O����P�� Y!���^7y8��O=L�!�ĄKv�l��	A�v���`�\�,t�'3��^8���ć�"�,Ks.�4ZR���.����zZ�T�I&&dX!cQ�SWo�"<���[���d
Eb��ҬiA��S�HC)%8ax2Y���t��V�}ǚ��p+˽6R������z�.�D؟�[�54�&|itĆO� ��׋�OJ�=E�t�**�~�#�,.����so̶8*!��X�`����_���.Вb�!�d�]x�D���E9y}��,�.���
O~5pA�-_�-[��B�n�	)7�
�HO�*�*ݸ��Kz8ISNU,!xh��S�? ^�X� �%�"���$J���C�1�S��y�*�;���W��򅫧ʁ��yRh��wpA���/��Q���N�M��Ob$��O�H���C��Ĵ���p2�2��xr#Y�6��d Z�4j�5BF��/�y���>q�<�CdP<�b;%��/�(O����+kFmIp�Y/i	P�ʐ�Py��!6Ύ���ƙ�.�V��B
�yҊ��O?�a�O|��a5�lz,]�p�8�O��O�`�G�n}��z�
"Ti�u�>!	�M �y�S�پR�=`�D-��E�>���D:}B�(2�bi�q��{8���ǁZ��y�M�_òD)��,{H9(����HO���;�P0�3HP�M��\�FP,�!�$�10����.�/t�p`�C3�!�ę�Rnh�"T �P�9Xu&ގ:R!�F�[�6�����o�x�rb��#C!�$�:2\���2�
�Vv�����C�jA��qӔ�G��<60� �ݡ��Z%L�&�0?�'��I��������a
@D�'\�9���f��!Ju"ps�lד��'�����m��w��aô��k�6$Q�'W��h,�Wh]:#	,ުi�'�p���@�j���ڎ6�B]�'����`�3T�n��f���hi�'�:��'oC�j� �vKK�[�~�
�'(���U&�V�������W�"�1
�'���u��z ��$ ����	�'O�1Z��	�#O�Q1D����j�O���L �|��ӆ�+j�"`+�b�'5�}�����N��7h�`��N7:j,!��A�f��"I�F7Hв�	�`
��D��J��%���k����yB�C�~��cʧ`|V�����y��)��NH7aƇ	�x-Z �ҲV".�����w�(@�LB��2����'ja~"%]�e�dXK�38p����6�yҍ��`�$�H�O���ab��V�yr��CM���(}���)ҧM�y�iK�}����Ǧ�@�:�Ba� �yb�Ԏ Z�LJ���.��]1���y��֡4�a�ȎS���I����O���韈E�O��]�y.�z��ۥSa8�hQ�S�v}x��*�S�OFP�ӆ�
d���H6'��^��@��>	���)N6Z�ղ�aL�Ddr�3�&C��	� �����l������lC��<t�G{�O�t�Dyb��'�th+@� 6 Iy�MD��yR�X�,���+|�fa�a���yrsv�(�)�� ����g�<�y�B@�E��EW�+���jGd�y�)�'@��m7IT�3`��a���:i�扄�#���:	�pj���̞������?)��Ԉ�ƩS����95�A�_u��o���O���6Ib�\�A�lB--V�4��':q W�G�6������#:Z<j�'Өi���S�zK�2� ܌tT}���?�Ic}�=Oz���`��C�z���]Ұ� �#4��;F�ӪFK�E����?@θ���>I��$!�S?1���D��z�B�&h6����B�b�<I�D[!�D@�B�T<dyz��F�'��x�# h�)���:������y"��C,);��<[� ��݊�y��?q��J�dL���4x䎤����df���f5[��a9TN�c��w�!D�� ��f�Z�jX��s�"W�2 S��	P}���ۉ.��,����_�t �7��*�!�D;1����!�vM��Ǯ���4�S�O�.	�֩P	f�H��F�%��'��MHP�Ա&q��E�3b�|��O
��ݴ�اu�6��=�B1j�c]�<}�`�@�#T�B�	�zQ4djtGZ�zA�5#5��:�<�˓s��:'�;+Q8# ƒ[`���hO�>Ej�㔬&��"7�[%�Z(���f�@j�'y.�Q`�K&�J� �I�eenq�/O��N�S�O-��h`H�32��yg��)�d#��yd�)Os�(��(n��"�|�'3a|�,�
V
�h���ڒ|u)�֍@���'���yb����T`�(q�!�t[�!��1O0�=�|
u���(YY���U� \ �Ǎs����$�`c.���l�1�<M#��R�i �Fx�'ےu� �g=������|R:��H>���%}�S�x������σԂA�C��e���^>~~dC�I���dag.#��Y�\�+�~㞀n��y�\���ON�ӒQ��uSWA� 
�'߈">A*O�7����d�nĺw����3��-X[�Y�ȓ?��W�.\j����)c���2�'��ɍ'���jƽ���)�L�W�nC䉷WK؄���[{���u�ۉT�\#>���T6fܒ�p�Q>I�&ܢ�Tx�!�D,?�^!�T���?�lIs'A3R�!�D�)/��Y��C�#n��!"�M�2o�az���8;p�� �T���"L�$R�'}��w̓ߘ'n�[���HG���+�pJpq�
�'�����ʎd:��ek��b�	�' ���"[$�L8IO
��R�'*LYg���U�9�R�0�Ȕ��'��� �F$cPh3�� n�	��'���Ղ׃>P�s��
r����'��p�!g��D���Q�̩����'V�	(#㖁�!)F��[���	�'�@�A���*�8��uƙ�'���'�H��&��z^��pM��t��[�'�bz����ڠb۲>T&�1�'���bRA�Q+�|2`�,:���(�';D} bY��5��f�e]h`a�'����a��VPP���U�+�'��Da��QB(H|*���O",��'���(�mH�Lh�ͱ�4e�]J�'`�\BA*Фl����ΚY[���'�rq6��)tq����#��M$�c�'/,�r�/yu���Ť\�7Ӿ�H�'��٠� �A�PL�/���H	�'�:0�l o���r��^�����'J��_3"��Q�A��^��,`	�'�ܬ��g1M�����1W��9	�'Ͳ1��'�O�V�S0a�&R� ��'񊙱to���4�[7O���!�'����w�^�FaV��s��5~l���'^��d��2c�X8.��Ԇʓ(/�uY�N��L��u���X<��6��d8`��sehāF�Y�aa4�ȓ}����"O�)%t�M1�LE"$��Ćȓ@Lȩ��^�$��	��a��1��g�蘐w��3v�Y��N��aIf���8$��`ڀW�R�2ȼ	\�=��+�^��!gEG�$�W9�)��^F(���K\�`��ETA�\�ȓK��9!�Kمt�1r�ډ[uH��S�? ���3
Ÿu��-��oċ3�xI"O�a:�M��jPA������"O��W��'/��eX�/����"O��y�/�S�҄: �ʶ*w�	�"O���Û 4x�*/T���w"OL�sĀ^�ps�P�.L�,aR��"O�|���@/ pblRf�A�!`�"Oz��3(�X<9��$:4�}R�"O@ء1ȅ��=9%�/r��*O�a��.ͷ/�e�^�R���'��� �N)�tt�Ğ*P�p4�
�'���p��!lKf��Ҋ��1� H
�'���2��	!���� �!�&��	�'��A;aÐ�E�!뙄oh��	�'�i2 �=`\x���(���/D����- U��$"�};�3��"D�����@����[Fb�-�#�.D��J[��lՠW-��6��mcS�'D�8�2���<1v�"�@��(,��b�#D��RD��6S�������N�v�96�,D���f�ȐQa�E���Y��3?D����+� �2e�1���:~�q�=D��fbC7~���I��C�H�b�V.0D�l8%D���%R�����РD.0D����+�VAh�m��PF�5rF�9D�h�G�D�[6Tظ��53j��g*D�(pK�Ter�
R���kYĉ�eH2D��&��fW`�X%�I�nÚ���
=D����B�$޼A*�H<�~� F�&D��xE�W d����$pjY�&9D�Īr(�#�Υ�Ba� bm���*D��ۆ���T�e�pkK�"��,D�Lz&Aˌd�L�zdȽl4���%D�(YaA�]_:ti���HĨd�"D���ˍ�<dȽbr�Z�z�8�J�l D�pcQ�\)B�:�qQ��4)־|pb�>D��j�EM�_�E��_��B�G1D���e挊b�jt��_
p�8�H0,4D����e�6l�]�#�[�E��ݒve5D�|*�Z?���JQʗ���M�#�-D��p��/���:#�׊'�ű#�(D�L:��[
P޴���c� ���T4D���g�4^7��1g�'�m��2D���&aA0_��2�e�m�H��7�$D�8Z��w��0�CY�ʤ�O$D�k�E�5���çX`��\�a� D�X�đ�y�+E��>T��\06�!D���.��XD�tb���0#P�!g�3D���eo^4D����*Ҕ>����/D����L*�e�$o��B�ݶ0�B䉸&b<L#v"Ab$��噧�xB��<r.�ua@M�z�p������n.JB�ɕ4V�3`j�u`x�2 %��zv0B�,"�@ˢ�7r	t9�1E�:B�I�4@�ԯ V�fed�7��C�	�c����P�'�����!��*D�L�I��e���J��T�?�$,�WC'D����ᄐx���z"�O..��i(��$D�<��OD$r�XU`'�<t�[�E#D��@��&g�P�r�z���Do5D�0��P���ˀ擸{�v�!�'D��C���;UNN�c�P�R�`Ul:D��R��by4P!���-^Q�b�,D��a�D1X����D�36]��P�)�d+�O� ƀ�q��1D��j�bP�XNb���	lx�Ē��-�	���f�.%D����ȅ2%��1����"\4�a!D�`�%�K+zHT��d�<�$��5�$D���7GV#.	�M��O�:�*� D� D�lV��#W��!��'ۜE�&p�'>D��c� ��� �҂�,G��")D��S6DPv<�@ǆ�!���0s�&D�P���>*��J��Ƶ:��s��8D�����-`n�)X�m�� ���(-8D� �kH�'��者��
���[�K5D��h�O�6\Cp"�5m�`ĨP�1D�4��A�Y �rS��D$��0D����۰_�ur��C�(`d�-D���W�l����1�S ���P@O*D�$ؓ� �"M�c�D�4
K�͡��'D��1���4Y{�պ���m�rq���%D�X�t�Î@X���'�Of ���6D�,�Ѥ�K6�pRփ�8(��a)D���Cǖ�z���k��ԯa/�����'D�\X0(�)u�^5��ҿF���+*D�{Ѣ�PIPa�n��[�`S�"6D�d��^�*�@XP��*"��ly�A7D�P���*�\�fiU/?������'D�`�f'YI4�$���WĀ�)$D�xKt�ɹ%8<[�
�DP��%$D�0���Z)v'u� ,�9&]8��"D�x��tk�	��C�9RU�0�� D��릂Ud�(��-K�`%PeK;D��	�F�e���U�ɬo���,;D�4Sa�̥
�ԁ��WF xA�#D�T�����`gh��,Ż4H=D��ʖM٥UW�����8hW�T�9D� �r%�:R�1@CG�]�
-�T�5D���燅w9p�J",�$sL��.4D��1G�@|iR ������%?D��1eG�&�m:���Nm��3��)D�,`q� 6R*��1Q�v��
��2D��8� ԁ`j��ÞC���e.D��(碂�qv��D�$5&>�CÃ9D��(�	Oô�����&}��:D���gO��#��}�'.A)b����5D�@�U&
a��<�p��TŲ(���&D�t�[-+���hrl�yS����)D��ID���B�e!ƍ��[1�$"q�"D�h��h�D�hJ��T�+B�qq?D���䪃�Fs�=zR��(:p>��1�>D��C�#.���gK�\?( ���?D�P��ٛS#���[��=� &��y��3 ����Q�*�-� N�,�y�E�}����r��ZX��e\��y�dX�.8��Zg�Ǳ7I��B��;�y�)B�2��)[����tn]x�.�y�lA K��h�FL�h%�-�m�;�yr�V�Dh��͙j�2��!���	l���O���(�o�m�
\#vM����+�'��K�L�.8�L�:�,���D��'��ӋSuޗ�a�d�z�N�B�<��غnx~-�W�LS� =k|�<i�k�-!;��b��
'2iX�/w�<���ֵHt�e���e��w��u�<�¯1�q�Y�(���ۄ�[s�<	��K>�N��k�)0��c`�Rs�<Ӆ�E��8�-�z��VLAd�<� "$[����. p0�Y�|�fi�V"O^h��e�<J���i��;��Cp"O�M�$n�
��� �B;Z��x�"O���h--�0!�2�@�<B.��*O�a�rǂ�r��2$�	!0PY
�'�J�#F�#RΕ��D��zձ�'�h�8���4U\��@�EC�@�P�9�'�6�q"�4S_�����0��t�	�'���JQ	��������.'�����'ז��� @�Ҹ��Ս*{L�0�'{�|�����sZ��� Ӊ:��tY�'?��#iB�1�Z�f�f^� N��D{����^�~�̥����t� !L��yi�:�< ��n��Yu����y%@*�t��'�"`�Z]�����yr��Q3�q)�	��n~�iR4E��y�
N�X��Q���w�࡫&�B��y����2�;g�B8r���v$P!�y��5,Ò�� ��>b�\)��P�y"�ΒF��� ).))�|��A��y�{G �Q�:ITVAeZ��yb,�X4�9Wg��@*������yR(
RB�D�_#�=��
�y���`d�͡4��<O^�B%D��y��@�7�xx00������-��y���ָ0G ��j���a��yR���6�I�CC��}�P��MS��yR(]+\�v��lZ�"���*��_��yBÀF�ؘS�I8��|{����y��E��PH��`֒$�\	@w� �y҈Q�$9�82d���0`wf�.�y��RXh�����ؚ`(�h�y�~��Q�q���	�'��y�.�9[����n�&28e��5�y�+T��]KCf�&tP���EJ��yr�ܩ�re��ɟ�l��ua����y�&5D6}��Ɣ�2\]`1����y�H�|b�D�Pș|�ԝ�QW��yR�pL̐��F�X�ibv�W �y�)�X6(��@���� :�KC�y2ڳs�A��y2R��%̀��y�'�P�)xЬ�3w,P�E���y�)�6?8�!���\�rO"aI���y�D�U�H���B[�|(��@5���yB͆�of@�z�GӢo�H�Eݠ�y¨YC�G�S+k��@��iL��y�ǚ�~��@E��7gF�"T���y�3L����醊�FP񆦉�yR�K�pK�0R�/���<���y��������%	\�!�nѩ�y�ڪj���K��L% ,Ƀ�ӗ�y��W9v@	�!��Z��\)�
ʤ�y���"C�H��еM�e����.�y��\��G�Ւ�r����y���D�P���N�� ۴�И�ybh��[�� �#�W�<�s��y��(VR�ZsD�U�)dD�y��B����K�`�J,S��H�y�ǂ:�8�sS�͢5ْIP'�yBm�Lh$�1�[}����O��y2��mq"��tC���SD_��y�NP�a5�p�7B��pb�!B3���y���;�VY�4��#ԌfjJ��ybK�Ou���w,���|��e!�y
� V�s3h�/X������X/g��c%"O��s��U~<�SV��:~Ҝ0"O����&\EA��ɜ	���"O�UТ���W�����8�h��"O��B+��q�d0x#�%n�2�@�"Ozh2I٤�d�de�/�l= �"O��H5�T�At�鲗��=c�N�`�>����
|�� � U4����h�s��sl@�*FN�<mt:)""[��q��nZ�]c��oOb��E�[2U�ȓT�V<�u�iu,�pE�.4!��|�fxƤ�UhP�Ã���ȓ8��eK7i��^��`J���nM$d�ȓ)��&lҴ{эЯg�6��7Ӽ�IS)��ZѢ�o�����'Ry����<.��xAV
 +����Ej�I��J$��{�m�<ft�ȓ ��d����jj�G��2�$ą�3f��
?a�
�A(ϳF�����}��I�dF�4��kãN�^�\��_f!��`&���Ҡ훂`�t �ȓ2���#�'1T�*� ƶ8uV���e�Ѝ��EL3�l��q��1@��)��Q��⃬]  �����V2X��ȓh�p���dѹd-d*���Ke�a�ȓI�DP�3/�80�µSԱ�ȓ[�\���Ə7p�u2$"C�>4
���i�&�T%ȸB� �W#G�(�zA��n�й6a�<İ�"��#�l��ȓ 
�Ir$	-\T0)��uBVm��`whYU�t� �P0�O��H��� =9�T�����t���L݀�ȓ]O> WI��&@�����Yӈ��ȓsc|��7)��1�ԽH��T+Xvņȓ�ҵ:�@ �R�%p!i����ȓN!�e�7 ��S�����	 �>Ub���}�<����?�4xƩS��`|��_<��"��J�|$�0�秕�[<$p�ȓu��I!�PI��[V�]�Jfh��ȓX1 ���0n�lD�����4U����~�FL�lS>�؝��*%I�`�ȓE���2��T ��)2Q�� j�`��e/bQiUa�<Ka�����H�Ly�ȓᎴ�)Y\Bn�Su!�Jc"|��?mX܈ ��s�KE#˒>]�H�ȓ�@����7.����f��	E�V���7U���C��")��m벩ӽGxx�ȓ0X`x�D�B>	�r,k������ȓ0�X�h�,|dR�@P�E'�$�� c���Q��h3��J ��Q&���}.��`�W�P嚕�d�ӛQ��E~2(Ɔ2�Q>�Q�����5J�H<��Є#(D���ј^8 ���a	20�Y�/����q@L�IqO�>�p�܍*+�q��-��A2�#3D�ڷN�5s<3�����Q�*}2���$0N���P
@�@�=��͈��_�x:����^�{LX	 �F�-������-d�e�6 Ñ�y�N�,��i�,��� ����O��q`ٜ����b�Hpd�����#�(�y&�vw`%�`�7z�.��!���~"�A�����=E�dB�=�rm�bJ��$IFl�
�y��Ѻf�pj�	�<T�������ēx�$		�9s�qk4�B"��L<j��Y�ȓh�9�'$�����9T����ވ�ȓ3�<�q��̇K���{���S�? V���C�l�\!����{K��7"O�l
�M3�,��#]!8���7"OȜp@h�=[lvp#P��,L�6�3�"OР3���/�`�q�.��5�v��"O"���Ӧe�ֹ:��X��M��"O�T�֯K�M�|�b�����з"OĠ2��2�Ȑ�6�]�Tc�$��"O�,H�����Kd�>V���"O��P��ˠf��S�ǕW_�Y�"O$�1��H�����ωs%(A�A"O8�c�ǛE&
���&�w/@`�5"O������9�� ��d޴e�z�+7"O�1�1�B�O>��C��s����"OvA�#�H�0&>�rE�D�.qJ"O�TKFD)uW)a`��9�Tl�"Ot=r��BV�ll��Cߗ$�<��"O���Q8n��1�r��l3a"Ol�+�0�v͘)�+s��M��"O���iAl4���I�y�V��&"O&��`W�]�$)*�Л1�(�!"O�@�V��'�p�Lޓ/�	2"O�=�ь�6nRh��R$n��lң"O��a��4Y1nu �OX�}� �ѱ"OP�I��*� i�����P5��"O�����l�h�7��K�i�"OXY���J�~Q��F%M7���"O�@���y�;����k<�a�"O ,[g��7��poY<w�I�g"O-���
v2������R1��I�"O�Hd�׶c:���Q�:��pF"O��;q(��LqJB�	�o�ЃF"O��z�یe����Ʊ�ޜ�A"O��Zp�74Z��3�'B�LY`�"Olh�!䛒-���0���k��ŢG"Ot���&7�,�X��P�2��H�4"O��r�������#E�xf�B�"Ox�kR�
�PF~UӠdU+'�Ԭ�c"OV8#	�  Pd��&V�]��s4"O,���+t�fPoL�6��pp""O$���$��y�	Ѵ� �nD
1"Opݩ�l�I
�)
�s�Z)�D"O\��JŇ�^��Rf�,q�h9q�"Op=��˂+ EP$)VdP�e0r"O8 ��w#l�ѳ$4t
X�#"OF`�� B�@�(����Ƿ+��%Q�'VX�C�(�ȟ��w���t �/��}= a�!4D�p�lƵj��3D�\�Ib<=zà7�Gn���Y�j֢|2d*޴q[�]Qs��lRZ=�A�<�� D�z�^yq��A4h"8(�N�-F����U�vx@��'�"}�'�V��`/�f`��į@�x�X݃
�'�4�bN�H?NL���q֤x��`ˣ-�"Q��cĥy��m Gm*,O")�"G@�1�t,AwnW�?ЊՑP�';��#�+��j��\�E�ٕ8��򧔕z}h$���dT�Z�ʑ(<���3.�TH�e��6IL��vM�P�6HJ��&��+$$��^u�h�|B��T��U�5]p4��L�<ɡ��&ѡ��]�u�BL�\�`!kӜ	����%]�.�<���O��r�C��?].�����q'�'$���ѭ<�DO /|����)P�n���#��P�O�ԊG��>\�
���->�<,){�lbtqҏ��/����剷 ��4В�^5"Up-Q���f/N�0"M�:Ty(S�̽#�xa�BT�b"������GU`񻀢U�R2�h��C/i��'�`��T�G?8W�X@��.{@�:�O�p��O���10AE��Y�1�#�P��'�
G�Q D��h!��(LS�}#ր�v(`��؍�t����g1�z��t%6�y��ʱ:<��F�F�zO
�(DM���PxB�M�? "�*�f
;ڒ�R��;}�	��i�Sg���c�H�C͌��w��z�(�5F�Y�'Y�p���>^���A�Ξ�����~�Zb�8~bNpӃ�R�,�T�r�/��c�R$�eg�+.�Q�S/�- F��ݰ>g-����ٔ��
~V���GU���<� ��,�]z¢?�
�a/U����'5i�|�ፘ�J��p���޹�ȓro�MQ�[��| a%��h	ȉ`W�ޗC���cA�P�5�f`�pl��PB��8�y7g�5��}Ӑ̟�u8�����Px�H�A0�{�A��P벍�C`=`�c�>q�h���+�*�Q����C5�3�� �xT���W�
5��QxB�N����	�N+���7�H'?cV��__�� N��C��ɨ J�	��I�Ɔ��ha������Yj���s��f�8�!h;+��'�K��p����H��l��<�ì`�,�g蘻��T�]�1��mڔ��p@�hPD�S�yR���U>!�%$t����ݾ=36��eR�]�8hg�Q�;v���c�#�S9>|���w�D���gЫPu�1@�9��Q�'ܚ�a'ńL�>���Ԅu	�I� �X'p^P���Ҋ}�Ta�YX��AB�EE�'��10B
��1���9����a� �	ӓPK�k�4��֮�A����C;�b�� �O~�����Jk�4���'�.���
�8w�<� bf�3?��z�yrF�>��J$�S
Y�B�K'.�!`L)��_>y{�l� �,�����.d�f4�T�3D�(�wkL�-�p@Q�Q�m$D$d2{��,�R��S�)���C@��|4$|��z��ɹ_�d�$�8f���+)D���G��}vx|K'L�7��|�F9|%�9�W��Ww�lH��ʆ�h��	l>޵8E�P�|�L�`T�	)����ѩ&�<����v�us��^���QʐMƎ��w��7VȘ��D�L��I�d�;Y*�P���ў�VdӱG|�0��.��H`�E��r�آ'Ͻc�B�ɱ^�@�F��.�L=]�����Z��4�?E�d�U�:� E�D����n������y"mG�Z~Ÿ��7(�p꟯�y� P< I[��@4B
�I j��ybI�=yBЩ��'�@�r�X �y��G�v��z�/��&佒�+�����hO���@Kt,ڊ<;�HR��|Jh���"O9�b�l`���O�"&a��D!\O2���R%T۞���El���O.8�%���#'��:�J7{�dX`��E�<��V�[��3�.SQެ���fYA�<!�j\�Gĩy2	Y.�)Qcj�P�<�FI�& � �1��%3�r�i�t�<yAi_��:��w"�pr��l�<��@^1i��A�늦��%�c�s�<9��FC��@9�K��wnI8�ʉv�<�@=c�YX#���=U�1@��^�<����1c��S&����p���r�<���$> ��[��dh�5
�,�P�<1�/��� ���N�QE֌!r�Kp�<c� M.Rp0gA��>H�e�m�x�<a�˜'S�@��I`!Hm�<IWBÃ%���*�Aً� �s��d�<��造0a��ä�M�L�)�G'_�<U�\��!K#b�=[��Q�<�'�ӼϺP��n�&�����Uj�<�S,�/*����'b�er�rgy�<��G�J{hm�5�R.^f$HҢ`�N�<�um�8{�
0'�ĶH�ɩ�VK�<�5�\�d�>*5�:3���Fl�K�<y�π6$�DY���;u�&����WE�<yD)N�G��ه�F�E�$l�|�<��I��u	��,��-y	�u�<��R�/ Ԓ@דc��hb��m�<i�E&e�8c��<��0VA�<���e@6��g
-FK<a ��	B�<��@
.V����`�(O�������e�<!֏ϿVp�8j�E*$p����Tb�<� (���E�9l�ȅh L� ([�"O�b���5|��&��h�S�"O���G�Q�vz�CD�ay��8�"O`I�"�!䠘��=l��7"O�:'#G�Pw�yZb�OP0�@"O"a��k���ɆςLHdQU"O:�	��Y�)�^�S	���y "O�̫��O8��a�jW?$�d2"O:�@�ܿ0���t�S0�ΰ��"O���a�(=�̼@�'^3`�2�c�"O:i�@Ur�r�"������"Oj�(���YZ1�v��'n�`��"O6M�u���O|2��&�8��"Ob�!MM��Bu��=����"O*̺s��+}^��
���</���� "O@IC�E�D�xv6�|11"O(�Hւɑs��Pӆe�u"O)�`&�ĵ�cJI"���i7"O&K&��+x
���\�4�fp�q"OYj�S�P���(�jƱyVa*�"O,�*Q��*|������[nEi2"OjW$<34x
� :Nr�d"O�l�eC�h��i�� �6��`"O2����T2�Ib�iD̔k�"O2]h���y*�J����� Y�"ON@�+
�1�B�R�Øz{����"O�	G��ba:�r�"�:4�h�@"Om�R	Y G��`���I��EiB"O|�*�L�-e2��â�mx�\�"O���*ĽZ=*�@ƃ�$'a�<��"O��@Qa��T���ՃDMn���'"O�Ej��]���0`�
1]H1ɷ"O41�a.�wz�3�MJh"�'� |�f��9t|zpjL�`�
�'�.�ѣ��Du�x����Z㔥y�'ш���.��N=���'^J4d��'�d�`�o�
I$��)غRt���'g�1󐅘���0�� &��'@�5�3�2ZŎ�;���++K�\��'�^��
$&3"�Q�-�� p���'[���0��	K��SF͚
����'GTE�p/N ��AfУ]P@�;�'o���G/����`�:T�ш�'���i_�\�I����WR|��'����H{jPˢ�M�E%�%x�'��%���5���
B�C�+,�@�'J|��XM$����J1p�,Ԣ�'e��gi�9��
f�lrd���'��	�"������9`�P�\�	�'ޜ p�圥!�����E3WLdL��'HTJ�'�2���� ��H�J��'�2�S6EK�"@T:�]�C'f��'�5`Q'S:W"�Y)B��<0�(2�'#��Y��nK�h���B=t�2�'�����<v���Ԁ˭�,Y#�'�h!�@��>>ou����L��0�'p��v�P�+����Bg0kw���'�85��U
ت�'U�h��5��'��)��h�5#�؈p��4l����'� C�$�[����u(M�Y�(�I�'�,��"AD����$S�W��e�
�'+
��k�~�X��jI�N6t	a
�'� y�O��Y���w�^�W�|�`�'���:�"6E�r��(F�LT3	��� ����Ok���c�� x����"Oz�� N�8(8�qfə�3DDdp�"OT88bNP%0�@p!�4X�2f"O\i�/ܺ9�P���q6�0S�"O|ɋ�(�h6N`���ޢw���˖"O�$10	�, Z�Ȳ\tNPA"O-Z�aW-%@���
*.h �c"O��` �ɹ-�b͚f,�f��9b"O��[�b��
Z�9qf��>�:���"OF!y&fПO�����Aѧ:�Y��"O����@�5*dc ��~p���"OD\8����K���FǇfv�C�"O��A���fk e˶�ҩ5\!B"O���ꗀZh�I���qa��7"O�pZ�dE~fE�(΄z`�(�"Ojt�׫ۙ�q27�V9m"!J�"O��uM�>�Y���4x"m�e"O$�;U#Q�~��Q�҃nk,�h!"O������v�i�撲3IP��#"O����R�0�h�G��b����"OfpA5�D2-<���+�'&��X�"O8yF�]@�$h�@*P�y���r"O�i��D��IS����j�"OT�96�(u�J%���ĽX�,�#q"O�E1�&�>1�>%���?[y����"O�ƙ
�@�0:�+�F�r��a�ȓH�h�ȂT`�B�.$!~Ą�xb$<�Ώ�w�d]�QA�������Q��)ই�5jy�Ň�zH��*~��� ��~X�T�RM_=L�m�ȓO���Q$W�rF�7MK�#E�Ň�I����w&��.Y��rb�8�����9Z@i��F�%����F�4ɺ���V���YǠȼKuFD������ą�e�I�#M:�m��DP�MZ�l�� �P���/����5��sID	����i���(�"ɛ�b��"�
���(��tHdA��5:��W�3Y8ن�^�j�����^h�����Y���(��;Y�A&�x(�3�W'�h�ȓLΜݨ�+�S�l�j��1]�����"0�5��\��r�(]�>�졆ȓt$����GM-@=Z�O���I�ȓ$@B��U�ȋ9z�N��+�!��B|�las��#_�x���M
ZI�ȓ#��	cN��ք�b �- ���ȓn��1��Ʃ
��
3BG&GK���ȓk�Υ�iF�񆸀M:/TPy��y��5 ֫cJ�X`�Y�@Q���ȓ�Eڑ��I��E�f�
�:)؇ȓ`����RQD`�N��>�ȓ�2$��FM�%n�XA냯
xq��mH�+7'
�*��pV�N H��a�ȓH� ��m�!4��7�
�İ�ȓV�ⵊ� "r��!S�����Hф�.,�l�K'�LȪ�H[:�!��[՚x8�f$7��B�Ȅ7��t�ȓt+^uF��2�|Ȫg�P06n����N�^4j��4�r�Y��}=��ȓ+�p��̐m�J��� �U�`}�ȓk�hY��&	&3�Z�;v�(��܆�K� Q�IGoE�M�#��~IF@�ȓF�y[��]7������Ï|_ �ȓ$�j�3׎^�x8f�C��]�;����S�? �!��I�N*�l�y�LpX�"O�D��F 2�F顂�9�vփj�<)CjO}n$�B�/��R%�(jgH�x�<���܅$�R��4��:Q8�(��	u�<A�
ۮ\=��zN�$�d�Р˂N�<��lǇ\�M�#��6/jlQ�p�<��|��@�	"�A �� t�<Ǎ�6A.�ђ&�j����q�<�c�H�l������
�T�,�Q�h�<Y�.Q��n]��k����4GVB�<���\2|\x抹{���Я
}�<-=���f�� #��q��� I��B䉮FnE!�c
mG��"GN��6�B�I�	��C��΂f䂝sS�In�B�I@x�۶� abi�U��:iB��@LU�� i���ʎ�ivC䉴P]���B�-(���X�"� ��B䉻|��M��@?-AziCp�H�G>�B�I�`����Q�Ϭ�ZͲD�F�&��B�	*l�P$qPB� 8��E�d�pC�I+ ́�2`��C�k(C�I
rIH�)TD��xy�d�%(1aPC��e�X,�$�M�А�e�R�>C�� ��9 Vm��I���sB"�#TC�I�����+Q�T����	vЄB�;b��-��S�)	�����V7w�B�I
Z�<�����p޾��K	�5��C�I,1�8�A�K�bj����F%uN�C䉨s��A�O�5����-'�B��R�S���I`�]���	V"Of���嗍s^h\�3AGc	șKS"O0 �(5��"�&[�k��Y�v"O�Z#%K��P5Qs�Y�=a�lIG"O ��Rd�0.J��r�C�HW��7"Oht�-�=s���(���xE�e3""Op}r�ٰ���@@��r]I"O"$���Er��yE�ʼ^�%K""O0�+rk΃x�i�'�Y�I�-�"O�(�f�TcH��hF�;D��i�"OBȺ3G��6B���֕���t"OZDz�dKT��6��c�J��R"O�� ��YY�Uh�	]՜��"O6���d<V	
uC��b���C"OH��K�6dD��g���z$R�"OL�c�N< H�L	��T��"O�T�A�7>�`��Q�[b�P�"O�}��퍚Nҝ���kd4D��"O���aL�%0�@A"
mv���"O�i:e�\�7Y��+B���:_���V"Ozuc�J5d�H��~���"O`�[��U +
�|���_<qx�٠6"OP C�^C
�l�!)J%����"O��pa�W�`��*����l�&�9�"O� ��,f3���'��uٔ4��"O�5�P�W4Z�@go��jT�� d"O8T��9,�*%Ir��^�P���"O�0 4 $Om m��Q�vLE"O
`�e��/E`I�� �eH��"O$l�ԎEn�@���xV
4D�8�#�q�EҤ.м$뜄ӂ 2D�TX�e�� ��P".�-\&1�ց-D�| �J ��귡�/sB��3�1D�,�B	�w>�� �M� ����m,D�\�TN� N|�
�*���/D�� �=��7��D+P�A*2qh�"O������Q8� ��C�r4@4"O�Dk��h�q	��	.G"O���X"]�D�x�a�$�#"O��[�韤%��]R�ڀiȉ#"Oh#�����%�τY�,��g"OtxEGq����� *}���� "O,Uȥ��,��J�!ʆE�"T0�"On���c��Jmk�Px�Fbr"O =�"DO�N���{6�S%E�p�Q�"O�Lbt�V�^)J��Bm4U��x4"O m�D�L�p5���p&^ ʐ�E"O����2H���F�~2Z� P"OJ�h7"]uɄ�9g(иi&"O,����#��EځÌ���Ȁ�>�D�F�V484�a�^U8�}����U���CM0&�(*2$�d���S5쑝=��"�'���ho��5¢"�f���yCQ���S�j�Mb.��}$$���o�6DH��ۖ�)�tlRV�BY�����0�ඬ�"��0��<�}�ЦQA�R$����pܐY���ay�$�Z��(�h��j�!�z�$&s\ ��'�ĽEy��i�[����'��x��D���� s�eEy2�OljP�e��f�h���ٚ'M�ݩ�℉w����9<����>��d�A,�%�0���)�5c͎l�ʤ؁ �&�.˓4:�㟌E��&X��ɷD�0��IAň��?��kP����Oɤ`4����Q�)����]�A[P$��a_:eRN��Uy����$�*�0|�"g B�P�O'�`���"�Zܓz1D�iٴ)sDI�����pJ(���A�X�9 �͢f� ���놴]d�'�*�����5%2�D2(Z'>��	S���Jc�	 h�Q��|j#mP�#+R}�q��2u
�kǋ�ퟠ1��)�'�6��GdW��H0p$ϮHN����O�O@�g�S:�(��\P�ҽk�5#��Jf�fE��<�����C���Q�p-s#D�O�fUS0�|2dHI���O?dH1���	��[���3Հ�r,O Ȋ��S(g" jBc�82&ey���h.�B �(OQ?�����D'l%!�!4l�A�ٙ�(O���I�|1@l@Qd��gF�r�n@���O�	���)�ĥP�)�z�W�_!�N�y��A�j]q�"�!zd�х�?,�����?*��"�1��C�ɡ7eP�7d�%B��#뇏j�C�I�L$\D�Èċ;��	�5��@�!�d�rR���4�
 풵�6a@�~Z!�DJ9fʺ0�a�%L��H�@��$�!��M�l�\LR�DS��LX)��R�!�� ���0��cd�I(��%�!�$L�dn�	���>j@L+��Z�R�!�ɈH�
�;�A�mQ`�@U�X�!��W,!�N�үS�$�9��j�!�DE;tؼ��
WG�T5�tK��y�!�d�]�r�z�(A�U�f�ժ�x!��Ó!ڼ�
�Ʌ�2%��$F�N!��1T$iu�Y�K� �3.ǆ['!�Dn#��0�΋5�B��a,��z!�d�0�ܰՋ��O��t�� �!��;�U�ש�%��y�&&�n�!��D�T�v���N8�B�u�!�D�+/B\l@�"����0A��F�!�DUtLP�d��[��\��iҢ�!��V/W��}�al�*$��ѹ��d�!�d_3t��6�_�z���9�E-=�!�D �H�Y�.�_o�|ȧ���!�dV�A]شiW�L�M=�yJˀu�!�$ۍ~�R`��A�f7�1x��G�cS!�� ��pT�Z�K�2�FmǗo�
�q�"O8d�F͞� ]¥pƫPx�"O��v��TSc+��o[�4��"O��rFųs�zdYK������"Ozx��H#�X�;u/��i��2C"O�T�����$���*A(��y�"OZ)��Q���5z��G�\��|�"Opđ���,�%��O7܉0"Ov��c���Vr֩�%o�'4��q�"O.8��/�*Qц�D�[�4E`�"O�ܪ���2>��$����?���("O<�8�b� 
��q	3���P6�H"O�=��߰v`J��@0V���U"O�سD�0R�x���H��h��"O^�Z4JB�Lh�7�M�@��P�d"OP���b���t3ee��Q"O$�tH�m��kƣ[#�����"O�u �LH74ڜ�
@c��S�����"Orp"�R	;!J����-[���"�"O���`N�i����&�\-CN�0R�"O ��ǔo�\,CwOPXG�	K�"O�m�
p�F\��D f.\��$"OB�de��B+��X��[�7(���"O8��p̃�`�t�rٳ2��#"O�A�eN'�H�SĐ#N��D��"O�@���]>4�ޅs���<S��"�"O. �pkN�{Ǯt�Tb��!<�ٶ"O�1tN��\bd�q ���"O�%���7oLeZ'��	'��8�w"ON��͈�5�XCR�@�4��L�A"O��إ�9r�R-���""O��RɜD!N��Q�8��(T"O<����2wJɢ���71Dt�"O���e�4�(�a�,�_�$Jv"O:���CY#j!������\��w"O� ���X+jp:Tc�̒$9T��CE"O���'�K �@ 
��B����W"O64Kb��%��,��A�R��Y�q"Ox�[���}߀�E$@	0���y "O��-HBM�d�W���SvP0"O~]�4�K�Utd�f�
�a���g"O	C���<@�ءA��wM̩�E"O
��Bθ<=@ 'a��~�ѣ"O>������� �c�@R����"OP����A�8��N�?����"O��k�6~��4t��A��"O���1a6�0�saI?7��	�1"O��� �V?�y��OUa�&�`�"O}P��H#<�15O+?��y�"O��2 J�F$��")��)Q�"OH�� ��G��;b-��� rr"O�%F��vY�1�Fm_�P�.���"O�;7�C;5ݮ�P�6<�t��"OX�+�iM$/�E�R��)$����"O���r={>"�"���:+��u"O���A�,��x4�:$h"O.��F�L�.��Y�OH�j���V"O���<"�@�@35�:�C�"O�X�v�j,ȉgBD=)�"]"O`�����|:J�I@�ʢeup�3�"Od� �䈺�蕃���\tR�Z�"O�1po��Hl��\_~(X�'DRZ�<�W K"!Gr-B�k��j�`LPZ�<��+F%��<H�#A�'ذ�!f@W�<� ��s�� �;��!k�"O�|�$�_w3�X��4`y��r�"O��@� @�t)dE#%vN�#�"Oxt�ӥQ�nMĵ���SU���"O��S���)e7�XpA'
LR�p�"Ob����R�T#*�qE�3	��"OJI���ԼP� ��2#Ul����"O �� k��s�N���Bʑ���8�"O�違�^�Yd�a8� �Y{漸�"O��% ?8��S�O�+i�|H�"O�cc@,�@�fdE;Cgt0�S"O��zq��^��`��GI
��"O8ik��_�N2�U� Dˍ	D�|��"O��# �qf:��Q�U �6�%"Oe�fF4p�qB��l,��sg"Ob� 5�F�e��P���·c 4��"Ol92b�t��ysT�ڈy%��xV"O�� f����1�!�	L�T1u"O���@�Siȱ��Ά�Va�"O�5�$�ըY��p� /2~ $��"O�-K�eO h#e��}�j`�U"Op�z�*�G�؛���O�Υ��"OD��@�5*�����Ɣ	d�D�f"O�-��횀M�<����A���ڳ"O��X��ׇ~g��&��8g�\�B"Oʁ�a@ޔ>� ś�*{!��Ўi�!��]D��V(I9i�^E*Cc�5O�!��:w� ����g�HX#�$@�	�!�˾QE<�����Mm tK.�!�ԂtlnA�riX�i�="��]�4�!��B
x��4(�́��u��Һ�!�$�S,��&��$�Q"!��6s!��3|X��7���t���C.'O!��j����DGc�	+!�K��!��ܖD���K�aI&Q��m�V�/4w!�dJI5x��5)�#��#��{k!�,e�\�С��-^ f���# 9;h!���� ��R7;��-s&���!���q+F�c��E�~e�ظ��y��|��H�hIS�JJ�>t6	`$����"OteP�eQe�D�G)R���:���D8�\�d�]1zK�j�c؊`S� =D�Yr�z���@E!�>z0�a��y�8C�� ��ĺ/Пr�%h+ː V�C�%הe�1kV�|>Ұ��)K0�`C�	%sx���C��#4�0�Gc	W��B�I�t�<c�Tdע���E�a�B䉒B�V�S��5.$� 0��P5��B�I0�*��+SX��R��0H�C�	�RH~�*� G�����O	���ȓe�fEBFI�r�Ƶ!PlT�K�\l���@�[�<�F��P	�<�����$�U�p�<g��`1�H�A7J��ȓW����拥g�0'��%Z��ȓlH�1+�cP���m��nК
����Zy����A]Ε���[;����>v��ȝ�s�<�kC�"���ȓ`�VM��b�j�X31��q6̄ȓn��YY)��E]��㐥S<nz �ȓM�0��QH�6qk4�ͺqd����3h���V=���Z�G̭xL`$�ȓj������_ht�2cA�+M�	�ȓX��P�	�4s,�����M
	��g$�,г�H�%���$S5N���S�? z�1��r렅B��=	����!"O���V��Ȝe��JM�_�b�x0"Or,"�܏�B�#A�a>aR�"On�i�ߒ�1k�IT*d~���W"O�1)2HI�A�|�*b�r�1�g"O�jTB�jJ�L�1�αl�1ʗ"O��R
L�V� =JQcR�R�`x��"Ovr�-X�M� �q�Aݼt���k�"O�$��H�+Ǹ��v��"���15"O(�rn�E��T�֊/~����"ONA��@>r��hsBi]�@���"O��s�EJ��dH�ƂL��9��"O���2`�\s�9h厰R���z�"O��ՠ�:���f���:$"O��X���k��@U��\�=P�"O
�A��1W�Wc	"�6��u"O�ĺ$�^#RĪ�W,f&� 
U"O� Y�
$;�8-pF��E����"O�Q9�@��"�ds1DJ�E2,���"Oj؇�V0��]���m!pM�"O�|���� ������e)�#�y�K�&K���RVė9O8zQb�ޚ�y��_,���)�'ְA�p�d.�1�y������I`L :ozbu�ɮ�yRܥ�]��C�db��J��yBh"2�l�9�j�+	��8�e]��y�(��B�P��'�!O|������y��,5B�8��DX'A�fF��y�BD�q���a�*�0%1!��
�y���0L���A�z���3�!�=�y"��E(���ϓ
c�e��̕��y�@�%8�lkG���x�NIP��yr�W����c�r=zI"�W�y�`�,� yI�h��<���\��y"�ք
�N�_.y�!O˨�y� R�����!ΐg2��tᗛ�yB�YT�HCu,ݺad �C�A'�y�j*[@��y��ԄD>0��L��y"ʌ&f4"�ԃt��I@� D��yҥ۲Kުy��i�s�Ddه.K��yr��S��L�X�lɰ[��^��y�� �9Tfщ0Q�3�"t�ݑ�y��+��p;7��17�����(�y�	[6��I�����(��f =ј'.b�� ��Eo�����o�D��@�с੐����h�b�C[p9b$�'�B�'8��Y'Ú>V^du�C)���P,��ěs/��7����9v�Ъj�8����W:D{��č:�^X���V�p�x9���Ǐ>�����끅���J@	<w:�
�C�bH�6��n�P�m���M����$S?����[قMY���\)q����'c�O���pp��V�Dܠ���2U�B�;�i3\OV|n:�M�O�A�a�ŮJy�
�U=�@�f^�NQ8��4�?����?ͧ[��h���?���MKT�Ä{l�JfƢB��iiJs��L�&�B�@��c7�m��@��Lm�S�?A��4�a`&�s)L�;�${`�L����Q�@1��Y����F�4�`�)�$,�S�y�Jհd�S��6:��}�J]�[�����O��'�j�2�����3sk׆>z�(!m��!�F�Ђ�G+3�b�'�T�'Y�,{���R6�%�5a�=<IhR�{B}�|<nQ�����4x�*	�p"�g�&\B�Ȗ"oO�|�g�'~j$��gչ���'���'�6��������s���AClР��;o����M #7���$υ*�f7���*[�<��˻x�LXȋ"�E��v���M	���;�ϒ}Ѵ�R���|i��P	O��u�c�1���Z7K�dѓ�|��A�F���k�n�7�޽���MS�W\.u��h$�x����%�<����%�����E�T�K�Ǹ� �I֟��XX��Zq��@u@�����mL
03T���e���|��g�T�)�<I)ء36�&�i��P�1�]>���v`D!I3$���O��$�O�)����O��$�O��5�ԨJ���Dj�$.X]�,�<L˜�������r�%Y���t��LGhQ�P1�F��N ��#��8v�)�Rb"�m��6ˋ���qd�ԸK^���\�V"<a���쟠"۴�d� ����II*":�
��ޯ=&qx��>q���?��Қ�ĭ�318��Q$��K�x�h��<��'a{�-]7Gd~����֔P$��֦ف1�f9o4�M��K��vL C��7��O��$�O����( ��! b�$Hp.��C�9��\C	�OV���OV%��n��|��Ɖ<~2QD��0�i�/z��9'	=��+��?p@4m&���<s������0*��ҩY�#*�`Q��..�D@�<��l���u4x�	?��'úh"�C��#1�'G���%G=g�>4Sa�r��,��?��4f�z7�A>L�]0���N~���	�����4:����'+.�RQ��W@��I�Y ��%������>����?���vK����?���M��	�)ڑ�0H6[E�,ڲ��3��*4>��҃�ݨbuD��SM9=��-�O��D��UAMz�<d��97Wp���O]�fg$ٴ��(tGbL�p�&��ًVA@M��r	λM��AB�mT7Gh���Cˈ�������'0@7Q������,z�>� ,*�&dۄiS�M��`	��
R�'�Ob"?A�&Z�L�z�ꒀ$�J���+iܓ.��Cv�ڒO �)�� 6흕�����b	d)���B�����>��� 
  ��   e  4       �+  f7  O?  �I  (U  j[  �a  h  ]n  �t  �z  &�  i�  ��  �  2�  ��  צ  �  Z�  ��  �  -�  ��  �  8�  ��  �  X�  ��  ��  � B	 �  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�rdFz�Q�`�'�@o�	�*�)�D���	�%��	�OP���,�2��AK�}fԠ�2�Sp1O)l��y�S�`l
)��S��fE �6�����B|*����;�	�D����&�!3��ѐ���c�� Y�~�b��}��?a�bW�W����q嚱xNCb/�Mx��A�Zy�X��A90��
P�T� H���4 ��ԥ�4H��`y� �+	B0�*G#*�D-�S�'q
:-�b�� @٥�'Wǂ1�ȓc�8�y0�n�&���@,t�^��vC��Ezʟ��'�(���,�B�qE�|���'�`��R��D �uN�i/�51�M*}b�>%>y�<��( :l.��1p��
T��CR(^�'���OZ��ڂl+�Y�͟�xd��a�?oI!�T*D,�=�.����� �Py"�)��m�f {� �!�\�t.<�y�I�$�b���ҧqED�X����d9�O0|�1�_����c�>n�����'��Iv��/|��  �ۃ/��d�@:X��B�I#c��Q;�½��2G.ԫ
��OZ�=yʜq���6���惕{¤����B+/;�	o��,&`��t�d�9��(5$���!�O�I��y21ORc?��Oô�i�O^�L(*Q�M�J��9�U�'8�d�[��M���ׂ |`�	p��<0�!���k��\�#i�/o
��v�ٰEr!�ę���4�����8AX'�eQ��E{*���r�m��F)��I���R��	C��'�ɧ� ��h��~�
 ��	M�Z��LkET�̅�	I���X�I�~�ր���8y2����8?�Íe6�@���j��yq*T�h0�@��EPN8�J�9%��<r�e(�F����'(
8 ҏH����@Ќ]�$�Х��	O�':�5��!:w\��ҕ�I�<!gB�<]xT�v%�
�\}��WF��$���"J m,B"-�V	�q-!D�Hh�d�J<U�uh�� ��:�J;�Or�q�" ?�1���G)Y�¥�ꉳ�BB�I�Ly���&U��T���ƀ5�t�D+�|�ў�)���؝�b����S�O5\Opb�PQʗ��\!h�{s6pd(���F{��	�-_z�śv���L���s�1��|b�xb藟qMCfO°wk:h㓣N3�yO�>.~��V�y�|���!Z��yb�+ �
rTh�p�p�S�9�y��H�Fp8�(��k=6������yBH�]�X#�Æ]EfD�`����yB*H�`D��ᓋ�*km�8�V���'�k:�)�)%N����A
q�İ�v�.s��Oʢ=�~J�J\G��yb�>Vr�P���s�<��AY�oBTA�a� І�Z�����hO?�	&��!�$Ɯ:& �iU�B�	.H���q5 ͡M��8sY7w;�C�Ɏ�J��4�Զ;X�AWꗚ�NC�%�
HgL<D�ipP@�-%NC�I.Nb졂ӡ��;���q�
יByC�I/^�L�p�_�	
�y�!`FC�Inڠ�:E�7.X��mqm�?���I�.�b��C��j�^���i(~|!�$ß{���˒&�2��Erԡ��-���^��H�����]�v������zB(�"O�x�֠�/~B���%�1�:Y��|�'ffD�&�z ���C<O�T�Q	��y�N��M�F��H�����)�#�y���FN:d�5%حv��@� ��Oj�~����0,8���61�:i�"��`�<�%������
5b�����SE�<�W*_4h0Ɯc�C�\�pHQ7�]@�<�ԃI*<��#3��E3�5��M|�<	��[ J]0��@	J!&�~�<ّ`_�`t&A�2�[AdLC�	C�<��D�FBJ���
b��\j�!])�?q#Ĩ�bT�O���d��lj S�
�z�2�+�7w���' D�܁�'&�Z����AΌ��KYE�'��aڷ哠D��r�/�Y�����!	�2�&��d5?y'�M^8��%JR8QhIp$�G�h�D���K�mE�� !���X��F�F�w!�D��l|x�� }��d��/R2e!�������"I��\�s��TW�R9Oδ�G�	�Z\��GܼR�p�iv"O�dAӈ�#)`����_)J�b�C��Is>��K<�m��BX0"��|�a�(D���Z8'N��H&ŀ�A
b�zT����x��]+ϼ(@Щ�� ꞡ�����y��J�)������:q��u�N��y�R�6X��p�Jo`��+�8�?y�O���]y*��b>�yEgP�mt"-�J�� ��E��H(<��4X��@kD^��#Qi�}Zq�O��	r���'�l�S�Y7�(�mح\>�\�瓐�b7��h��H�> j�!$BOȾ��$&Nqxí�N:$��.�=/@�ȓz��	�#4-��b�S�R>���S�? 4h��j��"�r��0"��!�'�IC�S�O�d�a� G�Q��R5�fǦ��"OH,�b�O3�D�@e�D-�`�2�>	�tD}���˦}5�m3a�ѥX :]���?q%�̆#���X�O�3�9j�b}�<�ǨĲ�r(j�I�?��0QaGx�'i����i���S���-�̘�f��<]򄙳&Vg�����΀5� b���Bb�9YS���J>a|r�|rI�=>lʱ��/u��Y1l�=�xR�'`��4O�Q�潫�@��@0� �����ȟ�mS�^�.��ć�4���O�)��ʆ�$Ԕѻf�W�>Hj�QpE�ܟ���2���`�� -�R�*Fc��GČ%����ē�(��Y�M�='�|��J&NH�f"O�i��e_24 �"Q���`k�04��D=}�1O��?�cJ�;IҰt��L=�<h�ڟ4���+�|h��g� �r�r�JU<��l���1��'�*ub��B/(����d
��C-�,�˓�(Oh�C&bsD0����x�|!T�$d !,O���yʟ,�'��a�EoD)2�
��L�(�dߓ�'(�P��P�8�0OĆSH]���'"<O����O� ��
�HP��*0��'��w�i�V��'`��>O����g?٥�C�:!H )�.��"�m��U�<�"��й�񨞂p���r���P}��)ҧN��[�E�lde��̇+[�L)��#P,�U�6�b����c�@%�4����%�qG�<��,�����i�`B�I�N8�)8�\�G������;8B�IOa6=�B-֧D![��Lx���=Y�{��x�-�C��xp��T�J�������M3�'O����Ӷ{eT��cM�
�4��'�T3P� :�B�/Ɲz��'�zuH �E(f� �;�0`�'sʉE�$4��:7 �,4ڽ��'�^�C�(�"DbT��l̲L�^,��'΄)zäT-m"h4�%�!?P`��'6��VA�<b,~D���"m��a�'�1[�*��GN�a�X��H�'0(�����4h���H�' Q�
�'�h%�r�]�,cl����rɒ։�d�<i����q�P����9O!RLh��Fb�<�F*�';�^	8` +�N1�E.�c�<��f���(c�.'B�4�ӣ��\�<�`�A=��HS/��Yx���&V\�<�1 T!�����jǈ~�lx�7`MN�<���=t�d���|/�ɂ���c�<�qȋ�m`�5S��&w�v*d(x�<�Ch ��R-���$n����b��x�<��B�:�*��,נ*��q��w�<QO�9"g�<����>�(g'Hu�<9�'�[�D�	S��cd]��IOq�<ٰ��4�kU�Q.�ʤ�w�<����,z �&&�i"f���*�v�<A�EӦ>�Bv!�Y�6�S��v�<�d�G�i֬�Z�J,ql�qK�[�<��m��^�@q+.yܢE9��V�<�GcO�"�~���4d�Й[�QR�<I��ϵ(�d\0���2r[d\���y�<����Z�j�
P0L-��"wDq�<𦑒
ʁb�FG�K1�Q���c�<i�L����	�(|���9w�S�<���-~�2`��Jp�4��E�<���&1�<R��$5z��B!�D�<���2Tqy%�^H�����j~�<� ��'�ε$�b�Gs~���"Oz-���L�]�"�Z�;v�3b"O�8`����0�"L{�bخqpP��"O������TKI2f4XZ�"O�hC�M�3 ��b�ɀ�c��&�'��P���Iٟ��џ��	���=M,ʓ�8[,C� �I��I���I����ǟ�I��T�	۟\�	�ǾI�d�Y`�<��"�� ���������	ޟ����h��������.<xs*�&�A8�a�7u�����I��������I��������I�0D�t8�J��S����P��`�	����ٟ���џP�������ߟ0�ɋJ���4���9Z�ͪ3�:��	ȟ�	����џ��	����۟P�I�Q*@p�UnR'�Fi���N�;����ß �	�$��۟��؟��	ܟ�	���=�r��(T0�e+���J�j,��ß��I����	���	����Iݟ<��)�h�h��K\|�0��B�������͟��Iɟ,������П���"o�"4J��"������!^4u��������l��ȟ\��ӟ�I˟��	/�qA�õrD4:�ҳ]M�)�Iٟ$��ԟ�����X������̟���!{�m�hT�|$��0�K;n����Ɵ�	���	<�Iӟ��	͟����;�v�
�m#�s��(�d����������\�	������4�?��b�V!����VP��� 2Z��#^�\��Cy���O��m�Cv���&��X�\ P��L�n�1Dn<}�i���'���/�9r잴Q�g�4 R}���Pi��7-�O4�R� ̪O����'���xR-�V��^X.��j����5@�Z����<I���7ڧqn����g��J����N��9r$Y�&�i��#�y"�����* {U	��3����&�j��
��M��'3�)�I,r�l]C7O|}����+OH*�ؐK�;-�8��0O��r�X��l�KO*��|���a�� b���f��$�5N���ϓ��6�d����s�m)�		�&%!僕m"���`��-%��Dx�\�������̓����:���;u��^^1�+�/�	�5l4p7�-(�c>aAW��,	���I�/����ƚ���1gĖ�sW&�'s����"~�yL���C�o�4�#�.��Γ7p��N"��ᦹEx��E��Q���Ym�0��7d�<_�Lp���?9ܴ�?�"ċw����'��쩷n�$����fح�D����]�k_h|IY�zjў�`y����6|��x�BXfv��6J̎������C8�J��P4��JB�K�=��Բ�Hc�z�[���	�Mϓ�ħ���.��@*q.V�ML�9��]�6�"�[��:"��'�2����7W�z)�f�$Hy~�"�M ⼰4�O�h�ҒU)R�8�'(�'x�6�Y�l��B/.�*(;��H�K6>�� �<���iӎ"<Q.O��D~�
�D��
�0t��N�]2 �剽K�@��%��m��ǿRQ��;R蛻	�8dI�O?����)B_c ┣ǈ� t��P4�Qؔ�*�'��]�d�����8zq��(Z��c흁1砅a���Ҧ��c?}�i��'�)S0oH>mK`�z�+S�dv����?O���M�r�i���E,d̒�'v���to��ZT��$g<���M�U�1�����W5��rF�x���{y��'�$�R4�6.�L���l˝����'�'�
6���1O�'�|��Ȣy��F���S �i�Odʓ�?�4�y����O�X��O[V���f������k��Jn����������Ĳ��9$$�O��׮��D#(�qW@�n	�U���OR�d�O2�D�O�	��0E��]��zٴ<��Jp�C���#�"��!����(��<Y��?�����4�ʓ<���C�~E��Dy�`{G���7m�)p�dW��$�����!=FNqJ��gy�kVO���j�x��U`g,K���'�r\��G�ĨD
j��ֶ��vh��l[����+m�|��E��b>]mz޽r�ML�{�=S� Y �Ez�A«�?!�4�y"T��	����� M� 4��>O�Mj!I؂v 0Y I�1?n���1O�-�၊��\k�;���<ͧ�?��f�nS ��Elr�!Z�b���O��d�O�Y���IV9�y��'=��q2� G!?�<�P��¬sh�'��Y��ݴW���O*�1X��r/�&f"8���#� &����?Y%�W4P��� ��3������"��v����?b�����6.�(�R5���?�˓���O?�I�*o�d���� ��A�"��r��牫�M�`�u�z�^#<�ӗK6:@H#�;S�͋��BdF�	ڦ���4�?�%̘�n�l���?��4���2�@�,��� E�$-(@���ܤ��4�B˓��'V��	��\�G	S�%J���!?�ֺi�(:�y��)��L¤ʥѫ�H�S"
"<�'���iD�)�	����a�Dy*��o,��H�˰Er�8FE�\�ɑa[0��,��)��E{��O�{tx`��LQf�jL��KgRW�d�'�'��6͑�U��\�T\���R�,�R�L��
��Db�#<�,ON�Dp�����I�dy��-�,^��$��:UĹ�nI'��ON�)%e�J�li	������3�5� �="��Զ*��9[&
�ZfQ�2OL��O��d�Oh���OD�?�ڑN��O����N�Q��	F��y�'R�}����7O2���O��OT3QI\�v9x8wːo˔�@�f�l�'&x6��Ʀ��ӊW��` pNi��mڛC��:���>��%�W�V�?."�¶�+��LY2�hO>�į<Y��/��.�2!R���!Y���*3/��<IO>��io&u��yB�O^���t���A��/Ř�"˟����`y��'1��<O�d�)�,�*����+m�(p�A��' E����}��JW��\��66�2h��DE�2Qr��I�HRIf��7j,�'�2Q�b>�~���J����{s$�;J͞�a �g���H�(m���l�<y.O6��4�.�r0�,KlJi2(V�}��EnǟP�F+5A�����d`�P;[�r�� g0?&i"Q��:w��nD����Bi̓�?�*O^�}b�@S�`f2I������r�f�;mE�����'���I}��צ��q@i� {l�Dӱ�W�6�pi�	ڦ͓���O����'a�����S��y�N��\"*�w���YJ�ZŨ5�y��x�� �%ĦU�ў����v�ۻT�|���4N78�v���'��'��6�LU1O�Q6���czn��T�٘r}m��'/���d�OD7m{�p�'���R�@_�L`�Q-P��V0��'� ��F*Xq���/���⟜L��_
Fb���	d�ظ��N�JKu�{q��$�O2��O&�$�O��������4L��rs��a�n�K�\�Z����?���i�Œ�'fr�xӦ�O�9��If�.id�!i E^)8���
�:O�0n��Me�iOBLR�N��y��'�LASĈ�-|M��j�E��0`���( Ϯ,1d��W��'����Iџ�	˟ �ɭ�$`�pc�xo���q�C�:�N�'�z7M���O���?�9O8h����/b"����퀵(�Ձ���gy�)g�NM1��n�8q&>Q��?�C�Dս���1����j�6�,A���J�5����0a�*)�&�;J>9-Of	sB&�J�����W���1eŢ��D�O��dV+jtfo�jyr,{�fH��8�$qX���y�f���G�W�s��O1oM�i>�@�O��l���M[��i\�z%�83X�c~�1MV�C�j�@F���y"�'�d�JE�Q"}V�I3�W�l��5F�1�j�↨E<7�*���R�y��'���'���'�R�)٠N�� ���U�)M�9p�k�.|�I��O�����1��w�����M{L>i0�7$���jW&�5vfB]1đ
��]�0��4[v���O0�y�v�L�yb�' f�GF�9�.� С��Y�f��݊�p@�h vў���ay��'�l�!��T!L{ϖ0xQ���'��'g�7���r1O�ʧ``�{�	��yJ^Q �������O���?	�4�yҜ���O'Z�w�
�"]ˤ���D�"8�!�՜s��5���9��$���["`ѤkdV�O��f�D�Hۆ�AeE��v�BTI�O��$�O��d�O1�&�'"�F�	���ReU���H� Ӄ>,���'���'ɧ�\�0��4�2�E&��n����3~�u�i��6�/o0��:OD��ҙ� ��r���sW�$���hc ԝ,�6Pb󏁕b;H�Γ��$�O"���Ov���Or��|R� �.f��x����c^Њ��A��OV"M��'9��O��d�'"�i���1��4B@�Χou�\�f#@(�4n�M���'��i>���?���g�PZ��	Qj�2r�+\�\�Hb�PBh�%#��q�n��&!l|%��'^��'�<Dbq��I�a��H��ϤY�4�'hB�'�"X�x�4z�A��?y�MZ�c�cֲ(`j�c���d�>Y��ig�7�C�D�'N)�WBɁ���ʴ(�+z��O.�pk /k �횑�,��'pU��
���O�z�n
"�
�"rrEr̘�D�O6�$�OP���O��}
��\���1�-_�O욄��nõa�Hh�����v�݇�y��',�7"�4������q��B��brLE�m�����Rٴ(���M��E��p��'��C�t�"�[EËvlb�ڗ���
�͘gf��d�(e�w��� �'g�Oƨ�� �f�tis��>]��@�O��o��Ojpc����@�Q<΍`t��x.�-�P�F(��џ�l��<yL|���?�u/����4Y!���&%�榙#"t�hkl~B�M�DuH𐓈X*ў8 ul
>B`�Xp�Er�-�g'�ß�'<�C��M����<�C,
+7XqHW�G���a���I?��4�O,ʓ�?iٴ�?��\u[ذ��	�y�����E0m�p�蓅M�<��
j���@w_���'�$a�AR�Нdgdɹ��+/"�$�7$u����\y�T�"~JGb1Pf @fL�,\l��C�^k̓7�ք�����Ц�%�P�W��s���Z1 �����CdR�<)/O6�ߦ��	��1K1����Ƀ|��`+���#M����+
H\�@�?���(��Sn�A\2">If+Ըgu��y3f�AN��wgZ�<6�á ��h�`P	:�p��#f��`!>"  �"����6pp$�Vc�'���S�*�6�B�A�t	n�"cd�9'��%�%◷F2=�֣G*�I�aMTd^���g��YQ���c�#�|��䚡jZ�]0T�L���BT�|�:�B.�����(FܕA��Q=)_h��(��P����٦��I���	�?u+3�V8G���;b&��g���1�a��ē�?��0ц,����?�����#c�֑��Z9.a�4)�4�l������)-�����4?������S7��� ���G=~�%��)�+��� ��i9��'s&I �'�b�'��v|�F �>4�`����^P����_ɦE�����Mk���?������x��'��u��I�h'��H��=]B�$Bd����O����O ��~���?��DV=RH0��DF0}�P����R��F�'���'�����e<�d�O������Bl�z�*yXD��� `��@%�lӺ�d�O��$�72���O��iʜ=�Li �oB�� �a�͈�.�� �n��b�dl�&��@h<�b�,�RE��KN�6�lPbiHK�� ���:�xRr�^	E���#"8.M����^�Q
�z��]�$�q'K�EO��yd���M�e�� 2:e�d97�U�}RB�;w�P�~��@��8�,�a�v�H�����#��g*�6J0W��,	C�¹��dц��h�R��O@���dң�mR��P\(X�D f�:- ��'BrJ�M��'
2E��u�,I��΀B���iCF}����ǧ�8h�ʰ2#b߱*m	�̒Ʀ�R�1ʓ`��	XTA *U4��������C�#Ղ]��IC��G�����o�!�M�#�e�'�|Q���?��i��o۲�"���Ā���13h[�K��ҟ@�Iɟ�F�/�F�,@ڧ.N%�n��b T>�xR�zӮ@2U�E-_���R6ni�
5j2��o�]y���+N�7-�O��Į|"E��?���Ͽ!� �� ʓ�Mp�H�����?���1���
t�r�y�$·8��P�S޷wj�dA.����5�<p����a�De�Vd��>AS�,��-PvB+6��a�H�+:nH�RJ<�N @V5�COA�\ 6b�T���&$��NdӜ�oZ����J`�T�L8���7�	� �X���h��?Yϓ'�ؕb%P��8� N�<,(��ɯ�HO���Oξ .R1��"x�Ъc������Iȟ��I�PX9sD/^ޟ��͟������1�+\Rڠ� eN;Kf�;DJ �R��⃀��?������ы�L>чΒH���
��[��ވ1�� m�����Iз)���QΔ�}&�p����	�H|����Z0�E2iK���Y4�U�)�3�DS7�1�g�/:�}�0�Ǯ{Y!�]��p�W�8J":��pN@3&M�ɩ�HO�#�$12���@�B��G��0��H�]�n #���#V!��d�O~���O�����?q���?�Ѩ�"t��ܪ���n�DXւ��&W�I�w�M>]���J�RJx��!c�B�\Fy2��8i��)&"�&�.y���O�=K�Sx�+B�ҝ������ `DyB` J�4�p-�\��A�����r�Cԛ�D{ӊ���<����$�<Q@���n� `V� '�d��F�R�<�"=8�v����ToF�Q�R���t��lӮ˓}��,6�i���'K��j@�&h�.�9D�%30�sq�'d�M��'W���>Q'l��Bb�<��Q�H���mɟp�j����ɷhM�@Y�ьKd>�I�n;ʓb�RE襭�-\(r�X֫\xd��ó.8$V~p�A���$=r`A�L����Q
�#
�.��O@���'Y�@!�ԵL4)Y�@�"g��ʰ�`�H��ן��?E�$&L�QXR��0��?u��M��x��s��|A�2H���S�8�i��g�Oʓ �,\H��iq��'��Ӕ����ɒc(Xe�5d�9'yJѡ�A��v���I���A�p:�(�t���sj�9�S��^>u�@K2F�@�D��Jzr�+}��h�)��������I��a�q�g�[d�����	?�"�4����M#��i�����9d�,qL�4������l-1O��d8<OX����W}��2�hP�Sʨ�'��#=�Ӏ����	�v
�;M��p���8�X����?��S�����Kǖ�?����?���7�N�(�$`:�?R�g��Z��D#	���ⲹi���s�
{1�*!zV)�y�_�s@E�� ��D�����7 q�2��L��K��ܺU1h� %Sc�ӠBʊtY�4��$�#��E�|Hb�"^+]T� ����O`���O��EE�Oq��ܟ�q�����{��~����AG�gq��D���<1E��`����v͕�B��ɐ�HO\�)�OPʓM� ��qdCQ���
u�J�t�b!��7Bz��h��?1��?Aa��B���O�瓖,�PQ�Cl�½��S`�paU$t5�d�U�� 	q��hVaC>'���;��.s/2jRE0c~!�v�֪ b���� ����K�1��ݺb�ٚ/�Hp�N��(OХ��cZwd��p��پ9@Uj�S�Y^��h��,o�̟D�'����Z�#@P����/ʸ�*R��<	!�I�;`�z�ׄx�� k�� %�1O��l�$�'K$\��f�|�$�O�lJ�I$��B�* ��yrM�O���I5�4���O�擄�TTs��9�DDq��T �"�R ��-�wbI�2�H8�2�3ơ)s���x-�t�ľ"����1�V )F��[G�]N`4��oȎ]��`!t��B�2!X�Ƀ7 h�HN�Ƀc���qOȱ��m�!kΜd�&C�	2v��jf �4���#��̍Ny0C�ɍ�M;�l�^�QR� D5�.�AI#��F625iQ�i�"�'��ӱj���ɌV����BFYL̝7�����I��p���p-��q�	Ē`�������k"MA�TG��ȁ�Z�	.�>w�JA�d���:M���X�AĴ/Թ�ě�
 uC����}���:4��.UKm걋�I�z�'��,j���?AJ~�L~� ��q5F͸)�N�4��Q��!����O��D݄-�N�r��'cP���&ax�%7ғ;��0Z%d� 3�ȅ�VΙ�\�|Hs�i�B�'�	���Tt�']"�'��w$vX���d��+��X4NND�hP�ʍ'��@5l��ꕎ��--J��1O�e�r/��X<�pf�d�@(S�/�X)�G�U���(�)��"&q���b'T���tK�=�$;pڳ�Z���ϟ�X�4�?I& [��?�}�'&I[�T�#'햾\�L��fӋ��{"�|2C_�rڒ�saA@ZW�J�.��$�Ϧ��4���|�����Ĕ�~1`� I�f��D`%��v�d��@�,=�6�$�Ot�d�O\�;�?�����E�Acf��˄z�dɲ�b	6v(�0�'$��d@7-�h����F� 2'��x�7@��3g�J��= ����������?A��E�AYf�1�͇w�B1��Ar�<YP�١0k�thv�V�W}�M*�)Lt�(��O)1d���9�	ӟ҃(��~�^�"`�3Z�H��Ў��H�	�f�����']��aZ���*i��l���O��h�㑃��D�w�É]ux�4�'I��ҕ8A6���aܬ[\�tц�$G&�BR(�g/�@��4T�
���q�')�c�E.�'�f�B!ʓt�(�0g����Ţ�'U�)��
\��`e��MΣ�nP
�'�x6M)4]����N'2q���
�N1OXq�lIϦ����O�L�''�U�r�ԡ8>�ċ�LP�wj�u���'��"��>���T>�u�]�anY18��XE�:k���O��H��)�8\4�@qg��"X*8x��`=_1��'�\p����ɧ�Ox8T3V�N�jܬ�s�(p���[�'�<a���%,X�@ԆZ.,|��
c����=VHL�S�Œ&�p2�7D��(fC��d�.u���L*~� 1"D��J���q?�I##.D-^)� �#D�P����c����d�)X�@#"D�t���ޚy�^yK'�.��=�E)-D���Ǉ:R�=�F����)+D�h�����\��Yhh��0���h_<!��ψp��(�ę5W������e�!򄌚*d�S�"4D�T�!���5�!��/%;*MCE&�nxP��p�!��O�F� YK��D�)�p�k���Z�!��6�ʒk�=X��J�n�a!��P���HiB�(��u�'�?	�!��2~�PQ���P��������f�!���m����+�D���_<Y!�[��P�@ˇ�,:��- �!�5pbj5Yw��\	~����F�!���q:ŧ_�E�*cC��$8�!�_�u5��H�܉7�p	4��r�!��Ωs����jK1_����T!�{�!�䌋�>�Ãj

���h��E2�!򄃂 ��p�vk�@oN-��E�*]�!�sC�	�̙QZبq %A�m!�D@���9��:Bz�X�c��!�d�S�~���E'2�����f�!��QB���eU�'H-�Si���!��Y�?�Raӄm�6&�K��B�!��C�^���梗�����M(v�!���F�<� )�![W$yQ"+�3)�!�$ &����DQ� CP}`QC!�!��C�nճ��g����Ä�H!�ė�w�@Qr�U�ijz�Y�L-!�DS0[�ȳ��YH�x����^�@D!�DD$qFiއ:����1C!�:zצ�)o��2 =���)4!���4@�MrS�Ɋ�Yåm��Q��3��� j�LpW�٪UqX��e�<���K*x��ǆ�K�D]1!*Io�'��YP�cȔ��]H"�zJ�CK�i1�N��`�3�!aV�0� �6Snꕓ$&{3�|n*C������f0�5����v�0�G+ݬ7��>�|��l�43ޕ᳎	�6���<� B���Ӛ0�z5
��E� }�-1K�!�܇�kVGԚ\�ԑ�b�̅E��|�b��&�D�ˉ�D9hf�]Zp5��hctӄj I@�_�|Pt8y��'��iap�Q1�:�	��^'"��Q.�
��$:FiŃ"��t���Ĕ�1�,?)��͋E��͚Ԋ�	��E1�-VI�'���2cBr�&M�̈́���5x�
��G�>1���W	Q��h�Kٲ!���zp��z�|�q�[�V;�,V�'.�R �F<<P,��W����Erh��=q�@&��<��O�}&4Wo�T�(A�a��e��	>��F8RDҒ�3QT���%��]��a�+Umy�2M5�	ނ��ԭ����L�!V�1�'�Za� J�!e��hO��%4ڗKW
��Hp��2pw����#v�|j�'��T�r���B�%`�%�'#VH��G�l~�DY����{/T\S��D�O��ӥ��~�V��d��+UWT�Z%I���q�`�T<El@�bG�)�A��'L&H�aT��o����c ON��L�,:�	2DC�+˜�B&�'It7MWAijpm�H$��ó�dXFy�	��?4X�ӥؠ��0ՆQ�z��ϓҘ'��0C�� �E	J,�)$q�TFtkZ��A�'@�|��J��y�=*�m�n׎�r��c�9��'Z��jl�fǮ��	�dZc��}K�) �?B�LK�&1))�%ȰΔ+^{��V�?����'���a J�VP����i��8�'���Sr�'�:7�B�UԼ��ܴOcv�I�ϕ-w,��%L	sJD|@�,�z�H�p���P�2�L�'TO�=���o�xxr�N�{VI�'U�@�}�������
)|���M�/�7�ى;z�Gy�X*r�d�B�G�E�2����Ta�� ϓ�~�S���uI�Ks�@�� �����7��t�0/{PQ��;ea��;���Y+��HH�@�xT�e��$�<����W�$���#�䅲�N��jʨI�"�1�	�	�c!��	a#�
U<�S��U2K��QL�����M�"�|�.��2w��I^���O��D��<�K��d���D���`6M���0�{Q��H5T�����CQ��t ØWكPK�=m\.m3�*O�Ų���?]^�5�AK��~�n8��'97͛�F�hH��'�-c� �a����Dy�nI��h�3G�gH�YԊůjh�U���~�꧟�l��8Z��b�ܥAa�0��E��QM�h���U�o�Q�\��ߔ�nZ�6Xu;$�_�^`��˙ �2�p��j`�堟��O����5W�y+c�[.x�V (�,Q)�$H'5m��R΄�pf�T)?�u.��*`
i�� �Iz�Ey�n�C���?q�s��а�Q�c��(�&7K���<(���F2P�lQ�*Y�MxZ���œ2Y�l%��a+�ـ�E]�0(��~�dH�q�Af����wk�O\�D�$]��bR�Y?7�1*��1>UQ���.B.Up�ŋ�ժ`#h C�	A	m"��%�I>��Q��[�����M���1�g0�Jܲ���.H �Ґ����Q�G]�n�Zi��+� E�ؐ��*�	s��|��z*��y���$�
	�t-�=�`�Z�ÆI�'kp�2������J�;����O�\�#ǈ;n���)�Õ�W�9�G�E̓�B	m��s�%�tex���49N��ݥ|�b�%c.{rf �Ek�~�n��C%��6�#o�4���c��8{����'�H�.��s�PTG�S�6i���tk�	�=�tl0��<t	��(J���7j@*{�X] d�pȧOj�=%?qP��7Ɋ8b����}.4U	w�A�|ᕤ��Q����JC�0���M���h��L�Rl���Mԅ�ڢ<i����u�Lb�c̞J���DD���9��5�G<b����׸}�<X���K�V��'v�l�s!��s-�C��.~!2��e�=�~���9�J�np��*Ӝ�5����5����*]�g�����a'{���UI�.��z"�H�:��q�c�<�3�Ʉ�	��\�q7"0����gc �3a�܊���"Ğ��4i֙"B��GyB.�o�ʘ���c0)a ��|dB��rV�<�A)}����R��X��1o|`x �:W���#��� �X���ɫ.�aEA�g���eO�N<���H�1��`�Ox	F��O���f�K�\\�'�))U>�K�"O�ݫ�O5,�90p���G;H}�P�i��ৎUG�.����@��EȖ�-d���lُ!�����r�,�5Lӕ�yb`�Bj�kS�Gi6�Ͳ���s�<IQ�)��񇥏�z�&A��[�	ƥ��.U����}�V �� �z���P K��qr*A|�<�IƐ! PQ�둓ow�jD�d;
5��	�H��I Cp�@�e!P3�n��W�@�wĶC�	,P����ٴ���"S̙�o�t7MG"=�0<���O���=�Uj.�ab�c�R�E���l؞L8F�H�z@��'�l�x�Ć���{�%�N��$��'Z�� QLD"8ҘP����?і���}�_�%��ic�TQ�π �h C�m��K��/�V��"O^�[v��#��a�l
lk\�Yv�U�%'X�5�?}��"�g}��'s2@I����Z�\��R����(Oh8��3�@H����|\��VV�����k/2ɪ�㗤aM��+fMk���'�p�]y�AF5_?$i�N+��qnZ.�BU��4yw��	d�~�`'D%!\A�sOI� ��C��'O��ڄ��=�X��÷v����R�Pa�fL0O_ڨ�+%)6`�sG4ʓ]{��õA �!����獧1Z��۱�Y<�����c�.�`G#5М�82ږ[9r�@p#?��ױaP��&�e���~�P��#S����d
Bv �RGA�$�4�p"�@\ؤ%3��($�C6���N�Nh8�LN�l8�H�'��L�B�,$����P��`ٌ��1R0��0�&ߧ�@��mu�y�`�f<j���~  �q�I�'I� P�egփF�(�R:����
>)i�Ye'[>ZV��p�4k剽,��i[a�Ӆ'�Э��GZ�"VB�<����G�2;eAԺ)ƹx�^�+�^����Q��S�Dx�%9�E�tM> �M_u	@��C�!�3�\eH��м;�	�%L��쎯IB�xD�UK�OH�'#D)��Z�ۀ��4��CG�D�O����i�j��"<WE�;,�%���~|L���D~"[�@�ȹ�ta�Z2ѱ'�̘22�6-)7ۮ6�ƣ�~R�O�p���$�?�gG��� ņK�6nG�'!؀@�+��Rm���Q)cv�z�(D;qzD�|�8d{�q�'� &!A#N�!0�RA�J�� �5��"A*��	>Qq��SC�'V�t	`-�+&/��@�3tm�ir`�X���G�Z���Ē�N�?arq�����ɗC�SE���U�W�|��5A�<�Q�;Q��
����-1D����M7j��4LAi��G\�(�Xt�OR�F��B�m�Dl01���F<��B��9?��(�h&Y���dj�x}a���2�� �'��*p�ىL&޹R"!G�=�X�Cݴ~E.5:���+w
�O�]hp.��nI˕n�VzPH�ӧ؃3t)3OϬٶ�R��^��&<:�I��rs��X�e�ȟ���b2�$�1�X�Hw�ʹ�?	7,F_�,�b�-7�*\٧�wyr����h)�tm��*\����G�(OpM�����!,�h�DG??ڑ��)��'J��"�)�Y�|"��n4z��݄m ^h` ��Y��:7�V�h�L��&ƨO�����3��nJ�r�"Q`b���n�Q�&#'3�&�)!#���'&<M�QF.��	�g��,up�xp�r��T��/�Ov���D?j6���
7\dj����P�$"�'n~�藬�5J�>����O"Hp��ߚ^���O"Ir��Ϻ	�]�@�ӏa8P� *�!?{��� gl`M)A��Kk��OM�N�v��ƴRD<����-��I�x!ueU��?9��&w����AǞ4�LCqyR�'�@y�h@MExB���=�(O�ų$�V0m�6��Vc$>��m@��N��'<J�ڂ���V��G�D�Ɉ	�-A􋞅(w3��ҩ$4���TI�2?�XF}rO�3m,�H�weޱ���ϔjNr!�k�5� �CU�;+8~L��P���Az�T�YN�$M�7,,�pөL�N��+ fD�o漩W$,wu����C�*����SHܨ����':2��Ŕ�W�@�c���o��$/�2�����wPj@�e�������:���Z-�?Q����:T�`)VL��۲
�p���	/1�PL�jմ޺,��סi���גxR�c��9�#�ڟf�(r��8��L� �k`��O� ����c���@�'v� �O*Q�����#�JM�.H�W��qB5#��@K�OZ��nN(��D�$OG�i�FU��f �T"bi�s��'rt���`D�-��G}"*��{'��z�w�dB+Џ-��Ri���xT�A6��G��^�®D[D�^���(S�::����� 7Ҡ]����	N<�ēU�R4�t�(p{bk	��}�aV���'�- �$���.��,"�,�5"��kgyՈ6~X�ڃ�@3X� ������`��}(5�� (����`�m�z�l��'Y���ď�1q�
�)�P9"m�M�,OĬ(��: e���3�C�-�0�e�I5�����Y��|@�S��Sgi>���x�<�G��N٠�ܡV�� dGN�pAƗ�qn�����=*e�D~r��+r>�ͻv�.�9��ȴwZ��g�*r����'��l�?E����� |���-��q��,A�xȉp�	/y�n ���I�Z���I(p��#dଚR�]�H� a�-��w���'=2��|�bZ�6�2 ��E�(��q�9x+z�0bl9-<a�Lֳ��I����*cF&���-Ad<9� ��o�ax���T�s`cǧobܛ �5��đ�]F��ugPW8�&n�;DQ����*@>TF|�5d�� ���q�;-��ɐu�B})��Q�i�m��KL6'�X[�&ķ"��y�@Ȅ�5�D>p%*�sA
Вf0x���ܬKAK�
7p���ߊTP�0�ȓ��h(@�$p�\0IƊuz"I��p����Q�Y�Nq�5XՆ��G�P�ȓ#:p@��aM�U�����E	A�
̄�ev�{����c�\�8'C�#bR��ȓ$�
�k���Bi�Ё�=S� e��S�? ��k�#0�uC�A�1>�<�"O��d�Krz�-�s�}�t�3"O�٩���+$�*����B����"O��t�ë=�4y;��ԝ2A��"O��!�n(��!��$0 ��"O�����V���U��P`��y��Ʀ*L�L���W�P}s�$��y�͟"mwY�@�&}@8Aq�JS��yB������O�!'vE�e*N��yr\�B��K ����`�$8r�'��!`�.^!%ܱ12��3k�~@�
�'B��D+U ���☎6�\�C�'���@����j��ѣa��D�A�'�hy12���Pe�c��atS�'�@@�H�3v��R�-s���0�' ����΄���!�BT0li�j�'��%�/Bh���b�Sj�x�'1>ܒf�@�q��R�Y� ��'��Q"�<�,�1�ΐ~�2$��'j$���
"�)� +"��uq�'z" ���FzMc�A�*Di�I�':�$7D/9n��f^?;���J�'f�*f�*l)��#�gכH���'� %���'D��XUE�^,`�'�j$��'��H��M�4�U�r�Y�'�P��LI4z
���aˆU�0l�'� `��d��]�N}�ӥ�;�����'_�	kQCH�&&���7�� �����'H (�+]�E��U��B�0;r��	�'�,�bצ[S�BM	F�ڵ"'J�'4��00�{����V�="��R
�'/�̛C�G6ߢ�1��&H,��'��}�R�ؤ@lZ�A����']Z����C�ia`aH֫LV%��'�d���N����{w��:Lm��'�н��%Y�q�����:wǤ�'��2b�kGZ`��+i���0	�'�2��ăE	!��B6!Z9��I`	�'�x���� �&-�*T�7���:	�'-��Ӭ	8|8�0E 3O��q�'�9*��:�6 ���Ǎ.�(���'|�{c���H�d$�"D��
�'D<i�6A��+ap��G¶^��
�'f��ƃ�1�Ũ�O]$	$�b
�'���	�ߖ��]��U8�< 	
�'t�r�lA4hY��� ���I��'�B�@�B6���g
��'�H��5�&��"�"hV����'��!w�_�76�
�bŊ[��r�'��m�ԯFRB^�)�CT��:�J�'%pA���D�zu�I�%�([�'���B\�0A´ ��)|��
�'>��(&�ן#����H$�N(	�'dNh@dNѢ'T��Ґ#��q�'?��*� &c }�0�fR8�
�'���ᏉN����G�[�.���'1J�r ŗ�^��l	�O���',�u� W�}�� c��r����'�N��f�,\��q@"�Ey� R�'#���JD�ٲu+���nN
���'<��3��;�(u
�c޼i�Z4�'�	b��S#Q� ���c�����'�%ad�_�}ݼ��k�8a}�D��'b��C�/%<�"J�$'������ �����p���j��<�U��"O�M�1&��J���#ri�9$N���"O6����6�\xb��o"�Pw"O``�-Ԃl�i��F_�J�;0"O�ѺG@�]y��(�IP����"O�<����t�p�t�ѽ?��P�"Ol�B+Q�L	�A��Q��"O(}���3tސ�u!�=�p��"O�Bv�	,�Yh�O	%4�ěs"O�e³����Q[�.;��2�'��O$ԛă��%Ȭ1'@�r��Ek#"O��E�-am�	H�l@A\T��"O��E�D�M#pmZ;*���"ONcFl_�3,ġ;2
��z(H+�"O�T�W��Ii>��/�c	$��&�'��*>�)I�M�)h�)@��r��ȓb�
���j&�"wh�M���ȓH<����
+�6	Г�Io��m��X�=�!$-+;��K0^�Ld<���m��5I�!�34����y-�Ɇ�J}Qh7,51�r1*̍C ���1�P��wr���Y�OC"���C�<!��־b�9!��&W+~·�]~�<)&�F��)���V R,�E �LQa�<i�IΪ�"�7���#�ppÔIP^�<餈ֺ|��
נrp[�l���5��ϸ�����,ȷ�jȬ�@��� ���8����ġ>�5c�('rd�gD�H��`�g�y�<9���~0�Mb�煆N�>P
�nt�<!�bƖHk�h�揜~nT"R͖r�<	%�������=�����F�<���Y-	02y��\�e�tt!h�<�w���W�6u�3��#t�M!uM�b�<Q�#Noj���L�1�j�e�]W�<��N^�*Z5��U�R�ub�B��%�"��a`8cVR	:�
�+~��B�I�&Kv͹�	�7!$-�7M��*M�B�_�l@��GS����8��B�I�B�4�GD��r����IPs�B䉭`*��bǭ��V\�|31��MP����e��Ӱ�_�.h$�k�$��@Q3��&D��p-�m�4`� �%�8���%D�P�$� �̱a��\?KF���s�0D�lS��H�2Zm�@c>9-�l9��.D�X�Dc�0l���҇�&A �<��i/D���g��.6X0�eˍ]�Z�1�1D�,z�%�u/$�9ƃ
X� ])�B;D���/R(�f��@'a�!�S�9D��A�W�����C��kS�� $�OJ�'�5�PiT'"�8�)�
F��"�'�>YYv�M�v	>y��'^�9+�|��'�ĘJ��}�Ph��N�#�\�'Lh$,��HQ�%�JT�R�'���r%\=1v�Q���%@�pU �'�$��E)y(�,!�!��2���'�MR� �dV�9�T卌r��\C�'��� Κ=Z*���П4�� ��'���"`A�}���$ND:&Z]2�'ސ�Eo���p�gcY5vht0!�'@�⤇��3-���	n�����'��}�r�H�� \CDJ�Nt��'/���!@בk ��G�ȷE��T��'rL��g�H�75$"w�S�)q���O �=E�d���="�"q��k�pM��E_(�y
� ��s�o;9n9�����9����"O�9��z��h�F]I�.�(�"O�D���O�� 4�ѣ	
H#�tZ�"OZxxЊX����"�#�.~�`��"O�PAB��TbP�Ԉ�7!h��&"O�� G	�7�P����2��P�E"O 隤�
z��#��6ob���"O<} &k��t�#HfD�x"O �+��K>\2Ľْ�]���U�t�'�O��z�)�N�y�(	.$�p��"O ��'v�x�P�\g���*��-�S��yB�	7!�A��17��i f�B$�yҍ�X�4!�a��c$A@���=�y�	���C���6aR �I�'�y򢌌Bάxs��o���P��ybJѷ �&@;톡��ӆg\��y��b���!�Iª&��q�u�E!�y�Eͨc���틦(�]���ͅ�y���"[��G��@�P�g*�y2��Q7j��A�����p΅��hO|��	�t�Q�ɒ71�U�T/:�!�D��9`�)�[�1v�`E�B�d!��^���L�⇕�jf((�K��!�$L<�Z�b��R8�PWk���!�dJ >�����E�x�(�� �h�!�dW�2�l9(`e���@��k�!�ۊ/��Ś��ǂP�vɻB�ۉ�!�dD#r�~!��_�`�zp+�!�E\��,Ac�^�5�d*�*��nT!�G)����m�3?����?U�!�d�
�:�C���X�P�DQ�t�!��P�"Zd�B�4�L�J�a��Q�!��Ny�d{@�O�p�I� 
:��� ����c�  Ȁ�ӈ���'
az��#%#�@��"�抝�2�Ё�y��«h�
���(��F��G�"�yR����r 
T�ű �"�q)��y2GY�T����W�����a�!�?�'��}�O�~�
�!�!�9�"����*�yBf[.i��H���SiVd����+�yoO�����M*6��LZ�$��yM,$��|��ʄ|�D���EϮ�y���*4�� �r!I$sg���ꊮ�y�@�tp���//rV���dm �y�(�0Zw��E��m��A���y��-�Tm�E�L�_�ޭ�ԥ���yR2)B�ȘgN�"iĨ��֐�yR-  ,�%���l��J�y�_?5�@�tk�"t���b�!�yR�ĉLt�J��_ vV�Yg�8�y"��΄��C��i�hs%%��yR�P��	���ã`bĈv�yrH�Ly��Q)Ʊ\m
HJ�FL�y2)8/`����FL�U7�`%��yҢR;%�$Y�⌵EMڡHBM���yr'S+.�^9�c��:s��4���y�A�tkh�Q4b�9t�̙���y� �V`t�Cu`�����S�K��yBD�,_@���S����Flı�y���9�}q�胾(�L��bLÄ�y�D�
s<��]$��]iRO��y�E.sN S���"��0��#��y�^�p��j <v8{! B��y"�/s\X�W�X f��ER��y
� X� e��**�⋾r�� �'"Ov�Qg�	��(0����9���J�"OV0���l+����K=6����U"OA�
�^!z��9E��`8�"O|�#�X�2 �8`T�إa�0�6"O 	��&��]��� BI�
�(8F"O�`�ҋ��m}(�J�����z5�D"Or�s���'l��2e\�,�ڦ"O��G�{A�A
�,t%['"O&�!� ��$��i̥��3�"O�y���<��b��Ý+�$4�"O�yPu�F� q���C3z�<���"O��[DF�\x�"H}�8Dʂ"O��HeE��+���b��� &�Aآ"O��1���n1z`o�#@	~p�"O�A�bCP�*!X�A�M�A�N�z1"O���� 4$"52�&^*@8�ӂ"O�s�Ô�f��5ɗI�{�e�!"O0���o683A��16��y�"O�\��h0)#�͇bA^m��"OT��p@<2eг@�4*�8`"O�<�DI:�X�B� 9p��i�"O����Oπ%���T��<i��8�"OEyfJ�e��4����-mT�}{�"OdZp��,�V%�Bo
����"O�=�gdF�k�4(��OU%:�,p"OtLs�* �Ld�AJ��f�\��"OZԹ ĵ [�)��(�Isg"Op5�τ�͠	�$�K<V�X�k�"O$���k�?nXH��뉤)�މH�"O@���lHo��+'��?�te�e*Oj}��i��M�v��&I>Z(�'k�H��!	�S	���
̺6`�U
�'��0��@����ԏ,�n�Z�'��@��/��9�����.2+l��'�V�*�$�*<��HSt�V&����'�6-3O�-�Y��K1�P!Y�'Ξ9�M�#=:(��BǕr~�,��'�R h�´xf�ђ���e��|�
�'�U�G��4+U�)IR�A�\Iճ�'�$�pK[� Ҽ0�Ҧ�/Xl���'��Hj� 
�0�27�L�U^����'��|��D��M����L�\�B�'���U0i���V��$Ii���'k&����r��y+��� lH���'���g�X	Z�ްK0HS$e�Y��'�p����pi3�b�{¹��'=01���(tL��B����k�'o��8wi��BM!�!J=
]"t`�'R�`BqFѼ@��E�lR9�� �'.�#��F�~X4T+���21A� Q�'b`� #�q87oŁ,����'� e�C,ޕM�)��**����
�'�P�j��bW�U㴯�,x�A
�'4��Cv��!�,�t�bA#�'�`���HͧU�~����A�d# \��'!�����O�)�nQ�Dl��Za8�b�'IhQcǒ�\34�YM`H�''r�C�*b�T�2n��Tr:��
�']p%�ƿIJ�=��m��w:y8
�'��]���Q�+������ȇc�`���'�,Ȩ���&��a�W�]�6��':�0��X(�����MۻK4�}x�'2�h�LJ��z��F#X�8���  DCg�@�0��5�GX��E g"O"h�D��\� �� lضw���"Oư�p�[�:����K^4kb���"OޙY4\�qoz)p҉��Xj��"O��X��͝/2����%�� �t"O�Ђ陼D!ظI��4M<��"O����Ĕ:{����&��4��\K"O�i2&СWæ	�.B�m>�)��"O ,#î��jv��{�B͎'
r���"OH	%h�:1���Z!]4�<�j�"ON�Jf�
Z�6A��F�C��w"OJ��e�c�L9 s�_�D��Q�U"O\���3��rQ��1y1@"Ob�wjH�Z����N�\I���*OV\�2�I(��{��PL��	�'��	�DA%%=�(�F �;� l��'�p3�cW;(�J|��Y.@����'�PT� #�* ���A�$���`	�'� 1�㌊w�� ������	�'=B�0%E�<],b� �C�;����'38\��NR<�.L3$�fD^��'Ҟ9�D ��u�e��c�m��'_i���I�d�8��R�ʤ^ඍ��'���z�Γ��*	2���]%j$
�'Ϯ�K�KS�~�d����ҝT�.���'�^�$J�qp]�$��G����'0���)	�N��%�smW8
h�'zp��m<#F��S֧C��:�'ܪ���bϤ@S��"�I�8��`#
�'LBTxW%ɰa�@�rR C
@|:�p
�'�Bbem��Y��"�"�@U��I�'�0�2M <�bŀN�D���'��{�&\�G��)��b�1�P=�	�'sD���iJ�XsDkδ7t=�	�'S)r�@̂``t��8���'�͡�I�)T�q��(�)|����'�v��u��H}�CK�"mQPZ�'���فf�;A��@Jd�x��8�
�')J��ƌ,� 1:r�G�A��'�ZV ��1p�U�I��ի��ߐ�yRH@VN��A�P�6(Uy�+�y�ώ�RL���@�a��Ń����yR��<�~5�q��(8���e��y��
h��z��,p���oS��y�bX�Zd��O�y�t�qį�y"g2$/�B��#d�6�ȠH�2�yr�$q���1-Z�n�����9�yM&vc�ȅ� �c�!#u*��y"��c4��BR'�f?����y"(�rv��g��^�Lq�ϯ�y�^�o�@��d�D�J ,S����y��֍A_:`�bd�Wڸ�P�I�9�y��@�S����rg��x� \��G[��yr�B!^3J���ejC<�2����y�-@:p�4u�E̗OHj�����y��ΝH��8���ρD�����y2�A ���@O��@�
��y�j�n��"�&6�j�x&��y2i�'
`����#B-��*͌�y���RC�ǯ2b�`�ץ�v'�A��v�f0��Q&T��3j�.5n�ȓC��I�v�i����cF��ƅ�ȓk�J�i��Q�/� �ec	�"p*���|T��+��P&~�D��L.q�̆�S�? ���𡏥^�pI)�@��t�W"Or���J�P��q���%my�Y��"OSRoW�7���@�	`����"On����n�Kҍ9�.ċ�IY��y�"�$ ���h��#?"�1rဝ�y2S�qw0�U��*�r1`T3�y�Po �d��cĂ9�f�h��Z��yk� ~`Qӷj���(��7n�7�y��+I���(J� �`'-��y"B�����$�0y˰��6e��yR��}$
���ۭs��\Ж&�yR�K:<�BQ86��j��!�vm��y�I��}��a�WƓ':����y�G �|ds�H��
����k��y��:1���� T4�����yB�T)ʴd�%�wڠ�2l� �y#�/
" ����}��,q'c�/�y�Q`$�j �D s�$TZ��_-�y�OP:� ���Ԛ`�%��`ً�y�����E8�(]�8�s����y�"V�.>�cB�@�t�I����y��6VH��R!U�w@t];Q	ۋ�y"��r��L��k&w��-��j��y.}D�(i�\�ؖ�I!�y�ŌR{`��6�ИP>bqB���3�yR�C-PN�irsE*@���j��J��y�P�A�йZ3k9g(�f�V��y�C�yD�	����9z�� ۘ�y�̅� m���㒆m��Đ��U��yfV�Y�<��C]�|�7!�y��U���"E��U&��@�I&�yB	̪o$�r�ާ}���iֈ���yU���ܲ@�~�f��K�>�y�F@�:�<m�"N�JC�E?�yr	�a�|,H$�;Q�"k��y�'T�EX��(��D6T ����ԏ�yW�����5���q!C$�y�@�<��E�E2R��h��y��E�, �1�����@STDkVgD��yr*N�)��yG@�9�U�&aW=�y��#a�$iؔa��0t�4��[��y��=F0Q�D-H5P�0I&���y��Ӻ�X��t�+�\�"�� ��y"-Ў6QЙ� ��x�x�Μ��y�FnJ`��l
 v:����>�y��J	e� �AӅ�}�
pJ�!��y�,T��-[V�$�x	���yb,C ��iN4)kb���y��.]AM��KU%��mBWf;�y�D��W�������d�� �����y���;B
"3���0a;����'�yҬ�%� 0���@a������S
�y� ��	���y�� �pՖ����y��ƁGj���ϔ5�e�a��yb+C�Ƞ��d�?�x���J[��y��[-K*�T��Ύ	��Z��à�y"l��k`dJE�L���9�͊$�y2�͢oX4�u�Yofp�#a�#�y'�o�0e� �aN�x5����y"� ������D�T�����%ӈ�yr��I���'Gr^I�J���y��kƴ�r�ƅ5������y�k�5jI+u���4�4���HG�y�D .Y,����%���U	��y
� ����D8�C�E�d��0�G"ONP`���_e�\P�cS�#S@	zd"ON���]�H[Z�x��ܘqb�0ˇ"O����}12�4X�(�x��"O0�s��ϋ^J�ʵƛll�Y�w"O$b�{�E�SG��	X�@c"O��k �8p*��Y�f�	o�8��"O
��ɕ�k�Ÿ�R 5➑�"O�;�\�l�ZQw���uҰd��"O�L�х�'��]��G�6Z�b�+"O�ͱ"� =i86�"�U>z0`��"O��bv��<&8�h��Ӣ`-�a�f"O������U45k��3�I�T"O��&KۀH���!^�PWhL;�"O�tRW��) !@:%��-u\�]q�"Ofh; ɛ6]���q��� I&0�"Oʅ;dA�k2zl�É��Y)^��"O*��W�Y�N���0D�S���K�"O8�	fMS<˖��u� �L�<���"O4,c�,*]�b8H��(@L���"OF`4�P6_�v�{Î2/��Y�"OZ})"�U��( 
E�
T�� F"OP�2K�2Q�ܻG/P;�JD��"O���[�j�P�@1vH�ɰ��ô�yR�4A��xآ�R!g�@�3e��yb�)2n0]Ð�R:t�(�E�I��y����K���� Z�qO�pxeF���y�� ;+��Ȃ!N�aո��D
��y�h��'[��AV�$)���1芌�y�H��
r�D,�/+���@B��y�M�� ke�=��ؒQ&���y�ʓ�oz���	�p���eW��yR�GsCN��wG[ü��2�B'�y���?l�i	S���٤�����yN�
��a���Yު��7�y�-Q����G����Z���y�JY���̺�	��M[4採�y�E@�l�tiB��]%3�p2�(C��yRŇ�-��K�mD|9B�f��y�+�T�$���L�yϾ���aǎ�y�-���ba�u�ʄ#iİ�yf�� cA�u`B8$�r!�4�H��y�i\)Z@��ÀX��������y�
�~)�f����Y��X��y�ƠWITE{i�6�X$G2�y�ȓWDl�&��B���� ��y����#���`�D�O�p��Y��y�oܡ� �+�L��N"|��� ��yb�X@	���@G"?U��bJ�yB.-`I`�F�[�9�zHc�a�=�y"�Ɍhq�`�/-s���Go@�y���:L����'�Ш!������y"��I�}���V8Ghܿ�y�l�(j�0�l�� �P5o_��yBD��9��DB� Ӡ��!�̋�yR�ȄJkj�P0�
rI�j6C���y���;��t�ceX8\ר,�U�4�y�菽#G�EYA�� ��j�)M	�y2"T�$8('�CJ dx#B��yR�DRm6}���U�h��qiǈGH�<�d́3c����ϙ�\#�U6�LN�<��ǜ:����O"��C�J�N�<�р��E'~��i��W���k�J�<9&o�7\xs� '*4*HSK�<� XP�@N+1��	Dm��u,^�
"O6�ypƝ�+�z܂�nԋ(����"O�dX���	R���y/�F�"d�B"O�������$���^�f�
�E"O��94�ҷIҀ0��-�D�@ȳ"O���G�ë��%��-�k�L��"O�QŊQ�N�zij^��eOJ�a!��-r���Y/ *����6LP�E!�u~*D�D6m�%`�̛�R�!�D�5nΜ�s�L*LkZ���
$�!��4+�H`q�L�2^YR��!��u[!�D�9Gc~0f�1*�� �hA�t�!�D�>XNˏku.A����!�dΈ?��p$�C� ^�����Y�.!�dڟJ!K�"�-B[~}��%��!�UT6zF��adF�=XC���"O� �7���|_<,�Ţ�=>B�qZ�"Oґ�&�����Q��z�B�"O
����^U��<;e ),mz4�g"O�x���L�aH(��/L�\�-{r"O<8:�M�2�*�aů�]���j�"OIs�T�uk��k���I�a�C"O���'Q m~}0��O�!<9�c"O�00㯞&w�z�̏�s<@x�"OJ�kDN�$X��U#æؘj�A�a"Onl�iD�!�d��GI-F����"O�}K��A�I-*��6�Jik�]Q�"Ox�9��Ӏ���S".Ѥw�Lq�"O�yy�K#� B�>I��j�Ck!�����L�W��|��i�/�%W!��@P��9�
�>���b�g�G;!�D�}�Jy�a����A�y�!��7>�xI�%	�J�Ph��E:%�!�VmV�qR�רQ�pi�3e��~�!�D��o����l�!+���k�K7\�!�F8!�>� ��ΆT�a�("�!򄍵7����c��&1��#7�!�ă�
�`��ԻD⵺ԩ�;g�!�D�>�4�hT��=v���Aj���!�03ݚ4�s/�'�,@Sv�C� _!�$	#W����B��,�v �i�I�!��;0�P���
T��!���$n�!�O�=��D��j.��d@�3g�!�d��_H��� �y�q�� }�!�J9�]y��|w֘р�\Y�!��Z
L%p��//vT�I�B�9Y!�䇘]����自TB)�޵4�!�$��*\d8G$�&��� �p!���JF]�"1G� y��͝�!�$
k�詁���@Y��d���	�!��.��I�&�m�0�����!�d�#njd�Q�B9(�Ҁq쓒!�5ond᠈Ĺ/dй���j`!�$��z�^1H�MJ�3�z=�q�ՓT[!���C��ᕎ�
�Z��S��">!��F� ��ФP�*��4�&']W-!��z�6a��0W��B��ת%�!��Vl@h�_X ��ANF%�!�A+yǖ��`F� L@4*�L�'!�dИB���Ҍ�&�u��k��y�!�DU�)��5��Ĉ �P��Í�w�!�� =|�P)�C˙&��캧,Ζ\�!�dV��
a��K�,��{�k�-!�$��V��k�b�=�\�1!�� �`j��S*~���EL��#AL-à"O��YѤ�P��h)qd�F���T"O��� �;[��P
ѐ�� 8�"OTU�"F�Js���ɮ��"O��c���zVq�.ޭQl8H6"O4D���#M�0Aː;�L9r�"O�ճR�^&v�9!L��]�|�g"OX���!��/�⁺�ȑ0w~��"O�m(�� 0k�~x���N���"OF)�MR� ��1�f��Ӧ��*O�(���Àkʴ!�c�a�J)C�'V]pr�Ni����@�^%W�~\��'s��3@Ǜ�q�`���U[>��'��)�A�n�f�0���8/�h	�'�0�J�@ 
�ɻ�j�)��z�'�x�&��2�����R��8p��'6V5��aԊ�t%���S@�"�'6�ٰ��$�a!wi8=d���'n�Á���S���k���:	�E)�'wvl1���lc��P�.�:�@�'���iΟI��X)�ȅ�P���������g�
�
��E�ʌGN���ȓy`ɐ�Bٸz` D	�^�W#�L�ȓw֦��r�:
�0�0���	I�ȱ�ȓ?8�q� +��p�lŁq��t�ȓ�8}(3�����M� p�d`��=���M�,��s�nE8>n�d��(��q�C��g���E��`����ȓ4�j�� �ڸ�dnW�R��t=`�k5��7ư �'-��p��ND�ĉ���'g�����/����M��H�W
��a���͌+	�	��WȈ9����;)����'t~L��>���c�=V��+Q&�<=)�� ]�uS��(��Q��D^<�ȓ �qP(�#,�)��EN�;|l��6�[uB�h]�,p$�c/�u�ȓ��:�%P�M��"D8I �y��;�ኀ�g� ̡ �H�ܩ�ȓ)��e�נ)�(p���(Nr܄�g�P���@:2i���u~rՄȓP�C��ڤ$�P���V�vTɄȓ)�X�m��,��&C�=X:�ȓ-�����+Sr� i�%��R�L�ȓ^�ڭ�1�PnDxз)�:(	�(�ȓ�������_��ɳ�%��[�����G���9�c,�J�c�i����}�ȓ1��hP��Ky��Tb�WS��F'�)�&F��n���˱r���ȓ�y���Α7��(�V�M�4Jń�;�<Z���Εbы4L�ȓJ��@1�`�C�����ޅb-j��{��b��	E�
��%���l��ȓ2����@ǱL%� j��[=7�����6b08����}�ܱ��<B������d`��� oV!R'�ܸ�1�ȓ}0ST����@"�(7
�����#�Ȑ���U�U��m�-�3�����x���!"��>�6�G�vꄇȓ ����ᑧL�P�wNPfr⨇���Q�	Ւ_)&`kC�_�������D`��5�3b��ȓdY<kQc��85N���i����N���
M�"�I�3�G
&b@���S�? $i귦��V.��ԃ��:  �g"O��R�
\�9�U�J�I)��[�"O�2���R�ļ���ֹ8 D��"O(�i�?�q� -C�W1��S"Op<c�"�K��M�w���"����"O����m�"�A¤��2芁`"O@r%�#T��1��[D!Ru"O|�+RfL+o�e
�Ӭ%j��"O�S��
�qY�	B��.E6��G"OFh9CC��Q����s��,G��A�"O�b��^8Aa���C��w²HR"O�,����j��$�6���Ё"O~��ŉK'E-
���T
,`��"O�diDN���G�J �Ԃ�"O��Q��zpa�e&L�]�vX��"O����o�
)��Ӳ��/"��i"O�$3����[(��ZV$�"8pU3�"Ol�C��0F��]!�"C Nȴ�Q"O(x[�m8H�&c}�x�ča�<��Vq<�%��G
M�<�4a�<���^Z���TE�~j萁��S�<���̵-V5	7/�s�,a��M�<�a1�\)�2�u�9Vb�T�<a�o׌�,AZ�&�>�E㧈K�<�G'K4D�,AC���a��㖥�~�<Y���\;r����-8�z��{�<Y֤�#W�\����8���z�<�R`��Q'*<
�˚B��lZeL�t�<q�Ɍ�A�d����&8l"��Vq�<� ��2l̘ ��,It����j�<9R#^Q���%@��RX��eC[p�<i��"C�����U&
�Z�cv*Mi�<сe�$txܽ��m!t�¡���GM�<鑪�T�S��QUb����L�<a��N�"]��IW��E��I�d�<�c�I�E��Tٗr1~�Z�^�<��΀�[(�����WT�U�FG�a�<Qs䈧4k���Go�e.AR�N�]�<�5�NB�B�Z�@s�����Hs�<Av`�=`��h�>'R�C�D�<A�̕�[�dP���H
�z��E�<��`��hӤћ��aՐ���NEG�<1�"��
�<9�H�خ	[��YA�<1�ސW���[�I����v�^h�<��لjܜ��J�#���!t�b�<q��]�2�q Oڇ-�&a��`�<��$S�*B��yǡPO�ʱK��a�<����5��j�/\�˓�_�<��F�>(��8I4z���SDM�^�<����'��N�6Bd����A[�<1���l��1�D1"�R�k@o�W�<	���Ka$(�#��vB��PCQ]�<�V�l<�k0���I�HT�c`�^�<��o�-���&��*; \��i	A�<�`�U�|�6�X�
��w$p����T�<"�� �I6/]#{+����*DN�<��K�&��2�F��@�'p�<�!��?�X�Y�菗nym�-Kn�<��![.%�f��F��JFhD�q��r�<3�,V��
%�քZp����
H�<��b
#H�lzW&�M��C��C�<��"��uP�I���ړ7��4��aFg�<I 	�(o�X�3M��	�n��-D�IA�Y�3Ϥi�H�nJLuQI&D�� �Lb��gک�&9/t�!"O�X��wft	��h *z2!"O�4[qC�O�)y'-Y$A�$"O `�Lc>𳅆�2Y�}�D"O<�#�+_Dm�ǅ]��NI�F"O�D&�P8	<$��c�&_|�<8�"O�����?1T����@�<?m�B�"O��Q/�"��� �Q�y;�"Ov9��B(0<�֍S�S��`"Oh�AրK�N�2���0IB�I�"Ob�{B�U:���0��"M�2�u"O����QM.4���(����`"O~��,`�.�%�E>k(�b�"Ox���b
�90,��(Q_��c�"O�d	bI_+,�l���;_e
l�#"OT8��V�t�B�c�F�N�`���"O1i�h�54�$Բ��߉Yy��2"O�-��� *l�����. ^0l�&"O��a����x���W��3f"O8�� /D�5�1�R)hqnp0@"O��s�S%Ƒ8Ca�9ol8)"Of	��(��=�s7�CaH<�"O�����б.���/�+J4I�!"O����F�٘1S���Rc��{�"ONE�B��4�&��"�qK��! "O6E�`#@�tf$����Dv.���"O���1��F]��X�$�2K����"O,��s�ٳs���d@�#=��0"OR!a1��(��T�D�=���"O�!�
E�Z�0h;B�×(�&HiE"OB��h�� ��S�
�7�V9q"O􈔤��<~�=z���.0����d"OJ!���E4 ��$A�AF.>�^��&"Oڐ���fp<�E���&�B}��"O�H���>�Q;�e>�P4�"O�U����%0Xp 2/"��[�"O�ӂ6��i��Awg,�Z�"O^�!bΗ�4W���A�D�Uȵ"O�0#G�۫:�	;�	 튡�"OLHb�̚t�"��2N�#�*)z�"O, ѣ�t��H�vl��Z�"�q�"O���BO�=T��Q��]�<hQ"OSt@�T��0��'+�Zy!�"O�bS�h�JA�2�^�}����"O�d8&J�'B9<q�
ɇ4�:`"Ob��\�	ކz"�<E�|Q�S"O�ŉ3���\�x��һ��I1"O~�PC�8Ar�(&��+��eP"O�0xGf!H�(�O�%R��z�"O �'FQ����s��;��dK%"OXA��/9?߸Y:��<�P"O�2bӠ$1�Ѫٿ<�-�@"O��2�d��1���3�� "O*5	�V�IƔ ��%�2H�"O�h���]�x8���k��0r"O�#�l��^�|�zG�<a�f���"Odq�d#Eؼ��W�e)�t)�"Or8c���(����1���t8a�"O�rB�H�I��ȱG��J}44��"Op`�2���'<i+���:Y�Pᨶ"O��)w�x-����'��� "O���#d�<&h,-���E�b�AA"O�,�&$�-AL~�ɡ��2�
�q3"OH�� 2�(B�fՈL|j�`A"O� ��ÔE�.r�����%%L�x�q"O����7"��3feoEP�z��'k���R�D�9��/��0v�y�=D���j�(�<颁 (,�Z��h;D�2��[�5�&}��-B�}�:@K� :D�Lڷ�!%È4ȁ�\ t+x�@�<D��
�K��3��M��J\CE4C�;D����`��;���a�Xc2ȕAa$8D�0
r+�)50�,H�h�+h�൒�%7D�|����1���IES�*�ӱ�!�	l�'��	= �t P�Oϻu�4�@�*�O��B�Ɂwah�S�Mϥ���4$�*_�B�ɬ$�$M��k�3��a�2m�.5��B�	��D��.�1+�A��/
�_Y�B�ɤ�X���$�h]��7ȦB�I�EE.� �G�^c���E��h0�B�I"1�R�p!�m^r�����nB��,,�n�0u��4�P�H�#c6B�	��]I"M�R">�'�u��C�I�8*s.��w�p�����_e�C�Ƀ>zp)	��9k��QCŜ�\bhB䉤C��<���\��Ƨ� �B�I��D�@�lZ2L|e���=]�HB�ɑ%���v�˥! j�PGG:0CZB䉞Qu8�3�+@�R�:��4�#r�XB�I?uz�u�������ev�B䉘Vj]9� P a�9���_�D�B䉉��R�?\x��`�L?.C�ɦ��'
?Q�8��V&VB�I�$n���Rdˬ'���2�� 
����<I�'��p @ǂ�#�xI��@�B��X���x���3c�Q�`^�^(y�C_��y��ke�����*D�>1�tj�5�yB��N�eq`�Ȕ6��#̈�y�`��6�v����Z>H�L{��5�y�iӊReY�$��8�hB�����y"�V8c�ZPX�I��.E:h�$�yB&�PY,�H�@
	�H��c[�y��ҝM��hP���p�J�H�"��y2b��-H��+�-Ѱ~��ԑ��y��ʙ'j��b��طK�h\�@)��y���4k~ 	�A�4hz10��1�y�M��ua@�#��
0(�]���@4�y��&*0���ᩅ)!IƠ�9��=1(O��I�r���r���XK�N�?a�C�?� �y��^��U�*֋�����'�HՒ�N(5f��"�QC�1�':T|�fM)&Wt僴ĎY̌�A�'`�Hү͌uڀ1iC��eu8��'�V�A�I˚c�����D�S���	�'l|µCɅ.@qCf��4���	�'J&�rgÓx|(qgG*)��a[	�'H�պiR�y� ��Hҵ��@�'D�t��o�<�����̢���'>�-pg��}d�@�ˈ��m��'��9f,�tE��"�2$�z�'P�� ��S�Q*F��	��Y��'��m�2�N�g�H ¥��Tg���',���x��)�/!<��H���xR�ҁdpT�Ԡ?̠��[��y��������5�	b�.Ѻ�y�jR�wӌ��' �xoP`��� ��y�@�Oe���������y"ÛW��e���0��ò�'�y
� ��K"�L(���E<n��܊�'j�D�AX��LZ�`S�i�6!�$�!B�T,�ф�	1C>t��J2Y!�d�Rc���2Cʘ=�"DV�;!�$�(8|�$e��&�ޜ��ԛF�!�Č�w9��!��ڮ0�zH��ߟI|!�$@�D��ԑ���7�P�;���_w!�
�(���u��8*���Z��
@h!���shf�귈��)꼱����8!���
-0�Y,� \�bf��2�!�D߅ ;�dp�ctV\QSP��!���D���9$aD$rE�	ڳ�[��!� |�(�`6C�u���;�/ƙp�!�D�;f��x�K11�h@�-J�x�!�d����oG����z�lB(=!�ƜN��Xh`뙿Gx��r�
:�O����2?UZ9H	��Yې�$Zu!�DG�/�Xi�a�#چX��N�:Q!�dW�J<�5�E�].onB!��,l7!�؟-`�\cQ)J�mba�DGMB!�$yw�5��I��`�	����!򤟆N?�,� �.��U�P�N�!�R�?��U�A3�Ne9%`�4�!�A$B(�4��@ĭ��9�4h�!�$S���$+�͚�~�>i$�@�!�'�X+@�p-���ރ/�!�D�C �@
DLz�� ���*/k!��13�d��:>ܹ&o/}O!�D�H8%Z���2xg(�%�ʜ@!�D��/�h�&	�t`Fi��
I"s?!�Dǲ}�mh$��o�� 	;]&!��Y�Q����J�[WŠ���J !��F�24Z�p�`ڽ6vx��J^�q!�D޴�]��K7Ig��D@5!򄁡KP`���R�Z�P)�A��!�K���s�"H�g�P���
ԶM!�D"5�����Р">����¬v8!�D��!K� ����%s�հ�מt$!���vi�X����E�Zq!�dзo���� �Z@f<
��R�!�D�S�J���h�R�u�$>!��;�~�Є-S7��L�b[�\�!�䛩��C�̓fFkQ'�D�!�dīO��M��J���䆚�o�!�D��2����ٰ]x4�q%�%P�!��� ���)��']A���#$ӡN�!�D�9{~�3�D�qh\�'A�&s�!�ǇK�~$��@;o�8��D`���!򄋒8��$A�(Q�u(dU8�.з"�!�$��(lx<��M�.t��01\H�!�D���)(�	��=T�PK���$Hr!���&e��)��݃hOܹ�$��U!�d�/_qGY�sX���	�n�!��7U�*İ�n��A��Q:&�>�!�D�r>�@�!C��>��9�T&��p�!�$�!�l[� עT�Ig��B!�d[z�e��دP{���5蛫, !��Φ!�&�ӅAt�(�5B1;�!��ɾl�����$߱_���@���!��^Ŝ��Wa��{��]q�C�*�!��<H��}adO4Q2}�d��( �!�>)��I�'�S/+�>�0�Ƚs�!�$�:���P�ŏ�4C�$z��C�/�!�W6c�A	��J\&��C� ġcL!�� (b%G��� �.��j Ńe"Or]Af�@�i
h�`T�
�/��@B"O�9�bA�i�" iq�I�z��"On$A���->��H�֏�"����"O��e*�$p��0 NK�|�bd"O�y�c�&Qz���d��19�"O����O������)��G�
�:0"O��j�������L6G�25��"OX����'�셲E�E��lS$"O�	�T@/vn�W����4Bw"Op@p��k��C�aA�K2�1��"OP�e�;F�d���o:�R�!�DPu�N�B �:I���U���!�G�9�lD�s,�'k���V�Y*�!�ĕ/vH��eM B�"X2���:^!���8#���1�F�� $���jU!��oP@�F�[�kpd@���9d�!��*E��\�׀idh��q���;!�DE,u 0S�J�Ml���s*�(H3!��[
�
�[��N&=�5*]�!�$��j
�jN9a�by���4!�D�B�T��Bʰ)�FW��!�d���$��E�8����}!��84K$�q�*�	�&���Gc!��ݙ*�<�;ńʯCϤ�3-���!�́F9|�bB���'ɊqX�A�CF!�䜥�*�C��U��ukӀ�p�!��d?��E�Z�z��� @�"r!��S��P����5T���2 �"�!�$Y32gj0����MS@$��;�!�D��@��!��h���-پ$�!�B�����zs���;��C�	M��	����9\�
ŭ �4~C�	�e�X8�a�������� 4S�B��jh���'#ů����Ă�4tB�Ɍ'x(p��/p�x&���HB�I1�X��Q�Ωq9���g֗t,�C�I���Ă�����I�T�*�B�	;k��H��B*� C�6ϪC䉾���ق`�mæ��FHЭ.M4B�	��:ᑲH��JfڌrG���DC�	>f���^�bB�(��_GC�ɱ!�ư���W+;��A���r`�B䉺=V�XG��3���@�-Z�B�Ɋ~A��WB̿����A6d�nB�I�@��#e��P������t� C䉞 q:��V>)��3��@��B䉇,l��c#�&GlhU���J���B�I�a!��RG!H�-����$	� �*B�	)L�bSG
�r+�M��Ɛ�P��C䉢[��x�Ц�<,*�=Kׄ�_�B�ɠI�ʗ�ּ �zQk �߸n�|B�I�X���C�@�1�N������F�pB��_j�y��K��<�Yr��g�PB�I�b���k(����\�lB�	;9��ɕ�Y�H�ҡ
�T4JB�	�5�̡��]T��kV��T�B�	5~��<�'���{=d$���R7d��C�I���zh�-=\�� �5&�C�	�y�%`T�	Vo�%*��˝dn�C�	<f�ı�DH�lʉ;QDɿ#KB�9�tŊ��߬}��p���ZF�C�ɠ�V�A��H؝�B@�b�2B�I�8l�5��7p���b�nŐX@C�)� ̠8�c3+H�,�U��$Ҍ*c"O���bD�\�̝ĊO<��
�"O�����,D5�{e�?�*9��"OZ�b�I�k��(a��<tɦq�"OXи�F*\���l�{�v�y�"O 0�υ!ڈyà�!�$i�"O�	�t�[ W�(۷�0��mj"O�@s�L+]&�1kV�նm��i0�"OХ��-�	��lje�D)	���C"O�4	��p �'O�Z�D�v"O�A03�]'��L��v��E�w"O�}��l8�iE-t�98"O
�J�HF/��$�(k��t"O�U�(\�ܴA�-��$6xrE"OU"��O�w��A��mJ� 7��*b"O�h��N�m�P9��J�/3�H��"O�8�B�)a���It�RP 郡"Ol�I�#Af������$[�AU"O��� &D��D�q*/q:�+4"O�����X7�;�W���F"O�P�B@��u~��zǁO�cV|[�"OP8���ǓU2��f��'.�R�R1"O�h��
�jc!�?V��$�"O��B��M���bbT�u���#�"OThأV�e�DM��ҏ;��� "O������6�:ucZ9Q0��`"Ot`#�O-I�B0�d��?3j96"Or�p��kQFI1���W�*��"On���d	!�> ��1�"O��(�̌�t���G	�H]�E"O65i�Z�DE�K���6a�Ѵ"O��w�޴m&m`J��`E�"O��#��4�BHz$g��>�\4ч"O p���ѦJ����pf�&*��C"O>P�پ{�Ld�ԪG�f�2�"O.�R�ؠ/l���G�vI��"Od y2ˁ�rejV�ٷf�^���"O,���R%g�Q�t&�A��'��� g�O�fu�p���$�	�'��`j!
D� �Tii�LL	6 U��')�	��J�%;�x�'M��{t�!9�'�:���I)"��8���wM�X�'�`Q���0�H�ZR��u�,A��'4@��(��@���3v��2�'��H�bb�*kc|��W�=ET�8�'�`�>g+.�z6N�5[���
�'Yj%+EjͲu��D�0�Ս3��uJ�'Z�:G�C�}Kt����C��!�ȓ!�P�s��k��8@�%T��܇�X�̄�#ȓ	�h�g��� ���5K\]Re�<!,��ZҪ3.m��.�@���
���
����ȓ<�0}I�%h��X"p�Ӗ��(�ȓY>�p�nC3gBv�:FL�w����z���kQ���"�V��$F楄�.0vx* /ҏrZ�q���E ��ȓ}֠��3���x޶H�� LxP��sǤx�Ƭ�#:����Ш�.BA�<��):�� K�"`ެ��GB�<�A/	�P	p�S�=��Q�S~�<�4k�* (�t�B��]�!��|�<�2��9���caHN4)|LPf��N�<95��?!�.l�V/D����EI�<��jI.u�z��5g2sm�9+�HK^�<� J\�wo��~uaP�NԔD�2y"OV�hJ^4V�����
,��"Or9���ՈK�Tz��۴2o�	�"O��`fB#:��B�,L
!^z�S�"O�-���+5�`l9!J6B@��X"O^e��]3�%yb�Q�U��H�"O���0/�bl���֣�E"O�]YU劚Ò���<s$��w"O��3d%K7	��+�C��($"ђe"Ot5�3i9Y�4;��Ҍ8�i�#"OX��H�D�X)�5jC�}yХ�F"O%P��Bb�T AO��bm��3�"O�!�1E�y�ZI��'��Wc2"O�q�0��`�xР`H�1ax� �"O�� E	S��1��t����"OrP�t�ZVɊa����Tѣ%"O,j�CM* c�X������"S"O��"��=���q�A�~��MB"O5k� x>5�W��:�V존"O����f;�Z͈y3���"O���eo�:uhB΍3*'n� "O�T{�^>9�,4k�K�'"^e��"OVɺtLE>pCX�4)� �e"O�Ib_�R�n�a��#��E"O	�CdN�"��\��/n3��"Of8a�m� E�P�bh�!�\�"O$!8���$wT��'E�<i��W"Of���k��fJ
��E %ļy�"ON�q#GPn��i(�d����x"Ot	�w�ўM�
ِ�� �~p�jP"O�]�k�7G�rIQ#D�8W�Ų�"O&T[aB��I���;�i�%p8>�Bq"O��
�%��D�2JP��"O��+����~Od%3��M�> htA"O��ǆŚH=�-�� �5H�s�"O��b$Ym�:��Ca�+��!�"O�}�'�.^��0k4�$&��!"O��s5IX6s%�� �?ljH�3"OH��$V�M\�R2/D�
�&]�R"O(36	�?nKZ�qu+Z!:�ȓv�*��q Ya���@6D@��J���*���#� �*��� W����ȓ!0��#N��G�L5�$C��/D��p��](V�e�!'�A�pl#D���c��,j�SD�H��=��/4D�t[��"v/&������w��њ�4D��
&�H�Z��t������r��0D�dr�޽U���ivmsxac!g+D����.�&G�0�*WG�1/rT�i�i)D� p!"U:3c�h��a..��p�%D�4Qsn��d�(p��/ЙC霼���$D��Ga�Caޡ�J�Db�q�G/D���D� �"�p��˗ah}��M,D�h1BB�:sl�2�̖��@��)D��� f̄�"S�u+ڸƥ*D�X���'wx(���Ͽ �$a�3D��`/H5hB�l�7Ǆyɱ/D�������=�^�a�Lʋ�XɃ�7D���DyôX��`�=BBp�w�4D��hP#�5�zY!�0UX4⑆1D��K��H�_He:�@�>+BRb�/D��C�͝>\S!ED�B;�ip'2D�������E�Ӌ8X��u��%D��#$ͩo��jO�A*��Yd�%D�� J�;� �d�ƍC��A�
ي"O
1jB�ʶo��p� S9�R	�"O� � $��ɠ�ϑQ��,Pa"Oڸ넇�d����C��,�4���"O̽���)p��2�aS3S�p)�'"O�8��j¬v"2��OG�L��!r6"O�u�f�[���6�liy'"O8�g��>A�q0�kH�2��q�"O ��b��a/�|���3Vq8���"O� "�OD N�	'�A;gb��"O�(H���R��
��\	�Fё�"ODxP�	2X�ypF)`���R"O"��N�x� ��f�&�Z�X�"O��hӶ�4� �z�H��"O��`���M���� �A �`��"O�]�DN�G*cC-R�zț�"Ob�G��xv9��˙���R"OL��С�E��T�֩>~�2�"Oέ		@tjddI�Q��Xk�"O|x�%V@
T		����"OL���M!�j��ǘ;o�ճe"O:aaa��9!YDM�$�R�S���90"O"h8@EW:)�r-2�L�|HR�"O�Y��I%(�2�`�#�D�9�"Oh�ZV L4tb��\}���ju"O�<�fC�n����S�P��ꕑ"O�����D�"Ծ��C����!"Ot`�*S�~�J�c�#9����"O�i(���Q�gc������"Odx�d���ʩk��)���9V"O4���Y�T�y��Ưs�D��"O��࡞�190��#H^R��� "O�)2X0|����@��sB�=��"O�h	$�O���E��""[d��"O&hɒN��$�����[H2��"O��#�}�Vl�Q�֙34�`Z"O�U�
�/I%��D)��V򅂓"O��b+6S�^X���u���s"O2��cؘ��঩۽}��TAT"O��*��� n�pda@��y��A�e"O�a�oG�V��8�U<q�f ڤ"O���g�Kz�a⤎�aҺ5ۤ"O��8S▶1��Pk!m��S�T�g"O��C7lQ�ܸ�yցf�*-�V"OB�3",K�L�ņ�b�$�)�"O.|��߯E��DЅϲ�Y�
O�6��t`����2$�VAáa�=�!�� %�\�����f���+�'V`2Op0�e��@���E<\�X�"O,a�%��+h�8�,��uLBd�#"O��d��G��YSqM�<"O��:e�^�q)��3��������1Ӓ�A3DvCva��u����F�Z��%�[*U|d�2��+ ����*�4iσӒ�RR��>P�$)��}^lіƂ�a��]*��2m�:���u���E�+z֔�F2?Slņ�k� 1H��Q��)�C�Y��$����}��ԙ:0�i4%�)M��I��m}t��`Y� 	$TA��h�9�ȓWa�(��aئ�.�
��V?9Y�!�ȓ��������d�^�{�HFV�U�ȓ&iX}�L^�TƼ�+�K���ȓy���g�ۗW��t��|.T��S�? ������6*�����M�z���"Or	�,�0:�����׉^�Ԛ�"O��j�M%�iq���[��4��"O$P�6ćt"d�T�D#3*^%��"O@���3C´��E$�\�y�"Oİ �E��xxQ�/r��$"O,q'�W�ڨ���J
*a�"O��R��W��N��P H����"OB�c`�ζAXd{2B:�"��"O���P�gh8�*V4�̥P�"O`�z7�R6Rj���@�(k�X��"O���oñT�T��`�0 ����"O:�sE�5I\�3.ޔ'Ҫ�"*O��"�Z9%o�4A�L.cL$
�'�����),d��`�o�Z���#�')br�Ջ7��Q�]�F�����'o��b�� r@Y�-�E��
�'�:Is�� �JDr����A��0H�'�P���f�0���`�]�4ڶ��'�8��(=,� �IA`uVQj�'�P�#�C���=�AK�/�:�'�j-R�ʅ�X�|��`��x�j�2�'ʦDj��~)r�Pw�F�jNFݙ�'�,��L��+��kݢHt `�'�ĸxaa�j@�<*��UoL���'qL�Y�:`!�䊥��!uJ���'�u[g���*U>�J%آsbd�
�'r�	��U)�
ݚ4Ŝ.X錘�	�'�~��w��PG��bcM2x\r�z�'�,b`-0Lۦ�B �mX�X�'\�9��O�?B�e�N�1>�i
�'�~ԉ�hI<f��8�b*A�.��1k
�'u21a%cА>�����i�Q����
�'�K�yU��b��1z2��Q�<)7ϙ�R PBE�PWH���(�M�<�� ��_�<�5*�kF(�y�oDL�<Q�&U�z�J�³�N�4Sz\��*c�<�7bpw�JA���o��|�#�j�'�y��/������9Yh�$�� Ǧ�yB�A� Q$4��f$R����=�y�[h���R
Q���b�%���ybcJ�8��Hxc�ĜE�v�t���yb�F�¬D�a�$+����f���y«��lj*��^�V����q�.�y"BŮL����֯�0(������y"I�#.;��UO�%F#��r$��y�HS�Z
�j��X�EB �����y�!B*/��%ZƩM�EUT������yRKS��`��@>�:�ie�N�y"�ό ��h{@�ȗ$���ӭ�%�y��d��S� ��^�k �K�y"�	o���qᙝ�������y�d�;K��-Z���R���yb!�Ho���5�	H�I1�T��y��^��|�"/H>M�R �7Ɗ��y�D[@@Q��gO,e�	*'OE8�y�eG�WRơBQ
�|���)�I���y��/�H�f���g?�샶X��y�̑<�j* ��*�|صEY��OL��ȢJ��h���	A�b8PEb�!�DV9ef�$ȠD�H���P��_J�!�DL-�\iQHO*��8�%G�!�$\"�$qcUN��2�0�O��_
!�D.h2��I�4�L��eKO9s�!�� ���Q�;�H��f�-D��5��"O�Aې� 	A�dFo��^�H��"O�(�jF�g���-�>���8b"O�,+�M�)�^M�'�7>��L�G"O$�F���]��B�����"O �T�Z>MN`D��g]����A�"O�Y2%֥5�$�w�E�-K�k%"O���V�6SB Dh��FK4`��p"O,�0F��8��y0�(l(L "Of		��S�;:9���]<Gufc�"OJ�d]V!���jD��3F"O8D�%eQ�G��xr�E�CR.�"O���(ݨ��9��٢,��% �"O\	��"�&���C�G�)!��8�"Oܬ�wn�br�wmȽYZ�q3"O�mpC_P~l4� B�2�L��D"O D�eҋ+�L��A���,���5"O��|Z�C5�ʻ���pn�v�<YEւn`8�U��*P��}�<a��ۭ S��vBH&(r"£�C�<���Y--n0a�$'��i��-~�<����n��K'��) "b�h�t�<�D>
�R����G*��e1�#�m�<��̜�4Az$%ٴ0&5��A�b�<��(J?�Y!W�I�Y�^�	�N�W�<I��3B���֠Md瞱��!V�<�3����\�֣_$~~,�4f�Q�<ˉ158hXpMY�eQ��@&R�<�cvj*F��7������Y�<�7Œ2Bh۰ʯ)r��`�U�<&�F
/A��S"���(��a����M�<q���@@#��N%fV1@�h�N�<	�"%��P3�J�5�FmM�<1��[ ܼP5�L9�j�`�J�<��]�u
��cJ̑~����M^P�<�&nM��ܠ���)0="e�E�<�OSo��ǋV�;Z�A��A�<��iIE|��:A�]�1�wh�|�<��9�r��� �-
�%�`^O�<���Jt��Z�oR53JXy�G�<�%F _���S6$�es,�@�<�ʂ!>D�떃��"��H���V�<��˞(V�;w��5fIq���~�<���6.�9[ ����a�łIs�<q�σ�%�������e��݋2�Wq�<�I��4�D���a>�`��r��l�<�� \G(��E��1pXӦG�r�<�FU$3m&z�I˩	�-�`�o�<aC� &4i&o�%S���áb�<����i�� k���<��$	g�<)2�K�~�U�KΜo3�@I�+�b�<�3�� c�ȷ����$=!��TJ�<��� $��q��gA�+��iz"��H�<	c4`帍!�
β_����wD�7�}{�n�����+�X����*[�Cl����n��\t�����.D��0n�S�����ʃ> ��3�.D���Q�1�4*D�jS0ݡ�-/D�P��S� ��T �"@�"�}p��-D�p�Q̉P�Xᔨʗ�>@ˑ�9D�����³:(����#+A\�T�7D��@#kS�n	P�;�,�5��l�5�5D�t�Ԏ�$a����a�ƕ�h�yS�>D��(�AA�m"� �8Z��A��*D��@"��8�8��w@8�J1K�+D�� �Q�,Ԋ��e��%�T�����"O.��W��?=��=���;$��T9�"OеC�KTK&L+��V	`�8���"O�)8��S�L򁐌Q��9�6"O���*�ؙv�^�q8L�RV"O��eL�=()v�cl�_��$"O|��ƇtaÄQ-�� �aQ!N�!�dϖ9m���ڋd��� �o�>|�!�Ă���(�Ҭ��)�`MQ�.Nf!�Kgzt0����������-��cQ!�d\�-� �Z�I�ɚ�"��!��5�L����>Zȶ	��aW�i�!�Z�� 0EK3��ݪ
H6Q�!�$��_�ܠ���|�R�K6�]&�!�ȫU&�Da�H�N峇���,`!�Ą�H�v�Ht��5��0�2�Z�t!��QR'L�$���FI�K!�ąu�$��R�����K���!��\�H�$R�	�P%���äs�!�����
`Μ&x�����'�!�_JP�ub��x��xa��>Kp!�$�T�uBBO� %��['g��m!�5\�l9B nq�V�G�<o!�DLX]�@#5���1�I��43�!�
;B{ب��M� ��p4�� a!��>*�Q�E�ݰ�V�����Xc!���+|a�c&���|x�D(4!�dT�7!"{�Ȕ37ڄ�z�$ԅL!�$�`J��y���8I�p��!�U'R�!�$H"&��Ip'_�k4b +q»Rc!�D�3UN��*��5*D(@䎴�!��PO����j�=�:��!BG�(v!��C�ldN4�wƙ/���;�y��&]Bm�������.�N裢J	$6J�3�΂"�y�o�<���B�!b�a��Ϯژ'`�Y�On8��P��C�$$�%��F�5��Cc3��hb� ��1�īߝi\4d�R��|)�
O��t�^�mgL�� ��0�����'��@C���lܓ@Tq�T`�T��c��S5Z��ȓKo�#R ��c$ΠPb�&`&0�'�F���e�S�O�z�Y�ςMٸx	 ��&|�zٲ
�'�`%#7o]2[�Q�玔3v��K�y�.T�u����7^� �!�L�2E�A�B�8]{�Bቯn��tI��44��f�0z���B�WH<i�jҵYh�#�f�4S������ _�<�b�I8��$9� �'�Xxf�W�<)�@1|������6"��u8-�g�<!�*F-]�H�ҫ-��@6�b�<YAf͗(ZxY�,)sF����ʕA�<��L�6u
 ���epbh��͏f�<q���+h3�������J��s5l`�<�m�,h��������$'X�<���M$g�"��ǎN%z�R�P��[�<)&D�N� U	gJ�&_ST((��M�<1`�͉&��`� �L�z\��f�Q�<��N�'
���REnP�$�v́��L�<��1�R=�$�^F(���O�<�!bX 9�,}kS�T�a�h�H�<aP��?QRdIT�Տ���yE-J�<A¡N28��sl[dxl���y�<��G� ��U욍0)���(�v�<�g�[�bo����LI�+�考u h�<�㏗.���AG d����B��b�<ٖ-ɽMDd����G<H��P�<�  ]k�
�ui�`�2O��	�L��"O��f��v���5���$Ţ"O��23�P�p��%���K.%�L@"O��P���;�R�vbF(݈\�"O���ƫ�:R�h�PBH�5X\U:�"Oິ���3�΄��lƘZ�h�"O. �S����mXrL*y�&	X"O�LJ��+��;�L�43�~�� "O|@@�(J�d}�17JY7C�@X"OR���ϕj�~8X£
k�b	3�"ObhpC	@V��	DD>��b�"Oܴ�I��D��"�U��A�"O��S0�7�E
����@���ȓY ����M��/p@=�сE$:V�݅�u0!��h�L��7�ҢB6��ȓ=G� A� ���$��'_9��J� �1"� y$��C�+P'|�*�ȓX�eQ`�>pn���� �@��T�ȓ8��hpĒ7 }�y�D�F0@����/x�]0���<<��JƂÖT��d�ȓf�䬸b 	|��M�@�M�3$�͆ȓ:��`!�+R [�d�p�+�\.݆ȓ7\�a��+Z
mKډ��HN�sQ����;�&y�W�"�N��F�H,Zڶ����%�%�B�9[ �� �ϩgxTمȓ޼�[@���b����S��` �مȓlL�v�A�2���Ď�=���ȓpY�9����="��������Ԅ�|��� 8b�6����{�����P�a��J�[}����/)�b̈́�Z4V)9�̖k�e�qc�Ӥd�ȓ@=22�иK��e��/Fg��Y�ȓ�V�`I$(�:����<0�y�ȓM��,Cf�}rP`���I>v/����zI#��آ�i�e$s���<�u�r��b�״�h�\t��� �ȼ�����Ƙ��"O��p	W�LC��H�d�9a*�;eH� �v	�$K�?��R�BS���'��!��; G�!��.�����'�d0P�߭*8A��	 8]hU��&�͊��9�r�c�E�����H�����1$�<ul���*-O,8�VOǎ#�t�3��Wm�\y�/�C��B�OCB�����̟�]k B�I?]�\!�JU��a%� >�ʓU�ZR$UZ� ����׽"S��Bu� ���m�H��E��#�:���m �B�ɿ�tu�v��P��(���*F���3�׆i�P+�i�(�JI)�$���'.����ż42������M��X���*԰]��ҙ-��HD��`O��BÎT �څ�"N%B�Q9�$��6�@	2�=O�ě�͔�4����%�F�t
��	��D9bC�
�X�Z �I%��ܳ�ˇ� X���q���Ga�]�pȐO�}ۅ�U~�>t�0�ȑ(���6?O^}��k	��<�-n��Y�!�}�6x��(���5�v�#��ʷqd=�$aU� �!���.J����Iǟ g�ӣ�H*?����ʞI�f�!`���?������?��#`a|z5�'���a�IԿ�B�����P� %"	�n�����̪HH�_
@�����&A�n��3$��X� �<j�`p:��F���O�����^��\y'HM�r�3��I����R���.���`�[�u��9RaK�
z�0��H�l�<E2a�����ৌC����f�R�I����o�)T1��uKy�|��ؼr�6��CX�V����֎�M���3�Bi�S4U
$T�S���1�B���Oٛ`�tC�ɚ�p��W�#��xyf�Y�`���Q�ƻH1d)c���f���[�(F��,�B�/O�L""ҫ[y��a�K�+�έY�'�м"F�Ҩ��dꍤ-̎�Z0����$3�A��J��t�l�� �]#��M�rџ����֮%��d蕄D�����4�{��Ť���� �"N>]2��g,$�&���@��w�}���ٻS2�0p�����?�֠��
��Xs��R��j"$��<��A�6��hb)ϩ Oh��.��h#�J���a��ղ��Hw���to�"p�<���S�? H1�@�(0Fp���iz�f�
��R���J���k��S 
�2EM�CyB�Q̬�⥈�%�$D�B��0?)FAA�@�ޔ�$��>���!AFEڶС�+<L[<	0P#ɽp�ԍ��x�T�ˌ�$�#t���PE�zp��0f�7%���jTN����O�D�6�^(D0����T.QX��jO	}���� ��J�����=�����+��0���Ad�3:��rOI���!�d׃��!��!�?*��&?�`'J��N�@�nƷ-��K 	2D��`�IX�]�.X��m�p�b"DB��Ř�zwB���G�%E��O��@��O~R�.e���Kۇ�v�ڷh���p?Q���=*�vh��� "`d#%�A�]�E����60P↷QU\�a��,ܼ���X�2�8d��>e�}1�f¼m6�����A�RY�1��K�6�u�1�ElU��kVFKW��`C�"r���v�Hx(<9B�\&`p�#�X�6W<]s�qy�i�b��H�$�.m���U������~�`&V�
p3�gЦN4���bp�<�VcŨ������rup�z����Å)��#O�rwt�b�&r�'��r�B�(�-I|H��)I/h��U��d�۷���
|(%f�Z� e�d0|hr�H�@�Pa`d��-2LO,2h��_���;@E�)Y��X��'�PY�W�J�R�t�� � EA�3!f 5V��
oAx�H�+�!�d�;#%dR�!�+e㔉�c����1O���C��碵;Bb&ڧC��ä� =����c�]�>T��ڎ)����4:��D�C��8����B�3!8m'�9k�H&u�Ć�<@������ �`��7� ����ȓp�N��ҧCW��h�ЋT�=��d�������-l���vB�y)L	��9f����	.t���b[4$2E�ȓ>s����!�� �э.\��ȓ&�X�#�ۥN�>|�DK�����ȓi�=��(��+r���t��Җ��ȓG���/�0�U2 ���B��'a6����P:�L����X���!z�!�CM����$͢\�V�3�n�!�d�sz4��Rꌳf�0��&��	W�����'#��=��>I�B��;���⬌*_/�!�i=D��b��^�-��Da5�H�:�����9D�)V�0�v�qB�2:��� 9D�,D`��a��� 	�(C��r�. D�ز�\xW�J���:!� �!D��选� P(�'��al�d�?D��9��d�ڬ��ոr�h@�0D��z��tV6�l+L/x2�q�0D����] (vU�g#��K��z�;D�t*��=�څ�"�8L���/%D��s1�@&I�0�áEʰBh�\��?D�Lyfe�2x����I%+/p}���!D�j���=��Q�bA6(m
�-?D�����.8�R��׬S���צ>D��+A����P��2 �)D���r
����i"T�X�:���1w�'D���dI%)���$����5�cO%D�|;�A�>\�������e�A��!"D�P���L�2q��(]�x����V�"D� 8UhBY-X��F�d+T�#��%D�8�a8^ y�A�q><��@"T����hJ���2#��>���"OXy��\�1��
ŨQ������"O��1a�MJg��3�ǘ�c�x�4"O݀%�ۜ"M������c6���"O����E�1�"�I����A�@�1�"O�Ւ�d̻����w�WE�8="4"O�e��gߚAjr�`w��a�Ȥ"O�
�(T�
�I���+2J�0e"O�q0k�<my T��+-d�գ�"O� �۷&�	`1;��F�	��	e"O�%:q��T�|�5ዩ �X��"O��a�n��h4�ŏ�(S8t�j�"OX�#bT.�p��m��l-� @"O�1b���3�����mK�6B��`"OV8Z�I�04	���6\�X�Ԭ�1"O��A�jR�6�M@g�w� ��"O�̠��~UR��vl[�)�$z�"O��!a�A�/>1P+X��HI��"Ox�����(�к��V)�䡩v"Or���O�K�NaB0g�$<���j�"ODe�!��3l�,�ڃ��<\V��kt"Oz|��[#~A��P�X���"O̅�pj �z�0@T�L�*�"O�0�Ŕ��~�"
Z����٧"Oj<A�:8$m���M-.�t!�"OʴpD�
�o�.�� �4���"O|�%N���-",��%�❂"Of��C$[�c+>�pu��E��,�"O^� ��Ԭ\P���7
�9�Lц"O�Y۶G%�*yaG+�	pPP�h�"OT!ƁQ:)�I@dI'r0��h�"O�lx�g_�p��c��43:,3g"O4��
7L� ��f`�:�!!3"O�Dk��N*m��qrO�4`N�iڵ"O��U΂�r��U�#.%U*���"O8��d��)����C��a�"O�	Ht�׶|f����N�^VH��"O�g ��P�0Q
�NR�L3f���"O.8��O^>�ҴP4G�,7�q2"O�Hb��DP6�Ӷ�D6S�2��"O�� �-"��A[�&焅9e"O�8��A�6V,��0�5>�H]��"OZu��a?.�v�:�BO7�6�"O��RrI���x( �dьUc"O�%Pc��.
���"��F>;��	A"O� �R��� �m��VNmH�"OB��0G�"&�l	�*�2zGt$"O�B��S���+���i7"O^�p�D�HJy	�ʰI$���A"O����&�� ���J�dU.X/8U�2"O�h*��4m#=���-[�}��"OjŰ�
��	�#�	q�U�"O6�25�U?_�v��sV~����"O e���.��cB��7p0@ɐ"OHe
�� �5Ж��),Zm@"O|�s��a:��K�a8���"O�̰��E�K���p��.w�~ĩq"O�=�j�4��Yb�
����"O伂�B�7Rc�ĳu�U)Aj`|�u"O`qB��wM�:G�Z3�"O��#���Jx��Q:D8R�8�$�h�<��'��1b 0,��`�/WM�<q�_�EDr�Q�
�g�<a��D�<a�)W7}�Ա�F��0n��B*A�<Q���+iTu@f/S��Rl��D�x�<����*<��ۗ�ůDd�,��-w�<��%E>
�`o�%#�z�I���t�<Y���`k�\�l�qRz�WMY_�<���N��+��+Vi
�(P~�<�ҼB�*i�L�2"�	�q�<!2�H�jȑq�I\�S!��qNEP�<���8�QQX�J�93��P�<���ٛ92ZP�Ү�nm��AEh�H�<� �%;2Ń�+�ntb�
I�5T4�D"OЭ*0��}KXU��Q
)��"O&�FB�
�b�
Ʀ�T��`�"O.���R&�̐��@)Р��"O�|�pM�sI��q���4�؄��"Of�5�*�(��
��-�"Om���C�([��K#�^�>��F"O��$ۉ�\\�E ��\�R�"OP��F]4F��v�5/��E�"O踳ÀC��p�#��2 ���g"Oz ���l��:���P�jm9B"O��q�ɯ>����r@�ku8�8�"O�$�#��aj��#HA�p��"O�����~ʘ5���޷*�Μ��"O�e0�C���ã�
L� (��"O�5��'�=82Z�T�T"���"O�y��ɗ	��SD� +n���"O8A�$�0rFh�'�T���"O�"��ڑF@�i�@�(w�Z�ّ"O�(�d�<Z��L`!��t��;�"ORpAv�ö����M61��3�"O����&�Q7�\��ɀ �N�j�"O��(�1�R����qƶ�R!"OHr5�)G[b�0����n��r"O��[SAQ�}S����\>:[� "OH���L�Q�(0P� �o$:���"O^U ���3G1�ȡsn��b�.��S"O����T����$���*�"O>E	p$V�?�y��߶Tz\��d"Oh�Y1�ؘyP�IYC��8j��Q�"O�]{4�V�?@�l �ϕ�[��X�"O
�8f���+<��g��Kx�CD"O0"gnJ:(�tX�d�wߢq�A"O�,y��D$-�(b�F:r�%J"O�%B�*� �bls���Hj�"O�9R*W�!�^-+���e$Y�"O �ʀ�C>��4�5�ä<�Q˔"O5S���{�jR����R��"O��C썠i��( RC��a}�A��"O�Dz0T�s@���5"UB���"O�`���8'�H��!�Q�l��"O|�3���0���8vO�<f&�5��"O�:���'{�:�J�LR�a�95"O�ɩ@��:e�� �
�	'����"O
��qgˍs���i��ϨC2"OTx�%Й#�������q"O�r&FS3>�b���*W��`-�yr�f�:����S��]��lA �yrDʍ0Ϫ�3�c�x2|�UI�8�yR�Yt`a�ń0x�يm���y"d�$CdTm��cO+��A��CR��yb�E�`��%�:)�� 򔫍��yIِ�8�!ǸV��$⣀_�yr�5\anm��ė�bh�f���y���Q-��r����2X
�F�;�yR���p�]is	���܉j'��=�yٳ8'���K��(���+S��y��8/�L{DC�-=:.�6�yB��2� ���#�� �F�ڤbϋ�yB�K�b���3�jV��|����>�y��PT��!p# LO�^��#� �y��v���.LE�l9��A��yBɔ�RE�UoՔ*� �u�^��yR��4�E��/�@%q�S��y
� ��0͘�ls�$HW��$X��0��"O�D�����Kl�E9���;X~0� b"O�Se��a�r�`gI
=k�0q�"O�8���	ژ���gH�[m~@C�"O��z⌛,�PS�FR�rt�u��"O���	�d/�L�!BOֶ�"O<�V
�L��tk޾H����"O4��V Ë?��,����(W�B}s"O�M+ J}�(�Su!QU|e�"O���4���/�:1���H/X0��"O�Ȑ��7��t��	�o8~D� "O��z*�W[4Y�(6�p"O���¸er�,��>����"OlH:e]������\�*����"O�hS3 W�@# ��:�&"O�	��\�uNEP�C�2��5"O����FL&p��H��L�5�V1��"O���'�>�pt���F�Z��#"O�\r������*Ԧ8�v�7"Oz�ˑ�(���ϼ�MP"O�(G�ڜz�]*�O�R��12�"O�(*$��'s��5���+h�"O���*����A���x,�0"O���S��0�!��T�P��g"O�ڂD�P���5�1x����"O�����>������V��5+�"O�� ��/�*E	��͝X���
�"Ob�h#�קN�^usfo���}��"O�t����PО�ì��)�j��`"O(�X�d�6�iT���T�Cv"O�\���#�.�1�R�s����"O���B�2i�8K��!~v2��A"O���$KE�j�p�D�(+`�0"O4� «,a�b��qh0S"O�LX��ƐԶ)x�ػUwd9D"O��ya�S�vO&!ס�;Ħ��S"O��U#�:HӴ\���	j�"OJ��$�J�XI�����96�6[�"ON`��^�)0���GIA��0E�"O�ā��.��%sc�;q�8�4"O }�lL)O �`±cE �����"OƑ��K:_�zISl�5H�٠ "O�5"bt<y��	�)\{�A+�"O~�
�'5��Ъ���$.,9�"OJ-��X
�� *V��j�X{"OR��!ɰa�ujH�K����f"O��('Mܪu'�-���0�����"O�h j�*	��]��ΐI� ��"O�I���4�L�E���Q�j��E"O� �r���o��	���]!O
 �Y�"Oнh2bPKLJ���o��A��k�"O�A��mV�s%�@� btnd{p"O��� ('��}�.P�Zhhy�"On��6�^;5�8���CPF6��"O�Qk@G� A>���ĂRK~�#�"O����Q�*)�l;bl�t2��2&"O�
r���&r$!GMK572���W"O��PaU(Y�$5r���j��	�"O��S)9qm�DI�5'��L"O���aMЙ^�v�����
c�p�r"Oa#���#�p=rvBŔs��<�"O4�qqDڌI?|�� �Da��9�ҘH���#�P�h��I3�(��$�����ce$��Y[��2��-W�����Gx��TÜ
��S6�
�9"J��cJ���$�2�(O�>� ȱ��̃�e�a�p+��Q�jx���i�}Dy���W&n���
M�^h��r x�<)�O=<���Nļk�^l�u�Q���H��}B�e���'3��=����&}��S�Q�vVVy'�t�%�)��":r@�D��,�<���K<��J7d�<E��'�DhE��Ο�]�(���e�"�MS�(�S�OD�ms(��7E���@�a����S�	��0|����B�r����h�f�:�H	X�h�d�2��O��I	B[�q��
&���8�L�056�O���a�,akn�!QHK�.\%���	�_����-"�D�#@_�,Ȝ扏I��$jq��S��"�e�2St�y��+''�@��Iv
�.?NbYp��DP��}�'{���#Q��jlyj���a�T����	e>�Ѐ"Ȏ`��`�"Ň�)Ծ����0�I5o�Q�������7JRN8�e	�eǂ��6�xb �R���	����2���U�`ʇ�S�zr���U��>a�&3�S�OD���əd�HaydڈҎ��ٴq�<�<E�4g��	̲֔�� Ff�����rQ��b	�'��E�@-%̝��ဳ7��!�>1��-�S�S }z���d��)'�����7_f�OL�������d*x�h�@D�w��"fĴxd�	�#Q�"}�ダN[Z�Y#��m�:py���Ц��I+�S�O:	d�Mx:���B$�$���'G���3��_��Pб倊2�|�	�'i�q��ެkz� �f�ɟ*�5��'��Mr��1άx��
���fC䉩}'��#c��75p��ܔ6UB�I�9j��jB�TQ�Ʈ�%}�C�IJJ��" ,ޛj�����܎1M~C䉔M/��!��en�Q����7��B䉽.�f(�i�� f�1ϔ��\C��:%���,9U�l�0ā�1n? C�	�4�����OӒ&������4O�DC�I���]���FH|R�D;5�pB�I�5�J �P&^����F ;�C�
Y8�h����5���"��)V �B�I�!h�hy��]� ŀE��H�fݪB�ɦi�l�`"��hxE��ޠ�TB�z�5���0P�ȤG	��C�I�6������e2���ؤp�C�Ʌc 0��e�4z���Kw�՚ڠC�I5PJ@��mR�d����9JXC�	�o)�))�NN X�`@ �-�PC�	�8u��H�T?Z���Фn��C�ɞqT�<�V(͓r�^�xU*O2	R�C�I;F�<q�en�5 @h�#2��C䉗b���;I��VzPq��M�|C�əJZ�����|�T��d͆�fC�	=Z�!�q�_&.xj�hʀR0C�I#��Y�ecڰyXr�((2RB�I<�f!��X�.֍؁�V�BHB�	+S�nhQW�9�! ��'oFB�#L�-B�
5i��a�JS%cA���@�L�[3���H�ٺ���*j !�d��i��I��恪,��I�IA�!���I���B��S�!�%��<x!�_�
�Y�BnΈa�e;�eS�+m!��{���ArJʐ)R�f�a!�$�mn�k�%5���^9�!�dP�# ��tn��I���I�!�$��r��-�V��k]��"�֙�!��8.�楹��B�1Z�|�H�4-�!�DPzN��kA��%k���ǡ׽g!�$ձd��K@�Z6D:D��r`kZ!�Ą2�9��O\�3rȡ�fE!�� ��E�e$�a��^:��ҵ"O\U��F�Y~�PO�#�
U�"O�0j��A:���1O��}C%"O�����
 m�AME��"	�"O�iqSaũq�@U���)x,�3�"O��6�P�.ABQbդ��|P�+"O�(҆_�Ъ�c��I�V"OT��6�1oy��ȌL�(��P"O��J��\�2k�MySВY�J쒧"O���'{f���M�7��@1�"O��;�� 9��Y�>�8E"O�	�`%�
[o����Vr��h"O>���ΓA��P�b�Rp0"O`�d!E[��+�E� 	��"OtP���t	��JE�P!yޘ��`"O�Ҧ�ڀС`� �5��舑"O���D�A"pU�`*�_Z����"O��E�b.�܈O�7<��@P0"Ol}��&��I�2��у0��� "O��c^�E E��SRh{���y���P�رRǆH�
U0`���?�yX28-HlpA���*�#���yb��.0}&�^�J"d8�J>�y"�_�\ �% BU���
����y2!��L2��`�\�ZQ0ԅ�kW$T�QJWC/��8w��qҌa�ȓ5��+�*Ј]����b_�hԚ�ȓ6/R;dB�]�zH)�,384B�I�v���0�"�>jV����G�"B�I�a����/S~rħV�B~8B䉸(~�u����)c� �Oc6tC��.k���ф�+h�:�{�*C�ywJC�	�`D 4s�(V�	�L�b"O��J�f��Av��f�I*:��|��"O6}�!����ȱ����9!ft=@R"O���/�<g���Ui�+a�4�"O�(�5jǂ^w>�2��)5J&4C�"O��{w�B3.Ȣ7�Ša��	��"O���TIٸ���!�,��V��"O"*N��N�A�!N�m��C�"O�y ���_��y�`@�%xc�"O}��̌,� �鄀ۄ+�dE�V"O�X��0�L��.�9��1��"O��@ ��M.�1��n�S����"O@ �� 4�ƴ�� E�bP��"O�ah�@�$o��ԫ��1��ij"Oz�a1"δ���
�ʜ��U2�"O�;���(�αS$iФF�.H�e"O��i�]�h�!��*J�d��p�c"O\@9������HKZ P�Bp�"O�� ' �����S+o��`"O} ��	%��d V���0}n@�3"O��C�C;HA��N+w�VQ��"O"l"�.�a6���5�L���Ԁ�"Ol���o�L]Jx`
��E��ؚ�"OxS��<J�-���ձ�l�hv"O�Ą���[E�L�"OPir�%�_��e�Q�CaP	��"O^P#q�|�r(Z�ˇ#l	rX� "ODqc�x�6���Z��4[�"O���ϔz3r[EG�[�P"O�7iJ�no�fj���.��"Ot�D�Ja�1�ө��5_ A�"O,\�@'=�����׭PD��bC"O� |Y���	]j���F�)b���"O�<�W��T����"zQ��؇"O$<j�/��]x���A�I
s"O.���Z��4˵C�;�BE��"O��r(��|-�F�èe��$ �"O�P����8����O̹�B 0"O�}��BŠ}v��8d��tB���"Of�A咝0tr�P�ְQnD(v"O�5	�O�D'ݣ6A�La*(Y�"O�9��@ (%������&Z@��"O�d�1����gڤudʵ4"O�4{���<Kv99v�фaSV���"O��Cv��)mEJ;o"H�z\��"O��Xe:f8���;]^�IS��N�<A�=>,<�2��C^���UN�<�chѨ-⨡Jce\�N����fW~�<��K�\���n�?�����y�<�dh��5b��F�Z�[v��	�w�<��!J3M[ h*wcaD%>� ��d�@�	�3^w�L��˝;��H����|8�,;V��]� �� 0̕��X�����IA��(;�#R�z⨇�$F~�[U��!2�4y��ИMd�@��1sv��Q��0W�v�@6fļQY�Նȓf�R%P..�b�v$۸F\���ȓVx ���a9H�Y���\x�]�ȓd��P����~�P bТp.q��``�B-�]��r7(��s����ȓ8�0���ݵV�J,�2
>$�Y�'��~�
K<LY� ��W	�x���O��y�M� >M�%�w_0ղEe��y2�b\�f.F2N�E����m��C�	�b"�}��ឍp��$��ή.7B�ɴ/�Z,��Ȣ��0x���<HB�	�C�8�@=-.d����Z�qe6B�I7�@|��cW�nq`dc&�����B��/u�����$0�.N�lA���[�<i�☒w;�}@4 �z�>8�Qd�[�<��G� ��ܑ%�;&����eW�<٧�� h��CWEm�r��C�S�<ٓˉo�Ly�Vn� �5Ȇj�i�<1�>]% �PO
�u�2U��A�d�<)����&c
�2摀��k "�d�<!�c�?�� % =�:<�g�{�<�u�Vv��R�E�Zv�����Q�<I��K�c���J��٢Akz���*VL�<���үJ7�Q�c
�w$b�����F�<���Q��R3B��*g0`����l�<A�FI�~�")��f��I;��$�Hi�<	��)CbI��O��U��Y���d�<�b吧� @S��i9�};�Qi�<yW�dt����C�x��Ass
�g�<�c��M�L+�!_9�ys��c�<a-��IX�8���=&�qc�
�c�<�tj=k�ĕ�w�D�<��fC�b�<�&k L�0ԀS�ӽq60��vBMT�<i��N�h��hQ���K>Ś'M�v�<a���
4��z��\32[ Pd(FW�<�V�J��L`����s���U�O�<��D�`��	��pڲ` �Yc�<��
Wސ�Y%B�7[V�Г��y�<� FZ!	�goM�:�����\q�<р�^�'��h�)8��zЍd�<ٱ�D�R�X[F[,da庑��]�<� �SV#�"�*��փ4��b"O
�����|�dEj���H.�DpV"O�E+��D�FR��Qh��\/�xd"O�@���K�(��0IR%�+h|J�"O24#���(g��  �=�L�p"O�dh�(*�re�\>k��"O��&�)�(�B��I�"O�%zV ��4���B�*H����C"O��1s�G�x�<s��Š�$I�d"O&UivE�8����"��T檬�"O~�B�����jݺ�p'"OV��r�b��-�f*�=�p�"O�$ V�̩�r��cD�[�PMj�"O$������l�X�BQ�{��4�'"Ov}3��;i��x��{u���"Ob P��m0ܘ���C�8N�9�"O�V՟�^��5�1y�PͰ�"O􅠇A�������1��"1"O���1�9st���%��"O�	j֍S�Tr��,�2�Yy�"Od�ńG8_ȴ��	~�y+�"O�0��H�
P�V��V�]�P<�3"OH�K��U�K�����l� �H(�"O�P3d�51D������ I��Q"O~�sΐ�[�1��A�0=���"O��5�K"5&�:��5`���"Ot��Ĩ	4p�X����h�tU��"O����   ��   d  �  �#  0.  V8  C  �N  {W  �]  4d  �k  �t  �{  ׁ  �  ]�  ��  ��  <�  �  ��  �  F�  ��  ��  �  T�  ��  ��  �  [�  ��  �  ��  �  ^ � f! �' �- �6 �< D �J �P W �^  `� u�	����ZviC�'lj\�0�Iz+��D��g�2T@���O�6�M���lc"�¥�V���E�q\I����:&p�\C�
4��ӛgή�#�_
�@�Xw_����O�N�r�O)<4`�MƐHhXi"!j|����CmX�|�|К1�],dD^��Ǐ�.3�qs�nݽ�Ն]�?�r۴p�z���J�����7Xúy�I�\��б�'���xRB�.8e��2��iӚ2@<ON���O����OB����m3�-A�M8��D���O ��ح$L�oXyB�'����f�Oar�'��i��G
T��� C��0�y`�'��'���'u��'<�\wK��p���j�eh��HtԆؓ���/?�64�JL.�	\�D�(Q�P� ��\{l(bo��<G��5�T���'��5�d��<��٨/+��RD>���1���Z�K͹y����*�?a��?���?����?q���i��#G� �K��@k�F�#V�ZHKu��O~�oZ �M�u�i��7��O<�oھp��<)�4;�@X�3앝w0$|�VM߼v{ʥ�耓+�8Q��iU6M�O@��{"�?+�H~\@ @�@���z4��	˱;��p =jX[��O@o���MC����T�OP�kgV�:rP1=dqЇ�s��7��
zJ� �tG=j�v�I�5�.�t�F szTlZ7�M�½i��xX׀N}
�/\�u:���u�$s�Zy��QvT�7MTڦ��۴^�E
��;�`�S���kt�� �2vA��s�ʹQ ��YQ ��&���2;�ypR�i�6m�Ԧ)���[�"h�(��������_6��$�]2f ��lN̜��4l�R�F��R�j�!�i͚E��L�����'��!�\�`������N�Y1�'�ON���O���ۦ%�O�"�J���a����7�9"�(�Z����O��D�OTY@p��^L���6!
�r��͛�xl@���(N����D�.ͦ��Ԁ�F�Q�dH��(�ѳ�@H�.�(��GT<{&�y����:^Ed�C"i��BKJQ�t��=uQ���S'�<rY�Hq�`�*	�p�{ዖ�\�������OB���O&�O:���O^˓�?�TNB�6��IpJ�H��Y�iF�?��q.^���������|ڦ�'���x��Q�s/��/��
���D�d!�0oß��j�w^V9�b
Z�x����?$������?)��ʡ�&aB#L�6H2V� 3IGi�� � id�$�Ou�
�B I�]v��c��4{��	�-�"�a��:]��9Ȱ��=\}Ƚ�M�V�' �� TЩ?p�9��	�+N��'z�8��rT�)%�'��� ��Y^"h��m��ؤ
� ���?Q���?�����Z��]qA��n��c'K<h{ў����M�G�i��'�=�։��dJ��x���
4%.\�W�q� �D�<Q�J�������?�����S���L ��Yq��Q�CI  $kpi��P;:�@T��8�"�A2�|z��mF<�+�DC?A�[6A1f4S�P�X\ 4K�,.,Z�:'��>
}3��7@��`�|WÏ�t��	�q�h��#�;����Ԩ�&7d�n���\�F���O��3����p؊���M�Ţ�
H�ۢ��$�S�O8����+�:u���2�h[�j#���'�R�mӘ�oZJ�i>5�my��[��� ke�àP��� ,s��}�ah�>���?Q,O�˧���I�u���g��Z2&��T��2I 4�:;-^-��eb@����"M*{��Fy���<沽�0���@� �6�L0d퐐��NX8>��JG�
Z� �2�	I!a�Z=FyR�գ(���%ȝ�W'��!��Z6������V�0ғ��'����M�>cs8]9`o����@�'���'�ў��<��L��	sp���	b�
��j�ɶ�M�Ƶi&�	�x���4�?�'����@�/jRN,@fB]�_�:�������O|��v>�m�8jn@�,y���!V j�<]�N�~_l��A�3=t����ߨ,N<�<��J)� ���ػ
d4!æ�ҵO���q`�:4�̓Faט3F�`�G��(n�	� �]���o���I�M�ļi��j��O.�ƅÁ �@���J?g��٦������?�}��\w�>9{���p�d��Lr�����?A*��Io�*��eB3��
A2�p$�иd��jٴ�?Qӹit��)�tM��	AY������M���J|�q��/`>$b�h�*.��9���?�����4���a��a|4��ɓ�\P��>��Gn�4^ ��`d��7�y'�^~2��O��x�dD�	�=�7-(tF,�@d� OX���O{���Չ�Bx%R��2Ce����O�4J��'��6�Wq�S^̧QG�a�r� �A�Z�a���4�$�P��^�I����Wy�	w�����#�,�1 �
�N�#?�$�')�v�'�6��OJ�Kf���1p��@VяUo6��G\�����fyB������'���'�	��5�7"Y�<�. �#)׮-�"	
(�MJJQ��H�=-�h���m�x�D�O�~��vm��~�2(��M�f��B�^�0��ƃ]d�)�Q/�-I,�I�jV	<�E&�(��S+mK>, 3F��AR� �"5�4��&n�
Q�$�r�q���'�P�:��٘�?���?�bh҅k��� ~,cAr�z!J��|�)�S{<6ujd��|w��*ׅ#����O�@o��M�M>��'��/Otģ�%�8�H#�"��@�@]
�oџ�	��'I�S�|r1��C���2Nя	)� �0Q��Mzw�[1I�Tɑ�
��8�V�:�j�9C�d�<9V
(Ah�{e��`h�#ѧ��~�8�� ��Z�����% x�B�aL>a�I
�����<b�y:���w���K�I#D�,r�ڟxb�4葞�Dx��Ҭ~�TE3�O��jЌ�yd�B��?qO>���?�/O��O�a��9^�Fxi��R-U,�� �O2�oȟx�ܴH�F]>툵�	'�M����?Y�^Ĵ9��l��w��I��L��?a�>.Jm���?ٞO�r� $َF��m���YHH`�� �iWέ.�r������=_p��땶A�2`���Dɮ ��5�cj�;��7-٨A�(Ȫ��� @�ѫ�$#kW���
�,*���3�& ,�O��3�'D2���Y"��^Z�tj�2*��x3pe4���O���Dv��$���Q�`g-&��O�=ͧ6-r! �'!3�*ܚ3�L��1nc����$ۧ!�|�D�OL�d�|�2$�+�?��)9<բ'��1����` �?��r�X�
$8Р!Y�$�3
^<�t��by�ȟ����H��8�����%\+@(Ӳ��Њ@oR}��Q'�S�,����E@^ �=�gmR3*�����KK�8#�0gW5v70�rF�I⟨F��9OLu��F�>,~D���A�5R��af"OZ�2��,,f�E�qf<3.8y��۟�8��dق*�IS���VzU��++�(lZ��T�'����C�O�B�'�R^��#����7�D9��`�I j��Q8���L�-� ��C%bܢ4�O��
?���O?�E$�'y�4*b��
+�p���l*�9	�AI�#~`	SE��V0(����%-�2cB6�hdY�K�U�K��q|�H�B�fӾ<�'uȈ����Ο�'��j�V�~�d��SK�V���'�"]�(�IA�'��$RA���S!L����(g���R���'�B7�Oզ�����M�-�>��|
�d��u��P�3���l�* ��&vn�r��D��?q���?��5����O<�dg>��rm��3�\�R��`5g-�qF^K�)�55�HۓJfڡBa꛵kJ�)K�nMP	�l�U(U�#��劥ӪC�a{d�?Oq&t�s���3�f�Y���)	>D���?����*e�*�	�f|��YD�(��|��/A��X�/,7âe �	�&=�h�$���ڴ�?Q)O*��7K�W�g�R���˖�<a�!��1 ���<���?���*0�f�B[�:S0�$mHl�J��K�ò��A�aS���� ������F�'������V5T��Qa4�L���F�l(��Rf�hP躲��.|h��R`�-*��u�|" 0�?�������;:Bt]�f�+`�6�T8V��J>Y���0=�)'u��+�!lu"3ʄM���hO�)�A"�߾d�$Ls��:|$)@�	�ON�E8�l ��i��O�����p�ډp����qƇ�D�a��j���4��K$�T>s�F����B�@A����=p�H�#b5#�*�D�L�SB��]��H�O=C��@^~�RRL6Vj�an�0cJ��5$�-%�������2�mT�1p������	���)5c��$���){��iq>iyb��7��l{ө��e��@ׅ0�	p���S29FJAjCC}���v&L��=A�-���o`��OJ�̛ۗ�Τ��1l�
eaE���}�I�h�ɬ ��iȒ����	̟���ݼ�&FG�r�
��Kȇ=r\��->�"�xl�P�u#��9;���Y�c>���T�*��"q��u��eِ34q�P�w�R��R=6X!R�U�؆� u�I�<1�Tiq�'���:fn�o���:�e�WCb�2�������B�'�ў3���,@��iqpK�?u��!��R�<I��=мzPfC�w�Fc!b	Gy>��|����KChɫ����;'D�1%	h�@v&��[7<���O����Oj���O��v>a5�۽p��!@��G�$�#`a--�*�7/�tI5G��%c�D�A,�G�Q� ���T�,��w�Ӛs�d��B2H#�`B�*ߛX�(�Y�	�+�°�'�E�c��m��I�B�=b��ݛ4G߬c�.Iӷ�IA�T!� �O���4ړ�O��T�U�*�q@d�70�%�'�'B1Ob�*�CԖK��<2��R �x낚|$mӀ��<�p�'"h���'��ݕf�ܚ���9vQL��7�2�'�
��'�b9��`�#(K�`4�ZaJ���V���@Y�8
 �ִAw:��C흩SZ@�?q��1[�Faطd(@Ȅ�G�
pD\
R�ȮO��)Fmȸ13��e�'FB����'�*PsR�;�����{s��0
�'���Y��[�ve�8��O4��<k	�iIR�`��ѣ ��*"�bӷDM���y��ۣ�i,��']哥u���I�erQT�X�|�@�KI61��5�	ȟ� �NِC���"`3	�9iW	��j�y	�v�t���U�&�����H��i&��$^��E�Y����v��1�M�g�>3z(��O?	�֦	�@.��Hg�_5^���ôh3?��Θ����Ij�O��[?;.���"�V(�۷�ħ�!��$J4m����8���i7��j�џ�+��I4�lpY�O �\�x�gA
kV�6-�O��D�O�%�ڬ;e����O>���O�睑K�
��$��Da�iJ��@�6T��E�7��D��o��Q��d� z�d0a���Kn�K�Z�ڈȕ�K6��y�F��2�\�$��+Fnʓ7f�"��8����]�����l~R��;�?����hO�����8� �EO+^
l�+�=D�4�!�4	�$+Ύ;X�x�O�<ad�i>��IMybk"JJ�ܪlV�VH�Q;w��>�6ዧ�P6,���'j��'��������|B�iP(~>�y;��[]�r�3�,��|��0��CV� �Ih&,Ӯ4����HR��<Õw�? M{�؆8f<�"!o�)K�L@���� ~�Uar��0��QI	_��z�gԎ	ғO��z�焘@㢍��cB*�M�Ѣ̛F5��'�b�d>�'=�Д�B��Dܙ;�'0?��P��	x̓,mTU�!��<Ri�x��(�e���%��;ڴ�?�+O�E�p��Ѧ5�	ԟ)ҨΪ!rz}�� <%�L��b̟��ɴ8���ΟH��*�����$��}�1Ѝ����M�$'D�rB�X��(�H���7H5ބ ��9ʓ0%r[���/����E��q\8��tk�7.&�!��
��ĉ������iB]Q%�|�C̄�?�`�ip�ɢUf<yi�E�)?�,�	��Q?(�O�?�# `?	w#ݮ6?B�[pJm��u�}��hO�iA���+RN��XZ���%�~�:�vL�O�4sb>O̉����!�I����O�܄R��'ݰ�qGL�-N���s�a��S��H��'�b&Q}��:d��E�r`8����t�Tez�FF�d��SpC��G�OI��g��>D�n�'�J����N�lIa@�M�]�~4y�O�n�]z\GY���M�,�S'�U�NP"�Ȇ*F#����� N�)§HQty��$}�ő�ߵVF�ą�M�4��!�,+����� ��G{"�'C�#=�,�v��%���n�AЏ&ț��'�2�'u��h���2�']R�'��N�?�$@ShׄO���#�?}�(����Ol}")��+v"i���y,����58�
_�M氘��a��c�>���ZP��|�<a��+�>}¦f�`�RM`��ݟ(�'�x����?��+A�nP��OY#Tnv�2p&�Y�`B�	�):2�#�Ԕ[v���C���˓,������'k��3��}�J�Ue��U�d7�� l�7��O����O�˓��b>��b�.���P�R�2�x�YEI��y�@�sH�=?U��c���`���$���Q�H"s��Mh��u�Sm�d�ဌ�k�JM��&?TGd�s����*���K؄zR!2�d�{JQ�f�oKB���Ֆz,��e��O&$m�HO�"<	����u"|�(�mҦhapH���Ig���񑁞�E�h��N6��%����4vg��]�$�b����Mk���?�c%�+|���v
�{�ڕQF�4�?A��iG�����?�O�H(�B\�J�����.1�hs�oXMdh�Q'�չ{���Y�/ԡ�ZAp�`�B�'^p�)��1L���p����*�Z��t,B2Z6�0)\D����+��B��Ȁ0����0G�|B㞒�?����$�?$3��k3E|�����[;zn�'���'�� A�ԥ2B�z�`HKل�ً�i>����=���9'��H�1n��	VyBn�(��6��O$���|
7 ��?0 @�L�!��DJ�V���X�:�?��Rb|vI��R_`�� ��K����Ƃ�l�aQΟ�IS�ڠ��F
A%B��@�C��T�j�|��Y��#�" ��������ѧ�40��:InD`��/�8'�m���v���rM\%��џ�E���' �]{�f�X�X�@�30�FTs�"Ot�PQ�ٺr�����e�H`s�I̟h����D�7�؁�%͡%lD�����*l���D��ǟ`[aMTD����̟�	�D�;B[��� F�n��D)H�`s��A3c���GjZ�Z$C%G@̧m�Z�
ց��<RVh��Zt2��Hb%���S:u��`��	ɼ����&�L��#ŮNE�4�_�j��7=����1R�d��Bh�&����'���'�L�(sݬXcs��%J���'E�t	S�F9X��"���_m@<����?it�i>}%�d��I�z� � I
5ڒ�A�hd�|��Fʟ@�	��D���?��	П�Χ@h�2o	
e�5�����1lӠ3��k�DN�^�<�$�!*���3��G��(O�Ȼ!�k��1��E�`����	P+��˄h]�3CVTB�F�:{�4)	�咧{�>-qЂ)�R�{� ��u�_2\�+gF�'���"��'���[�'	�� �f{��#�۞kD�	���'���*�K�X���ҴeV�g?��YI>)C�i�2S�Dx�C��I̟�z)��%�2�hq��)< �M�c���(�I�aiƨ������ɦ��:�dƱT|y��E5�y�
	�0�X&�_�>�:��ƌ�m�ĩ��+a��u9gO�-P̊�F�_�O�H`2�x�ʡr���hW0��$��!s��wӎ��'�p��%�����W� �U����?������i%?�B)?K�|�vAD2��m@��Gk̓�hO哔�Mcᎌe��UI�!�"LS2
�Y��X����˔"�M���?�-����O�O��t*O;`RJ�0���z^�p9���O2��V�TȮ<��Ǉ�s���¯O�ST�ԉESen����̉�Q�^0��䛌-E  �e5F�5E�DW*T�DY���B�� �4���	6��'d�>A�/�:�b�,Y����`$�4��p��p���3�G�cД!������E��1ڧ=�Z�k�d�@c����æG�68�۴�?����?�!�$�������?���?a�w�����tF�9q3"��KW�I��Z�
���9fn���K�t�g̓3) qs�˴-���R&Ȥ-v���Y	 ����b�":x�8J1d�ȩ
j�*O� %І�8�36\t��'*�ɣm0���O<�=�@`�F�0�s�D�t�i�	@%�yb��6�0paN�68PcD�ؿ��$�{���$�'��	p�%1aOF7f��p+��K��l�
3s�~4�	ğ`��� ;Yw��'x�i�3v�x!���B�<�豠CEu�9�g��}O��Bf�T؞J���Y��&[l�<����(;;�̰�b�}#p���UX�ʃ�A/p�N=���/�\I�,Uן<��^�'}��yV+h�5� S���-��/D�@��F �u1�����P�3��	.�$�ަ��IZy��,k�6M<ʂ�E�{\�⨜X�Y�~���<����?Q�O�jP�Ď#S�Ć��5<dm12���D˖�j�\�'�V�ː(��H�'��s�'�R��ѝ7��p�冈�
H��*�3`�Йa���(�%3�NS�q��8;��Ą-��Q�|��Ą�?�f�i���DN㤏W�|`1�%oI�p'�D{��$J
T�r�A�&ݮ�&���ƒI��OҢ=�'D�&��*�؝�cKl_�C�5�掭�M(O�,A��IЦ�����D�Oq
!���'���׮��M3�l�E�$+e�TH��'�2�iЮ� C"�^�է�,�Bo���[���*r`�0I�G�f~�B��g�@��}ΖHj�P�@�\�֙�t`�%G�R�`���u�,��[��od,�����S�Oo��ò�X�QSQ�"&%��
�'6l)C�Dg���Jѣ/���Bl�O��
�`��N�
�I�`:37T�9$�ic��'"����j�9��'���'�b8�v�j4)�x�6���O^?u֩�P`C9q�r����'�t!��v�3�3�|�Ƨ�"4��w)K:%~@L��Q��qD\$k����2��X̧Y�\$+)O.��1.SA��"�K�.�ȱ���r�^�m�П�V���T�|�'^���:ږ�A�|��,�_0��)�'m)��
�52��А�
�/� ��/O6an� �M�J>�����.O
%�䌂)J�ŒG��@J�[�$��7�O��$�O������D�O�擒l��t�1�<�Fq:�޹�Fp����������L�<S"7�Q�}8�e4�?�I���ԚR�!�a�l`뛞m.�����N�mڟ6)��r +!�b$�|RK��� � �<��<����(~D���?i��d)�@ĉ��Y��x{�/ܢ H0��	v�x�h�X�`�=�"|yQ�W�<T
�&����4�?�-O���3%Dt�4�'r�y!�M�ml6��f&��1ⅪC�'��F�jw�'��	��Wj���� @>�'�.���@�2�Щ(�&�C��Ó.e�0�gH��i�Z���dC�Cy"��hۑx*�{�e4O<�c�'�r���-�ܤ��aР�[J܂W�ҒO�����H9�4C$�ʇL��܋%�g���<���T>��: �	�RI��rA���U�-Y�0��vyR�'�26M)���|��aʜ#!b�*|N��� 	NCh@���?Q�A�)=� �'
�+h@R!��4��L$:B�D�ؘ<�5�:%��0���`8%m@'B.�a@�ms0Ԕ(E哒6O��ڤ,@�%I$�0��\��$I�|�	�MK�����'z��5�<T��h��0�3%�2A[��HÔ|�'iaz����,����#`�;<��zHF��hO`��TA}r�IY�?�.�-�1yJ�B7E��Uu�����B�K���I�O����Oʓs\������Q@�`pI>¤<
���<l�������6������+��O��'�~��רֱ�m��$f�,@P�S�K���;RgЛN���J��O��'~ }aj@)5nű�OĐQ�"M���D_�!���'����]
v���WRd�d� 5��C�I�ZѪaӗ��g`l��!
4�����O�Gzʟʓ)����Ą9��8�i�&2�����8}M��'�b�'K�)�Ӗ&� UB!��-7ʩyg�6z=���J^">`��q!VL8�-���_���O.tbEL�b_d)�B�ֵL�V�{���
PT)��*k���Ս��}�H�?I`�\\�6��u�@��,�e�y��	��`�Iq������'Ņ�6�$ݛc+�f�I��'�1O�d+�^�M�l$xG�G�:,PԐ|��>�(O�5c��A�S,\��] &�Ɍ$~�����&��$�<a���?��xDFA񥄗q��B���9ޔɃD���t�p#)I�.�E�\
hџ|Z�Fϖ���1ۄE	���aH~Ӡ��e/+�S�1Q�dDBF�=�?)�����X�`�S��	vq~t2�ʍ��'d��'r����@$>D@S!��PK&X��i>�A��_&�a�"S�������cyP�Ixy�獊M��S��S>e�I�k�	;���gJ���䤒�#X���锢Tz"je_:P|��C�'���O�բ6̅$d���0k��:nFh��O��_3_i@0�/�J�Xq1�j=��1�ԼJ0�L(�$��!#�#,���;S�M�IF���'m� �����LE�5�%�	/>]�S�"O�x��%�N���
'/�|R>K0�̟����*?��L��(��Seo��s�>�n�<�';���Q>�<��B�U�vDh�h�_.y9�JEY�|s���ɚ9��hB���[H}c�mȴ�b�` �$LOX�A���=$�F�p��TFj�A�'�T@B����y����c���l�цC �,!�$Jv�q"�ʜ)a�ř1� +`��I#�HO>��
��R�~E{4��_�T�Ƌ ʐ�#�4�?)���?�(O1��)u�a�����Rx����+Mp�.)�r`��hX����'`���L�,]:2��A�
)�I�`�C��P�$�_�Xy(5��;;Ԙ�+��Z��٣�NɈH��,����O|�mZ��MC�ҡ>�;2Nh8��Y���P�d�d�$C�I�kP$|)V�@�, h�dL |�O���'�剕:b�(۴��iР�ড�!A ��%o!��'����$I\��*@?z�P9�7� c�ax�G��O���9;�mz��<�v�P�'Z�����ј'(�Y�%��L�KD&�8�D��'�\eha ۂOD�:�D	h\~����F4��F`��'�8kr�\�u$ܖ��a��\7L�'����?��H� *� yG.�.m
����	�_�Z���s�ʵ��*��?E��[>g��)h�Ǐ�t;2��U���E���;��<��Ђj>�'�h���ԳGzB�2V ��.&f(�'��J��?���)y������~Zjp�rjǄb�ȵ�5�1D��bGG��(���@�^��myAi=��^�>u�%��aSdT�cAL�L��D@Q`�Ob���J�<�e�ր�?����?����ę#kt�8Q�͟�9k����次��#�s� ���+IZ��b,7�3扙A^��Xӎ�|�`̡cIYx��eA���a�Ɉ�F���M6�3��&���Aa �� �t(V�h0�6?i�P䟨�I`�'����`*��DY���&4ct@�["O
�+�#�?����p��,�"��dX�����?Q�'5@%� I!�=�e;b��%P��i"՗'��5?O�M@���6���\0���;L\�����Y2]Q��8`�����b)0���?��#Hae�^fsri�A��>�'	�^x�'Y) S�`�`��<A̰D|"�іL,�Sfb��."�l����,w&QAL�?ٶA��h���bV.�-�ў�
���OF�d �$8F��
tÌ�l��*���#?���0?� ���5��q�'ghw�q:�QXx���(O�)k#��8jm�W��\U�pS�l3Q��͟D��ߟH�O1�<�'>"#�O;x��D��/)v`p5�(K���wmRAsp��q���d�i�d)�Ϋh@Pb>����B�m��X��_7.�peKg�v�d��OD�K!$��.�-DV�7MSV����g�M�T2�Y�-�Ƒ��dΊ}���cw�\I8�0O�؇�'5�������;Sҩ�r�H	|$xau	r/vh�ȓP�D��
�>
�9�g����?�� ^����q"M����`S���  �1N��ݟt��q�q�F���h�	��<�	�?��,.����d�6̮�0!)��-��|��ĉ�.%����LH������o�deԈ$I��O�S2�׊@�d�4��s"�M��#%%���G�P�C.�xAդ]'+6��'q��i�X�L�~`�;)�&�8PHťj\�9�Dሥy�0��'ҋHڟ���R�'L�䅚>z�!�H�d������oE���<-�0ae��XT.qk���v?��d�|�����'���"u�ޔ+���*\:b��3�Z�t��b��������џ��� #^w�b�'�󉋌q�V�:C�T��f��t�F(���)Th��"�[q؞�:GͫMb��ÊEк0"��N���#bfZ�*�zhXۓ~G���Ƀ_�F���>kh�Z���)D��I��d�'��̂��� �h�n��`�k�4Ov�=	\5��(Ҭ�N�ʐ��@ �l���M����2.Pf�O�9���Ү�8=A��s
B�4�ĩ:!�'�Z5���'�2�'bv�
a(X�+#�=��,N �
��B��+����q�Y5X�z�/<bv�(j�nD��(O�J�GT.H��h��	�V:(B��*c(p�A����ɴ���&Y$5�q�ό*T��R�.2�D�*U��'�1��ݪď�F\r̘1� *6�U��_�$�Ih�����&�[1%=t�	b��{�|�����<�ӏO�Q����掄9I�%C�c`y���9�6�O��$�|�0鄴�?���n' ��E/�pC�0�g� &Ԝ���V�Xs�� �K� I�ǀ]@ \b�)M�J*���/73�(���<>v	��y���z4:X6,!��]�r�:`���j�*��*jܗO�$���!��dC�k� 뮬!�'����?��O�OTb2O� n���ڂS�@Iz���H�F�@"O��hg�T�5ظ$i��*�TqF�D�O6�Dz�O�pl���2���ɢ������'���'W��x�.�6�R�'�r�'��֝��b��"9(��&��Y�f�ȣF����z�6$Y��W>^���O�B��!�t���;�е�J� ��!!�R}�����Q#�.ڡH�27�]�&*�|���Q� t��G󼋡���2(��L��vP�&)'}ba���?1��?ɍ<�����݆&��ؙ�11.�A�O�y�w �$|I �G"3)�y8P�O,�Ez�O��R��yC.�c(�����VDոl���%C���O6���OP���?�����4�޺`�����e9+[\-�T�W3C�u �CªK:����C��|rx�'�
S�Gy2@B,UZ1�R!�3x�89�vO�K�x+����sB���9_��� �O��F�Gyr	��?9Un ���HSl�c�:,�P̨�?Q��$%�`.��9������r'T�����<R�Q�"�%�F�:�m����}�'�h7�O<�8r�U�i�r�'7���.5���%5�������R� �(o��'r m�5�͌-�p)�'>hqTd��'�#M���
��R�s�HB���sװ������#Lݠ$&^�Wf"���A�|��,F�e<T2#d�	~x���Y~��xXSF;,H�O�hX�'�J�?��b�&w����
$%��|��e5D����C�Y`ո��U���:'�=�$0��|��T�h��^�����P/>zd��ǵ<)��?a����ĩ|�ɟF���
��f���ʭsvQ�W��̓�?��O��S�'<�N$���
x��؀	9�?1�4�ē8� $FB4�8���͹F ��SDbB�9��'���w�H��I���S۟@ϓV�����b��d/�i�+۱\y����U�Mk��!}p%)���y"Ʌ�������3�?�Xa2���3%�^�J�#�KW�5h"%��'
r���Z���s��Iϟ���͓$��X8��"�ڼ�Si�a:=K�hH������<�d8���<)�nknz�-�'J%
��%
F���Ph�4����'\���?�&��?��ȟ����?m�	�jD�F$M�a*΄:% �,��{��oL�����l���C��@�c#�x���]��u��P�UI(]k@��vp�'� �M�'	v	����?��w�d�'2��O_V=���=d��] �ƞ_���%�!O��D�2���'K��]��Γwx��m��Y�J��4�'NЩ���1�\3Z`�=��4�yr#4y�F�}ӚMB��Oh�]�?���Kd��(�� +g��ě�ǣ���ܴgN�k�'��h���?!���?��'8��I�Oe�ɱ-�]A"�=L���-DD3�40�,����$��?1o����,O��Û�1�	��6e$��ʂd ���"ORe(C��|p~ �b�V��4���i&r�|B�~�/O�'7��Qt��4�~���[�J��|��X�(%��F{��Ov�1�hB�s�]{n]�%�q��)��<ʓ.Ql,KT)�aK��ſF9Gz"�'�����+�>[�و��iBb���'��9P����5{�Ol$h�
�'���B�eu���q��!v�PIK	�'a�1�2�T�x�"�j�`�x�K�'}��c�`�@��)��kC�\�B�R�'D��:.w��PJ�FI��9
�'�p�T߯=4	�w	R�i�2%r	�'QP�B�`�h���q��q	�'QJU��j_'n���a �%=�M�����O>�D�O&���O�P�e��_^�*ch��)����]������џ8�������@�����A$ւ�&�'�/GL,��Ƅ��M���?����?���?9��?����?a���9�n\	�`O�L|X�J%͛��'D��'n�'6��'$R�'T��~��
�G�<F���а6-�OJ�D�Ob�d�O��D�ON�D�O\�dX3He�e"��ĵ��ũUIԏV#�mZ����	���؟��IϟT�	�ɾL�=xy�W)_=�hAY��٦��I����I�0�Iן����(�Iҟhi!��5se YfʷK4ƌ�ɛ�M���?���?����?����?���?1f�+q��h���u{�Yb�Z�
F���'6��'���'��'"�'�2A� isf}�V!@�Oqx|;��E�p�6�O ���O���O����O����O
�D�,0���䋱"��иpaM[v%lZٟh��ӟ��	��`�Iٟ��I՟��Zpڤ��73��@A�Z��a�ش�?���?����?Q��?9���?1��F�@��A�G��@U/M�6�!q�i���'���'_B�'A"�'���'Ӕ<r�ӥG�ƈ���\/F2�I (x����?�,O:#~� �,"5�&�G	U��I���M!�d̓��Os�7Mu���V���f>WO�&u�T���M̦�Xڴ�y�Y��&?��g"�����D&�6�]� �j���9e��I�o���������E{�O��Ą7 �H,�&%ڮX-����?lX��$����41т��<	� R<;≜�r��j���'z~�=Bt��{}�)�imZ�<a/���BR��^�p����H#͌��S�P�e�_f�9?�'��	Zw�x��/ap��K�� @e>\����!��˓���O��}�F�6U�4Kخ"�]2�Ӂt� ��	�M[��t~�p����S�3x��#��@�N.QHӄ�;4[�5�I��M�ǹi2C�i��F���H�n�%0Q<-	����
�Chn��G�D�eነ�&��̟�'U1�X���i�0��C��	5�I�Q�p��42O���<���4��|��(&
^)2N�k��[�
��1��a�0�IR�O|��&���Th�	 �i)LhP\�HS L$,;�O���GP:x���=�I>H��}�!!>$�G�$I�Z �ѻnN���A0h��3��0h�"�8.���<Y1��8,��P��G:>N�A�3���#�"�#��O-T�+���� |��
ܜg�tq)ݻ���Aàs��eM�+�:mj"���o��[dӂ[���Y�/С,��9���"g�L)� ��;Y(�G㎗�yR����I��@C��BE
��Z�ҩ���\�{˂�x���*�d�B3.F��X�ȓ�z���KƔ7��±&	@Q0�O����͓-��H@P�լy/T� ���$T �L9�9}��.>;'���1� GDP��=X�z�S3CM:����N� bF($_r��{t��`�'l���)@�6�ػ��C	,��@(�� �z�:����8.t�(����Y��DRT�&LbR���q%IM#O��02A(Ėm7�%P3�ڋ����4.C��?��?a�����2����"��'�^,�Q�])5��ڥ ʆn�@-#��'��'�'�B��7`pP��O�Q�V� 0W���f�ҭֈ	�w�<D�\q��S�I�OT��0�:,O�=nK�����NN�,a���	�' d�R�@���a'�?q������#/��@`�+b��W�-ԍ�! l�ZP�!�%E��m�3�5ܴ�b�ٕ3�)9��
3 '���@K�0b��I�a��YL�TӢCߤ:��|��@��-mN�(FF*x�ˤ�S�_�J� f�*_�Z]`1gߥL�eR�d��'��[o)�����"|���I2���w�8}0��@]��rf�A��͹T��n��p��D�G$,=�5�b�>y�W���(�I!����I�p���h�,�˧ń�Bh����D��3�~�O���'|7��Ŧm�	ٺ�v�S9�$ �
�k���Z?����h�� 9#K��B�c��O�I��,��'�ў�S��~r(�>:���QƂ(ƭze��%��˓LӞ�)��iC2�'C�;�1�	�qA��*cI��z��Ȑ3����T��?����4~����H)~{Lpyߴn�X��cL�f�O�Us� H���p�ŊFԤp��O��iD��W�4�4C	����:��e	��ŗq�x��'Ae�q ��]2lzj )P��N�x��'�a���X�F�f���<ҧ �V5�F�:k�D���k�/S��O���>lO�l�D���=�@����.��S������3��di��#�Y!� �t@i� �0n�.�?Q���?��Y������?���? nfޱ �F�	l���aR�_���ɇ��D�	�'l�"H<	"u.
K����͑���3;���ep�,t:�Ƅ�3�,9`�]`=������!!o�t�/G���I�52�V 0�-���`�Y�=�&��W� �^��-9BN�
L��Wz����M��'�������?i��P���V�`��Pb�C�<	fC�*/e�;Ff�u6����N�`0�	>ғ2�V�'T�I�_%�D9���8e�X�Z�D��d���5Tƽ�I���I�H1��p��k>Y��g�亙`Q��%}av�)���%}}�ջqKU/a^��ƛ"��䣌�DVi�z�	# �0ނH0��]�ǀ
u�� �f�8�!'P���O��1�i�ER�_�|�¬��
�;�� c1O���ڴ�?*O���$��b���Ŭ�n1���\~c����"O�	{��Ŵ#/~X3v���ZRf��G�>��i��\�8C�a�M���?��4Y;����훌0q�����~@�5���'S�qa��'r�';V)H�c�H�Ar�KEE�2&��_1��Q �l��l1�C�0AѢ=�U$V��(O�	��M�Dl���-z�~�P��ہ<��Y����ft�D��f���HR��(O,��E�'�������|Հu0�Ƀ,S��%&_X���O⟢}���@=7��8k4#M�)���X�'�F����'vn�'Hb!�]�``�\�eǠ<Cb �wH�V�'�Z>���ԟ�lZ�My�I�!HԵu	�)#0�L5���Κ�b��/��a��OY�T:��r���O`�*K|�D��j9�®@7a�@%d�e}bN�Ec�8 �I�_��J�U���`�F@�OO�5is�T� ~4���CO��"�2���ş�ش�?)K?uh�X?���7T`y�ք�g2D�p�/}2�'�a{���8�q�F�(��*������O�mگ�M���O�PFJ��H�-z�*�Cu� 8�6��Ox�������Ov�D�O|��A8�yW�K�Z��H��!X9wW6t�Hx<�6I��yZIkD��@	�(+I|�ը�U��ʓ\�;B��!�,���ġL�e�g�M�3w�31+G@*2b�hy�ʧbd��H�nňSy�Ε�N̪(�hF{B���׍X<\��,O��V�'�h7m����nݺ��l��� �8��C&�*!��6z
>���%Ϥ1�,�y�+G):u���HO�I�O,��M�d+��!'����O�>���V��E�<�   P�II4�|��ɜ�G9 �
O��D�7$�X� ��G�n%2q���y��̮'���37왴?�,�������yb��2y�J8�W�F*/ p��B�
<�y��U!���yU�U	@$��l��y�&ALjX)��x\�}!���yF���f��T��{�$�˦G�+�yB��)b�.��P�8{�$���H�'�yT�,�^Tis��K��[��y���>�\�Iw�ĺ�"�B�)���y�Ɣj�Z �X� ƀ��#���y2�����[�y#n��SL�y�R/7M8H뒅B�F�+Ƃ�@u�B��B�`*d�ԢV�4a$m�zF�B��
w��Y��g�,���.ޘ4��C�I.,R���ƭCE�=�3/��C�%��9p�.P欑�W�͜49�C�b�&�pr�m��ICNJ�"hC剝B>b�s /5w���򖂍�`�!�D�j:�j��d��(S&�5�!�D�$vp�����0R&|�j�E��4�!�C:8�j�	��М�T��ɤ�!�\5n\N����1����dC�UX!���Xd<�����p�0cc�$6�!�d]*8�y�Vd�v�l��%']�ԡ�#�'oD1O?�6i����� \�12N(���L)-�C�ɞB�i�IڢP�~�����{8�dY�>��=*E��o��#����tl�ţQ�;-y��,lO|8�'gE ���f�it�R��'=�z�8p,ƣw�8�{�'�`-�f��w�d9����d�dL��{" Y3T5(U�v�Q4q��|
���"y�0�0���m��ŮHa�<�C�Rn��c����vT�XP&�+3��iu�9e/L��fʤF��ODM)��P�|T@`o$,�%�2"Oْ-�AcjPP���$)��b��/��YB�����R��'���	��ڶ#����b�3��؉	�ղ)F�W��m�t��KQ���eOi�Yq�<'pĸ�ªO�<1e���.�0P�	�@Z � �IybM\&�
y�dcA�)R-�q@K&�>�T�،V�pQ��L�r=ĥ�<D�<rSV)��H����}�L�1�K��2h~�JO�[�X�g�����<i�b��n�s�J9�# �>�b���ϮZ�ZPXp�g����V�P��%Xq���n��eI怀6p�C5�Z��y�Gԙx@Ppu	�0S�����O�s�(�<eS6@�"�:q�)1�q��산x�����"  TӅ�04�D��N�3X:����#ğ7r�QjQ�f�8��c�
L3T�!���'�px�wn˱[<�������ֱY��鰣R�<�|2ѧ�y��F8 ��M��Qrِ�
N"55v�{�(ٷM� �07MX/&��:˟z!�1�p�I�Q� "k̀f�|Тf,�8����dŊ:�����e���#v���JL�W��h/ʼ��h��eX��s��E�y����Xu���U	q��� Ea��	��Fz2��9	X2"JE�NTl���/�o`��  �V[���&)W�8�I�-�]ʔ�{�'�h1����SFlP� >��Iڴf[��aҪI�L��{4��&F��6��!����|�1AC��1@g�*A�������\�*��ȓ:w�yX �G� έi*M�e�,�Ӄ�\}n� 1�Ȉ .C}��#A����aM<YG�7�` ����8��tX���˓m�������n���
�� �\�p)��17T�挝-F��aH�ω�����$,aI�P�'+C d��!"oĥ/h��ta���2!X���e�q9�7�>����P˘eZ<C�e����c�^8L3"�Z�'�j�J3j��H��|�3bT%��$ݴXmJњ���i}\��t�� �F���ԭ|���kL�,��PX�a/ٶ�ɲ���!��%*ٛ��
�B�������6V�L�!BR�J��z��ZƊA3eY?�`2eW#ܘ'p@+mܼvBY�$]�`�1	�%��:�B�lLX<��\������ɪ~��$��j�)�UJ�L�����I�u1
��G,�!1ܩ�GN@�}j�=I�����3��t��3�_Do��cM�f�rD(�t�v ���.�y
� R-�P�ԁi�ѩ�K�8h�6OL��표Y������GlV%�@��*m���W�<T��	Q�ʛ0��B�I�2�:YF*T�JQç��a���'�����&N�|���O��A�ڠ
���ir*O��f�Z��'j�y��j�1oz��
ɘ#@�l�T�p@D��'�0p�{�&r�O5A�N	YB7D�����4c�D�R6mΨ
�t�bqe5D���0R����f��Pؒ�ybB-D�tj��=b�L!�+	F�x��<D�R��ՠH��,C� E�m
�qR8D�$���I�n��*W��]}%C�8D�����Z�,�t59�j4,y�@
��6D�Pu�O3$Y�yb���P���:^�!��Â!�0`T��?B��i��OD1@�!�Ҋ'��iJ@���h��#�$�!򄕺�l�j$��|�
��W�=�!�X�ĸ0�LZ��53���!򤙁��|{ҥ�k�d�z�A�h!�d�r1,u���2.����1ɍg!򤖞�"�ˁ,?Az�uz�jמ!F!�R�]?^|�HW�A��p�ș"<^!�� <��᱀�%~����g�y=!�ƀW`�(�UN�u���<�!�D� slLq�tHΣS=P���K�o�!� 9���w��EJ�@u��3E�!�䉽u.�@�S͋	~��&֚r�!�б;X���f��2�<�a���yx!��<���T�tԑ��� |!�D�%�4+R�TXvz���A	Wg!�d&p���$��x���1$��3[S!�d��P�jEb�����ҥ�DΧ_@!�dA1p};��B5I����$\�-K!�$Ve�l�p&N*fL\��D� 8H!�
R�*�(���OB�)P#��!�54>�0"�n�'6��6��>xB�I9�̲2�YP� �C�:�B�� z�D����/6_����eN#n�xB�ɧG:���G�Ի4�`��O�F�BB�ɉ���p)�������1�
C�t���)�K���]놆�$ �C�ɓ!(F�	h�A�)�T��;-�B�I�}D�u�酹X~� *�h!s�C�I�Y�<P C�)M�\��eE)>tC�	�I[�oL4H�u;B���"C�	�ePL��2�D�i��u���D��$C�I.Ue�!At����+(O�i��B�ɺ�@�`c�¯kgn �@d�w��B��`��|��E۱h.�U��M.B��=h:��	S E24B�cR"#/BB�	/1�P�X��O>��	���%2.B�I�v_TՓeEX��;ᘋz�B�	�G,�l"��J����Z�'{�C�<h�Qk��Ѯ&~ZAA�f�4B��h�<�"�%'�VU��fA�pQC䉨>���Av��K����ܞ!�C�	�0E���L��N�gH�$hƨB�-�ȉ"�6<Y$���DzB�	���B��=�ܻ�I�Jg4B�	��4��Iâ�$�V%�B�I�Q�D���Όa�T�Q��C�I�l�	@�L5H�����58�C�II-�Qz3�ƶc��Xu ���B�	�	����f�Ӑ**zPtH�Z�C䉈u�HƑ�i�
Щ�qݦ]��S�? ZU����/y�v\ٷ�D�[0v�`"O:�`��)+��H�bC�3m-�\�2"OQ������t˥bʯ��p��"O�9��FǢ��q�tv���"Op$Q��ܐ{�"��N�71��q�"O�\�H}�	 �m�^��t�#"O��8�꘾}�hQ�썵6a��"@"OHE� ̀�_?�q��K!6kls�"O���E�&��8�IRSR t��"O�$H"��/j\���3&�^G�TX�"O� ��N̈:Q���Ee��n"�}3�"Oj�I��ۡx�b�c'S�B����"O,dKD��{�K5kJ	�<Q�"O��c׉�#u��Yd�ǀL�,�s�"OVā�	�'C���v��kbz��"O&y���G�ܞ�p�1����"O4Ԩa�)�$@���?��5rD"O�@f���y>⁪�b��P��"ON\30+��)Q�"�k�l�Q�"O�;Gb�)q����59��#"O�d{4!�G����� �0�H�ȇ"On%�MT�Yv��(@�P~Z9z "O��S���:V\|cA^�	}��q"O���ұf��L�(��Ae���"OnDٲ�өL[�(kP(Ԍ�$��"O%��@)���G�4xY�"Ox�)Ba�|�{%O ^�Ε�'"O\�j�!��T�8� �V��%�"O����,Uf���#
��U�0"OD�* F @�b����D�D�bv"O��k,	D_H-	RD��ZPp�"O�	hE蓍bcJ��TB�*�z$��"OBE�児��!"D!�R� ���"O~��G�@�|�|�/՘>���S@"OpyA�p�t�q)k(�"ON�	F��S�dD�[�.�p�� "O�Ipj�#�dIa0@I>v�Nm@�"O�4	b��
��Zѯ�Gi�M3r"O�\�S`> ��͒�	34��"O��A�(�
!�bm�6�@�.6*��$"O��h��#���P�L�5kvH�[�"O2LZ��ˆ<L�$���X�f:x�"O���ǡK����`Ԥ2?hi�"O�!RѤ��"jp�	�('�x���"O��Y�$[r㴉C7����t"O�b4˄o���8IG�	���s"O��B�%��^� �K`+/b����s"O�x*!��/�*��tj��ȍ �"O|4Ⲫ��	0�;��B<ݼm�U"O���B)G�O:PX� ���\p{�"O�|�����t$*v�	h�X鈂"OF	�(j� L��┘8.���"O����+�Đ ��$u Z�*g"O$QG�8O�D��E�ās����"O�#�h��-juBf[�u��0�t"O��
�CݑP��c�2y����Q"O�آG)�>mPY1�F7��0��"O>�ҥͼu74�P��@�b}	t"O�)���Q+�V�C��K�@�ȐP�"O`T���\>2���
dƕ�{����"On�Y�L��= �DY����}r�"Ot���n�͢��C#k� K�"O�%#¶U]�ʡ�.�~��"On�b7Q�PD� �e��O:�Z4"O� ���A ��O��a �O60N���"O|9Q���a�.��oF�K4�q��"O>�yD$��~�ҎJ`:� �2"O��0a��&X|!3�#ֱ�x�"O���pɄ�`�}ˡ"��_>>�A
O�}��Ⴙ/��� �� e"��2�yҪB%>����!�5y��E@�ޠ�y
Tj�R�R��F�tt"�/��y2�O�A� �8�
ؔFK��ԇ��y�� 
"�0b�G%?�~ѩ����y��]R�3�a�:�|L����y��;�l�+@)��ڞ�@w%�9�y���w�@u�憔�x�.�7o��yRJ�����jS#k�f��DO��y2$O�2nV��%_�ay�{uj��y�P1tǢ԰�j1�H8��b���y�_����ֈޟJ�b�����yR�
�g�5�ЄʺHU΄QE�;�yrO�J�HpRJԄ2.2�2呝�y(�~\�Y����PQ"�'�y�@U����2��h�|��ių�y�G
%�Z���IO,.q�-(��O�y��f���W��4۴ �t�H��y����PN
S�"+B�������y�e�?U�}�B��R7xH��+��y�	�D� Dct�N13)���$
I��y�@0J����*
�'��D�Z�yb@\0%���	���10x�cUV��yr��?BU6��A�(6�uҕLQ��yB��c��A��D*��ůX �y�K��]^"�iFB ���GD��y���$,�
W��iJB�B��y���{����d�C��~��PI��y���;d|;p�!�iu%[��y�CS�;V�x֭� �h��ⓒ�y� �&y?�Y��#���{��Ԏ�hO���F'B�`T��OV.TD��#�
�"!�d�v�t�#JB5T����3 FpjFGa؟����!`����!��A~q#�&=<O���%��7C��?}hP������Pqe��_=�9�ȓ{�}�qO�S�������^x�'���ש�;}p
p#�/�n"}�D@O?&	���&I2WҀ�6�l�<��Xj��R��1���a���9p����M�6-}�����L>�%���t���õ$��G�p۶Ji(<�荚N�Xx�ɒ+�\��F�.=���`���W�-���݀9����ě�>�9gE%#IJ����ʆ��x2�5]%*�'Jے�𠡗4>eV��BB�*!��P���G�f���'�^E0�٦?��mȶ�Y�Dָ|"�OVٔe��"I,p�B.śh�`9��k-�S"�v]��胺QJ�E��%�-w�4B�ɪY�d�ۤmN�d�1��'z|���B��-���­`a�2��b��'��H"�ӓ�>	8��B��jt�� "�I �a���;W�.M� ��D�(���+7��e����*��y�*ƞS>��P���HK>�-J�����ɣO.Ui�#ʢo���`����D�v����MَI(� �JP)P��C�ɑRw�؃�j�	N!
��#���SB �K�3��:T�(Q>��Q�A�8�ƨb�/�h�`�Gh<D���5K��y	~����z|���3��?sDi���ϸ��V��>�&4�}&�EN����8Y4ҏl$�� %�� ��]�pn�����D~Ar�ۢش	��ά,���KG��p=Y�F%�nd�R%�8l�%ES~8�0��EZ�ؚ�S��$-9�ŲW隓fꌸ�+��PnE�Հw!���1��qA+**Y uS�g�6��Բ� �<{��ؘ%���@�Q>9I��H��=�0�
���0��=D�\i�@�8��Ԃ�5{`�mkb˵6��`U�Ơ�?��˖6���>�O� �t*�te<���>~X2���O�u(��7�<���k����@�˲yS,q���<���E.f�v����ӛu�d�� �ªj�џ�a����4���l��BM��x ��ԐQ+�1z����y"��-$|��r��Cά�*��Y���d�!F\8�2��ӄo�  r��ĸ�)�-�X�C��b�j��b YǊ��둬,$ؓO���が�<I�K?,u�[��Kx7V��Ǆ�k���H�[�nL`cc@ۘhn��A�W�l�4���Q����4萠p���P�<��EB�À��?m��#C��3��	�A�@$D�Ի`.?}�T�i,A�N�!���<Qծ]�D�:➢|Zu��)[���+g �	t8�7��@�<�Ѯ�`���F,�%p,�Đ'O�0��Œ#G,O��e�O"OǬ���/�?A����'̼�a�R|p��	1�֢/���C'�߰_",d�OZU0���E�:ıO�8
�0�!�'�,��)��8��'$�e	P �B�bԛVeͥ�V���'d �A� �0d�Y��B.0}b$���)��>yd���$OP�#�P-`����.�r�<q  �S!6��g�5(�}��EG� Q8j#?�&���`џ�������CE�l�`��K6\O�Q�3
�_~�h�[�V��!]$.�T@i!Ʉ:B�Vl�Q`%�O6���g�#;�`�T�*	~��R���$�n��'a�a�P�"���E�����T��%�@��'H�!�E�\��)�.�-$��x�deI�P��)O��!�Ń�]�$�E�,O �Z`f̵x4�I��6�Iд"ODmIӄ1�8���gʮ*�TkdMĶt�(��OH����h�'W�Yp��=��c�K��7�j0
�?u��Pt��8i+�)}^�$qEU)\��B �Z�V0���Q�T���	�CF݉��}>DлV(��n��\)�C_�����=�Dѭ�<q�'y��[�슲#�M���
`���

�'Xt�AT��J@. /X��+�MGqyB �@<`D�'��a!��~�Ӧh޽�6�]�^�zAzA��<E"�	��$D��[׎�3SW ��E�v���sf�Z}�x���Y��H�s�ԭi�Ɖ����|��=%bB��KI3o��a�L	��0=ᡬ��w����E�x��(ې`^�vs���lA�%�Ÿ��M��k3O�+KeXfN���<a�i��}6����W7sS`ѐe �q�I3�`Вa(j�2Z��V�u�|��'G��$Q'R{���G$F�i�C�\�B�	�+�f���@�Ac|�a1��4K���ֲi�PJ4`�|�����T?1�n߼K�,�/����@�P�I���ц\bh<�A��l%���c��txd4QE ������y"��
B����d�R����X��Lo��2Rg�`����r��l�N��> *����'N���
K���B��t��1ࠁ#5S���4�|AA�^�z�5r��'�H<�[
�l�+x�.9!H>	�#%8U��H��b��~r�id�(۫)[� ��Nd�H��D?H	���%m�, ����',�D���^.}' �	0��y �'����s
 ?���	^gV���엉>@.T�uD�TpC�ɊR��=��
�'x���'��n��*Aaͳ��D
A��F�%��RQ\�J�RW(]��B��k4<OJ�PS M�H_B��c�UE��h���6�*Q8f�ޗH�Ĩ؁�<�I��T��J>=��ꤍ�F�p4��Vz*�'fp5��F.:����'�܀���?	En
��� ������,u��	�'R>1p��\���0�\�1"�#W���#����<����<������>�&"J�_NB=)�
��2f�l�3�ph<i�JN�w��xP�T$� �7�q�Z���^1X�� h���0�ORb�<�& �� ����c®I˸�!$1<O���gҎ	K��%,�/�|��kL�C���	�d����L�<)g�ݏps�BvŎ�V�2M��`�}̓8�ƍѪ;e���f�}�O�X��*ȿ	��!�%g�}�Q��'N��Bgm�2%؀I�S��<y�Ե��4V�,Q����S�O�L�q�㞳&�<(@4ǁ)l�ꙸ�"O��"�ݣ/HP�	����f�|�2����&M�8��	�Pl�H�\%&}�,Z3CM*]Ql��$��h����f� ���S�ItX����cԝj��(4��)7%�rPN	"��Rꪜ���;ړ/��L��B�B��qJ1@�<4I�
�8b0�"Oڜ�p%@�z����H�V�"݀A�'�r0�W���O?]��˸2i"�qr�\�7�*�K��<9�oJM9���pW�^�v�xg�St~���=����'��3&�Pd��R�B�Y7d��!�1r�tq %���M,��s��G,{�9�'�ԝ�rB
�3I:m���#�$-����)iT�%����%���@��Y�i���F�<6��?�:�XG�[>T� ,��Cy"k�.yPb��|R����(7����H^71p��rM~�<!�GBO�5(�E^&!)�(IV�I<L�& +	�=l%H�H3��Y�tH��W-&����}�$R��9qh��Hq�63<idI0e@!��@��0���?=�d����1�џ�ƀ�/{���>јCM��A��F 4f;� �QO3D����&N0YG���f_�	Q�h �o�<��׻=!&E�<E�d��&L���vH0^�¬�r��/�y�n�}:I���A�ĀX���=��-āZ��,,OBtp��&Qh�}2f��+��Is�'GBur���K����!�!uа�A��2O�zC�I�i7���eB�58B�1AnJ�I�4�?��b�)W�Jչ3 ���� !4NX�M6 �"O������ ������<���qqT�l�ׇ�
�ا(�ҌJ�b�	��2�JQ�V�時@"O(�j�iXr��Q�.W�mXg�|�&8����D^�y�Xixªϝk��J�N-iN��LN�9+Z8	��efA���"�vaq��54��3��2f@$��K�1a�({T�$O�06�IO�p��C�&�R����Gl�C䉉	~VMy����J���A C�ɖ @���'n�b�`��$CĴ]VB�I!{xL���]|@���n�B�	 A�j�M�+wކ*���2��C�	�&��4�5�w�
|�2E��-FC�	0Ɩ4Q�$S�/��ݐb��	(C�	|����0H�6=镠�7��B�	��~}��ܑbQX�2��4S?�B䉚t�␳��� .�$%#ȗ���C�	+sb hqʇ%��8�hX#��C�ɴq��} ��+"�L�	X5(�C�I�J~H��Q(iƒ��ѧQ�Q(�B�&`~��� E7#rl@�@�(:xpB�	�2�tJԃԂ.~P���"Pi�B�?kܝ�H�1qE8,bb0�B�ɾ6.l�k������D��m�C�	�3�����U�ک�e� 9KB��_:|3�/����Q�E>C��2{-4�;"�ʓB�RY�BN�-`C�I:W�b|٢FU�aĊ�3	�(C�I�p� C+��?���1��(6i(C�	+D��)�EU/,
lDa!�M!�B�	�r0��gˊ�b�-{3��C,�B��	Ii
����"q��e�Q�)I�B� }�V�i���'Pnt�zR	�(;XC�R�aP��)f���ر(�C�$C�I!]H㶬ݫ%�8�juA; )C䉫N	0�X�	�L�,�9��� C�$8*���'�P�t�!r��N�e�FC�ɵa�d��U&H�C|L�Z��;? C�ɛ9�M��\
ZPs���w!�	_6ʜ"�cé-T.d�G�ΌJd!�D���b$�dLO)E.,v��!F_!�� ֍��R�wZH���?��q�"O��,6Z���fW�t���C�"O���Q@
h�{CdE�S��x"&"O~|#�� 2�� �Cлj��9	�"O�2�$�v�1���]�`��0""O4P2��#/�zm(Dl9��g"O�%����`�A�4B6�Y�"O��e
ũ.P��Uc3�x	d"O@J&gL�;6|8$ė4,��+�"Oʔa�j�$&�2ą\��Xp"Ot��)�b��Xr�C��L�֑3�"Or!�FE�6��Q��'�!%�x��"O��2�!O�=`���쐢D��mЦ"O|DhQ��/�"�Z��Od�~�i�'�r�YR����vK��	lS�'�����2YW�!�.T�.�	�'d�U�ª��-��j�f�&��=��'�t���:�|A�SJ��:�|,2�'08�K��C<>�����?L6���'+������ Fř7I��Ѯl�'0��B1Q�sfH֡.�֐C�'(���2ظ�$n��ق�'JU�V�V,1��𣢘�A^ء�'��<[�J�E�4-���:�88h	�'�\4).��{*�,:�b��,K���'��j���a��U����
����'�*��wEPbYP�KCϑ,G&,��'���e�=pF"��r"��l}S�'��	��ӱ7�J�� ?zB�"�'���J%傛T��i�C�T�c��Ԙ�'� i�q$�$(�1 c��$]����'?�ţ���H&�J���\�4K�'��;�1�:*��Z�B�0���'�cpJ�R`rQ	�ϔCM�Q��'��a���!�=�`���C����'CPU�cc��K�"�q5�W;z�R�'7�� {m�L�ԃѨ#r(�
�'0<kGo�@�~)�t�	eC�y�	�'\> ��nY�Z�� !���c��}#�'��% '������ Xި �'b��#%�Y�(�t��_�'$�1��'&�Q���s}���o�9"�y��'&h��b��?JP6PW��R�lP�'�A �jP�
*2��6d��"#�! �'�6P��t( ����i�' �(�$6���{�F�6_Z$��'��ma�:����׹|.1��'#�q�Ŭ��ik�R"���	�'c�uPr��14�(�@��xdr	�'�8|�k�,|/P�b�B�7���P	�'�����DC����jK%R�h�'�Ls���	~���B��
��p�'6ك�5�XxR�n%u6��'��T�?�r}"�$�"} ��b�'�^Ĩ��Ԯ���戌z"Ap�'k֨�� ��mjLu��M�uG�BJ�d����F^|���[�w����aW� �����>��/GY+�(X�AP�U>�Mc�d�q�<��N}�l�ƈV�AG�D�Cf�<��T�e�Q��3�"%�)C`�<٦�����3A ���v�)bN�a�<�4�%��|H�J��E_P�1���Q�<�
�~Ę�	�=�B(�P��e�<��d�20���"E
9	���r0gc�<� ��9w��3`�"M�b�T+�8�3C"O�I Bʕ"s+�4�`�J��YI#"O��ҧʈK�� ��Qu����"O�� �@�T�u@�m�&]
~�ۆ"O�1�ф�TбK��qb�<2�"O�����hX�����b�dѡ3"O����Y����Ȓ?9ל��B"On��&*E�P���F
�t`��"O.=�k �:! (/}f@�"O$Q[��W G`f��$ɯ]B
��4"OH�2�'���X�eEA�仅"O�����I�|�i�I[�1��P"O�T�f�.gzPd��	�0���"O`A�t�"<�B����B� �S"O���s�Q�{P��P�a%.x5��"O����Â�rp4a·v�5;�"OH!�a�T�Za�Y3�EK�r�I��"O���tE9oʴA�S� 6���"O�Ix6��2 ~fP��c�6��s"Oh���h�#�60D��$w��I�D"O�u�f�
�������,��%(�"O�`g�E}�>�Х��=�*�ۣ"O�R4�ʅu�֭Y4a�p�����"OX5�4���(��oQ3�]�"O��q�� ^�st�̯7w~M8d"O DqSፗ'"�	��knl,�&"OH@sR�$R���
ИZQ
Q�"O~�(Rf��APj�;�*M�F��,X�"O:A0vA͐<xڐӒ) ׌�"�"O<�CD��;b�v5�T��/o*d�D"OTZ�C1N eH�eәU�-R"O�;�����R��S��a"@��"O���N��(dP�7�`�h�"O��ce:1��]r'쒕GG���"O��ȇp#)@c�� ��X�C"O$�Q���D��Ģ��с`gP%"Ovi{��L3x0�;�(
 g �(�"O�]�w�Ê�@k���Y=�L��"O�uS�Z�'Be2�F�`��"O�H 
Ӑ� ����?�q�"O���E,��\��҃\��(�"O �b�W�	x(� G���B"O�E�e�eȤA��%�,��)h "O�1j��Ǔv*����n�� ݸ��$"O��z�lT�ҥk�N�:rX���"O����_],��e�V�&��h�"O�p��e5 f
�E�: @���"O�F�ˈnipC��_�-�#�"O};�U�-u��8��~!|�!�$>P*��#ʚZ���:��J(]M!�$� |s0��S�~Ub��K1&D!����tt�}x�7n�&01eA�CX!�䁱`��Ӗ�~��Ȁ�"�-1�!򄚱+ "�J��E�d����I�!�	�'k6��.&�(L�#��!��<����J�0���Nұ�!򄜃�0Ċ��˔T���;m���!�ީwм�*���iMn�ˡ��k�!��"_@xm��ǂ
�����
/�!�dɳQ20(���֎m~�5[A�ʳ;�!�d��V�֘�%7jM���R�)�!�č#��!�Р�h��XB�7^!�d/F���x�D�5�*�
�!� a�!�D�>N�00᷏\1�q2���{!�� p5�
�2c�Z%h���@�X��"O��g�KeKD�U#s�=�P"O�)�AA�P��X�_�_X�(3�"OH؋R�X�m�T �D_�]A>�i�"O��f��l�$0�<t*ՠ�"O<������	�j��&�? ���#c"Ox��sD�$��
�R�FװiAt"O���fOG.1վEӠM�,'���"O̠U�O��i���	��Q"O��y��ûF�� ��L
E�"a�2"O��s�J؆�d�/Px�� �r"O���7Sq^�s��43�h�9�"O���@ �R�Ȍ��
�Xhv�0"O�%�5�2 ��Bbڱo �;�"O@�pkQ�� ٚ�&I[��v"O��Y�E㨥�tX���'"OD ��Q5�Δ�c��5�x�R"O @��Fȱ
,����B�-n��ۑ"Ofa�c޻*m�Izȃ1 pD��"O�7&��8 q�0�P
@햕3�"O�"ǩW%�h���$?��Ẓ"O>�+)]�}�VjG/u�F�Q""O�D��D�g<˒	�Ś�"O�l���Y+�F�`�AD�b^�8�"O�\�#@C�pvʘ�O�4����"O��B��c�d%Y�S�t��pw"OV��SN�)N���0�/έb���{�"OVI���,!��pe!O8U@�L��"O*|p�G�W�Heq`�&� "OB�"��A�r�25��$}����"O���QM�$<>�ѱ�b� %g�D�"O$�Yvi�l��܃�d��c�����"O|���B�j�,�rAFN�ba�"OLEµ&R�t;��SB�h�8#"O�Y�,U�V�Qx ��,ĺ��"O>�1�E0^�5�DAף9a�d35"O�[�~y�uбO��w�,P�D"O����+W;L�f.�OlRPb�"O^���L[?���aN��uI""O@\83 �-p�\C��49L�ku"OZ���O�<?�PW�!Sᆜ[ "Oƭ���:5�^4��Ɂ>(Иe�V"O�Y��$Ӳp����i�N9��"O@�U���WD���e*8*fѹG"O��⧧�r����RKQ+����"O���P��.�A��ڵh�i��"ONe����I<��S��F	�Ɣ�'"OZ�V�G0DrⰪ�#�
�D"O2�����;\W� �RI
O��	�"O� I����:� .���y""O���Q�Z�zR���mG�2J�M�"OZԂ����4hڈ��,T4�`rV"ObDbd?����ҧ�86�h"O�d�bm�@�q�]�R5�qJF"O���`������(Q�z0�u"Oq��̉i��Q�)��q�b��"O�i��* �Q�����T
R�~y�"O����6�Ҽ
pbY�Q(���y��L� pY��30M�2(��yB)B�eܺ�H@�����AQ��yҋEHpVA;B��i3�mQ᪏�yR)?A����M؜fCX�+���y�Ɔ/gCQ ���W� qd]��y�e�W"��yS���R��sp���y
� (�Ys���jW�A@M�H���U"OTʀ��)���ū^�(]��"O�ih4��(]�,1���U趽�G"O�QF	�q�zm����{�} �"OD|Zrk��g����)�>F��4�S"O� �b�K�eqBI�.!x��"Ofy	�G��\6��s�I�	o�	��"OpL���p����?�R(�0�љC�!�v���s� 0B��<�!��� ��9���_4N�G �!��DgK����C�Y.|�F�D�!��,$/��S��G�|�м��N�!�D�����@���-�t	�f��!�F��TP�k�U&�d��_@!�ŽZ�� Q�ϻ=7D4�`	U4!��Y�)Kȼze&J�NMX!)Q!���v��!Iw��-aqΈꥤ��-!��4�b�Ƨl��a��)Z�!�Dj����u��Z�"�S�!�d�2� <s�FI�G���R�!gG!�dP�y%xc6ņ�M#$�C1$͍lA!�H�F�A�0Î���+�!��U�*�DH؁Ξ|�����f!�d�J�D9�T#\�6�rp�E���/�!�DR��H���P� ��ϛ�!�R�L)�%S�^-�aB�K�8@� d��Ӫ��"J03
�LcpJJ�m�M�G"O,`AA??>����@�iSR�Y7"OR��d�5R�b�Ih\�h�8�"OP乃/"0�`�ږ^6�L}j�"O��y��գ���@�jP$ '"O��g��l������5^p�Ц"O�H',Y�E�Vy��GQ:F`�z�"O��R�F��O�j�9'�C!xAD�D"OH{�M�7��Dէ@�a��"O���@�o8��`9J�R�"O� �ǃN^�a��7�r�9�"O�����ܺ+�����u���6"O(��s�ޙq�e��@��U��9H�"O.̢�튮J��z�M�ĺb"O�I�2L8�(� ��@�Vq"O�i`�ڣW�x�r��5�M9�"O��F�$}�n�z$\��x}��"OP���ץO�h�P�&{B��"O�a�d�J9j������|��"O�$A��҉��<�i�0P
a�"O=Cuj?^�p(���TcR���g"OX�������F�7G�d@"OH�Ku��z2���wH�l>\�)�"OB8���ٖe�T���F!z�@"O�U���׹ib�  ����+�"OfP��!ڸ�bx�C
�-LS��X�"OH;��d0�����м@:Щ��'�!�H2^�Ds珉��1H��@z!�D��܁�e�I�uU����E�$t!�d� �H#��E�D����[!��Qc$�3!ޣr�J��aGj�!�$����u�4�*!zX�s�N,L�!�2_�ܻ���r����DG�!�$Z%0�9��ޓQ9N��E�J�R�!��h4�!�$�S�YHR��K�&!��A5��As�c�2,aʉ
�'xd��
�3k|�����Y�ـ�'���x&*�61I*!�V�Y�c�֨��� zD��(�. ��k_;f4$`��(�S��yRk�,
�tI��ܯIM\Œ����yr�ճ1^F�
��� �5�yBC��	@����?�`�Q�ݰ�y��U�n�(Ѻ�Y�
l� �O�y�B^S�Ƚ�����i N��y�L�lP�,12�Ӊx��hK#N��y��g�T��N��w�r��#E�yr��+�	r7a](l��D�L(�y��A!� ��6k�.�H� ��y2���6iF�¿��Pm�*�y��2��AK� F���=c��2�y� .�t���p��A���y2ֲ_����P�}�0���[?�ymI��A�����9��� �y��ٙu9��b�!��s�������y�԰FB���#F>n#VdA��O(�y��P!��c�K	X��(�A��y�!n36����I�8<f��yBŜ�kN�����M���udؠ�y���9y4r]�K����Z�jC��yRO�	GH��&��tj�$H�y"$X2_��ؕn�8�ʴѓ�ފ�yR��6�p1閥F� �y�4���y��I�F���Y�%�w�Eڃ���ybeG	F{7mH(s �}y�:�y��E�`�\���x����7���yR����XT�oU�i�J �g��y��
=��x�$��&3cN� �!�Đ�1�.x��Ѷ��xbm��T�!��V0�i#��	����>�!���҈`���_�9�Gܨ})!�]�q����@���bWl��H�
=�!�dǌ04�+���3?EYrs������)��<9�"�*OV>����D��*SE\v�<��LT�z��LS�Nr���n�<�TCW�E�Bek�A.Pd���P�Qa�<9�GP�&ĨD
���-`���kaU^�<Qwę)Ty� yS��[ܔ2��W�<��-H%`�8#��"I�X�2�Y�<��m�M߬��
�$#~���i�O�<�aj��f�P�2 ���?��K�M�<Y�C�v���!��'1��⃠�I�<!���2x�ͩ�.�9m:�R$UI�<�4/ċh l��V��O"����eG}yb�'O��Q̎�>��t�� <$|����O�=X#�P�x:!�2�$���g"O�X+W�I�@�Rc�	F�3A�� D{����ԂTs��-��%�(j�!�$c�Ё� ���^��&�^�!�!�$ܓ ��ʱc�	y��c�(Q�!�$ɂPָ�yf�C���E��G%�!�̝{ڐ9a���GY�aKw�ٲ4B!�D�ZOp��FڭfC2�[4�קh@!��=3�FD��I%nMZ�iT(!�$��t9P5 �'鬁����!d!�L�P��MJ�F�"!�E�N�QT!�d�4�T�s����,����E3?!��#����d�%Q��!3%��F�!�D�yCv���C1ly�݋ ��}!�ɊP�j�����&f (w͔#v!�d؈&<V�hY�~GEc6mG@j!��4�:9����p0���ըvQ!�X� �HS�`@80+��5�'a|
� Ă���`[wF3�v���"O����'"nmKF��������"O�e����av%��b
�}p��3"Oĵ���F�Q[��r���Ued��"O�P90�����5�KS�6R44S"O�10΁8Z�H,J$?H(���"Oܭ�um��aލb#M��]��[�"O�%��� Sb����_�j�&�)�"O֌R�`>4�3����@�"Ox�(�	۽J=����ш*w~]`�"O((�m�W-ri���ɐ�2���"O��""����~a�Uj�&V��"O� �B 2)�h��#��F��Lap"Onp+��D�"���aIF-��0�P"O<K���V��
��Հq�؀4"OĝhЎ��v"� �E���J%"O�A���T�24��%���Э��"OpqK��/M~|�d�x��pɱ"O�͂VA��8��u��(M�p �"O�1���ڒw�B���g.}q�"O��z5�3T:~����_�U��"O�3��J98�X<#����Sd�I �"O)��#�"���8����fR�v"O|���V6+τ@���1yC2p�U"O����JL�U� �g Z�����"O�3�B�IV8�t�K��|Is"O�-�5��5��]ᠯ˸�r��"O�qQ����h�-5T� E`�"O$��B�%�ޭ[���,;���(�"OD���*�`�h} ���p��@��"O�U�+ޤ�nE��c�%�F���"OHP��^�W=�0(�blaD�Q��!��X�q�V��C�8N((��BK1!�dN���T����h&����c�3�!�DA���5脮4"�����)�!�d�2瘴
��:w
4ݱ���#S�!��ƓPA�� n��j^�8 ��Q�i�!�D̈́u���7�B�gS�@ q�N !��1 I��B�KJ�I*!K��sf!��"����5�ٯpߌ�cP��*n!��J	aM�|���$og$��t�/=!򄁊[; ��N�fh:wi50$!��T:��j�BѱQ����畡�!�DC�l�YT�=l�&��'���!�ğ[X}ju�Y�W�T� r�R"	�!�D��;�p�C'����E��d�!�$;:MDqғD�0.�"%j֥��-�!�V,p�A�ϖ&.�}�"_�m�!�K
, �����ȗ=��T)��Z,DG!�.}q�"������ۆ3�!��
�n��2+в��i��+ʓ0�!�D�'m�<A�b4Ґ�2'�4#�!�LaP܈ٗl�PȜ��G��j�!�O3)-Kƨ���8��Ӗ�ly��'x��Xg�&P�)6\J�(p�
�'@|�$J��FH䆿>�A[
�'%����ө! ��b%#^�7���!	�'.lX׉B1p�V�5��Y��	�'Ԍ��!�R�U�Ĭ���"�~�R�'N��@Y�n�\Ap�mG<��$��'&��{�kļL����Ed�(��'nFx��@��B|�,)5\��'�	A�ƒ�R3���1�� &����'lj�i�T�h��]���I�<���� ~m2e���~�����4/��D"O(���V㐙"��:�W"O"�A���5Px8�b��o�P"O|C�G�;MR�:�@֮;�N,p�"O�%����nٞ��ѯ�={��B"O�e2�A�1?��]�LC�*�|X/�ybφ�Q<$�ӗ�B_�*܂F�[��y��վ%U�`Q1�,U���H1C�
�yBHȒc7�@�˜�L�� �@�^�y�͏�%7n�ц��;Iyx��`� �ybKّn��a��K!?	Ψ{����yrڎ;*�C0E�B�6u	�;�y⧖�^��Ȋ�`E�9D6E�1��y� *s�r����83�"��kU�y�F?b�v9ö/&3�����yB"�M�yҊǤ���c�-�y��]�M��|h�nJ��@��*�y�"O�z�Й+��� )� *2���y���U\���c�� �!ʕ�yR��[Eve!�D_+y�jUB����y�F�.�\9k�6x��5A����y�W�D6��e	�t��t���W �y�+��0��_:fz��@�� �y�@
`L���]�q�ǀW�y2%�� �(��qB�=[in}��bZ5�yr� p�����/��]{��[�	�)�yb
ǥ`|@l�n�',@���yb� �*Y|���/ �jE9V����yҭ��2���:���{�4��N���y"��84��"��Y<q���:��� �y�%�ĉ��[@6��p�H��y��_(--Qvi�?�T��I��y�@բ>֐�%0J���.�y�I�.[\Je���tk4NH)�ybOӶp�9tƁ��в�K��yrƙ8��ܫ�QFH]������y���d�^��BLԄf�<5�!���yR�(W���c�'�0^���%l�}�ȓ-8�@2�l�$ZQ��z�Α{"��c��-q����%���"�R�%Z�,�ȓ0����"c�?qm<���O�XP��x�.𳡊	0Y�>�"	B=l�(8���H�rnK`$��=2��!��"��4��ېH�<��+̴z6؅ȓu����KX	_�l�S��͹�4Յ�5����O_4z�]��')],��ȓ8� �X�y̌���ٌ`Φe�ȓ$ኤ(PAN|�ӑ��� ��x�b%Z�J� � ����_2�$�ȓG]�����7A%���	R����ȓ����bM�*2n���Á1��}�ȓ5�$�&#^V� t1d��Uf~��&c��b���*k���Q��0C���ȓ7Y�8���_5�ꄉ�#�z��ȓ9�Ձ�c��p��y�L%b�,1�ȓ6A|e�J�Ti�#B�)��5�ȓ.Q ��*��]�� �dT�,����?��|@�ϑQN� B뛿Y�$���]��0��E6W3.��5(K0ZN ���F���q�Ӓ��4P�m	��\��+���i����-l�-�p��&�E�ȓ7&֌˶��7_���{CD�c�*Є�#Kp�ң��N�̫��)�f��ȓZ�r`��d�?Z	H[��R%-/Ȇ�S�? *1iЭ�s0i 5�7Twb�"O�\��l�8�n(� ��
Ci���"O�i d:V��HB�G�%{�p�˓"Ol0����6P\܅���0Z����@"OH�sfF�n؀5�&�
!܂�"O5�!
�'� ��l�0G�|���"OnX��L7FZ��X��\�R�!"O@)�5�+~���ĉU��z""O���V�K���D
 ��Lȴ"O2%@�#B�YՌI�Fȋ�W��T(@"OZ �w�Tq����Λ �V���"Ox�zR���%���I���:�I��y�� �9��%%;V(�f��)�yr��]� �i�B�.grf�ڰ�yb�Jc`�B�+G�=��C��yr��r��@ǃ�)%����$���y��@ Wtn��(�j��BE� �yRb��b��0�$^��y�Ɔ�HA�,��n��V��y�ɅJIR�0����͊G�P��y��%_\�: �U6{~�"����y��R�����"�@�R�y�/ƦA�ニ�e��� �ܫ�y"@�Z9$h��a��`ۈd0�
��y��V"r�`Xc2��.� f���y���pF�9 �I�
(lД���y��KLqQ!'a�4%�%��h��y�43iޜwa�0hN�����y2HO�aI�aQs�ޘ#��{��y�È0�b�x.�&KF���T�yr͒+n�hq��E@����$�y�&��f�!�!��7t� �m��y�*)�%��m�>k��a3�Z�y�_�C^ �P�g$u휅�� ���y���) &�����m�}1�$Ծ�yr��-�4	3�P�fĖ�)�y����FQ�"̳C�>�3Sg��c!�D��3Ȗȓ�� �<ճ��1_�!��Îl�a"�k͕>��9@c�	�E�!���0�Q+�h�FFu�w��X!���?����b�O�����Ho
!�ĕ ?��T�E'�/-�F��f��0�!�dݺ*8�Њ��F�z�0�D��=�!�D��x!�PBf		8��m*�)�j4!�����=��̏S��M��O�d3!�O?�B�ᱠ��~x"��r���E@!����0ieR2/\P��/+'!�=�������)��I�:!�˥t�`Axvg����`mE4-"!��8!�P ��z�Ty#��3W
!�D��̀�uɑx��ݩЊ�{!�D��!V|���ٴQj0[�jF�g�!��X>2Ϭ8�pE_&]\񂇩F�!�d���,]8���$`�9�+޺�!�D�g6�Ӥ�:$;�2��.>�!�dٰRf� ���Io*���t�$H�!��M�� �q/ �"��O41�!�dC-oH��ע�$}vJUd흔�!�D .uJJ���<y���R�V�!�d	�Ry����S�2n�E
Ӂ�
�!�d޵,l��"�GZ�M�S��v�!��A�D:e��6	R^�Q�)�I�!�W$D�0�j�π/zU�  �4W�!�$���HHb�o�tr�/Pq��� ����F��T�V���..��I��"O��c���#\�BL���'Sj�b"O�p`g�
_�b��"r�p"ObDzq�@;z�P����3R�@�"O&��!�!o��0A�䈅Pƽ�P"O�mhuk��?��M�bë���k6"O"U�a�)f�ܴr�(���"O@���� `~$pta��64v"OƸA��� �Ń�
Z�'�� S"OΠ�ՙ3#T���/� ��"O�i�ק�.fL��G/TI��Eh�"O�xaǂ#R�jUNO2|tqG"O�-��Nc)"����E�dd�CS"O�ҕ� >*]�1�ƨ+gh��5"O|�R��#�8)]�yR0\a�"O��$O�OkH���$Y%�p�"O�8
a�U�uA0Őb��"(�1�"O�P��"z>�dx��2����"O�����F�+�!r5��;~�m�"O��j �����"�:u(&@��"Oԩ t��Q	�ա!A�.����r"Oа��$
�A���G�=����"Oм�*c ��5..]��G"O�b�=k��0l;rKf$��"OP�x�(Ɩg-���D��b�Q�"OX���L�k R�#��E���W"O� )C�̝��,㣪Ѻ@�٩�"O�l�2��;oi`�q��k��A�"O���I���@�k�¶
=\�r�"O�I�5��s�d�5��#@*d	�"O^A(t��0 �!H�#'����"O���A��b5��H��W�@���"O��􌟸�D���H��=��	�"Oz,`������L�#吚""܁��"Ox�cB��
(2$��ʉ��h�"O�jG��@�JabƌZ�E#A"O�}�1I��C���r�\�(�Us"O4�BfP�\`�A�L��	Eh"O�H�癄"��B�k^c5�;t"O,�y�Aw8 �h7$
�.zl�a"O|�ShB�x��С��U)ʐ��"OҕHuk	��2��V�CY��"ON�t�>aiCQ�B\��V"O�V'�.:����#둂:/�i9�"Of�3¡�;���j���2�"O$)�v┖&M\t[�Imz`yT"OH%aa�h\zy��b� 7�!�"O�u�EJKMv��b�3�}0e"O@�r!�ָR9�"��J	�}k�"O�HCQJW~�i[5@�D���"O�J�^�f�b�"/�I��-�p"ON�����'����g�����I�"O\��qa�''��&��4�`��"O��X�)A�RQ8�!cP���HC"O
��h�;O�As�	�d�����"O0`*1��.�69�1$�$a���p�"O�����!�,�hGm_h9���"O� Hs��Y�&�ҶKբH,498#"O��pqL��R�>mc��K>$��"O��{��6	iĥ��l� R���#"O@X�g
)�b�B"*X�T놽�"OF`0ʐ�܊�)�hR�[rZ�p"O�����$M0a��>a\�0�"O�ꆪ��Y)��;���A`�r�"O� �������l1t�#�� "O�Xj�$U`�+�Ĕ�B�ƹ�&"Ot�(Q�.^�ȕ����p�`%"O�<�#�خ{U��!��7���"OD�*�/G�p��pScR�a��Ӥ"O�r�o�Mw���D�@�|�z�"O���+D?8��@
#��N�\�!"O`eإM�b�Yyp�_*3h���"OZLB�-�9_�lٴ*�8/�9�"O��x�� �7p�h��̘5�N��"O|�o[7ǂݓnƹ�*ĺ�"O����逻A�
y�$,H jR촠�"O�\
`8�^����:P@��"O&�q�"�5�LY:����tL�%ʃ"Op�	F$�:s0S��:W6X|�"O����
l���2e����"ON�0�"E%zE���+�r�%"O�Q��F�04|��Ǘf�j�H�"On�s�#�����k�OQ�Z��z�"OL��#B�(��L�N>R P�"O`��FC>%a�X`�	fA�HJa"O"q� )H�>���ɼ�ī"O���&��B�(�{���bX�Xv"O�$!��ŷ2{�c�i_+i�@[�"O~�iG��5��w&\�
@�V���<��
O*���ͤZ���#�R�<�� Ǽm"�Yv̈\(�h�FNj�<�c��*~8pA0��"\e�t�#�b�<�ĉ� E�`<d�� ��YS�u�<���1:�
�a�,,x��Q��o�<��fY.�HؓAF��>h��Xw�<�`@	s^`�F�K�P(9 �]i�<�ĩ�� �yP��tF|���)Gf�<VR�,
���S��pHQe�<�BG�FX<ԉp�Xr0�a3��[`�<A�G0�����,� a�C�Y�<��U�L��,��FS�=�di���R�<A��Y�v��Uzv����@dm�Y�<� ` x�2�5&��P�LMV�<iw�ՠR(�4��̚+�p)�e�y�<���O��Q����"���%��w�<�� I**�� �ݦ[���/�J�<�����`����Z��<�)�hH�<QP)�h��AJ�@8��!A�<�)�JCf�� �L���:2�F�<��gZ&XN}���x8�s7E�X�<9D��F
�S7O�>�Rآ6#�_�<����J��T�Ѩ�Ϧ��6�B�<9�(�f� 	)�H�Ez�4��+@�<�M�!6���C���Z��q��}�<i`�W46��E��Q\ebd�O�<��
9LlH5*�I@��|o)�I�<�` ֙^j<�R��B�8��NG�<i���*q�01���uAq�/D�,�b!�O|8��mG@�����/D����OJX�J�
� �z��G�,D����g�g�Ha(��s�`�p�7D�� �*;@�s�Փ;P��a�7D�<
�c�6����kA�"�����c7D��RV�-!v�1�A�+��0T�!D�����F��l��K��2�DIk3e D��8#H�f���§䉟	��� �g<D�h�""��T��@A��P3�]br':D�[ -��'�`$�d��Q�\�Ѱ-8D�� T��X�� ��F�Y��;�"O��&i��m+�`JE�~@)1"O�(	�NO5L0d��Ź"w" �%"OV��/�Ω��5tn&�{p"O~Uc� ѯI��(����Ȋ�@�"Oh0hnCA�y���͞]tpC�"O��#��L�A^:U�3.޼d�d�t"OR��ݽJ��pGL�-�L�`�"O�ݑT��" d�����g�ک�"OVDj��։_��p1* :N�\A9'"O����ۇ%�n}s`�
-�X1�"O�p�%Tל�C5`�1N�
H��"O����$~!���EԳ]�Fh�V"O�@�q�	$��m�ADB�z��p"O���4G�5j�:��6<p`�T"O.�{$͚2[z=���N(Da"O��:aH,c!���B�;~H�p"O(��#��6�
���c�<�=(�"O��x���7��|�0��^V���"Oz]k񌈑7�2�Y��O�6��	j!"O���*��^��p�ao�'ɲA13"O��@�;s����c�E!NP��a�"O�����M��:E�J�dD*u�C"O���#� �Mȸ!�IQ$"O*̋U�],E0���e���4Ӈ"OP1�bK�F����ԂN=��)��"O��"� ިE�ECQ���}���"O�Eq"��NLN�����6�Ȩ�C"Oz�R��{6��+2�A$�	;"O���c�lH$�'O#���"O
�SD���� lHs��3΅��"O��[ׁ -2|4P���׌5IҘ`�"O�5�W���A�������
�l:�"O8����3�ԍ;V���Q�"O�2`Y�	�vƉ&Ȱ(*Q"O~���d��r6UYs"��S�"O�tI�iș|0��_���
�"O��*�e�N����N�J�f���"Oƈ֧��q��s��^m�%��"O �7��E��`.�JYtt{�"O��p�CU1e��X2vqXEL��y⏛H�$ rk�V�65V�ބ�y� B�m��l:�昦N�� U���y�H��Uˤ!��M�C�<�ce���ybA�u�Ta"�K�6C�Tɝ��yb-�>;���Qs%©~x��y��yR��wK�M#挅�$�"19��Q
�y�B�l��� TQe�Yu�߷�y�E��4]@�%�ƬWc�<����ybX�(0�Ճ!%� � ��yr���`٠%iw��B�:M��jA0�y)
�a^V�Ȕ��Af���*�y�҂v��p���͏%�dU0�A��yB$?E�ؕY���,���aܸ�y��9*�Y@��!O� iЃR��y�댦T�rd�c�$?X�X�]+�y��B�?�(P@�Z�:o�*3Nٷ�y�-@?*��ѳaC0��Ā*_��y�+a:�9� "�Fd�$�R>�y�NґqX�=��)ޮ`k�K��y��V9/�ږ�89�hѫS�y�X1V�	���!�\)A��yRmQ�U#�0)��:�~P�@C�yB%F$?��p��/��U�@��,�y
� �]��y�ҡ�,�)*�����"O�
��
G�0= "*�,�<��"O�e��*C;6z�����<�&��"OFQ���3���@��'4(F<g"O
�	����@9%�D
�	J�"O�D[e&� ��ȪQ��. �"O@��&n�\���s3�����a"Oqh k�gb��lq����"O�A�@�{����.��'�h�R�"O��p��S��T!���sWJ�Q"O&suKVc���,��c��;�"O����[���3,���6�1Q"O����@�)`�ZX[F��i���	R"O\"T/��vpެق)W�YIz�"O�X��.�'��r��ЕC�H��"O�Q��1;\��㇄�F(�8"4"O�b�N�/K�U�QfYOĤ��"O�%���~��]2��(�h���"O��Q�S����*�% >!J�"O�9X5�XTd�@u��/)���@"O<�2`� ��eq��_G�$�S"OP�T��s���֍�	;(@�zP"O��5䚗l�dY�dM�.$�-�"O�tʢ���f�0�@%���(Db��"Ol�;E��b�})V�R�]2Ԡ�S"O�H���T�,9��E��"�ѐ�"O�8����$l�v�e�%p� ��"O8�⁩3q����4KD�I�P{�"Obi�d�G/���G��`��l��"OtQ�s�#qѮI�2��qt�� t"O�$�1 ��xB��K��F&䥨�"O����@�_�huY�*�%\$qc"Oƨ a�U>�p�i�\*Hq�E"O�x�����gH�!�� �%"O�ѣ҄�|�P �D���y$d��"O�Ce��$kf4���\��Т�"Ov��󤘐"2N�3�OO Ӓ<
�"Op(��� �b ���"O���U'z�R���m��E�:)�q"O�(B��ͬ<��m�%��Գ�"O�X�텞@�X����3���"O����O� ���+��Ȣw�3�"O�9�T�I �R$+�.>�2��"OTE�G����q  *
�Y��1�P"O��#��E�F@ZP����~J�+W"O�``r`�z�u�BI7 �4tb!"Opp��ˉI�6��)�/#!.q�"O|��vK�#@�����A��1"O�\+��Y2�!P�ړ}[t؊�"OEcp�X&*C�� N�B��j&"OD|�G�B$��"���.��@��"Oz��a�_�	Or��̪*n~��"O��EA_�'�����@ԟl_��S"Ox�ڦDCPp��A�K[Ql��"Oب�t�����3�䙘.X�E�v"O����h�i�N=�G���BUt*�"O���?H����7<��V"O*���	�k���RR
^,}�r"Oj�1e�2_��8�g��~'��i�"OҐt�B.�bhɧ���}���ؐ"O��BF\`�AK��z���1"O$�fiQ� "�\�����"O��u��*9MÑ虊B�f"O��뷨T�6�젢$H-0�~a��"O� ��;1ئP��!�']�:�6h(w"O��sせ�'�����eBe�E"O�]�To�R����
=&^�J�"O:c�E
P�p��F><hH�"OL�F�ߖQ{X$k%�q����"O��	 ���(�����>q�͊�"O�}��P*R��W��U
2Pz�"O� �m&X]�MBӭ�){�|�pR"OP��V�z�HQ���.P߲��2"O>��*T�fU�M�5%̧)ct�""Ox 2'<\t@���YZ�̨e"O�3��'���ئ+����
"O$T�҄Ʀ"~��!��薌��"O��2dE�-x�3�_�>�dh�"O�]��͔Ϭ�U�U�
ф"O
q���`��^D��#@"O��r.VDu�Ą
V؂�"O�9!2bUHl�h&��?��"Oũs,�qk�X���7kZ���"OX��"c�+��Z#
�yc$]�"Ox${� �l�zظ��>	F�8ا"O�����[p�zƊ˯LtL��"OnQ�k�^MI���d<(��`"Ov�cD��;؂h�s�ϒ=�PG"O���� �"ϒ<��&�hR�"O`���j�<G���`�Cu
j�"O�Ā��H4wƜ�ۘx	�-�A"OМ ��dR�����Ge���t"O֭x�LW�kĬcJ�1{D�"O�(4�L5!�*�kp���_�]!�"O�U�0ƃ[�| �IC_�� "O��`#�͋Y	��!�����F"Ot�p�G�#�T]�I��M��5�"O�p�E�g��YE�G�l��U"O���ԬӟMj��z1���"T�A"O, �� ߅2_&( ���'����"O>��#�x}��3l��r4<���"O`�u�HI@�1��8B�p�4"O<vAU;%U��ժ��!
�"O��#��9�؈;銭I_*���"OĜ*GN� ,�z�m��pG�y��"Of�bS�Sn>�a4lҽ.�ZUR�"O��2T�W�g�����JQ�$�pLd"O� V�?%�J �@��&��*`"OXI�2�Q�=����V�O������"O�� �ǣ�@i�ʖ�;��p+�"Oj�xaiNl�F��RjM�aN|�G"O���D�P:}�.ɱiޭu�T�R"O8E�p� # �t�S��q�2MsE"O.8b�L�E��P���oZ�f�����=�z1�ԗX]�D1D����ȓ<�4F�A"u�ĺ����F����Xm���@�s%������I�ه�\ �aqӍZ)(�b��1h��J��ȓ1�(�xE@�"���e)Ѽ{�.T��F<��kr�9 � �yq����l-�ȓ��0����9�,t��K�_X��4��3�(f)��O�I�Vx��;��$a�`.��"�@)8�T]��6�Љ�b9n:�11`h�,zu�͆ȓN��5���H�?>H�`��T�:���s�&̓M�FŜu0��G�XcLp��,�hI�`�,]��`U%˺JFl��g�h��@Ԝ7*��A&��5٠���S�? ��p���r����>���&"OVE�bⓟJ����C��t��5r6"OD�5�1���S�$Ê]a�"O	���b��PcOȧ,�
Q�"O�:����:Q��rD!�>����R"O�80VQqH�ˡ���Mt��Q�"ON�A���g�HP2T�~��"OR��(��O�j���B�+|��"O ��=T��"*��9��!"O���3)X�r�m*S��~��B�"O
�Y�h�
v����䫜�_�N Z�"OI�	�=p ����MHi,���"O 0B�F�1dI�s�g^�B�R�"OT ��H	<x�YCMȨ7$�ay7"O�QI�&O"p���b�'��k�"O6�{����81"A�v�ژ�r"O�`QE��8`00C`�R}��w"O�� _�!
�����TR"Om(�"/f�E t�"`�i�"OL����
�p��r��Πn0��%"OT� VfQj��y#Y�7܆��A"O�t�s	�,�X�92�l�(-�&"Ov8z�gҕ$�R���O6����4"O��XւN�+�lH5�ףbLf�r�"O�S��	->+��9A6���"O0��UNE�P�p)����aK�"O����kĒ.:����>����!"O������C���������"O��/V�Lq"b&<��T��"OpPs"�]}��E��"�0�[W"O��%���"Q�D�W�V��"O��8�,$d����ql\�S"Oh�1���//�!�"�ԣ{-(�ڴ"O�I�� �,=&����K�]&�i�"OЕ�G���J��p�N5,��Ȳ�"O���㇜Z��A����0�VL��"O6q(4
��-���51\	�&"Ov$i1"�6���m�( �J""O�Yxe,�O��<�q�(܈��$"O\��cU7{�5�gL�e�l�I�"O�h#�h��^*���h�9%~p��S"OTa���֢d�֥Y�QgQ����"O^I���Q�U� ��%bx�`"O��+�䓪e4�J�N�%N�,��"O���V�D
(S� �*"�"O �Y���aX2�R��V�L�쁐�"O�Q�g&<E��):GN�1(���rc"O4Y	3ǲB�B�
�R!k�|t�Q"O�P ����0��J�<o�����"O�y%MC�<a`�H�m���"O�|Iug��|6�pF�Q�^�!$"O,� �
�v� P ���=���2q"OX���%1mzpѢ�؍a�n9��"O^�P�A�zrٛ���J��}"D"ON���f@1Oh"���+�/����"OD,z�h	�u6���5jڐ&~@�0"O^��%���oVp�A�ԻOg\Q�t"O���t-��ѐq���2H��"OL)������A��"V.&��"Oh�Ä�Q8�yP̖���3"O��zSf�f�:���HR	 ��I
�"O$)E+�C:d����R�F~�}��"OL�)Al�O��ui�H�.oB�"O|*7hT�q�Yz�+�KH)#�"O� NЀ 	����X�*H�b�q��"O����B��.}����o�+1�h��"ORti���-0���a�S�~�d%�P"O ۦ����Sc�C�|�΁�"O��� ��-['�����"x�d9��"O8mi%)�3<��l�bdݔ6m�(�"O�i�jW(<_��cT�T�I�q"O��:��.Sb����ΡS|aU"O>	�u���\��I��"�;k�ź�"O�(�S ��.�L�(���wj�W"O��*�R���〠0j|�u�q"O.�D/H0��9���k{�xb"O��b��C�[(�:�C�ot��P"Ov�$��Bd6���!`;�\ӓ"OpT�E͐*Q��e�]�d2��3�"O4ɸT`���d0���+)�e�"O����	uP;f��@M*�P�"O�(�F��J� ���F�<TԞ5"O�)���$}$v��$8�6�6"O޼c���8!$�r3C�lj��"O>͡$�{,>=��"_g	�-`4"O"����!�Z�*Q���6�  �p"O�xY�J,���o�,�:�(�"O��'E�����s&G\r�tU�"O��7��Q����P%0�|H�e"Op%8#��jA�hyգ/+�J�Q�"OB4���L�N��u�vlΰ%�Ρ��"O<�!�.��~`C"�U�Z��S"Oq��l�:7����K�uX4E�e"OD(A#Z�4
���ÖQJ~1��"O��pV���o��=B���M=���a"O����3&�,Y�!>|�H�n.D���d�ܑ_4 ���]���E #J5D�P+w�E%u����i����&D�`�a� -		Q�,U8;g����.D�H�s)�غ��"֐L�Ҹ{r D�X�d��[*� NӁ�x9C�<D�H��S�mt��k��>*l��d9D���0L�sH%�'Ȁ0cTbA�"�3D�l�1���B4-I�Ȟ{��aX��1D�x��`������^�6ut��$�/D��Q�,�c�\CA��,M� )�L9D� Hre�%y���)���8Fa�,z��"D��!FN�&�k��+l"tl�ak4D�`���)Sؐ��W:�v�h��>D�(AC���~�BI؂퀉C�f�X",=D��y� ������$E"�hC@�<》g��h�lŨCv� v�{�<�PM]6BHE걪[.H9�'�[v�<���U�	�(�*"��8ŚH^>�C�Ɋ[MB��Kaz�j�鑒�>B�	-#y�i
�)�?>t<|s��eHC�I�C?��ؔ��-_,�'Z>.S�C����*�7"t�d Cd�*|�NC�'~X�<i����/Y
�� W7C�	.}Q���n$���#�*h!C�	@��Y��L[o�53U�ޭ�$B�	8eiR�:�xr���� v�C�I%22��.D��5��8��C�	ǌ,��KKG�@ԤԜG��C��y7��B�)O�r%SG&ԟcR�C䉢 9�kv#'���ۡT)<#�C䉈��@pb$\ْ�c��;�rPh�"Oڨ�r�@���!�d�F)n�8C"O� �ː��"]��5C�b��U���c"O�չ �H^(0����\��"O�H�� G�|M�`�J9i��j!"OL���F�C�����\�nb��ѡ"OH�P!�Z|\" ���*s��SA"O0M��E�,?^��u�Х0i(Lsc"O2A��$�:A>�$ö���NT���"O�X`̃�q�0�GVP�EӴ"O�|�acқs6��Q������pr�"O�i�B�3V:�	ڷ儶82}$"O�uڲ��s��E�;9��Y��"O�JbaZ0zB,��(P�J��"O��
�J. �h�j�Na.���t"O��*�ݸ����2 
���"OS����\�VN��l��Z�"O��bd�B�)G��`W�߭�%K�"Oਲ਼	C(|Kl�*Uh�*�"�j�"OZ%���"�T�)t��6N��"O��c��Ԕ2-(tȕ�F�dV0��"O�uPlR)J�J4ÃoA*AH��@"O��� �'1y��qAͶ*G�%��"O�Y�c/��9�`�x&��.0<p�5"ON�҄�GePV�j�kQ.h7�$�"O�U���>	��ȡV�_CL�b"O��3t� A ��©�iBt�r�"O 쑂BI�atҴԧ�:)�}(S"O��i7��ĬE0@BE�0�p"O����X�>��{&�i؃e"O�\0'M�,��!�»,�Թ�"O~(�����Z�P���(����"ORE�m	�aP6��e�A���"OtظA$T(+ozF@߿VJ(1'"O��C�G�|c4�����y[�@�#"O2�FR$��ES�#n�P	�D�<�E�F?Z"LCDW��Xp�*Ru�<��ɖ"B ����_�)��Z���r�<I4eζ �
�9W��"�D���y�<�g �.EZ^-p�)�]�HxK�Z�<&E��Xa�����T��b1��D�<��"ר*�pAp⫊�Rj݄ȓ<��<�GΘ-
m��M݈$���ȓc`�=���&%�Ta�I�>6xQ��0�n=�h�3���&Fp �\��L��AE�_�Q-~��D�7�����u0��c��� �v�3'B x[���ȓ���a��8�P+�JĻU �Q��e���alJ�A �"p��1o���ȓ@�*ź�,g��@�ƈ@�Ly�@�ȓ"�-�A�3t.T�u/��6��ȓm[J}P �ܧPz QA��� ��c��2�Ƣ	k��!C0~V���ȓuP�ph��3_\6iZ���(u�����
e�x��,g*(Zŉ�<�5���쉫ӅO��13�O�B��ՆȓW�R�ɇ�^%���{���ȓ~��@��@�z�"� ė[%����7>V�3fE�Sj �¤OI�Zu�`��h���el(�k
�6l��y\���V�T�elP��@�m�ȓ9h\%�T�;JN=��I�G���1XP�-�p�	h`�	��)�ȓ�9�BE[z�v���I�4x�ȓ�f�R�	�V�P�����݇�#^.�Ï�>��d�S��
'9���S�? NԈ��L�Q�����T2D0�P�"Or��5�	�G��v�ۇe6HS�"O^�"�Ëb%:�i@�A!�8�"O��`��7��T������|�5"O\Ī��+�:��c�İB�X�yq"O<�Ƨ%N5�-��¿����"O�y� ��	k^�Q�[��l�D"O@3%�j��1, m����"O��&�T�a0�l�46�)wE�p�<��A5inC��D.�����T�<a&B7_�p� �'�le9��Y�<���6e��)��x��q�p�I[�<�El��O������qX��T��Z�<�cgؔ{_vL�"��7��I{�T�<�2�W�(��@b���- ����G�<�J��2P�({�dh��G�<���Z�5B(��!�ŉx�` 1�B�<Q�T������p����{�<y @4t�|q��__�Z�(Zq�<yF��8�v�����=y(dȡ��p�<�RlK	�����[9[��(1#�h�<wĐ �f1���Y2u�~|���b�<AD -*v��pB.cn�0�$�E�<	��K�1f�i��$(��GGZ�<�"�:q�����ɥ"�� ��@BY�<ٕ�u`d嗤D\�
5B/T���O� Ԥ�7��zI(e���(D���2N�	,��󄛐", %#�C:D���

�'����'�Z#$�I�8D�du�9I+@��%��a�q��)D�$����v�"���p��@o=D��F֚Ĉ�������5D����c��o@�*��eYUum>D�4�q���5aEM}<u��(D��P��.e�,�#͊26c8i�u�2D���D�������>��S!1D��(���d޺舒��;��\1�E$D�(�E�#.��O�$�ܛ�$D����̆}�^I[�bd*��w�=D� �g�;@`t�JB+b�����D0D�,��I�s���XP�][��%y5�/D�D8&ʎ$�cs�Y;%�	yR(-D�hѢB' �r@	Č#&z�S�0D�x�t��2�$��A,F�>�Д�/D�\��fa�1���9W��PAq�9D�,�4͍Y��ڐ�W	��H�5D�8'OR�U�������\�,5D�ĩVD�8�L��n��`�޹:ª4D�Qd�Q?f���b)V8�}��%7D�< 6�ȋ{�$�Qe4h��Ҁ'D�� �"�5+�0��
�t����k%D�Lˀ*Ɗ\ߐ�aծ�L����L8D�ܡ��ΧT� q�I�/b�� ���6D� *e�C�`8(�g$ج4LaJ�6D�,���ܒ}�,�4��r��7�>D�d�U�����r�f��3UH���`;D�ؙU/�2����C֭?T!��D�<Q��2:F<��$� 9��u��z�<#d^=(�����Y~Ԝ�pj�w�<�����ۤ'��!QDL�O<x��m�&-C�9*�}�5oL�q����X5��iB�3&��!)U��M����9⥃_�w���9�GQH�����A�Q;�cL;AV�+�EҶ��S�? D��$�$(6|0u��:(�(��"OD{�j�M)�8h'I%u�<�3"O��X�C�|`,T1��z�R�8�"O4�p�֧����� ��}jQ"O̔C��kY>]�%`RvFI�"O���JVks`��C̛n�a�a"O$�x�bG�P��"�$�X��"O�MB�E\�k�Tq`�'��}�8�)�"O@{g&�*	��,�7�5E���p"O4��&
��Y5z�yg�02] &"O<��
�'N��	���Z8�E"O.	�F��k��+�ř�"�f�rS"Oj���|��h��A�aƱ$"O��9��Y&�%��(��H�|�"OH�fPUKdYPGݏ栈�"OD�� iF�Z9	������"O8�����8�hH0��* ���1"O�L��
4��b�gI*P51�"O��
���� ����:\u��"O��k���0KC�U�?G`>��"O� �'ES�'%ƴ8��/_� �D"O�8�b�]o׊���@	�=��ѷ"OZ����L�pF���en�<��|y�"O\�@N�y��}�L6�F�b'"O��R�I�J
E�%�\�Yv�)P"Od(��j�nd��١1b���"O|=3��08����K!rY����"O��`V����@}�A,�q@*��ȓc��Q�� =j<���L�!!@jl�ȓT�&�K���_k�5��_�c��E�ȓrg�Q:�얗��0ao� {ĝ�ȓ7�l9 �!��a�H�9�-,�H��X���Ё"
�Pӱ��GH�d�ȓg�"U "�S/@���*�e�
p�!�D�!;�v@0���1�t�
Ei@�=�!�Ҥ@��`��ȝx�8d��H�!�&z�J�k�
�q�y�%B��!�Ě>`����Z9����͉j�!�D��o\DqI��4���V�K0nB!�D�&1IR���I����Ga˵W!�d�0&
6�3䘍+l ��M�g�!�䝯U4\��⠌�h����B�!�R�|�D)�G�[=,Yȝ3B�27�!�WF����I��t{U��*H�!�d,
}���(�?b�e��[z!��*�^ҷ��D^��С�W�9�!�$�(N!��e �*/�V��eg\#c�!�dI� �ސ� ��M���q��=!�#}�� ��+?ŪQ�CG}!��2��za KC���t�^�(�!��	}t��/͒ؠ���+�*\!�� =�F� �j�Qpv�Sf�W�,�!���\_�D(vN�+-È�S��F1�!��l�倂�W��8k����6�!�$�5f�S�� �D��G'c�!��K I]r��"�kt�6ɗES!�dɬAFT���͡3t���슇$!�䑦<�fA������X��FA
(q!���@���9c�Z�p������F1q
!��o��壴��/s�G`��~!�N�p���Z&��P���9!��$똱�!Q�I�>m��'ƠmL!�
99 �+�-�8��h��#!�D�04�H�A+��O_��SUd�%'!�� *����)r_l�8�$ъ6C�y`"O���#j���� �-bX��c�"OD�6�
�*��s��Re��
�"O (IUG��*B:\�u��4*0���"O��`�� /�>mڦ�њZ��(�"O��x� Q1X��)��'F��%��"O`3��D�d5j���eC�p�|y"OH9�hZ�	2�x�F���	��"O���Q&ޤae��pE��s���P1"Od���gE;{��aE�u�&�@�"O��K &��H)4��P%4s*qSP"On�"�@K�2�)I���W���"O x�l���Ȁ��Y�#�ݺb"O�����T�T\�����[&�bW"O؀Sa�J[�Ҕ#f-���R'"Ov$kP�ʼ'���!���
����5"Ov���CH1q^�1CD�%~<�x��"O�ĹY�̘3��Ǝ�.�)A/
�y�L#Y5�у�BX�e�|�Q�C�y�B�+�$ě�d͛�N�Cd���y��6KM��p �	{T *��,�yR���i{���(N`i���y�+�|4,��V$ڸ#t"���&�yrdݩ,a t���ǈƆ�k��y"���M��E#�^�H�`- ��yK��1��q4-�/#�p�Tצ�y2Ł�0���0O�2K��2����y�Ⱦ'��Qi�,� �����]4�y�`N0����q`I?U��Z��y���Pf��c�'l�X� ���yR똕%7� �s��T��L����>�y
�����(EiM����O��y� 5��{d���qp���!�y�ǜ�
�ڄ�<wNvYj�bZ�yRg�,;�*%A6B�/FN��8�y��_5MЍ�Bn;D�8 5�C��y���;3�PP�1��<b�Uϭ�y�%�$*����A�}bTpZ�b��y�cߝy��e�A���:�J�-£�y�`U�k��Q���'�D��"��y����H�+���E uዴ�y��na�$țR������J��R�'��L1�A��%2t���B�uެ���'+�HS��R��-A���l���'����R��$����@	k�ds�'�*�b5�[x6�:��.f�fe��'�hlh����z��3�F6CX0C�'Ԗ��C�En9����� ��'*Dʤ48x5�$�2^>��'�dX;R�v��1�Ѫ�tu��'�zC��R/�p�ǌ��l�:�' ��ɇb�|f�b�W8u�~�
�'ZB�f)��K�$@�Ć�`?$5�	�'����%���M�����-p�c	�'J��+��7C��3�e�(w4���'�d0��G�f�R�v���
�'�0�I`�B%a<�aΟbQ�
�'h�l�W�W�S�L\H�D8,�E*
�'��i` ��B<�ݙ��O�p�P	�'༥�dN� Bx�1�G��G�\��'ղp1Wϊ)�`��eP�Cqj=A�'�"d��O	�J&�����=�6<��'�@=1��=V4� $�յ_�|t��' {��#RD����c�7*"�) ��� �)(c��Mzѫ�!5-:֌��"O4�R���+xB �%��'+Jmxu"O���1e��V�z�N@58tX�"OLy���/��4Nʮx.,�8�"O����Y�9bmx��%zG>9	�"O>�Ģ��-����K#5h�j�"O�Q���W��Q�I͠}p���"O�q��	�(*��� �����}@d"OfuZ���w�Hi��	/�"���"O�pb���'5I���lF7�:qq4�'�'�T�R��})PT��D��6�  j	�'{�!!T +�욶ֶ1�xX	�'c���˖�N\����W5uز�i�'����be(�z�;5�s��b�O΢=E�$�E�k����M-Q��Q��5�yr���u��x�B��$z(*�3g���yb ��rh�q�V��p�`��
���y2/�#O���;�o^��&d��hԻ�yR��y��A���J$��''�yrnƀJ���sEC&���Z�y�L���h��ߩ1)�hr&BD����.���P����J�H���ض�13SN)kQ�K�:�!��<xZ9Ԉ��L?l�&(�!Ot!��;P{��A�ɰƚ%��M�$yW�zr�P�)�Ty��R� D�#�ܦ}p!��ج{p�M0@�̙_)^a�wB��!��D*Ϥ�3��,iB��S�U�J�!�da�=8�#�_&�1�9Uc!򄜙xN���S��ȁ3��in��dA�,�@�J�$���9��	]��p0�'La~��M,2l׻<�6 {楏+�y"�* ��`r�P�3Ҍ\#�N>�yr��#? թt�
�6�&�"� ��L���OdʡStͅH�Du�2kȫk}� Z�'u2�u�B#94���1J
9�]��'�r,��.K�4Rf)�P� 0.�VH�'5@����MQV=ۖe�s, q��'�d��e�M	��m_j<��	�_,|#<q3�SIF^�[VOP4{�ԕ�pU�<Y�̅#�
����ӭ3)��u-�J�<a�%�@v����({#������`�<!W�I8ڤ}�c�4��]D�<Y��W+nV(ۣ.!B�� tʊAh<Ad �C�ę��$��n�~�c&���y�
KS�.���#@�Yha����<�y�@6	��j�k��U%`}�$��!�yR� 8��9��R����Sǌ�y"(n�LYyQ+;8R`���y���rM�2�Y�8-BA�7*��y"�Т[���P��2iͲ�o)�yrbTz������<8�j qΈ�yr�,7�=��͇=2\�I1�ԛ�y���@����O��.���J�OF�y
׆Tg��:��ǭ;��������y"�D8�h�!�I^�.�'����y���:�V�;�J�F �q��+Y��MsOn=r�U>l��B�#C���"O����NJ�"���C��B�<@8�"O�L3�m�Z�$y�?4��``�"O4����9y�D��W#+�����"O����@N���k^�Jt)��3�S��y�%�-��Yҕ��5�2���y� Ӡ^O�AH��܊{�DL�D��y�*U�$�<QO~�'G�����
W��G.W)D���� ��'聹���K�^>qB|��q������@��=I�ٕ�̺��؞D���.� v�X9&�\�rh��B��N9��ȓ��ub1e[�X� ׌@�v���'��5�)ʧ:|V�	f��9_lQ���(KG|̅�����"�NzT�G��5�vD�<���ٰ�i��(���B�`�jԄ�	l�C��혇��q���ךH��uK����K�E���t�ʙ�>���?Q�g��nt<h��-Zk0*ф��yB�f]�hJ0��P9>�9�囱�y�g��tr5��A%E��M8�䂣�y�����H�,d���w�1�䓶0>��"B96�XҤJ�-V������E�<�qn��B݂��ϒX�V�˥��F�<I.P�t4{F	�Z�F�����D�<��Iن�̠��F�UV� 3��f�<�t�ǭ8@���)����Gd�<)%��-F� ���@��S� ��wcM`�<!W Q��q3�"��vJ�]�I���I��Iҧ��h�J����^9U~C�I?�0�ңG9�,Q D�+C6B��&j���3h�	��-�.�m&B�I<ž$Jc�ԑz��	�S��456B�	�p�@m:�OB�Xd�F��3G��� w]Q��}�Q7a���Ao��4u�X�3jI@�<�`�ךI�|L#�	�E��-�#��<1 J�{?Y�����R�p˕"�b����5�z�#`\��x��)"與�M�z�*Qi�/Mʌ���B�؜@��-ı�e㞠�Z)[d�m��L�ȓxv�=�1�� �6����9��L����pÅє�V� �c6Y܀��ȓcT���G7�h 8����
�dt��0>��ʰ�Ϯg\�P��b�݆�i3~=��"5|�E����zy�ȓ0� ��뗓%,)�SlK9"�\Ňȓ4d��Pn2
V8h17�̸@v"<�ȓk������L�`�ʹS���67�p��(�=� ��g�b�� �ͩ3�h���r�h�#��v�������$��\�=A�2LOj������ �R/Ê��ɑ
O6m�9hs�CWB�q�.����͔g�!�Ě/ :����#�+�TyITH�i8!��0b��x��ڷ��)3M��+?!��P� ]�YK jT: �PD�+C$w �'�ў�>����֭O�(��	�6j8=S�j6D�p�G�/(�髣%K�9�%�4D�|�ԃL�U	F��6e�ؠ�� D�L�Ra��B�|�c掸X�9�'�?D�4�V ���zuiK�D.}a��?D�(B���Eqp��C�
�8%(9D�4p.Ԭa}b��AD
�E�8�t(7D���+G�'B�M���ۻ\<�u{�g4D�����U�h�<��E���HF�<`F�$D��+��6E��R (e�����/D������6�t5�Tm�%>)�!,D�t�B�2[���ٴ�Sk<�6�)D���B���[��dBё;x����"D��Ҵ#��G��
D�z�\9�� D���7�V�M�-�d�C�T��$�?D�В�n�.z$�0FD�?8cN��"+3D��g떅]5����Vu$�J�
&D�$�D怗/&��1擿s����%D�� �8�ȓ�~���	�HD�e"O�h�R͕�6��z�_�>�Sq"O�M �5X|E�43&�z
�'����Ȥ�֨	�Οzv�y��'"�
�dޜ3Wtٙ�e��rS����'X�r�+�I�i���	m�zѨ�'��o_~4"M!3� �`�X�'ۺh�iR�1�h�(�@ʄ����'�x�vk�����S�_�	1�1p�'(��a�[�h�a�V&�n�9��'���+�0d�@����n3�m��'��Ԫ�d$\U�4JG�O�|�
�'X�K����H���YSG؞Ay���'��pA �$�0 rrj��fe�a��'D�=ڱa�3�N�CSgN�c�9��'UZ�Aר8���g�Ւ]MV�X�'Y"A3�!eN��g��Z/D���'⠡�)�I���� ��:��)@�'�� �JӞ%[�u�#P �ڜ�
�'q�) 4n�b2���)����
�''���LE�)�D�Q�-���	�'�8���R�H�y�
�ˬ�	�'&�h[���V"8 ��(t��-J�'Pj0�B[�D���)טh����'�Pp�PnAr�e VL'�h�'��i�킕;;|�%�ߵ\�z�#�'���C�CC���)r�MB�X`
h@
�'�԰a��2RT���f߲E����	�'V�\5 ̹����6o�`"��*D�$�犏6�>4�0� \Y `)D����/|��D����=6d"`+D�PT�[����Q�n�>���x�O6D�8
�]��b�[&J
|N�إ�3D�l3�ۡgg���v�;	$����1D�y�q���q�k�+�6��GF1D�p���.TU���s:�𽢡 +D�����U�<��ԛ���*�&ѐ�o4D�x��_	|���P�/�6��a`E?D���'P����G��B��e?D���D�	v[|\1	ZWXp谍>D��Ь;}"8ڇ"��n�F�"�,)D� �P���i�� SH'Rj�H$�"D��C&��)]ؐ��Z�#5VI��
 D�Db�J��``�u��d���ڵ�m!D�8��%į����!臰PB~X�.*D����*VV�P�3g��.�P"'D�X�Q.͝e�b#�כD~���(D���p��) � "S�3�lIx�i'D��P ��n�8xJ�mGg��4*D���G�&$Ќ���#G�~ǘ91��)D� ���U�X���1ժĖhg,lp�
,D�"M?]2��Q"̟�)�Dp��+?D�L���5*���S�[�4Z.�j��/D���g/NZ��)ٷ���p ���!D��J��E�(������4�&;D�@;���/l�q�ӌ�8)�,�m>D�����*93R!�6��+O�*Īi>D�� ' �%p�
ܨ��W�`0�%�(D�܂�C� ����aFJ�@9,s�$D�tr���R�*���������-D��&I��g�� ���x)��+D��jTJE74���0�K�=ixR)D�\�Q)o�d䳠DD�f���*!D�,��C��'f��OC<�z�8s�)D�� "��Wί1.���A�%z��xӑ"O��i)@�G��IC��?��t�7"O��#)��t����>uʬ�W"O(�S�͈.�%�1���g�vQ�"O��`�O!
D
��5��N��g"O�)��+p=�4�U�� :F�aCE"Oy�f�S�E����d/W7�b�"O�$m̈́T����d�4��W"O�%���ҥu��������u"O�YPwϗ#r���_�-l����"O�kG�:A�a�LY���P"Op�ۥ?���12@X.8A yA�"O4@�1%��@]O�:h�5HS"O������5tZ=�Rm	"D
N49q"O�d�0aF�*5(���+�FS����"O��0��Z�2Ơh�
K�l9�%S�"O0`�a��0�XR�+_�l+nȡe"O�� ��Yn�5�a�ƾ_uN@@�"Oʩ���It��p���j�ac"O`T�]�O�>�c���?8�nL0%"OĩRe7y�41S��C^t�!�"O�qKp΍7asz�bq���>��1#�"ODU��L	���Ь�6���{$"O	��ɍ+A�@�!�"v���"O�q8��\& &�$�'�0s�d@�"OL-����D�4L`į* ��)��"O�����&����LM�>�PL w"O(�r�<���R����г`"O�5�3���0�*,i�ꕥj}Q�"O$�c�A���ڤV��x�"O.H�D Q1@�>���g!g���P"Ov��@����3��'F[*���"O�Xi6!ʄR{r�2Fg������"O�p����O��@9 Ź�.���"O@��"H� _���1N 1�ҝ�S"O�d @�^��$*�2�P;�"O6����]l Bu�4���P"OTȩB��myv`�v-�(m�!�q"O��z����#��QB�G�u�
"O8�P�!�pٸ0���V���U��"O�ex&�sm���u�6��u"OR�"��4uC'��:a���"OpCt�����!�S�PH-��"O��Z���(��R2�тm�u�V"O���2-�0�Aط(Ц2���C"O5ó
:͚�r�'�>Q��� �"Of���'�*TDY��M90�f��"O�017,�R�A	P��7mfh�u"O� �e�b��P��7d�a�`"O�D"�*V.�b���C5AlU�"O�=Ze܋.���A�U":5Z�!R"OHٸ En���#R�T�*�Y�g"O��� ���A�,c��� r����"Or��� 6LD�R�rn��k�"O�=[�럧��<{7�8=Qr��"Oؽ�#�	K�x�*͸D~�Xd"O�@ 3$@�e�du���%_����"O0�Ҡ�2|ε�
W�l�&�3E"O���b,�f��UkEgR��jm�6"OДI&L�g>r��F�L�D�/�y���&Qg��xsIĨ!=P���g7�yB�;)x؄�U�>gr�Q&o�y�a�-Hz  �kZ�YL��1&��y��,{�Rؓ@c9N�@�еg���y
� V$��n�mz��f�U	$�8�"OR�+��ܳt7�H:�(H�D��*�"O�G��6`>��0H�:,�vH�"Oz�2�$�R��a��7#����"Ox��h_0�t����	eЎdB"O
D�u`�(%h��E. �c��H� "O�C�$�`8#���:�"�`�"Ot�K��[��KT�"O�l|�"O^��E��%V���c��BC�(��"O�1��M�)z���hҙ��q�"O~x��\5	�<�a�g�!.�\�"O����m�8a�EA�ux�!�"O�	����+�(����YUXpbp"O��si4t%. R�-݌K�@�"O8T�3���2&NH�d悓U4.�c�"O�jce�9:<.,)�")���F"O�!��Ȉ$�AÇEϨ�"O-j�b�)��!�Eh���"Oh0���j����CĹτ�C�"O4M�Tχ%K��iҥ�N2��+G"O6�)���
�j� �',�z�@"O��iZ��H9 !��u�^-���N�yR,W&:�r�%���r1��"�/���y�aьb��QC��f�q ���*�y�Đ?B��R�� ^ �\��P<�y��^B@�2�aZ�Of��� A��y���i�(}x�牨GG���KC�y���/��H!�T1E��J�-���y���.����4	!ha3dC��y���+�H7��J.ĕX�hǸ�y"ÇW*J�hVU�E%b����yBiE�@��D��<>H�9�#���y�DA�Y腓amJ�� ��æ��y�/�ν�b ��{� ���yr��"���v.��@8������y�c4D�v�*U/,&��a�H��y�7lͨ6�]63�`0�'Ë��y�CF�w砸(0�?-n�5�6/�y��:��#+U�(����H�"�y���?z4�Ib�ټs3p�-D�ա	�'~)�s��O��K���u�̅Q�'K�x�W Ɋ�,��g��]@�'y갱�&����c&�U&]�v��'��U�*W2&󪼩U�H)'��@�'Ġ����%�0�jpMǳn���p�'z,� �N�qJU.�:9����	�'��p�`D2_�`M�3眐-Rf�+	�'��l�%��Bb&�"o��)�'P�k)��9��(8$�º2�9��'j��ǝ>���da��b��E�'<�!���W�8�@���_Z�k�'C�IC̖&ǜ�ðj ���	�'�(�Ȁ��,]��X��JAu<lp��'�L��b'u��D�h.u���1�'�8iKԔ#��ز�ՔC��\#�'�&D�j@�J�{Ҋ�DMX�'- ��W�BL�:��E.�F�q�'�j��wʊ�):\)�.1 ����'O\�v�ٓ)pPMBD̞+q���
�'q�TpIb���_'6%��
�'���[��C8�E���)�줪�'�0��0���(�!F�SE|q�'�� �cM'����ր�Iƹ��'��u� �:p����5�6LnxA��� ���Bf�	+�b�+Ew��8U"O�e#D�2Jfx��gkY�YE�e1�"OT�C�A����
 J܍\X	T"O�9�:%��vҋ;�:��"O�,��΄' ��5y΅�ݼQ	D"O�:d�+lZ(���;<�F*�"O���e�(>���$,���8S"O^EpB�E�VtuY!Ι�`܊��"O>Xc6MDf�����^�VH�"O�%h��W�jϰuqd���uê��"O��:' �	f[uj��<�2ܳP"O�P���Η@�| PDH�9p��Q"O�QPG�V�e$���qc��8j���"O�L���F/{�~��C`Ix]�m0�"O�!�D uj� ��ZXv(s�"Oh��
�;�p{�I�^�j�iR"O�|�2h��d��1�C#��hr<� "O���#Oq����̣:� a!�'Fb��f����xa�ʌ3hx�R�'�8l�4ʏ�y8�ĢTY"�)�'�,a3.O� �R�2C�P�#����'n�}s��?Gа���>�M�'$X�
0�H,U��2�j��q�+�'���B��/O��B�?����
�'�@}�U)���VɈ�
ڋKzlX�
�'L`@�c'[��x�1H6�F��
�'�N���̩StJU	&���	�'�ds$-N"@"лF�4	oh�h	�'�K�Uad��p��Bo7Plp�'�� bR��6V��bc���dt��1�'MJX��� T�+s�K���!z�'yx�8Q��=j�!����@��'�`I�ਉ>HDɷ��+U�ݩ�'ObТ��U;J8x�wf�Q��t��'�(�ֆ��9h��;�UQk�(��'W��Z8I;T)ޓ^�h1�q�8�y��R�`�L9e�.L]~ �n���yBEّ*�,��G���0�ls�lC�y�H *���b��_>)Ln���y �.Vh��EGW�l�z���Ċ0�y�%�,+�&�Pi�����T��Pxb�7���):� ��F+��M��u���i��%BD�Bq�۔2�|���UP�%�v��"B쌐bm�ȓ @%��>(�Y��DP|��%��
T�F�8�"9A��X�H(\��ȓYF`PBl�%�X���Lt�l��=2��P�!W),R����NY뾀�ȓe�a�A�P#%�F|0���d�|�ȓM�v�����=�-��ǁ*kT -��ϨYX�@ѴH���b���E����ȓ~u�mkӊ�X�;�%L�x��q����l�7��,t��D��� =v8ͅȓ>f�V�>���U��'�^I�ȓR�P| $ �,)��aѢI G|`8�ȓ�hu�⨟�Zs ٕh��f����zy�1)�O�15j���a�DT���ȓ<�r���ޢTXd5����1~�"T�ȓg�4pAfX�Q����+Ү\�襄�Lv�{vfB�j���Z�x����ys,Hq���~Z@�B�n��%z��ȓ$u�e�C$R�}���O;�dD���R$���� �0����1.R��ȓ <��"�`�l�����␄�S�? ����l�q� �L^�dA�,o͒����s��K��M��$V/�7�R`P�%D���"%ւ�Nq�Ɗ�����H�Of!�pn&Kb� ��9k��5@D-j՚��%w��䚓@��ă�.¢r �v���k���P�i�`h`�̌��yƅ�,�,CtN�Z5��JT���'�\�ZUʀ�3)r�@A%9ʧj��a<t!4@Th�gf�!�ȓQ�"24��0|�l)�#m��"C�Gz�����<��Pa�����*��
k�a��ĸ�� c!��71;dQ�'�3c� ��q�]$H�u;�C��}z�cf�:�az�.b��!�n
S�~�´�M��0<1UNQ�q\��F�T%bԑpw	�1+8��E#�?2!�P��75��S�:�C���&�-����'L����-obS�(,鞼����Z��Cw!فx�N��g�&/�B��|T�"g�׫Pd�SKƥb�ΘI���tl��ae��'�hD�,�IJL̓v���C���|�qYc��5Έ���	�#��E"#���-�/=A��8BX��B@8�!����k�Y�q"����ՐV��y��]=M�.	:��҅)L�����5k�,��7霧D
�aҀ�H�"�B��B��|�h�A���b�(�#�^h<yǣӴ(��P��.��2E�%�OS�<���$�Ttq�D� D�.Y Ò�,��@���	�!Oq�S�P�G0��;�h	�:�!���%��h�%��h/,QWgQ�6��e3��PTdI�ւ�wx��?��vŧ�ēm���"�N�C}2X�	d�����`�����w�ȡ�B�!T�P�#r��{r@8
�oݩF'
 :U��8'_ҥ��'��\Js���T\�E�Qb2������y\ �qCIB�s%���6�O�6�T��'8������
�v$���, �
T�3O�u��̸}�� �M���!�i:��!7O��f�=�P�U7k���pc	�u��	 ��\cx�Ŋc(�!3�I����({H���''�U5��g�Zd2CJ�a!R):��Wldx ���4�̕b��T!����2l* �Au�xr��+�q���[�%��	0�%ھ��> 
�5y4���&�%KQ`QsC�'(U�Ue��D��d�ąA�3:nL��EߔS��5��ɷ{:K��P��Y S�1���B��*G���h�(��r�6��bPN@��M��R�pa��Pj3��@�c�&EHP��O =�"�ךl����'ؑ!.�c�i]L�b�T��0[��D�Ej�$2t�D�7��c?�X�t����eϴ$� P�d��Y�B��
B��p��Y1����j�y����Q$�$$��#�^��a�7(�~��A��1O\� ��[�ֱ�bn��*��`P�'T���@�ˉ-��*����Z�Q�h��`2�]Kŋ(V�V1����<��%�$��X��dF��U�A	��wp��E{rf	;:Qz$�!��;g�b@bcd�9f��	B5�DX+Q��x�$[	l!�$&*o0,�AEޅHA��S�CK�x�DQ�E�tX�w9����`��*n?h��	����~2��r9D�8�ϟalr 1P.�P�(!6�S~B��
��q[��䘦3��U"1.�[+4����ana"�M1LeX}I�AR#`�\���/�.( ��D�E&C����@"��!��Q5!�RB�	xؠ@����~��8��<N,B�I�Fx�I�Ga۝R�d��(H�(~�C��� O��=h*���+���C�4]�Ҩ��(�2����.GLC��sG�̊��:t����4C�ɷ0�X�1�M	��b'�ߢ|�C䉓[����bM 7=~��ȳ	{�B�#,�hJ $B�]йsG��8�B�	��4p�ЂE�*����/á)��C��8�>)*"�[�`�*0�H��B�	�9J��GO[�NIp�� #�"�rB��	�1�b� XPٰ��]�C��'3zl���
�2���h^8P[~C�Ɏ$��	$�˿h��$��Z�`ÔB�I�*%@�8qJUB=�pq��y]B�	S@ <��Z�#^���\,C�ɽw��: ��l�敋��˦02JB�I)N��RE�/e�Y��\_�NB�)� (�`�G'�t�@���4��*&"O�@r��Q "Ȧ	�%̀�$�\@�"O��2d��A"F��+�\�"O����!ֵ0#�Q1BC	�=��yr�"O*m�e��$yx�t� �#��Y@d"OF�r��V�8�asGYF̶�"O�h���}梴:�EE�Zo�3�"OZ�˵n������;=^����"O�L�7I!.���`�b�<�)�"O�4���}B
(r����$�9��"Ov���m����P���A �xp"OЄ��#EL?�����<���"O|[�,�-��0���0WȨQ�"O܄S����gy�!c�j�A�T��t"O��2Psy�!�����b�"O|)�F
�PKL�{��m��0�"O.��N��2��f�b��V"OhP�cF/r�)���p�Y"O��QOӓ�r�j��Y3`h�3�"O|�FN�<��`����k��"O��s��\��(s�B�=��3w"O�I�Q/��'~*@�
��� R"OIXףLy-:e�&D#?�yc@"O`��≋'p�|�ɐ�����Ӆ"O�A��e�(+w2U������E"O������+����GM��x�"O�|�t�#ͨ�{�H�? �a'"O*��O�cT"�2'�j�b  `"OB(0��_�|=b�d�M��P�"O�X =d�8D�cd�/U�%��"O���d:g���I�N��� 1"O��+E��/q����H���R@"O��f��;�6Pxp'_4)�2Ys�"OFـ�`�1 ��%̎M�´�'"O� Rꚹb�H�k���6��	P�"O* ڡ����d��-�=}��A�!"O�}�����,,)'ԃ^pl��"Of�+ ��Z�1p`(UT�T"ODH�@A� �	�ζVP�۠"OT- ѣ�*$)���1	�_/4y"OhX5k�\G@)
0CG�sRX1"O����S"0/}�Sdֈ^�u�W"O"#ŉ��X������O3D�h��3"O����EJ#s�R�Y5�?�b���"O�8Je��� �Tq!m�+G>����"Ou(�O�uZ�yꇬ��Xh�"O2A�p!�-O�
�k�mX5[��b$"O�\�����X�;�
p��ܚ�"O(�"�8)�Q����E�4�	�'bQB�#�\1�5��$\�b���'���!}���Z�bI��<1�'T�S�(�?"f�ݻK�m��0�'��س5�^�C�\�&��=Y�Y�'��h���/\�붣�Z�d �	�'Q@��嬎�q���V��$� ���'c(H��G�)���Ŝ�����'�j��6�E��K��s(�8BLGH�<9UF�5[��S�����'��E�<�6l4��!ՃS�2���Mu�<�?Y��HrM!�,4��ȓ*�j���l
�L����Aʉ �̅ȓ!�d��(�7u�	r�/J��`�ȓ(%�����'�^4���
�[���ȓ[�h1���qG<�@	6dbf��S�? ���H�<4�2���`����B"OP8���V�9 �ʵ�rd�c"O��A�Aޥ����A�T�q+"O��J���!|܂UAx	� Ϳ�yB [�(�2�0 �:��TDH�y�H�5G��
a�nY�|���&�yB��`E���pD�*Z
Th3̅=�y�
8� @��̝:\<11b�B��yR��mn�ĐF/Z W�X18����y�`�r�,Q��V(�	�K\#�y"�E.]$J��� �[Ƃqp�ƹ�y�.�.	B��D�G=D�<�8�F���yR�C�-�ԵxV�G��,���Y��y2@Ž6�4T��j_A����C$���y�&�rǦ<��D; `2܀��M%�yb�[*P���"�ϗ�y��Pl��y��S9�Z��R�t�tWN���y�A�<0^~9����o���r��Z��y���\��	h��[W9+V��y�$
��y����8�N `���yB�L�L`B�&H
4<�3�ό��yBlX��o�*O��EI䤘��y2��7p" �Ǡ8` P�#G�0�y2��*s9�����jWQY�\��y�d,+���bi]�gR� 2���yb�G�op���ҧ"M����R�E�y�L���P�5AR�|3���Py�GĎ/.:�0G(_�Z@���]�<ya K�	�`�¨f���b_p�<9���
B���A똠
y�-hc�l�<��i�%E%0�SA5Xz`:��S�<q�G](#��y��D�01^��7�P�<)�� �1b���#m\4F� s�d�<��@O<iJ�)��Θ�^�:��T)�a�<�E1Y���R��]���'��_�<y&#��.��J"�ײ5����n�Q�<aga��c�����gʱ}lV�9�.�S�<�fD�v7F��*�3`锌�!gLI�<A��S��z�±D�qT\a�ÞI�<���1zm��W�U�Xq���^G�<) g� %-<��@��f���1��G�<���~��:�Ɗ���u�  �<�BO�$<�K�`X*[��]�ZA>B�t��g�3~�@Q���%��C�I�a|*���(¶3�ʼ����iyVC�	�< �P��D��H�0z䊞�K]0C�ə3m�ň�E�;I��D1�\O�C�Ɋf��Y�s*��$SN ���L��B�	E��q`��D<D��D)�B�e�����e���1$��o�B�� _�<���^ ұ�g`Ğ*v`B�I)<P|1I���	~Ϧ%8�'���y ^�f+�`�	Fp�D #��y�F�*'`X�x4h�_� �8���yB�G�Y,�l��� ,d}cSO#�y��/�J IB�U�uXl(��Y%�y���3ͮ�+��׊�2�bcߊ�y⤔�/`ډAD��5u
Q�%O[�yb@g=������>5A��HՋ��y��)MR��aK[�>�<�;��$�y2��*�b��0
�cc��`Ņ�y�k�3yۦ�ˇ
R����
��y	����[u& ����>]�~��$$�5jvmͶv4((�%ǹIv����S�? ��P��<i٬�{T(_+�(�@�"O�hP&��5�H���H4d���!"O���B�"^X�h��ݖ{�8��"Ojl����0N��,¡E�7
���[�"O�1)q̊�h�B��)O��Ӈ#^�Ũ�Ba��s���I�.֖�`�
-	Yz ��1D��ʖ(Ok��@B�ߢJ<]�S"�Oh����&�%��Ɍ|	��p&C�*����.�:{���D�Q���aoP����L3����*P�K���@	6�yr�J��|c��JJ�r�y��K�ո';��z���`��"�[��(��4X7�@�Q�c׏��B��N�!�D>[��9�fI�$6j����V����e�߁h��Y
p3O�-K��3?Q-��j����U�X��Bfj�d�<��߭����l�Nz� q�#:c��
�/�$�����M`���W�>z�U���+ �`R�:O
��s��w�pa������jJ�^��{!%̓!1D���"O��`JA5D���i$$��\���/�&yx����^�!K4�jp��M�Ob>Eb�)�\��6�Z��VE��'���ѐ�W�V�}@�MR�k���s*��
F`�#%Y�t�.���Jۿ�ħ�1On �a�6x�͒�M;w�84W�'�E�� ��)Ѓ��(��:���&\~���9#���Q.@��ԅ��^a� �����}�|�J�C%�#>��L�G���{'o�-W"�\�T �#(��D���r���{S��,|(�Lq�<!E.�:��}K�Ƈ)7T�7.�:�y�/]9l���hU��������cG�;§@�q�&Nס_�v��c
=g�d�ȓ�LaoF�~�����2��Q@���p@��,έ$�2� ��Y��OY�ژ'��81q�^/0��� H.g�41
�f�<	2̐��z �
��&h�"]�m���J# ߰��qn�e�j9�ӓ}�ي�AʹK�4A9E��
H4Ez��ȇ=�|�p��L����`��"��p؃�������A&�R��GU.xB�It�r����
'mԑ��4z�V6M��3��
Q�=�H���	��(��Ik��sCn��g܈<��BB+ �f�j�<�!�E<t�������(CVp���#�B�;��J�{~Ʃr���$6�� �O_���s5�.v�ub֤�%QZ��0����$�!V�5m"�	�4?>�W'A8�r���bݳ&Q�H)3��?ss���	>m�N�zQ.B.7@�qS�C���HO~����] �y�5f	�k!l�y�F��Ꙙ� "qN�D��M&0�2a�]c�<��O ��B�O
�(Y�B٦�����^�}jQ� �!��p`�.4���\c��5��hZ[9�H��g(?|���'w�9a%<��\�F`�֊
 �^�U��ٻ,L'l��9�͙���)^bb>㞰!1dT��,`��&R��Q��+�O��+ ��2-���v�-~�(��D�
�A -F�i�0��� ǈ1�B���'�5����ZY�4��!�/�.�C��D�?Dft�e��)J�}�ˇ�	���1z
��Z*@m����#���&C�I4\q����h�Qj�	/�"牧��yZ�J��ΐ��o�5^#~2���2=�E��i8���fǛ�!��%_}���Q)׸I��AP�f��p�@[ê
�\�����'��X�`�<�619��	.�\@��h١$$&b��P��1 Ә��5�"5�h�0O��"@ÈV[�$����4p�"Of����?8�r(;�D	�P/�lҦ"Oz=9g�_�pJz(���B<YL	K�"O���/Ӧ8Ul�iu�M�k�!g"O69֨�:JR=���B�`UEA�"O.��A��Q���Ϊr:���"O�5+-�.��0���DJĊ�"O�@�ӄ�6�Mx��VM�^	�U"O��bq�ލ9h�t�[]q�s�"O�� F��#wz
��W�i���c"O���Ԅ�M{�M���}�;�"O�餀�y�P!�s��f�d�"O±0 DD;G1�%X���@��[!"O,(V�љ�`Id*��{���yF"O̡1��� qTE�ǃs��P�"O� �;q/��,D�$ce�}j$<A�"O.�a���TJ���ė�Xζ!��"O�H�KL/Ti��p�F�L����0"Ot���!�;I�Uk�H�L��5U"O����0`H:d���c&�s!��(IqRHBĦ!)Ҭ�'
���!�dG9�$Ub���r���ć	�!��7D�\�Hē��:q�A�3L�!�D�$G:���D���"W�.+�!�t>��!h3'��T��O !�!�J�i��m�G�"�����0�!��0�Z-� �S
{���A�N�~�!�$���< ���~�@�Q�
�-X!�d�'�b��l�Z��Da逡q]!�$�2o�&%��B֠��i8�cʗf�!��g@B�z� A�n/\���*_�!�>$��x$Ƹ<9&8�bU�X�!�$�&7����!�1��M������!�#!MD�����N����*%!�$ձXUP�:�#����l��o�x!�d��l}3Ck@=p�Bqq�'\�Hr!�΅?]H�(3�ҧUI�E��!t!��7��z�fӆ�0P(@��cc!�O2:l�Ƃ���LBů��^!�DZ�y�¼�k��nHd��.�G!��
P�a�F�ܽk��QQ�3G!���nDu�3A1>�0���.6@!�$~��ti0����01���y
�'Y��� J�@~�PQ�g�	-l!#
�'��u෠ͭRa�����"����
�'��0%� ��W��eP
�'���@�-R<f��92@�]���S	�'�|�(0^!9p%@�Ɏ�@��#�'�r5y��\�8�ቱnϾi�,� 
�'���r��O[
4Kf����WN�<�"+J.v8�	�"�d���ч�H�<�0,;mbPP�ᭁ8z��`c�<���7¡:�쌍>��9��`_�<�e"�qٞ0�1!Wm�<�e�V�<��C�*R,j��G��"&�9��řh�<�AO����� 3��*c]���Q|�<��,ȷA��!�
�Tq���Yb�<قGݩY��i�o��0L��dNd�<�E���%)�E ��[3�"=�"C䉭��a�"�
�m�m��Cb'jB�ɭZ_n��F�]`������FB�ɓm}&)�̉�^��f�K�D�XB�I)��)�qX#�^���	q�`C�I0�}��YO�젳�Ec�4C�I-2e�֥�@U p�$�U��B�
]�X)&E	X��9CӤ04B��qnz1"�M8n
u0��U �&B�I:Y�\�V�E nʈ|����&1�B�ɬ"C�l��&�?03�,��L�Z��C䉬s#J07ݞg:J%F��+��C�ɞ_"xqz1��9!.`CA��l�0B䉋�VpR�|y>(ӒM!�
B�ɿ`a��8�"	S�,+�JZ�1�C�Ʌ_�����NڧR����$WQtC�� $�pT���]CA ��`�]�?��B�ɫz4��Qυ�!࡙�[�B��#��DK'�W�R�^8�$A�aǄB�`N���5.��`�Q#}9!�$��^�*�D�Qb�4��a��"O� >�x��2J�X��F�r�X"O���GƔ\��=�U�ֹ�Ea"O �bb��� ��F»"	�]�w"O�AHviV�r������*"�d�U"Oh5�� .^O�[�&S�K�n�ٵ"OT�r"`^%���4�Q�
�L82�"O"1�P�a���UH�Qi� ��"O`�ZT#��fԈ��W�VKs���"OXȫ��	�d�� y¦�-<Q���"Oh�h%�C�}ب��$�$DY��"OvuA�?v� ���▒9G��G"O����D;T���W�iYJI9�"O���Q�a��q+��7�(�"O��(�nt�B���+[�T5�b"O�ݨr�߀4��|p2�G�gǬ���"O�m� ��cvj�����Wʚe��"O�d0�N�$y=8hu�)��\��"O�h1.�;g&�0a�Z"2�x��R"OЀ:���Q=�H�)H�2���"OP�(�(~�j���GY�(�]["Oh1�I�o�lR��]@�ި��"O$A��K�m��\ش0��"O�y�v`̅'�؁��G�[�6�"�"O�`R��$:AL�+�!�S�L���"O�]Wh�f��Y�f��
���d"OmH�jӧ^ɐ�
�Kǉ`�>ݘ�"O�!��j-l
~��C��m� �"O��x�c��3�^ ʷ�&@z�F"Op-pԨW��v�o˝IF椈!"O�1#�OI(��,���i��"O�xPR�� (�qE��gR`2"O޴���H5u^�)���F�ıB"O���kÏrW����T!@H��{�"O~�"*H\�Z�qA%�Q!�Z$"O�i��
]�&2�)dd�LB�(��"O8�p5k?+
D���	�l ���"O�,��=-h��J5��"ON�{�g4z݈�a�BK"7��Y�"O�����0!hmǏ�3�2�1r"O���V���eՂT{q��$2"O�����?���{�kހFOB�y�"OlhP1��l.���ʝ�+�8�"O|+'�0U\�-I`/,����"Oz�K%cM�&�jA򑍈����"O2P��l�*�@���"O��҂V�|���������6"OR@�W+U>X]pa���P�/�T�@"O�u�ޥ�ԥ�$'G�n�P0@"O8�	�f,i�@4 ��-U�ř�
Oʸ (��*����v-�"�x�`�&�=�~�.G6��'��	��"��'Q���&��+~��!�"cW#)� �� e�?ns���J<���|�A�G�Kd>4�aa�*424Y�&e|�T�#?a����0|z�k׳�:�!�V�=4�� �C8G�t�'zj����ȟ�F�M�Fe>#4ΙDS��±Ǌ
��Dܳ��9�C�U�)�'k\ҵ�W_|b}���G�p���]�z!���i!�S��yb)N.���X��Z�o���kDM�q�P���.��۶*��c�ۤKO�=�������U�Sta�Td��Y�@�#pKO��&,�������]�?�%A��������$˟A�
Pˣ+
��$�r���M�#��@igA<}��i�1[K̔г�Ď+*qcv���3Jt�	�=�J��Q��Y�Og���ħd��b�W'�ޤ��-gJPY2�`��/�|�x��m�vŰ�lI��0|�E�A]��8�dO�h��U�I _���5�m��m+M]��H9ç.Z��Ѳ#�!7ݚ%�cٞ��E�t��2�F![�� r������|֧���[�8���& �RN��s!�K1;��Q��-��m��a\�م�3� (9���_9��M�PjB�,+��;3��3o>���'���Č`�g?�O�NB�KOe[BQ!U�*	5���`�b�&��	�3�
ԣ�*G2����ÈMt�O��� B3�)�IA�w��U�g�v��y2� �>�'��}:����3ƚ����~��.I<O��I�X#6��?E��H31����/[�e%����+�?�C�9��������1"�P�z"L��.b8|���S�+��+��	]�Ot�i%��U�����5���^V!��%�̌p#��+e`��u'��L�!��+��������X�!�d	=B�`!ۉ1ɤu�$J�r�!��V�[3��1��]� v(��䀎D!�ā�q>�Bw �]dYÑEG�?!�$�?A��:p���\�T�ڃb!�$�#pbE���B���Kvcʴ+!�䖠\0N��l�Y����%iJ<V,!�\�m��YYp��<9����!򤘚c���˩J���%G�4G!�R�xF�X� I�C^��!��hS!�d\�a����kX.M>����i�x&!���|�Y �{= ��$��5�!�D:>ɸэ�H5($:C���5!��q��$	�o�'SqD���!�䁴H|.Y�c"�� 4�1���[�!�A�2���5&U=ED !��I&:�!��I+(����dOY�&V����a̚C�!��E'T)H�ɠ�ڞLV��ѡƅ0�!�d	�M�@��G�]�5:�aH�o�4�!��3iL�a��\#*$.4����/�!򤁤I�T����'gҌ��lVlq!���ARCC	�<�Z���GY!����9bT�Q&\�L
ӨJW!����������4֤`kt��6Q!�d4Wt�Z�:9߮����ҏ=<!��38Dv�sp��Q��5�f)T��!�d�gf��x M���	$h�!#�!��:dl�)��O�P�Nl�$%S=r�!�d�z���ࠜ9,��L:�"T?��򤂇"P��R�K�L �a��A��y�(v��%k񉔁{G��R�l�ybKO���y(�.�?&"��Bu��(�yR`�^�X��3e3,Ӿ�D���yR��%:�d �I�mb��È���y�-+%" 3J�h��P�C�y�
��_b�bq�\���|{�#��y�׮J�$�P��|����di��yB� /�p<Iï��l��T`D̏2�ybj�5��!y�̟�,n�d$���y�(е�a�#鐯3]�pl
�yr���gT\y�p�T�yu�0�d��yB����h�U�D�FY�s�܇�y�H#~�L��DbM�4��H�b`��y��ݴ!p�y�3L�9�gF��y�-�/l�r#f��<���0���?�yb���uU�d���߲*q�Eʡ�yhL����rA��h����-B-�y¯R�b �f�B�o�Ȕ�dC���yr�)a���D�~T�4Q��y�͘�p��!q"�)InV��T
�%�yҊ
��Hفq��-G�� 4��y2�DeF���镅A�ݩ����y� PE�$�ڐ�?N&!�cN̈́�yRGIc�����������)�yr��r���+U��jq�Ǫ�y
� ���%d��(�b!���9W"O`IQ���d�����:q���W"O
�ە�ˌk��-�P�@�P�Z"O�@P�m�%v�0�h��EX�"O����ʈ6���bҴj�^�a"O�����Ύ,��l�R�V��^|��"O��H�A�b��I*��6z)����"O*ܣ�,ېLO4%�!�I�JI ��G"O�Q!@u]©�b�/���%"O<��4@2��SA�?&� A�"O (9 �:r��`�@P.���b�"O���D�w�<[�.�o��10P"O<���.T?4�bU;��I�s��b1"OF�9di�=@��m��	 ��i�"O��K��,.��#������K�"OvpV��C���9�iC���"O.�g��C��|!B�
�'s��;�"Op�B$%#b�k&S4�S"O�$��E�;Yj�%�2���"O��`�ڞ��sD�9SF%i"O�D��i�i�JA�!D��q�0d�`"OR�a�,B'h�|̡��
+���E"O	�a�q�!AE�8c�쪓"O��F�܇YV���R#Vc��R�"OJ����~1*����^�fjZy{!"Oʹ���" ܨ7aA&����t"O��%e��7- 8�v/�Aj� "OHia���m�N���jLX�k�"O�R��܌V5V�
tN��\1X��"O"\���L%���Ԯ�!+��a�"O*@�p�C�q�����F)�l2D���e�{!b����
�C��%D���&��j����X
s\�I�8D�t�V��D��ey��I�p��+,D�T*@%Y�B���'�F m�^-a'+D��ˀ��"E��iD�q4.eZ�*D�<�"��=$���C�Bd6��ʷ$&D���'ʭr��Q{ǊA�Fu���4�$D����e��3�t��ç66cʅ �$%D�p�%R�
�8��&��#ӠA��(D���A�8��͊�;7�( /2D�8�5!S�Tׄ�k2��~^!���.D�T�v�F!l�u���,S�F9 O+D�p�Q� �y?�){D茅?h2�A�*D�$q��T&Te!�ʍ (����&D����I�#F�}(Q�J�i��(�M9D�<2�aMo2�����G'4��I*D� ���0ec<�3�	 �*!c��,D���[)�r�˅�`I>!�re>D��PTG 	2���Q#�<�k@`<D�d�g�� NQ�MT���X�!<D��y�@�&W�8�ǀO��1X�$;D�4��j��m��X[lϑ2{n����7D����$e�,�B��Ȗs�nY��#;D�����2_�(@n� u��E+D�hT'��l����&� 6����	+D�L��A�y����jǉX/^��d$D�h�'S9	��ۡhĠF���{4�#D��B�L�l�hU�\�@�	S�.D�̫�ɓ�^��t��\�!Ql]X�*O4��V�|@bŮ(sR��3"O���Q�p�4��W���5"Oth�#,X t� ǎvu�Q"Oz-jdKE;~ �&^�Q�H��w"O� �M`p�@b�l�`��0
�h%�u"Ox\#��J�S@�e��F�^Q�u��"O�����o�&�q'&�3��YW"O��kW-	4���p儥`O�M�Q"O6����ŚQ�hsF�67���"Ot��� �t8ѓ%�"BTv�h�"O��;"h���M�7��%/T�1j�"O��ペ�ss�����ЭGI�dB�"O`YAD��:n���Wc�W>N���"O\d��kɝ ĺ�*��6�EF2D��:D��oGDP�� �]���S�I/D� �ƏQ$�`���<S�Nt�$-D�؀���(	
��xW�V�FAN4�w!D�p�T�Kj�4�*Ӓ�0�c'I;D�4�3��S`�p�#.�(R��qp&�#D�N� =@k�$+s��S&D�:G�*B�'�	7$S� ���i��H��C�ɫ.*��ِ�G�U��l@�'�*v<�B�ɼT�p y�5z��H��P?YwjB�*�L����[mEx�H¦�u?6B�I�e�$�q�*E�)0L�����Ӎ��P,��j�"?�N\B�E�1�����Ĉ��eO���ؙQO7�@��L�\Y�f]pI�=�V/TE'� ���hbB��>/��}�*ܾ|~ A��q�,!b�ʞb�֜�r��:"e�ȓWtX�Eӕ+���aN�Eq����{]�ŹS,��=p+�'�9m�,Q�ȓ*]T5�ʺ�4 �5M�9�ȓu̍Z�AW�}gh�����gDzE�ȓf�����e�W�H��S0;@���t�B�HviO�,j��:��� ��Շ�'��:I�8���X�ĺBD�ȓv��$aׯM4.��� �+E��d�ȓ�)���4W��Up�N8��̄ȓ�Z�0��P 2XPeJ��5�ȓI�
���E�/��K��J�(ҞL�ȓZ������TZ�!����=y�@�ȓjb��k��G��F1Zl�� 0z$��b���BS�W;��J� �]s�<�ȓj�*���
D�\���D�V��]��/�E�Bߵe��y0�]�WG"�ȓd��s��º8,vu`%+\4A�&�ȓ/eL�8r�[��L�k�l�����'��Q�b� 2,��E�v�|���'&�<��J�	@L
v-G�:��|`
�'�L�Jeg�*�	jr�ֳ4�� ��'��T!�(ԡ,L�Hr&K��X�'��� �-)�ygaZ;��H�'`��v:�taejH�c�b �'F	*B��^����L
c-�X��'N�A�k�5Ċ�aY%UEnu9�'�&��PE�&K��h	�uV�)��'��l"���TM ��`�
q��$��'x�)V�*��hK��`�j��"O�xp��^��d� a҆b-R �"O����
��� � F�AyV�0=!���z� �pJH$	U���3��8!�䝣#�K� ҌD��tB�b!�d�q'Xp2���E�X�cv��\�!�$ɶ]P�R��$N�3ҧk�!�DD4!JԩRQ߷2)��'%��zl!��ЍN\򣊀JB���#ģ,�!�$�~ �P٢�Z%H��a\ �!�� ��bB�I,[���b��[d"OL�Al�:c�m8TH/K �"O���fBh�Y(�7.��#�"O�$�����&>���f�(~2��Y�"O8DP�AU�D�>��3Ő!N$�t"O6�`g�ѩo��j�Ŗ[I�a�"Oȼ#A��ڮ�	B�V2: `�`"O��ق�)�����N�Ƀ"OL,@�h��3vܼ9�C5#u*�(�"O�]*�F�NA�C`��*W�	v"O0�PpI]�`Pt��J	 B:&�`R"O��J�)U���гÉ�=P4��"O����:V���	aÈ-�0�q"Orl��
�Q"P��VAf����g"OFQ��ʀ�����/�h`I���O2R'�/�M+ϓ�M0J��f��@FJ�C��Y:X�;�(�U��7D&�R�.�%wN� j�*\�.}	�r��1��a�G^0_g��37�W���P�I�{,��D��B��!JXw��	� ���'��|x�^�$�4O	�:
.lJߴ�j�4!��`%�h&Eۂj���z#$���
%!0}��'w��O�9��Ãh��-���tG�Ӧu%���ݴ�.O�]S���am�52�^]-��M�T��;PZF(��/O:�䓙
��Ѹ�⑏
���z��D�-�DH��"۽�} ��%Ր��RlI�,Zy"c�ɷ	���hs�[�H��C��|!�h��fY����)LY�ͣ��[�C�����	��'7�@������eX��KC/ž m�-Q�!۞P^ұ�O��$�O>�O�˧��D˅*n�l����7=`���,ғa2!�dUl;����]� <HQP�l��0#V�i޴S6�F�'Ҷ7mA�;��o���'A�\�vءf@Пa&��BW"؎ֲD�s?}��'"6� ��D'�����
?c��{�$׍�\���ZU�)`o��NU���#Щ#��$�>a�l� ���q��1��Ḱ,I�@�L4�`"XϺ{�OW'hˈ���)$���
�GLE�'��	�ɟ�M�i�"���h4}�b���75����%F�|��˓���O>�iz�(r	N�<���s�L*0>pu��I즁�۴������^�	FL��F��4mW4%l8X���-+ɛv�'�i>!��\�^�Bu��Rt����ڒ^�����}��HV�i���Z���"�[f�?u�S�D+�.�rK��9s�-��d��eh�}Z�J9M����p<l�)h��ܠ)xr��U�^��Hcޙ�q."U��|x �K[�^d��L���?�7�i�ʓe��D���߹q%�۲�Vm�QfO5n�8���L��?��D�<�Н>��+��D����
�m{�9 CO~ܓ8қ�Ck�v����5���?������a'm�$wX4�6��_,�0*���d����M�	ϓ�MK�HCYh��䉑(�Ȩ;c�ҿ.p��8��\��Y��ς:(��K�B�s-�A��B���lt4q���4F�ѳK�P`��S� ;5H�	O	�""`ݱ�e'����c�((���s��f��)$��"r�pQ��',N7-{�	�����T��)Z�2$H�Q�6�r����&���'%�yS��5��`8�Ë�LenȰS"
�]$�4h޴��*O�đ1�E��oچ%�����?$ܠ!��E�Cwt���O��1p�J��Д��kφTpU��
�vPPp�çC%b�Ce��W�J��S�I�2�Q��P���p�a�Im�0M�C���$���e۾@麬�T�^�?q�aqG�'1Q�y��O�m�7U��a�BU�sf�%�UI��&~~�ޟ��'����?�m�5F}4�ѐß,$v�)r��!��B���՘עR�t��"S� ����G�P11���|��`ݍ�IN�I���#�O   ��   �  }  �  W  �'  �0  �7  *>  }D  �J  Q  IW  �]  �c  j  Vp  �v  �|  �  a�  ��  �  *�  m�  ��  �  ��  ��  Z�  �  K�  {�  !�  d�  ��  D�   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ��N~��\	?Cv@ӎҿF��(8`����y�DG�|�mYDG1E�>-��'��y"	�*]�MYԤG,Czr��v���y�M��ۗU�~L�S�Q���(O�pD{��D�� o ���G̿%�v�K#�^��y2'�q�
�1N	�%uJ%Qq���y�ԆE��,F��H���[�y"�C�@�h&��5F��8wFU4�yb���B��|�g�Q{I� �&.Ҡ�y�a�3���C�'Ǩv���p�7�y2�" =��9��H�vVXt��kA�w�t˓��S��?i0A�x6n�ڡ��L���˶�t�<ѕ�צ2(=����j��{Ro{�<yF7BX"ɓ6*��P���Ã�Ju��'���%�B)ct��և
?��q��>D���%,]>d�h���K�S�z5���1D����`@����yge5R��P��,D�,�a��Q,�|KAI�
Ԏ��a�+D��c�����0
 e��0�|9�4B,D�Lx�U��� iL]LifQ�@}�
��'��|r��=z�t3�e�rC,�Д����y�#Ɔ_��,�!eO�ky��2�G��y��Ӓ0j����֘jЎ	h�/˘'�ўb>� mI���"��M�'� �o��'"O���U͉�P A�sFQ
0��!�"O@�B�¾?l~�ѷ�ΝpƂ�l4D�h�P�K�:B�`�e�$"*�
%D�\ɐ��y{�yc�F���M�H$LO��{�{��C�R��x�"�"D�|�y3
[��y/C-�n�Z��ȱ<M�9��+	%�yjE�R�e� ��Q���K~F�C�-,���7��>f�y����3H�C�I>�0��A�W!���'�A�A�LC�I(B��r
�.Ml�+d���P�X7M1���҉@�0�Lqɇj�0:��%��'(D����оPX���G�@���:&*%D�� "$�v*���#K6���e�.D�|�֧YM'Ĝ���J�x�,�(�H!D���F��p�@�h�u�2��W�?D��"�)/˶(S҂ܩL�52?D� ��DT�l��c��4�J	h�:D��X��W0\�l"��5��8�@6D��p�Y�\fp��7=ƺ��'D�,��,G.��� �_4;�h�Cv"8D���`қ1�D��1��m�Vr�M7D�HBwf�u�\ �[�^�dy�ƶ� �
�U��Q�5l��kf�j��t��W�`� 6��{s0T�6����⩄ȓ=�����"HغT�R�6�X��G;���c/H?52�*�%<;��L�ȓ!$l
g���p"���.@��	v����6% "��OŶ�$��`�f�!�+'D��5��2H��)��B�L�怣<�'�.}�U��&?�������!CG�W��D�R�C��C䉱]��Cď\�a��U)P%l��O����G�U�������;��Q�re��7��z�d�9I������8�	�dJ�K�!�\2y
�PB�O�U̤Q�����'��D)�)�S+��!�i�(X�܈��d֫w"C�ɺ:g:���	� ?��Q�ĆF���L��'U?j���
x��	
�ÝI�����(��T�2��8`�V��� ���{Y!�$�;R�d�/P�l�@�2SD��$3Q�,D{*���mCX��y4j�17x���HH<�$kԒW��6&�$.x0��|�<��G�:4Lm�T���PC�3�h��<Y�ϵ"L,�`Ҁ
F `cfH[x��p=	��yW�U��)U.q��I][�<A� ��yDA��D�I�`,�LLY�<�L�"
mN$Z�K��%��)jf��R�<a�ɚ��i;�d��X{H1J�g�V�<�C�V��h�ǩ�O��h�WP�<	c�2a�p35dU�8�4��H�<���X����0ݳW�Pܓ�M�ϓ0dx�Ч��1�V�I� V;ڤ�ȓ{ez���Ö�uVH�R�H�/��ćȓ#X�r�ʋ�W]zcܢ����M�ȸ�T!@�#����Q+���)�`B���f���.Z�6��a�'�YFy�𩃣E~�;p��S}h�f�Z!����)�wӳmV�Y�a�!�P�xk��"�P
��$�"-]�Y�!��q���I ���3b,�%|�:��ȓo�4�8��NP8�@@ c��t���f��6(��jP��X�Eܴ�ȓ��j�M5sn2i�II�$��a�he�`�W&}�R��e�O�܅�S�? b���H0��q�$�7I>9;�"O�Tb��ۨ,�D��;�N���"O�TC'��by� -<����q"O���)F�����,
�{v*�Z4"O��:㋦o�ja�d
<pf\T��"OZ��V��Frġ��K�O�\��"O ����W��8�é J��p�"O�<⶯B24UZ7O�i����'�I�R��x"D�2Y�(SN��x���&���yң�x���(^m��(�a�_��u�8�8�I�Þ��g
\XW!���*X�\����:���z7G&rn!�Ow��ĚF�=+���ӕ��(�O��=%>���Nɪx�����!D�!�:D�x[U�>s^A����.ZǤM�be&D�L[�.��B���� �D�8AdK�n&D��a%���j��X��+vu�y���#D��2p�@�Jۅ�;ռQ�A�!�y"a�� �J�B�3�X�ж��+�y��ܠ�B��O�$�ZUQV���y+A:/$�5@�H͹�qQPD���yr�ŏ;b�i�%���0Qh�8�y������W�T�s�j��IT��y�l�9�q���W�f���!�L;�yMX'(��\�G�$�:�&��yR��� D4cC����az����yr��;Zd"݌U���Հˁ�y���+�XH�E��I>晘Uŉ��y2��WM����

oӢ���n���yb�ЩX��(�0m�QH��bUJV��y�!ֆs�V;��*ۘU����yҍ=zE� !a�7K�����O>�y�9ܾ\����:pN��x���5�yB��'uS�@J�F;cFd �ea�4�yC]>�T)�k�(��)�q���y��ZY��A��a�����,��y�_�۸���̑4,���p����y2� �&�`���3� �7#��y� e;��$ȃ�
=$���!ڀ�yB�Z�u�l�p䒊�^r@J���y�L�:-��q��T�q���'*[��y"��7U�$���Au��Bn���y��2Pe��`��qȸ�v���y�撺)���K�pX��6*��y��VU��q�Ҧn4��q��y����-
!]�es���0j_;�yr�ɣG^E�`�O�p�52Ǎ�%�yE��'�D�C�셹W�ԑ��
��yE��'^��}�U�UkA��y"b�x�|�A���LX5Ċ��y�a���H���~j2� B�yR �$ln�дG6t����FD�yRBD�C��e�v,��ã�ʋ�yr"G�%���[�M�h�T���T �yR�ī>�������j���h �yR�7���h��g ԟ�y�D�P7A�(Y�
�+A`��X�'X�k�@��|����T*�>j�t[�'���K���6`vi�A�Cgm
���'/��H�bO� ���"Z�l�lѣ�'�Ȉ0#M�w���0�@�V0�0�'~��cFmFV�JɒSz&�3�'I:q���m���ؑ��G����'m���̙c���ʄo�>�<	��� r���^�k/i�c�ڶj�f�;�"OV���. ?��ɕ�۪:�jT"O2�!�g�� ��92���	$$��s"O�L8p�u�����l1���2"O�%C���\a��̴)�)��'�r�'.B�'F�'���'�B�'�fU�'�O{��P��[��1+F�'�r�''��'E��'���'��'��1����*��dCأD�⠢�'��'b�'�2�o�������X��!�l��r���2NT�3�ӟ ���0�I��,�IӟD�I��8��џ�`�� /�Qj��J?n= 1�mʟ��I���I��Iޟ������ȟȩ�ݦ���RbE�7����I͟�	�D�����I����	ן���ϟ(""�B���2Ŕ{�~����$��Ο��I�T�	ӟ��	۟��	�� �Z�@:��k�@�$���!��(�������������ߟ$�I��Ĩ����SE/#����afFҟ��Iǟ��	ȟ8��ΟX��ޟ���П� V�F�v��9Eh�z�tԘ����h��ğ$�	̟����`�	џ��I�PR'��k6F�kA�E�t����nY������������	�@��ӟ4����2e��1b���6�	!��E(5�ٟ��ڟ|�	ş��	����l�I۟,���(6I^Ve�Ǡ�z�Dߟ|��ߟ�����������I��M����?�"�6SF��g�����:�*[)����\�����ĆȦ���ӈkkJ��f�ZO
a饠�]u<�;����4����!SO�H���{o�JR��M���=���ݴ���K�=T�YrBG<���&o7��;��iM`�9�쟜b2Bb����\y��#CGQ�g˰o�)��]�c5@��4�d�<y���(y��&�H�(�`
(~��]�6���en�M3�'��)擏B	|�lZ�<�B�������媵�qn��<	�!�A�.(81�P��hO��O���@Lɍ8�T�3���0�x��6O����*d�������'}���E�B��⁅G�ph���m}�icӠoZ�<��O�����>bЅD�N%2�j�g��b��K��"T�5擪N�;V�e���@j��	��� K��Iiy�𧈟�R�_z���c
f`�"�J$&{�D�̦AaK,?���i#�O�)�-,��	��Hz��ҋpt�Ц��ڴ�?	���M��O�Hz�݉u�HS�B�s6>�ѵ�)d�t`��vY!��ޛ���e�+d�F���ޝQ�!�[�x����H2�6=�u�ɋU����g)�	.��h�p��&R̸ۤŪ�9w�Z(��ꊻ�f����́A��-��O�%�Z#͕*T� Mr���O���/K,(��#f��!������B���t�Ȟ<�u��D�6�F��Q쁱:�u�U"3=��D{�@�4>�v�0�Q�b_4�:�MF�hw��ϓ;����a+�d�8l�#�W����PE]�7�ہʌ-;���(M�d![��Qz��U`aJڷ9�b�24��_eD��v+_�܍{��"Y����V���˔9=,���s�ڋ�tу2g�#:Ք)���ؾ6�ͨ��8"_~��Ο/����߁ �1C�d�-r^<Lـ$�"?�\�Cd��k0| cdB̋,6>(���Q���?	���?YtV?M���v9T����n�*��1��"��҅���N3���-�2� 1��?u�RkN�Z�1O�I�C�;T� �1��K�<� �oX! �Ru�#�D��֌��v���1sx�}�&
�-Rr��R��q��;o���*�+F#���#�a�L����s��nz��Y���	qy"�z���e�_,kX�{�k���xB�'O �X�R����0f��a�h�=��������&�DlZ4W|��ӯ�D�|��� �z|x������P��a������|�&#Ls8�re�bd2$���0^��V/� ��YU ���i��m�+/�4}Dy���qxr�� 0w�I�5c�(x����W��y���M�������*׆2�O���'� 6�
 zF���@�!�U:����j��i��Y�|�	N�S����`V
x[ M�z���C�O���0<�����
1�HX'�	h ��w���W��^����`y�����'�?Q.�.��
V���#���ϼ3�l f����OL�������LF�mJ���')�VC��L�Q�	I�0=
T�܁�d�r�LL�f�Q��s�J��5o�)�$�{��@�Q�rE��uQi�F��u���^nȀs���J�Oƌs��'�N7�y�'Ӷq �]&y��|뷊׬"��?����]CF�^�,1��]�QJd�'�ў��1��j�Ti��1GA�!ۥ�۵	���X�FMj�U���Ie��@��b���'�q�Y7J��K���y��ިB���8�h��YՊ���͑�gH0	���M����v�e�� \�\�D�p!�Dڈ�C�+y��rF	�9	c�&D+r2�F���/N�Q@M�$������C�,���d�?��i�7��O�"~�	�c$Y�"�>�ʰb��E���I����	x�����$A|�@4BR5�#<�����?��	m�Nh F��,HZ��gۯ�����ʟ���&���U����?����?��r���O��I��B��@'n���B��P����#��]�S��8)@�H�5��I�6�� �yf�1~�r�sAC��q��dy7�πzj�B4��-,��s�A�^V,��O�m���h�S�? L�#F�:^�&�H�IT�EP�)ʠ�O����'���|��'��_��Q�n���Vt0%j�j����1�'D��:6ʈ#)�p�	3��4*��`�,F�HO���O�����e�i�Z��Յ]�eC��jC:����'w��'dң�"���'^R��!)Z�e�BhIX��ECV���aH��@�5<�
�s��W/t�Ԕ��Fz{�ᲈ��;����ӳF ��Ç��P��e��'8@�E��$K�8-Ո��vq����<;R�'5�u@���n*�ȹ��J�j���M������U��}�Z��J�AB�� ++J��L� �S/j�!�_�� �6�P}�Ġ���d���Φ]�ش���>\�N�l�՟��m��N�|#�1��ٚW�d@Y��T�����'�b�'�h��fȔ4jA���o��G��pAo�d�FE��T�T�˲ L�ΉicV4�(O�ɂ�D��!���E\�-@��Z�`*2�0�D]��,��e��R~Y��,�1Q���VN'��F1PR�g�Խ�~:`�����A _>.R��iŭ�<I���>#d�#"L�!��P;
�h�z~"�i>�O<yTn�?)�B�h@�:,[4ѹ�eJy̓�?��V.&�bg٨� usC�Q_ڈ�ȓs��D��)G�	����J�Lj�M��N���`E�%}`��� ؟
b�}�ȓ88��2B�Z�u�fdZ�G� {Tl�ȓ0�pd��?RډX�� s2�|�ȓ ��(����'D���IK�sO�ȓA����fD�XT�@����v����P`Ĥ�� Ύb��Aؔ��?��%��BD��3�,��,�C���|u	�ȓ_���k�.T�
[���E���PU���U!X�YYԔ��Q.�k����R"O�2���6������&겄�5"OJ�3�l�Kg�}kC�Eޮ<�"O� �
H��p�u���Ќe�g"O����-��J� ~��dp"O���U	N-qa�0{��@�`����"O�<�4��9;�P8AC��%A8�q�"O�x@��Y�W���ѣ��)&أ"O�Q*�G����Fթq���;&"O��X��|��9�dl��o���@"O�90���(S
�	p��.�����"O�L�bn�{"��#�gQ�T|���"OP���i���֘�� hV\h2"OJ�2��P�:��7o@13�Y��"O
]�d҇|%Z<�B�ȾW"H�yD"Ol���"W�w��u;�9�(1��"O�ir%�Ͱa�� ���[�� �A�"OH}*����1� q��Yj#"O�0��N0I�PSǢ�]պ��"O,�y��I�FIN�b	 7(dW�'Q�oӡq��t��OķvF4bSn&D��Y�
i\�i{a&�/J����a�<٣啹P?�OQ>���'L1o/����-C1m���5�)D�T��
0j9th�d@�-\����#�4�Đ�8(���'©��E�*|�{2�K(W�Bh�	��P�d
��_�{�ș2�Γe>\!��x�:��c��	3Y�=��I�7
��H3J@�C�����">��V�A�`B�!�H�pY?	�����8��[�)�0fX6�)D��"3
B�U҄kF��]���QD't��U-]�&$�-��<�B� 7���Il�}�b,Ý}a�Dss�*|��B�!5�:�Z�Z�_�He[iY���P7�S�U;����D�U�du$,Fx�A�,%L� H��H�O~h"�F����>!�N��l��P��8��h�CM6>��=�2oɪ)op��琭f��e��l�"a�Ęg��hCFE�&��\Gz��ʩN6n�2Vj�� �&d���M�'1��R�a�A^l��p��Is���2��)�NL�v*a�V}��_��-YW썸@mTB���f��.�d7�s��Z�g��/Zq	͎-�\�0
,D���ရ?���1�m�6A�J��v#�i���G��>#_�l��D)���g�'RFyk�#�$o�|�i�AO
X���
�GC�}�6�Ks�? ��0����
�L��n�M9t�6$L/3�
M�d�DMX�Xꕁ*O>�rs��(@@D�N(�=2qC��נ���c���S3�r���]�p"c��#�ZB�	�#�mzt��Q�%���ABb�ɆǾQ*�N";J�# ���ȟ��yq,�,r�Kd��6>�4	Z"O���e*	(E��R&�}��t�Ԭ�&��lځ��ų�GB�n��g�'%* �����Pκ�bF��((�d	
�T��+U	ؼhE�Q6
� 	�Μ��
�}����R,�8%# �t�'�8�W��9ȞAC5��5"�V�Q��$�3'u�0c�((Fq�B̨|�W�ҨȢMȢs��H�O�<i�ŤO�h��E�UH�����L�@	�Mܴ�[��hy��i5'����w�z>�L����pL�C䉑tA��!����"��D�P�z�|�w�y��
�1Ǔ?��Xs7�D?G������7�1���6��xa�i�����jax��C�[cޢh��"O�|��b�&B-;�r�����>�{C�S�.l�$�u͘�:7ⱺ X)>�C�	�nnZ��
wS����.B�F&�6�]�9�4�"~n�����!瑶[r�b�Q��B�I�)z�i�Iöjh�����I������TAg�'��!�*4,z��䌕$�M��	��8�6��O���&���	����	؊<����"O� ٦OF�B�R:�Îfڨ�鉞 �m�#�"ҧqx����1�� rk�(31����{��Eáɳ4B�p��u�xm��(�t {�N�v�)�����˧Pm�X"�^�[yH��`*O@���&���S�׋Z��)�_�� F��j��I�ua�L�WD9I����F�&���$OPe�I\��	G/�v~񛖫��4ܸ�+'� �v�!��\�l��-ڃ��5a�l$�n��}A�I�+B��J�O�p(�`r�O�"�b�ӆ�(�x�7�@��'����E��;�F@(aM�t�M{�Oܻ2
R)��A��g�M�r���.��x�0��m������lr�	�.�3tyP���	�WyKP� i�	>{.�5"
ӓu���rU�C�Q�.��jلd�ቋr�ڍ�(O�˴F���4��Y���Cԩ�%`H�'��L�4ӿ���bR�T9*"�ON0s���I~2�0V#|���(��(���%�>MzE�y�<�����6�0c��ct(�y}�)ǠY��=�$�'��c>�D����̮;��3�#�.�tH�䯇�7!��܎F�~���1���P��(>L��iT��u1��w�i���ɟ�O �!��-�ąK��]EL��K4�'��i!&�<�`�q�>ɢg�(��U���� `�<D�&A�:�>q�V�J���|r�%j�����.���b������D�P����'��Y�����#O���Χf� a�@�E�0q�*F���ȓdW�MH��u���E��� �HvˤT� 9R���<i�*�O�S*��Ͽ+fFI�e��Aap� 2ņ���LF؟h�TĜ�.\��`ƍ��� JV0h(��4��$H�]d@���-%��1�;s�ĹFx�
P/M�Ԙ0T��[�B�R�K���Ozhx�Δ�
��$�k��`�6�x3M��4$�aJ���?0Y)�bS�wS-HG��za|#ۛD�t	P2���7.$AA$��6��D��Y�L�s�q��Њ��]�*:�h�4���`gD�,-�a�$��/h�zs"O�LQ�#��.�`"�jVK�����4u���V���	E-~��'(f���4���	�Y���@�a�e�TQ�cΰ}_a���3h3l����]*�`3�A�R����Ц��l���I
Z}��',;T-Gx�KÈ,0F���hL�h��t�0"����OFe�5ʗ�<�äQ����U猿;�xPp6,��:��?������I������&.��s*��Q���o6pSa0O֍0��D��<ͧ`SH���P��ư��JZ�J�F���x���3(���#EJ�C�|���:y3��
�zҤ�;����g�i�aQEݥ$p�[�GK������m)�O�,æ&�o��]!#�5�)�ٟ������<QW����/����sD@�46T:㮆�&ޔ��t� �c�ҥ���97��5���D���^��][Æ[�R6P���\��	�p%a|
� ���!�:�J�2�A
�H,� rS���Q�M҈�Bfi�[��#|"�O�`!H���00*r�[Ղ9LN��	�'����vωt���$u���x�[(,w��I�m�@PӇ����g��EK�EϐH�9s����RɄ��,�M�2��fcP�9����n�+A�ݺ"S�`j2U��X��Dɠa�L��	@�y�ŋ!�P;/"a{2(_�8�$h��O`������#F-)<� @"O�`�HB)����ct��M����)�T$
�F!�'1
0��;K�IX f2���ȓ<�2�х�c*��TI�%�v��%�?��'�F��'�z ��bMv�$�)�H�w�8p�
�'"�T�V!�07�u�S�B�d)�ش
\*%�N�a|�k]%g��T	q@Y�B�l13F���=�R��&F(]�w5O|<X4�Ҍ/T�ʆ��A��p"O��"�B�w;�;@��#uB�2���^(�2<AA`5�BHd!�5B����b�B�$%*��ȓ#Y8��e��	�ҽz�o�>�p�l�2>,ء�}���i��m�1�/}t;`��ob�� �'p�Y*���p������/qWt�@�O~��ѧGD��ʧ�1+~�j�e��"�� !�O
lQ�<�6�C8K�~=b�엡n��|b��}�<��Ϙ�[�"�:¬G4T�@H�d�'j&|�a� �.�y�K�7��	�a
\�s[�L�ȓiӰ@Cd��&��zgOA;V��n�B�����s�|�16�ë��h2>��/D��b����<B���$�,�ԥ�>���	�_�$%���3$��F�Ϲf�ي��I�!3���dճB��]z��iI ���+)�,t+���H�z�k
�'3��ZE���Z*�� r⍨>!��ۉ�dξyԬ���)X�O����^9K-vE�e@z2!�D Pd���#ƥVy�ܫ�d�"����<��c�"~nZ2����ۥl�z���!�%yjrC��}R�i6�Ьh�IH��,T�YE�D�p�'��xp����8�cY%V���r	�
l�L��>O$a���[�	�y�
�d�@=Ag"O" :�i�Vo��&C�, ɠ�9��1ѐ��iCJpֈ��*�����Kb�'�!�#-K�|��E?p��ݛ��a���m٬/\c�"~n��v�\��-ܷ$W ��ǅ�5X�&C�IO� [t��.*ޱ���>k˓z䩇�I�sp܁Z�ʂFS��	ш�-��B�9E��Ds�M����
"��!��B�=\[��z�MʀE�8ѳ&�*:��B�I<ix̥2@���ExA���f�lC�ɸa�lJC	ʹe9�Q����/7ZC䉻aG�-�'�Ş��uz�I�ItB�.Җ=9'���v�����kd�C��0W$�!1d�Gn���04�@ 2r�C��;UP���
ޫ&'r���J��C�	|8 �]<���y@ �-e�B��>�M�s�T�~&��#�܉NC�	��D8��� ��$�Ċ�*N(B�	�Q�N�rdc��/����G��X�XB䉊"\�ҳ�J'MȰ� nʁ"�dB�C���@!�8<�� �"�9w�FB�ɐ2�ę��"A/����A牛w�ZB䉜*n\1���FH� 
�[HB�I.#�B���w���QGE�:B�	�5�iÄ�M(JV����T!�B��Qܰ͹sKVkrP�T�?^�HC䉦xF���͙�d�\pkwE�i
C䉙GV��we��)�|��q�;!�B䉖yH�a�VkR;2 쀲�ë �dB�ɝ��dz7`�0(Z��fA�a�\B�)� :����1y�-�WoI�p|��"O(�Y��>,I�Xp���|��`;�"O��C�Oܢ:����⯀�F����P"O��Q� #K�����-R�q��"O�%��N	�1�ⱑK�$5Aj���"O&B儏�Y�D�q�LP&DF÷"O�L���#��d`�,�Ƹ���"O��-E*@N�B�L@�F���"O�T�@���X�$ey�k�1�B�*R"O����J���K�:q��r"O��1��vB���-��u0D���ע�3�Z���,�d��0D�,���	���a��A(k|��� D��	�)�98��*#�ʘ h�L��3D����d�P<����-f���)bh0D�ܰpA�9!4$�d*Z�o|ʰ��`"D�D�2M��H����}�8��=D��P�o]�$#��Bª4u��A��6D�(��*��x�֩c%�2`�~S'�)D��p��ì*`���锗/(B����#D��f*FCb�����ӞA���I�"D� ) �ՏT�8R����
�S4� D��!Viϲȶ��%�̴~����S�<D��ʴG(	� �削�þD�CN/D������>�6���O ����f�.D�����M$���˓�@*pY�� ��-D�L��h�E�ᛔ��S?�)�d(D����NT�mZ��#'��
r�l�RP0D���6���8�F���2z�Vx��!D���qЕibĕ*R`��ewT�Í!D�Ȩ2�נ
vfI�����8�J��p�$D��Z�kJ�������SnX�c
$D�8�Pb\�C{0�A���T7>�� #D��z"F� B)�p&�[/=p�K!D�P
@L���P2�,�,d� x#h1D�|�E��?�>I�UȀ�/��SV.D�  �� ml$i��Z*,.$i)�*Oj@#W@�	pW�L�B�[Y|���"O�!�Rk݄d�qق(�&
{5a�"ORT��)�p�h]Ƞ�O�z�2A"Ob!��S�V� ���F�5c�!"Ops�)�U��X��O�vC���&"O A�@��!�$�(w�ߓo&�LB�"O�TB`���}��K�R!0��"Ol�8��r�V�1��эod��"O>��s!YE!.�1�c��g��"O��з��0�bȨCYSZ0�j�"O8p�hC�T���т�
I]<��"O�92�@J�)��d�-Ax���"OJ���^$^tx� c�_*	�"O�x3��B�A���y�7PhL�"O�`
vk�r��xd�P9r08��"O>D`�Q�D�G��#S
(K"OP�qՁ� ~ߘ����y�ĝS�"O�"�C�-Wl�*S��4P��"O�����4~�t$��O�<��\ �"OX���?;�-� l
�0�vmq�"OH�rM	�hf|%�d�G�a����R�xR�)�ӋZ��U�.n yɣ�߁+�C�?E2�|�s�L6f�	�r��)X9C�I�-��i@�P�:쪤���N�MU�B�	<X GoU�I|.�:��ʾWLB��O�v��C���ΕB�B�2x*B�	_�Z�r�
��h@S�eM�C�)� �]b�p!�P�R���u�ms�"O�����c0���c�@��֤3�"O��)�@�>��%0�����"O�бABD� J<�qu��$6�6�(�"O��c��=P�i�@N�S.�к"O�L�L�u��ҷ��rV*��'��� ㅘ�p4X�/W.X4� �dJ.D�Hj�Z,"쐤�p+.Y�����+D�Ph7��4F X�y$�O��P�+D�1b�ʋb �!囌%r��+�=D�@Ic� s�:CX�3Z`I"�L;D��CԈM0<�fX��e��)�x���9D�h
o A�8��G	?"Z���!D��h���']b�Qh��6�L�'�!��$'�T#p�Ŕ��`B���c!�$��<��Q�0�³4��Dä�<z!�d^�qE��{���
lŐASDƮr<!�d�?z$I"�����+��r3!�$IbX��M�`�H&
�%&!�ė!�� rksfy�
�6no!�$L�^��9ƨ�
������'B!���^�<#ǧ�/��% �iJ1�!��Z��4I�D�*���8�!��
�<- �(O�<p~T��čB�!�d.
b��K Y�m^@l!�g�"�!�DЂc�����n8B�J�Ɵ�q�!�dR�\�`c��u+�U[VǽE !�$F
7��9Y�e� <v�3��,!�$	`e�����E�U*j<�a,Ȓ`!�&̄�`��M&-FLS��^!�$��`0����F�\�ɹ���)x�!��(8�n��^ ���7�!�A�"��m� Р�-���D:@�!�$ F��P���4?���Z��J�D!�� )h�`c�x���R�ꝼ~�!�d�K��XC�E�V�F��Ê׭2!�$��'���kcS7I�fTX�i˽p�!�d�}�����x�ԑ0h�CT!��;: �15*�t��I��ᑛt?�y��I�.q�����V�c�N�>\�ZB�	�m��µ�;1�jQ*�[��HB䉈 ��B�9#�`��E�)M\C�	[;Jhj�f�� �v*T�_��B�I#j�.y��'�p����Q&os�C䉌��̀(�d�`�c��{�B�Ib�B����{%A�a�ܼ�*���'���*�y.(���K�(�����'������UA�u���64q���'J��l̏*��5�����A�>|�"O�@ץH�4����2g`��$6�S��4}���EFؗ{\x�3NK�ZNC�I�&����y���E
�k�O���Ĉ"f��ԛ��Ʀj�`-��㙃o��}r��� ��Cò�Z�`=wN�x�a$D���T�a�|a��f�����"'D��Bc�I��igc�kZ�:��"D�T�Q�(���-�/KJq��H D�+ Y��H��&�S�<A;�A?D�lt�b�$B3��3D�*ՉW%9D� ƺ�zWG�scV C
+D�,x#F�rUn���.�@�0�kU�,D���7�F�g,�i{ ���]E{q%*D�03Q�N�=8���a�<	b�x �L;D� w Յ~]@��g�<X~���'$<D�� �Mႎ�:.%H��V�R�Pf"OP�s���C���[��]�t����"O� (�k /9�T��C�j�bY��"OT�"A�T(6��MIgY�K��i�"Oh= ��=�� ��o�7��X�'�Ib����@�a*�Q�`��Np��k��$�!�\)d"���(�7o������j�!�d�[2Z���`��X�Z�	��A+r!��!j���v��P���Pǋ�e!��FH�Xs�L<�������Va!�Ϭ �ReJW�ӟ5|��.D�!���Q��p�@�7^S��e$��g�!�V�Y,��j7QR�K�l1~�!�dVPu@M�� ?o�&��bL�M�!��u�ޱ��������y�!��'�hA�IL->���D���y�!�$B�-#�ٺfC4X���oo�!�<M}���`ڗ'�ʩ{��6!�䀖O3�,����.	�6��Խ[N!��~-���O��E�G�� E=!�gi�QB>zv��7
f;!�DҦ܎`"�`އ	 ��7OW!�$��5^���o�V��h3��b8!��Y3 �qB u�q�V �J !�=}� �zt��!�>DY��ܲ!�DJ;L������8]���C��S>y!�d#]*8��������`���!�D�~촄"!Oׇ~�b,��}!�d��
�����D�t��7�Љ!�K�uX�jWe� /�����ˉR�!�d^���)��)��m��xB�;�!��׫W��=k�Ȫ�F@�R��:o�!򄐀t�|!�NT�dnd�ڔHF#;�!�d�)ŠC�FSF�������
�!�dH5n<����"����ʈ?�!��k_
钴�<�扐G�]�G3!��ɾjb�l�!R��ʐ�W�o(!�d[m}����L�D2/
'c!�$9>�PREmB�5}�E��9st!�D�&=���+f�׃J���#-�6q�!�٩vĀ�qT �64��O�8`g!��2B$��gD	����3�2�!�N���a�N�T�F�ǆC��:6J�xk���X��B��ѳ'�C䉩>�*4K���sa�T���н}�tC�	t�h��̖�q3�xQ`�J�\C�	�=!��9�N�3l�
7�9w� C�ɖl�pZ�E͈t �=`'=j�B�	�H����@4Si>Vpˠ-* "Ov\S�d�y0�$�� ګRH<�1"OƬR��84Z4��j�K�l��"O�-��'ǳ9Q4��pd�%A1��5"OL��s���!R*ïD@|C"O!�`K	ک����T��2 "O8�pG��
g���P�!)"O4�W��!JY�=Bdo��Q�t"O�ڶ��#�8��c�I
r�"TZ4"O@Ę���<2 4ɂD˺d��b"O��s��۞O���B��U�Ġ�"OL�JW�H:�M
�#pǔ�	"O6 {���xl�Hc���R�p�"O:� dD�o��%��� �-��4�"O�d3�i��0Pe=�d0�"O6
E��H��1�B�&��W"O� |ՑQM��;� ��\�?j0���"O�D��b\�0i3Q�VAD5��"O栋�5OAn��fM,K�kD"OJ쫒J{� ]��Ѷo1Nd�R"Opڀ�.��dq�gEJd�9�"O��� 	*�[�3'�a���"O$)7�R$�
�Ic,Ir�pkd"O(��Џ�&h�僇�*n���"O���CI��+�p�a�J_�|@�	�S"OX�zѪB1vB-�a���7?~HI�"O�U	�(���R �V�i&�Ua&"O0�k�	�i"ɚb�"o�R�� "O�H���Q
w8�R�&��IB��Ѡ"O|iwi[�aN���`��)2�(�d"O6Ԡ���1$��Cvc��!�{�"O���ګI��#��^3,��$�"O�L� .�(�(SЦ���~�k�"O��1@�B�]@4�c�βM��<j�"OX8����RD. �s��'�5�P"O$y9ਝ
a�����A�t"�"O83��/�D	���3	�4L`�"O�����NRl��p��hY"0�U"On�KWL8ofL�䋏�u�e�"O�:@*�x�����e{�"O��)%�I,F�ވB3��L����"O���N�/O�E�c&�3;ؾ���"O�q�eFK��,M�af�W7��"O�q�Č��q�%f��U�A�g"O��aj�߸����N�uC||��"O�i �X'�̥@�%5��(�6"O�I���]j0��Q����9��ȲC"O�h c@��^u:Sjŝj@�:�"O�`+-@,�2�a4ꛂ>"p�V"O����*���;V�=\|�b"O��
����P1u�2>3h��"O�y�v8���p��q-j���"ODG
�
'w��F苒1/Ry�"O�ej�HD�=לMA�G�XpB9��"O:M� 
�],������"��dP�"O�%J�-6���+�@�
�T�0T"O�aA"��j0ҏT�>�>  �"OL��jˤvЬ�aN�,Sv0;5"O:D����H��s,��y��E�"O,�ć�&��Q��<Y��,A�"OJ�q���0	`ā��LhQ��"O�uP�.��n����L�:Q��1�"O(��"!������
�Z��E@�"Ov���%F7������K�P�6�ڑ"O�����YL���.R�n�*L��"O��c�֘"j�S L��	� �1"O$l�Q�^�/)�I��^��"OhŋA�҈i�u��X�"O8��aL;L�����FM�)�,P�"O<�c�OW2`�f�cE@̀	~�(rf"OQ�e�� >>�J����X*�s�"O��ԆR�G��ԧʹ|�
+0"O���ዂ1馬�'�*�}	�"O(�A3�/j0Ї+r��s"O���tMʭ�0��N9M�H]�"O�"�2'H��8�/S$�:�pR"ON�r5E2Z " 9@���~|*"O�h*Š y_T��ǡR1|Xi�"O�͓c��/8��P0�S�2@�pbT"O��A�fP�;`, �kЭAׄ=R"O� �hq�'ʚk#���T�I#^�h�"O ��LɣKD�:�J,��"O��� ӎ8�v�S� E�(�!"B"Ob9ːL�!+����/�nyhb"OJ��EK�q�puI�.�[�=�s"O�e��Mܖ1:��8cmĝ=�~�R"O
�"ף�L��)S�Ų��z�*ONI�vo֒.H�q$�7Oz,2
�'��t;U�ڦ Fȼ�U�˾q�d�2	�'���0�I�'���!KU�����':���dΑ*qZ�q�[l�T��'�p�����G؀��i�	]��%��'ވ�"�A�qP��)��I�|��'wai�ʓ�y��0��������'�r�A�O7c�¨[V-�}j��2�'kNY`c
�;tF��5`Z�w���h�'�Нy��ۜC��i$Eݭ e��8�'����2��nj����-D��
�'���j�!�DJ&m 		.XQ
�'�z���V�<E����
7>��'����E�ME� �1K�n�0���'� �r1���V��`���l�&E��'zPi�� ���-3��@�a���'2��@�!jV�5�_�8h9�G�<�I
	�*�rsC[�P.=��C}�<	�![
�xI�.\�|H �Bȃw�<Q ,Y�1.�I���#4�2��Vt�<�$�ɫ"��: �	�֤��i�l�<Q�&��h�k�O�h1�XX���q�<уf��]!�b��P��ׄ�j�<Yp-[�}0.���@�tPLEb7�Mg�<EI#��J� T�.���d�i�<2 ��HXp4áh��W���� f�<�$�^�l1P�i� ����iJ}�<Q.Rs~`��a�hM���{�<�q*̎Ph�Ys�B��0�X�j�z�<�R��;el�j��Q�'�0Mآ��u�<�m�;#q:���xLt-p�`�o�<ٲ*� R`e��\<h(���OU�<�HE*C���n�0�X�#�JP�<	ek��żu�&HM)��� QM�w�<	���i��!���I$"l�t�c	Ew�<�2���(��9"�ϊ7'i�-���u�<a��F#X`�F�ƶDA����X�<)��^�I�(�z�MX���J�m	V�<ႭÄNQ�P����e92�Bq�MU�<	据NV�1!� �(�$
p�Az�<Q��	6"�⼻'/W8Z0-U/y�<CC�2-ReiQ��q�J�:�Ȟ�<Ʉ�vT�:��[�G��AR��[B�<�#����In��L@��K�{�<��ё+��-!# 5 V"ma�u�<��dP�tQ��B!��2@}n�@���r�<«��m� �
�ė6��{��	l�<�s虅i���@e�ʴh.5q'	l�<AЊD#l$�9��ícV�� �LPk�<)�n��T�V��;䱱�ÔB�<Y���I����PJ�[7dD�eH|�<F-C���uzG��
�2��功{�<�U�.���Pa�*N0��C
v�<�#�3gk��#c�l�*��.E]�<�s�I�,�"�R MōOfV���Y�<y��E�!4���E���v��XōHN�<��*������9o@�0�UF�<� ���F���pFb)A��
�0=llʓ"O���J-8���џW:����"O�@r�Ͳ[t� ��� d����"O��3�@/;�r���-��S`	ks"Oź� �j��>8:�R"OȌs/�r}�%�� 	P���"O�<�GO
d����A�|;չ"O��*���v@��� ����}��"O����:����	<t�H�9�"OP%c��N�Q$�L���߫.f�mc"O�}��DG�n�^���G�^RNt�"O�`	��N8�a�ǆ?a1���"O���#S�(l>��5�<���'3�}A	] ��p��΢p��0�''1!d	�ږ��J�
QB6��'�R��!�Z@��2�0s����'L�A��Q<cD"�Pd�0�'���,��KD����gЉX��i(�'�LlqҠ2_!�iö���V���K�'�v�eȐ,E �R��K]D,��'|A*Ra��)��)�V
H���	�'�`��ϬZ����d�"A�:�	�'��Yb�f���hD� 䏀UԵ	�'��5xB�E�nL;�!ǇвMb�'aty�c�^���Kx@����'̪̂�Π]� ���dZduj���'�\eq� ��R3�� ��G(nH"-��'C�3s���c�	�cX|��'0B4Q�V�B�0��LY#kI����'ݴD���_`��А�@Z�4*8�	�'2}p��C9l���e�<M^�	�'��zb�!g��<��L�����{�'��B�*���"ҧ5� }H�'Jd,�����<в�f�O14%�B�'B�ذ�n�K��KG�N�/gp[�'UF��@�ܦOB�)���OH!1�'�&	�$ԭ/i�|R�]>ܺت�'�/3�a`1�%=���c+��y��P3j1���&�	����HP�J��y���#D�t��%�
�lB��y��I�lQc��L�Ԟ�G�О�yR�ȘN���H3F	�TQ���y2�C�9�4QC�f\&?��1j&o^��y���0b�0pj��LF����p��y�!_)2X��K��j�D�#�?�yb��Xr���cZ�LعS�ɜ�y��>jX`���5���wN���yb��cA����.����"A���yr�>5x&�3ĭ�#ܹY2���yɓ{Ĳ�@�7s/ع	Ugԣ�yҍ\����tlG6sW�`�T#]��y�`��2(n�p6��>_sV ���ǭ�y��1i����*ٞSb��Ku����y¡ΪBF�y�4Ea8l�6�!�d���b�@���O���0 ��N�!���
�p"0�+��ѐ��J!��J�f��XI�%é	 �{.�N!�đ�~+�]S7)��#�^	�Ƌ��7!��C�vE|�j�M��0�:�)�P
p3!��ߋ?���У�
�e*��r�jL!�dү7qX\�)�%<w� �d��:=!��UO��r�)I�n4��k֥'}!�Ċ���� ����P��M[�hޣ{z!�W 3`jR7�+��34���Y!�� �}���<w�8!�����N��c"O>Q{ə��@a@̎!�^@1"ONģ�#�!T��bE
�d3	I�"O��K�.Z�ն�Z�k�z4�ؑ�"O�iA-�3��Aɏ&R.x �g"OZ��0O���P���Aְ�"O@$�уZ�C��� �Jf5�ɓ�"Or9�6��;�t8���2f2���"OnL�s�چ�����8�u�""O�ف��]5: y�ˈ_��9E"ON��P�]*�!�����9�У "OL�� 
�laR5Cs*I�T��J�"O��2�.��Ļ��V�)Az��"O�q�#`P�/�W�Ӌ0@�)X�"O���C�>z����&�8+rpQW"O��h���Um,�S��_�6��S"O�=k�)�?ED�8sE��3t��"O������+��A��c� Z�Â"O��7ȧK��h�߬V�u� �7D���B�T�Fv���d��8WZ���i5D�L�Ł�-Wi�$�$�]1g1q3�3D��)�'K�[��§�Z;Vv<��n2D��{�o�"�U�@�Wu���@0D��A�DN�9���D� �%�f-D��A�*)�\3BH�'h
��f*D�|��F "l@�١O�-�����2D���#i�t��Z֯�x[�����2D����R6qeʰ���\�N�~��E�6D��G-�5y��Չ���])TT�"#6D�0�!̈�$`�����?E<i�4D��%�P|�J�Q��-p5)7/'D�dp6�T�e
Lx)ʏ1]8����*D�D2�o�57� �P�N�t�����*D���p��B��i0Wm�`>�A�H*D�,*��S�T7n�R��Mk�,��,D�0����3w��-�jF�}���a6D����iY�,��\+oè^o�耄�4D�t��F��6��P8Ҡ̓O:�0I� 2D��iT'W�a�ܘb�IJ�f�bA� J.D���'�� s
���
�%HN12L/D�,�C.2�x%�8yz��++D����̕ 7?��q�4!
"T��a3D����o�*�"�o���<�t�#D��z�-A��'F�8&�p���"D��11���s:���_��J]��E"D�!�� .t�nP�c��C��5D�(�Ҍ�?�6h�$���ƌxg�4D���"T�rn��ſL��ȗ�7D�P0�ݙ$���Ƅ�hvp��0D���#�=&;��	c ��X��%�c.D��c���8�Q�"�_�etN( �-D��0�+�"
_H �bL�9$m`u�Ec*D��Xwn�?*w 㙹q\CGD;D��RT��^쐅薯��Dq(xum=D�(Pe���/8�@!�μv����B:D���e�D1�5�c�u�y��,-D�肧�C�P���� %�)'���a*D��+4ɇ`L�n�*�x]PS�,D���V��t�����A�8�v¶�*D�����ʚF�D���F�^JNj�k;D��B�ތ3E�<�0n/e�Xa��M7D�8��1k{� ����;?�`y��
+D�� �@�# ���UE5�$����6D���E͕pp�s��@��t 5D�� �9(�8�<L9c'��)�����"O<�ȕ���uVԵ(�E\;�8�{�"O�����4;! ��C^+T�:!5"O.|@�1��� #C6}�N�q"O�ԫ�o�Uo���ցH�R��9"O����oG7n1��a�FЏl�d-j�"OX�q��\t|�4�^ R�80K�"O�Qc��3���Q
^�" ��٢"O����iHT�R�r�B[wd���"Ol����8z�T	{�BُN^f�R�"O����(�����NM��Q%"O����ϯ4t�q����5@�"Ol����=Dn|L�NR1z�h�"O^d��GU����qlޗB:�]��"OR<K �Ċ �BT�W�F�#̱g"Or����ŖZ�D�4�6?��9s"O����T9;/pu�%M	-�X��q"Oڑ�r X=n�m�7l�JH"O(�i�G�5=���'wOօ�A"Oܱ�F��^��tP�$����T"O���D�U���h
$E2�`�Z�<Y�EG�8�9���[�~A:�mR�<��N�^��yE��_?�ЗML�<Q&/�+\�u+��I��@��O�<	��X¨P�&�J�}:v��W|�<����Y��m��(�0q2D8�%�v�<���O<!��]�U.�.";&ɋ��Mi�<)�#R�%���AJP-;`�k���J�<AA�����iP1B�>p�4D�H�<��d�&�4r�m@�ڱ�$�JH�<�-G"�z)�b�+g��f I�<1vi�e��ybDƛ��Lp'MF�<i�L���'JχJ�CfB��<�JVϘm���S;&����o_z�<	��+X�6@Zd�I�f�K'H�^�<��⟴��t�j��4� 595,PY�<���-2l x���I)�<E $ |�<ab��|8Ҕ�e��$E��@�RdV}�<	�M���̺T�H�c�P��`��x�<)���p��K�:����+�t�<� Y-{�DS�b\��>0��v�<�`�4e�`�c%+�C��˶�PK�<�Ǫ�<V�pY�G�w��A�TN�<�Q^`}$��⊄�0
�Y�j�I�<I��� �� �7	�	`U��-]�<�$FP�&Y�ԺR�H�d�V,a�`�X�<F��S�Z�"a�j���(P��U�<�p�W>���A��Q%{#0�(cb�R�<���d3ب� ʵi�(��aDT�<A�B�<N� z�%�U>Ҝ��@�S�<	F@�9bH�3A�qb�f�<a�_!���x�ƚ<�L4p���H�<��K�*��y���}ͦ(��eH�<	5��I�\���φI�����P@�<��E��9`���]�؀X�<Yש%�l��#֢��r�D�L�<Y�#Q�U����jG65�	��EZE�<��`�) Bhh��F��s��A0C�^C�<�E��b�qA���SmL
��d�<Q"�ı
bl̺�ɚ2ih|���U_�<)�B�T.L��d�8���f�<Qp�Px�
Ma�
9�䠸S��d�<�/�4 ���]|�\�&�G�<ՍL�y��#�.V�Y�.�`�h�[�<� �u��h�I��e[�J��l����"O��9�I$Gb��Q	α�|:"ORU�7d�^Z��A�
��Q����"O:�����A�~�YSCB(TL2e��"O@���L�%G�Q�4 ˰M.���"O��3����u���oT,�5"O8S�ȁ6!b��5�T~�P"Op$XfAO�'�R}�d��g���P"O��I��%3B޹�����q���C�"O"��fŻZp�T陱0+ Sp"OF�Hd�I�Hy+�ʒ10*�y�F"O���C8P����1�ۆe���2"O�5� �>��8F��Wg���"OT��a�]�W�E��(��C��A�"O:�ǅ�	-ll�PοfH,��E"OrMZ倉4\��sR`J({W$@�P"OTEC��K*{  �O��+8�9��"O�i�$�����r/�5%�H�"O���S
2�ջh����;S"Oh ��N�2g�JY�q��& ��a"O<T��(Y���`��z��<�"O\��ɒ����wH���"O��I6%�"i�t2�^%�ܝ��"O�E�ri�8@��t��W"�Xɳ$"OJ�sQK-t(Y�@�	�G��i5"O�y���|F@�32���o��k"OX�Yyp�y�v^7{����Vh�<!�� �r4�iƱ �.����c�<��z�Z�`dm�y��`WH�<	T�R?A�v!��L��d��y�<��`��j����[���&\r�<G��9G;�hS��k�&=H@�W�<��G�z�8��D��(�ҁ���H�<i�ŀ�/����b���;aX���C�B�<���W*"|c�-�=W|�]�'��g�<�HK:b%� (��I��y���|�<I2�-X�ๅ�ךd�#�ɏT�<)��N�S�BaZ�OŠo��ҧ�N�<�r���	�� [��XI�Å�DI�<��"x�D�`cIK}_qkG�B�<y֪Y�( �b�N�<��eõ��|�<�W��-A��y#`�'Jʁ�sH�x�<���O�Xࠂ�/`�|x�ār�<Y�.�(�lԈ��30�����k�<�!��_��`Q�[�B����g�<���K�r���oެfR@��p�a�<��@��3%JǧR^��U"WE�<��Oѐ_��:dH�%'�|��\�<��1�p���'�h�C�,@Y�<��N n.�`Wl?/�E{�"~�<���L=�4�Ӈ�N�t�x�r��z�<���̃?�l�j�7|�aR���r�<�T�N>+2,y �͍�_(�!� �n�<�#� ad�tz0e��8NP�f�a�<�#\.u�]�Ƌ�v^���FX�<�D���#Ϫ��!4=$}����V�<��@�bkl F�ʍE��-aƃ�H�<I�^)yAfDA���lX�؀j�C�<1"��i����,ūh� ���D�<	g@M���9��-���P�s�}�<�*O6{z��{��S�7Q�x9l�]�<�Gˎn�ũ��%_Ɗ����N�<!��%�=�&��4 �7$VH�<ᑈD��R�+���HJ�X�AC�<� �h��A�5���UM����m��"O����b �!:�������(""O�� /�p7��@�� Q��!"O��[�/�)b�P��F�9d��ȧ"O:���-^,8f:�8���&Th%�"On�Z�\�1p���%��r]�<$"O��q��{۲��Reʨ)S�Y �"Or�{�GQ.1���4%�9�}`!"O
H�f�=�ڀ�pƍ �m�E"O�ܰ3F�7!��9#E�<�����"O"�J��Evv�*棍�#gҵ��"O:�pM�1�X�cE��%��"OZl��/ ����倳M��*�"O��7n��C���I"��k�"O����W�n���v?
�h�"O����OF�n�$��-���e"O� ����R�zm��Gٴ:ۀ���"O!��I�]���s�9�&a�"O�Ա�I۞0�܌����%D?8Tk�"O�H��б&��U0�`�M2�-�"O�p`r�¢ �X�!���r:LBg"O���4JJ�kc�!��GZ�}X�T:�"Odus�Lʁ[�F�F��KKN�C"O����9a5+!o("��F"O<���+i�+˕3T"�r�"O�}Bϝ$I�Y'JA�6�؈Q"O��˖��5�@p"d��y:L���"O��E�Ѕ,����'�-�``1"O�L����@�ά�F��I�9v"O�%R�� 6b 0Ħ�38b��7"O���teF�2QƸ�%�yu:4��"O,H� 
�	D�(
�䎄fFj䉥"Oy�c�L�6LK��c_,��b"O�FH�"�:���3]�����"O|A8�쎩+�����(F� ̌Q""O��h�'J�F�$�1�$
:y�8� "O�p���.R`i�,,:_���t"O�H!ׇ� ^���vLؾ.Y�� 4"O��˳�B�T�<B��28&�a2"O9
W����E.1pu{U"O��C� �H4` 	wfTFx8�"O���%�N�h�fA�t�
 [�݉"O&����9{��y#$B)&q ��1"O؉y�M(`��9���X=���:�"O�����;3���,Y����"O�i�r`L�"H1��Y2!����"O8��P@ Do\)h��$f@�P"O� ɒ�
>@��$ �!ɌN�bp"O��$a��j�.�9 o	����1�yR��i#��D"	9o��H��%�yB�B	Z{vR�/�6`m��y�64.�0S$χ�<��<��'��y��˵r��HÜ�a�"t������y��U��Ep��W c	��;����yR-�.`�B��W�"hY����y�(M-1��E�sĈ�Bb�t�j�y"�-qV4{!�-8���Iq�	��y"&�P��ْE��,4�@�`��y���P��-k��F�Lj��y�3nY�Ѩ�E��vq�ӯ@��y��AS�rlk��'0��K$��	�y�,]�-U�@�D)P#)(a���&�y�A]�v;4�s.I%#2<ɂ+��y"�A]�l�1 'N5j����y
� Nd"S�����db�߂
�l��"O^ib5��;�ts�
�-;�L!�`"O�Th�F�+u,4U�%@�	!�"OlΛ )|:����0кP#"O =*��J�BN`d
5ėQ��Q��"O�Y�.??^T(jQ#�-n<���U"O%#ƭ�g�c��΢O��؀"O�yZe�)ў��n��L�B���"O4Q��K�'���(�E�����"Ol�	�
C�&H
�B��+W֞x��"O�<i�Ɏ�q���P�(Ɍ�r"O�u�-D�w�j��@��!O�ɨ"O�@9R���	�'zf�3�"OH09�jI=XCt��K̿=��D"O����+=W�̛PJdڢ �A"O��se�W
0Բm����ʝ)2"O�%9f-ǱqK���s�Kp]b��`"O�ā��'�J��q�]�QC`�HW"Or����..jp��%�,8>�K�'�EHg�0w~�ˢΙ�����'�╊ �C�Ca*ț�"O��Si�.y(�-�&�!g&LxВ"Od�p�O&j8��D[4n(��"Oz)K��Ci���k��D�R�4�v"OD`"���'z=��e��j X�"Oj�`���;BԸ�b��"H�rq�R"O\`1�+U�U݄����	p�켸�"O@�X�嘡7U���V��W���!"Oh5����>��@��ɶU�$�8"O��1��B�G�0�!��ߵ�H��F"O�4:V#Y v(i(�)��<���1D"OJ��W ϩc��BG�4��}�"O|@f��R��,��[-|���"O��Y�Ή)~�
y�(G�P�Y$"OV��E͙3VܹU�ȜC�^�K�"OZa��h��sÂ��G�����@0"O�b�)Or� )&�V�$�P�R"O�8ৌ�,#�����/]����"O��[%.�/�v�{T�7_(i"O��7�C~�J"�<��S"O ��� �I>^�Qv#vKA��"O4�����(S��E�
w0v���"O4,A�W�6J�X��A�.
���"OP�4@�%�l���ۧ�>�Sf"O i�6�ɻ'i����ڳO<�Z�"O��bPG�^A9A�8E��\�%"O�	��M�����#�Q��a�"OT��­Z6��){���m-��"O��� w��03��q$�@�"OpК!�В�$Z�ew8���E���y��`ش́���?t=:YB2LE-�y��i ���c���q�W>�y�'�ʪ0@h �f!�8"�VX�5I5D�tI4��o�P�jǯ͙/��1��4D�(�Ș.P ���̞�C?>�h��2D�<J��68�������#�"�$D�$K�g��� ��A��6r����"D�P`ގ�2�1m�"A��*��6D�{D�<��B�J1r��y��i"D�,S�	нi�d2�-S�r�ҁ��;D�ԋ�F�� �9I�-�(�#9D��A���R��C�Ϋj0���ӊ:D�L��ǵ�!���N�uF8�ѧ�<D� :�oO2[ �Q*T��k48�Pa9D�� �0�`�^��+V
����"O�t0V�ų�8y�ө���-A"O�{sI��W�̼����
/EF];v"O����HW^�,�I#�����P"O���'!A~ެ�$��&�����"OL����ɨ��f٬��"O���o�N��<��/�.$Q$"O�5�%�[&F��� _�j��x�"O��f�0K�> :�	]9����T"O�,�k)C��iq��r���Ȇ"O^�"&f�2]z��8 ˎ23�� �"O�����G:z���ק��/�4��"OJɉs�ۘ)p�� ���!�P�*�"OFE�� ٥B�B��'7�$T1�"OtA����R�P�a�2�H�2S"Ob�z4bQ%S��؛�ޟm�li��"O8��j *C >����@�(-f%��"O0%�櫓�\�]�#�X��$I"O���͊b���EL 1��Xi�"O���L$�K���H��z"Ot3�Z&5�c��@����"O�� ),�l�gG�B���a�"O��7 ]�y��}CE�N9G��ܳ'"OL���gS�x	�`�b��4s�I�"O|� �͜.�R��R�F�V����"O�rJ�w�����S�^O�\��"O�1�(ɟ*8Lb2G�:f<viӲ"OP�``�^�k�P���FG?7���"OfQ��ƚ9�:��û9*�yQ"O�e���!I�<x�f�7fhl�w"O(���kO
B�1�æ9;a���6"O�A���%�PL�g摆FF��c"O�}��Dr�n$	�$�=�*C"O��1�� �D��3�Y4�<�&"OD5�MX��b�-�A��"O�@f�02V� �H(V���"OL]葧Ws�@@
���I�"O�����W;@�p��^\x��4"O�Ӥ(��s��!a�ԲB���`"O@d���F�t�a��ꃀA��QV"O��3�)#>�B���i7��l��"Ob��q�\
FJ��g�05�nYi�"Oj��`a�+T�(� ��D� m�s"OH���C3���3�Q*���W"Od�x�@٨s��a B:aP @�#"O�Y�RhՏ\4by��oΐy�I��"O�HP�ǫ��-(�n� D�Lk�"O��̑�P���$g���"O����.
�CU��ZB��,/`naV"OČ vg '8���p퉉TP�r"OP���N�F��A�)�}a�"O����?~�� {A�"~���� "O�+�n�5(�Q��C �*�(B"O¤b��߁#4�q֯3r��s"O�m�
�R�@�� NUTр�C�"OX����R��HAcF�\*ʢQ��"OH:�a(3��܉�޵I"X��"O��p��g���[�lL.G��t�"O�����9LMs�n��X�,�"O�	 �fB���X�nd�6"O��5L�ۘA��-P70bj��c"Oe�P�[pQ����X�zM�4Zp"O`����<k��A�&B�P���ۓ"OtL�weR((�p��B&L1y��)(�"O� ���v��tWZ�X�$�$r�n���"O��@��,s~��`��̮�J�"O�,[&� �]�RO	6�v��a"O��ɴ�<Lޠ�G�W�N�zś�"O�k��P�x�ƕ�g��?���R0"O�D��%����%(����P"O�e�g �/[R��b�ǆ!�"`1"Oe�sjPHR�2SX,P�"O�t�7���8�����n�: ���"OR���H��8-��Н"�"O�s�	��`B,�c,��i��� �"O��Q���+xY�|q�k��:Ɋ"Oн�U��+YB0��֧K<.�|H "O�q2��23^�3���(H�"O:����7_��H�nœgzX�2""O^=ѱ~��%�d�"0aHx`�"O���� 
"j��rk�38S��k�"O��;#(��d��Y�� %PMF�e"O�9�jݓR�0qIG
f6����"ON��6씥7�Y�v'^-7"O������I�4fߑ�H��"O i���#����&FIs�"Os����w,H!��"0l�aB"Oh��A�!Dc<�걃�+l r��Q"O�@�NX2$�4hZS�ãu�P��'"Oh5�G�J4�v5��f���Q�"O �7l��@���$�BhkQ"OPA ��!��Y��hB�wd�� $"OH�#�rϪtY���zr@ۖ"O:\�7�HyV����Z�/gt�x�*O���`�]�hph�0�:�;�'8H[�b���{g$
.%+|�;�'e�e��t���і	U�.��X�'nDM�Rd� r ^�S�ƙ*�x�p�'26�"'�V��#Ц�+vg��K�'yR��f��{
�3䎚�s>��';nX����BC�p �E
g����'c"Њ����ue�(�� _�`1�'V�Ra�2D�q�"�P�[S�(�'���{�j�-4Z���^�U�.���'�����P�^��>e:M�'�2Q���L�.�^�3��Ȗ^��
�'�#�ǚ�Ԯ��у5Pl��	�'�N�I� N##��A	�-G��a	�'qp5�"�K#��E{G��J��{�'x��cg�����K�b�����'��-r�/
+��趆N�-���'P���G�e����um���D���'��,�R �$5���� �����Z�<��b:�Nh�eC��U��|�<���ƂA�d%Y����3����C�|�<��$IG��������`̀2��z�<�3�ҏm��,; g�`��!dc�R�<�E`�XD��k̕FE��Dy�<q���!"�UW� 6pͨe�K�<i��F4& ��0+�*V���p0�A`�<A�dA�sX�!�j�%ǚ,P'�X�<���*b��Q㧫E/�pRC`�^�<���DrQg�b��b%�]�<a�-�/�h���]qj$��MB�<��й��*�K=6��K�V�<���ʃl�
��/�]�Ha[�GJR�<���T3DZBa1���"����a�C�<Y���.^���2�'I+#��k$��A�<� N p�+��6P��h�E� t�"O���SN�^wh�%�e��y�"ON�:��ڨKvh�qGV4D� X��"O��sL�(<��h#D-�g�Z+w"O��9�`
�_�L���2h��ɓ"OH<xQ/�jnP���jH���2�"O�8�����vHl9��?��ź$"OZ9{��ٛV�6a�@�;(��M��"O��8 ��j`q�J�zM�%"O��@aX7� A����L��"O��d�F��D���F���F"O�r#LC����bA+Ռf2�)��"O0Y���${^�M�A%wȂ���"O��3f��h~xq�0�9JZ���6"O��s�Ń\T
�ӆ�;4��c"O�iZ��~%J��lM,38�`)�"O�,Hя��yn���7�.,�՛�"OD����|0h@�?��7"O���eU2nTks(�T��jf"O�,ɥ��<F눬(X�S���#V"O�$���ܠc�A�a��<�RM�A"OXHÔn�,h�DY�q�D#�����"ORl`&�S*gX E`b*�4	�����"O��C�?O�52�T)zt��"O�=��f�x� Q��خKqFaa�"O��#�lјj䜻W��[�1�"O��zs��JVp�`)��fN�IU"O�<K���^�5�iA6�z�"Op4�@�,O>�٢G	m��y5"O�� �3z̓� ��L�V���"O
 z�`��1���+�6d�3"O��(���7&hȂ� "��H""Ot�"��Ц-�40��4���Y�"O����l�*l�ؓĚkaJA�R"O��`v�G�@����<B��2�"O�����K3x����V�K]�Ԫ�"O@���%��O��9� ��DS�D9�"O ���dۺG��|���S����%"O�a�Re��	n���SD�N����c"O.�3�G^U���0��&Q���k�"Ov��KG�lJ,�@a�w�blCr"O�Ѹ����v��o�W����"O�:�I�#�L��N�*g����P"OűR�ۨ\�t�03������"O��;�&-Q�<�
��)n�
�E"O���D
A2~����[,I�h���"O(��V?3���ȡ*כ Ahuc�"O��As@��%+�Z�C�,=+� c "OP%���R�l����aL�d6e��"O��jUC�.��YB��M=Q
LA�0"Oj�B��Ip�lP�Q�B�\~u��"O�uI�R*8q�l��(F�i��t��"O���СW�c�$(��ڨ��%[�"O���P�A�o��Ȁ4
$
n� X�"O�퐠f��U��B���)�0�a�"O0�X��I�v�Na�OC L��X$"O�i��f��l'�a����gݤ�{�"O(��AT6t� �g�{�60��"O��1�m�S�ʕ@��ןQ����"Ol-�����R��fL�C�X��"O�H����v���%��d��"Oڥ�p��9t�渻�iޅ�\�P"Or}`pJ�qA��*I�~Z�(Z�"O��H���j��� /I?lo�,Q�"O� �5@���%WMT�@7�-��"O&#��j4�{�,�>\��"O�9 �Bқg�b�����T��)�"O��ktA�;(ɮHk�K5eo���1"O�tb���J\�5�1��_~����"O:��a��H�7�� 5����'l������a�`�a�`�IeV���'�깒�
�gE�ᨆ��E����'L��23NJ0iYL��e�V=)O`��'Ʈ�x�}
f!SeG2n�JH �'�*�8�\(x����Ɛ�a)td	�'�'�v������{��!�'�`��� �sAʌ�-�`���'���%׳�&)Y���6s�`|�'������|h.�%$�X�|�H�'��SEJ�%6q�U�X8J�\t��'R��q��"$�n� ΐ�kq�a�'�p�p��x�� ht�B�.6���	�'���S&��5h���/~��T�	�'o� ���pG�90OU�p�$�H
�'����j��8�I��N��1��'ܔ*2(�l�؈6����d�	�'�]:�&�"f�iA%�)}-���'���*	����Ⱦs���
�'24-�ƍ�	��� fr�����'���s+%K`���j/Y�P��' �F!Tv�v瓂x���'! �Xt��+[��qO�4id^��
�'L��۔� �\������[|�dC�'����!N�5�Lܪ��Ii� �X�'�&�dn�� i�B�*Oo�c�'��i��˹z����*^�F;�,�
�'"��PD��[����'�,kxb�'�H!�7CÉi�D��ʄq�+�'�(x�`�U8Ȳ�[E��o �ٲ�'��-�6eO4�|h��_�dݬ+�'�а�A�EH����b���	�'��ԙ����&-����
	�'Ű$�k]+o~HA���m�� �'�ƑS#��t�&$a�鐶G����'�u�@���?���2�C�	�0��'ìᑓ ݤ4�� b�χp�d3�'�-@$
YSc@Y�AmS4a��'\.A��F�T��p�LƺX(@!��'�ts�(½p
 ���5L┙��'�����ˀ1^��B�L�>�ι�
�'_H���`�P�Js�ĩ
��	�'P���-;+|I`��^#k���
�'��Ȑ�=/0�A鎷e�~љ�' ��T�[�Fa8$m�XUԘ�'�NԩT`�1JX�DH,M	4	��'B�{�)P�I9��a�H4�J�R
�'��b� �!-�>��"N�0%���
�'"~hڥ
��*�P|x�+H�!����	�'a�Eq�̘�U��4����-���',T`���a�@����y�U��'y�Y�WI#��������[�'��@���]s�j�CܟF���
�'�����&ձ,��yS���w7Ԭ�	�'4�C ��;b0h�d��[jN�+	�'�z�U��0ҳ#W4T���I�%i�\�AE$0�����Jm�ȓ%f@�D��h�ĩ+�Ϗ�gl����7�@�	���}��s��=a��؇�S�? �)U+tMjh)�l[� ܂y:q"O6pb1��%̘�pM�T!x�"O&��g�1�p!��J�6��"O<���r�PX�0ʔ�S튤��"O�!�b�`�� ���z�ji�"O��1"6_8
���LÏ>ٖ�J#"O.������p�bA�E�4kT"O�l��I� (���{0��e�Hqv"O�р�`S�OO^``3��;f� �P�"O��(TaY:#l!�cXw�4��"O���%�A��u ڙ=��(%"O�i�ЫG�-�P;j�
I�� 6"OR8�m@.,���Y�I�V�Np�"O��D#,< ��@�E����i0"O��B��>7T���=6��z5"O���t�٠E_�t�UO&@p���"OT�[5`���(rf̩B$�"OjŘ7���M�8�G�ܵ�r"O��#�[��[�bP�|��#�"O�X�q�ϊ�� O�W�jh1�"Oވ��ʞc���BD�N���F"O ��"�q�p�D̓8.��L�'"Oȁ��̝;D�xj����v�	@"O�A��J��XPL9���V�w��X��"O� � �:��MC�K�I��I5"O$��Nԍ`N@;&nɽB� �a�"O��� ��p#��$��x�$���"O�,�ϓ	>��p�#Y&�~���"OP��A�^~�1�ݕr�xx��"OV�X6��"{ږU)��U��\�i�"O�)�e�2�Zq�� �)N��F"Op�?�j��ݮd�ZJ"O��o�)�
D瀶K� 
"O���gk)#x�����O�0��"O�Z���}���ٰ�v�&�)�"O<q��)�cw���shT-3{���"O��K�,�wn�P�C��8���"O��i��9]�yT&Q'���"O�H
c��,\�V��HCE"OXq��:@�,MA�L��@�x�"O�!@Uǜ�"p� jȚ�ti�t"Oj�M�y��삇FT)��LaQ"O�0B3\�<�(�0�����Acb"O��1#��w�~$Aa��$pNT�2"O2y���<]�#%��D��Pu"O>LcVN�7OP���D�.+�l��"Ov�c��V}�鑂ջY"v$�7"O�E�e,P����� L�b8��"O�ق���\���F���7�̔�E"O8TJR�ܻ0���L p�f(��"O���L�.:�$���	ߐ���"O�21�	N�>�n��pl�%�"OP�ס0!�@�M��Y�"O=����{�p���)K�<�!"OtU�' W����ʁ
��db�ԣp"O�d���4=a���&jZ�RQڑ�s"O�X�SÑ�9R�b��Qhm��"O&��D疸B����$OئA�}��"O������I��=� !\<1���1"O��"Po��zRPd*�� ���x"O�jA�O>��٨/�pX��*O�Qz�ܓ��t0�A�$.��-@�'�
�A���^�6�˦��-j
)B�'� !�o�)LD� �)X�pX��� ��a��%�d����T"O�X��k "�}�3"`�hk�"OPS���B
���F(ƢE:�q�!"Ov��.��+�عZ��8)L,z�"O�Xe(�8$a���I���B"O��c�G,L3�ôC��D�^�+S"O�-igERT�|��a	�o�r��"O��W�4n^r�A�y0ܠ�"OD��Rj�CS2}�с��SZ��9�"O�̙���f�b�CF@ոK�C&"O
��aI�'!��A��1?.L,��"O ���\�1�tCE,�9�v"O�X��`<5J�*O%茥w"ON���o�kJ�e��R`�s�"OD� Ν�;]��k��&o�(��"O8j&��'RzU"����g���A"O�m#�M!J�M��O��B��"OT�	n<]1&�F[�
1Z�"O���h
�l���˫Um
�AD"O��U	�r��<�,C�:j5�6"O$E�Ƈ�b�K��*�P )�"O��#d��TL|�-�^�b�!2"O�H`���ku~���f#3����"O.�D�Z	v+h%r�e�e٤0��"O�Q��Ą;K��c�% 0�B�"O|�!$M3 ��܋�E��\�A`"O��Q��G�@�� d!K��Ų�"O���d��mT���H�Vn���"O��K�)M��]�G?k��tr"O���@͆/(	�CA�=�hD;!"O~�"��&*pͫ%�F�[��l�q"O ���ЕLk���f�ך=� �"Of�	Ȇ�Lܬp�ӄ��w���"O�����VETk�a	!��e2 "O�S��B�UR�a��T#�`��"O�M��KC���Q�Յs�5�"Op k!`ԥP�0��-��Y�����"O�����6vf��KQ�/�LV\}�<����	�d������1�J\� ��C�ɽo�\�@�_�x}8S��#w��C�ɑk�jݹ�N�&muh�Z�l��q0�C䉙m�� ��;|8	�D�E0&�B�?,]� cFԢ]�jU����=m�B�:6B�;��,eZ��jՃߍgr�B䉥HP���^9��Z�$�)��B䉸Rg��C úH����\�|�C�I�]���Ka�� �b��; C�	�_�p���b��!��2��6~|�C��>,N(-;�@�?`���+�jәN��C䉧B
�JGoL2L��tpg�vfB�I-�&�3�bN2g�� jUś�B��	2<<�`��
h�(�3lٜ3�C�ɮY�FA���ʒbӴ` "��d��C�I/qz4�0�B.s�P���"r�C�	ZI�0��/��y����C�	��`-9T�� %/��ɵɊ�3��C�	�+�,E�>Z�r����ʃP�2B�2fk`@��o�L���a�I�R��B�I�8Lt���H�,���b/�  $B�I4Q�R�I��o��&ʙ�iB�	�!/�q�bQz��6F?C;�C䉛?y
����R7:�V<��M�Z��C�I�i4+�o�(qDZ��T-�PC�	�|&q��i�a�4�y'(T�cu^C�)� H�1�g�D�6�y��=X����"O�آ���_�����O�O���"O�蓴��4̾s��F*��m�"O���0���-�U��&���h&"O�}j�,E'�V	��`Y%��9K�"O�QY�-�;Nީ+��b�P}�"O�aQ֫H����3(T��A�u"O�&Z)�Zu�S`�?YX" *"O.yJ���B �Xj0�!:�5�"O4���mZ�%��cD�<6|]��"O�]�F���_wLi"��
�"O*�@c�R"<4x�fn����1"O��k�Ο�_{�$�V)̭,�~y�"O� �� ?>�q3
�茌Kc"OP�&��qa�X��W��eh"Ot���	�=HU
A�# X�3�R�Js"O쭐��^]#��G�n��"O�)�&e��d�� tA�aϒ�H"OW� 2���0BLIt.��A�mi�<Y��ڀi�̣��&<7�lIa�Yp�<�B �0`j�JN� U�qH@r�<1�Xk� ]�cD՞ �Z�k�<)[聸6,Y��<FF���8�ȓb�l� 4OJ-TPB8�u��4:=���ȓ �4�圮'`��b�&/RY��9�V��f!�)Fu�tk��F q������i�2��b\fM��_�/�T�ȓB��]8��X	2Q~%�d��#Zk6�ȓ��=���_�-�㎡p��ȓ?��x�FO2;���)B�:�E�ȓ@7���3l}�j Y��¸^����ȓy��=*�C	�H#f��WF��v��ȓC�H�I�o�{]ش�,P-������H��Bl4�ٲ�ȧm�LA�ȓ��]zGC�_����/{���LA����In�ŀ��ܺz��X��R6��v@9~�B8c5�80��	�����1f,]�&TL�׆�>����ȓ)C�Q�� ��pP�����\��ŇȓtAJx0c�CI��3�G[s%��ȓ9����L�'&�\s�m1 �TЅȓ�Nqpa�L>�^azc�ɯF�vm�ȓ?b��B�X�Wn@�ã��Iʾ؇�&H����[�z��H+vM,quJ	�ȓQf�M��"�6�"]��%J�hфȓ3�J��g@��t��w�j��ȓnU�� �Q�]%��[!�)�ze�ȓV.��I�����iC�",��ȓ����g�۪$�İ�C�~���ȓ/*���(97����M4h�p��B���0F��rA���3X�`��q�A��k�u����bF�������<�`/s�A����0}쐆ȓR�����'��+V,0�U�B̈́�Wm.�q�,
�v�s#��SQ�A��I���@T��Q��aC�-,Vq�ȓoq�ɊZ0>w��lG�'�J�;p"�v\�I��;Qh���
�'8B ��=/��i F:P��tQ�'�tSsFWG&qykDW�<
�'��4 �H�g��T�(	�'�%3��1�@ �$�0~�H[�'d�l����(51+� |���a�'|\�%:4���AIFZ�Dc��� ��R0���m�v.��I�����"O�tB���y�v���?���ۤ"O��9 ��<IFdۆ��?{r.��"O���AĹ+%�0yE"̍S� ""O�]Ε!9#2(�ۇYA�ȱ�"O�Eq*�x!�u�ֆ)n!��[a"O\��N��7��U��B����@"O<sw��#��ћ�e��iY@"Oz��
��K�I�@e�&Q�$�@�"O����+ɼl�V�y�c\�D���"O(��B��Hav	X��zh"O����]�K$�8�j �.i��"O�ap��Ш�Pk'�D�M�8i��"OBT"���'.�*m�w������"O��`�^�!܈�������"O`��ϬV��A�4n�R��<��"O8�ѡBO#tZ,I��d�]�"O�� W�[�k��u��\@=�h34"O����
�y�p���"4�X�A"O�$@���m׶�Ɂ�،d'ʐp�"O�œQ�F�,`@��	�|눝
�"O6ABH@B*�h	&m���r"O4x���:e"�\
�%W�Q֢��p"OV��s�.B�B
�E���y"O�ԉc��9u�(�CR8ydx�j�"O��zG� y\���"�8,�L@8�"OI���<S�4}�����\�i""O �@��=w3�ݓ�O�d����"O�kF���C0����;t�*)�2"O���"��^���#�m���	��"OL(�Q&�|մ�8�b� }E��s"OFݳ���00�⑰p\��+�"O�-�⎘;;
e�tAY�g�\,�w"O����ҙ5Y�(s@�{���҇"O��"*B�FYY��`ݬ�CQ"O����E6 P�J0�P�Eڼ "OV0�vė=P&As��֨m"�p�"O�%����}Ќ����-cA��1W"OF *r���8)�ᚈm�`�$"O�8B����ՋG+�X4p��"Oq���ȟM+ƨ`�IM�$�Q&"O܅sb�ZF��S���vӶ=�"ODh	P�,Z1�+��ŝt��YC�;O������2cF�1�_��ZTq��IT���"�`R�L�#��`�VC�ɷ��H�ᫎ�~\�7W�=%(C��'�<ت��ʉ"�d@�ƀW�I>:C�I3aN�al��5��R��8DAJC�I<5^D�a�\���Iw��:ьC䉇`�lʴ�	�,Q��^l�B��=p��<2��G�8[��C��:Z2����g�UW,�m:t�C�I�&��9q�7_�0��"ؔ8uJC�IM1��P
�.~��X��?d.VC�ɞ4�$�0Ӄ	�>I�*U�zC�I�x����#�}\y)W�P�=�LC�ɵq���!��X�1l����:jC�  3�X��b_��+©tN�B�I?Qa�X����o�*X�w�� �`C��T������Q�^�����;�B��7(���T��U�B�K2�ͼ��B䉩^YRT���j �(r�ϭ�B�I�x�$9�M� �μ�UJ
)�B�I�9�Z�#�a��0� ;�g��&fB�	$@$`�򆉆N�$A�V'�/ņC�)� ����T�w��3�C��+[v���"O4�B��/L�L�S��K�TF8Uqc�'�N�C��#���Am
̉3� }^苁 
�w�B�	>��H`�D�4�}��3;�'k��r��f?r����	�ԎF�m���	�%�T,!�����4i��^�:�L$^�|9+ �ߎYZ�ɲa[r�B6��|�bTX	(4��ꕮC �X"�C���x�T[���������*^�0x}�B@�l��8���>�O�k���+fL4��7W� �v�����ApAl5kt�D�2�?	���G4*fޱ��-'��uf�=D��z�����ڄ���5%p4A6M�<a���R����aDضb�X�G�dl~��H�A"�hk�L@:[f.���'��Â��,�����b�Pl�p��
2*`A�RO�M+�pHu�����,��D�6C�k�$�"�~���d��"�$hq�%�4�)�3$��)��D9��44zrIK��X�:H`����/�OV��0n��u[%Cɀ�b����>�\3�`��m��A#���n���O(��*EgӘoe����È,X�x�I
�'�r��w���M��d�����D�LW;�Dt�t̎7�dd�@k
�B�z�G��we�t&�&���ˊ�3=H����U�m�M��鱵��=r����K�JT�d(��_B,�k���(q��IĤO�Q���Պ v�dn�"D�Z����Q��,Z$NŮX'�0���ԃ3|杈�.ӂ@~��)	��5" `�
n� 18��*�O �PqJ
�$e��J��I�x�җ�$_��l"qB՗D�L�eH�w�H���ߟ&�C2c�9Q���ăL#YlYb"O\�L�{Z�0�O1%s@��f�AB�"x�W�� K��,+§oL	��t�`�y��I�M��8b.Q�f��HF�!D��P�hȚ���z5��m&�]��B] ���QI/QL�D��B&'��X��H�Q��p&.�V��N�4P�F�	��=\Ox�;R�>Tz���"X;w*���,����	��nH9�X��@S�i��rYO��|�G���HX��
�йG��߸'�Ԑ�b�,9�� h�����l�6�L9a!���3W� ��v�Y�a�����A�=�FC���� 壉��1���'a�h1hࠌ�W1���_0yW�AZ�V ���ݓ�wG�b�����K�B^dִ�I`d1D���dM��
��P���c۴	�Ҩ�:K��q�`��r�ua-Z2+�<��$�\&�Q�dq�ORQ|���D�O+/�%��'"\O A�c�	x����P�H�M>d�W������BE0&��y��}\t	q	La8� ���5x5I�AF�4-T��� 3�	/@y0i'��H��5��Y�u�����|��4hf@6O�8T p��%�y�攓ru��"L��F�V=@�dT�:i@aǇ�)�$UZ�UKN)���(gq�.�)GKn�kr�J�F����[�!򄞠NTXJ��I���P��I`�V^ O\@r�O���L��� & Q�DS�'Z�\�*B&Y|� ��
�;09;
ߓR��S�� \�L���&Xv��H� �p=@��#�ם]'�~��8A�Ph��l��:9��-���O�)��E�r�:�Ƞ�S(MB �C���<���{f@l�B䉞.p�Is���n�-rS�O>zՄ���4Vxx��x���'<��1L�+�f�'�����	�'�D��)e�y�6-_�-t�y[	�'&ʜ�m�6��IV�ɏ Gj�I�'���j�&]ɴ�xfE�3��}S�'�N�k D�)t�� U�[�%p����'����0�:��	���@��B,`�'��i�q�ی\�n1���Q�E�	�'Ќ ��\�ZɘK?Kԕ��[�\�p�*V�KWri����?4�x��'�Zx�K*=��[�(�9_1<܇ȓ|��{��X�DɆ$��"]�i~F��ȓF
���r+�;���bO�4���;����	��X)F�����s����ȓص�ף�{ʆ8����3A�҉��7L��� Uh�0�E���=��ȓ � bD��D�����[Zz�ȓ�}oȲ6��aҁ�X�	N�Ѕ�,�~�c����=��uR�G�P|x��S�? ��)5�7+�L{5�\�z��9�"ONP����U;Z`��ۧPbց�"O�y�E/�=[������F}�U��9���pC@7��ik�i�pvH)��w1z݊�JF�~��{�H�9-(p�����M�p�n��`�E<M"��V�<�AO.a�\��a^B,T��`�n�<YN_	��42֡8A�(���A�<��B��&q�a��nFxe~�l�A�<�2RlW�b#US&��6*
t�<����:JN�X ��:^�vy�"O>H���$QgL���-�;N�"��'"O�=��-E�6�����d)�"O�mj%��Mx4
QKR�M�(�1"OZ�jf�!/2jh�
ըx���"Oz�)g�ͫMC��bl� ^� ��"OP2!RO:m�%��A(���r"O����B�7��XQ�2�p�bN{�<�����P/N��q9}"�q�Hr�<��D�g�f|J��O�#~��)W�n�<�#
D�#�}S[0��� Do�<�竒�B\3�Df��p���yrk��m��Q�S�ŻU��X�(�ȓL̵`$��0pQ�S�n��ް��ȓ1D��ж$U���i���F<P����ȓ-�����Ю�R ̞<w���ȓHax�K@�9��	�  ѽi�v���$9r�Ksn��7&�!"�ȾN���@w��00"D�o �-r1�ݎ0C`D�ȓ7(Ԅ[�nW* ����PnA
.�i�ȓ{����c��g�
9�f�څf˾؅ȓ|J��a�&O����*�$����x��ӧ�K�>���K��)d&H�ȓ����!C%b�PQsep4�ȓt��5 �^�;��Q���Mxj*��ȓ:@jV�	;^vxأ�j�	?�"x��O=&�S5��-;�$�Ce���6��ȓQ�L��4J����C�ʬ3�|B��2�d�� ���}S�E�t��C�ɹ�F��6���5�xY���6�FB�I
Z����d�`����K>�B�ɂf(�0ؤ@�3&ԝR�+F�O."B�I������P*S7���<sj4B�ɮ;�4d���L�DY����vB�	88Հ�#��YRd��e��v�C�I )�H�2��F�g�t��p��$0��B�I�+O�����-a�N��dX
`�$S	�g�Ksc�
[��9�@�R�V�뉖o}�5����U=f�)��1T	R�	  �!���9 ��@�F$F��鱊�-c�1O����*��a�f��!"�'vJ�.O��q�f��'(�|�ȓ�)А �=F0F4wA�v��E�����=G1�$лR��?�' 2���cZ�}	�e"q����	�'ݤP@��>\���A���.0���v"
Wx�̓��w���퉷X�V�d.L�R���V�Q�<�����օb��/N�$m�6��G�t�nM
(zD��%�7ݸ���B>	��ˊ��r�p�D�3U+��%��p��c�@����%"2p]E�D12����"'�%�\q���Q��yRC ^�
`a���(�~\BM�� >�5�U��%���I�u�j�Y��L<9����3͚��-�"ވ����vH<��kT6p�i���I�y��)s�B�B�LyCЅ��,ٷ�Λ�p=qBk�ۂ4������QpH�qX�q��O?YJ��Pj�6`Kn%C��P�~M�G
Կ.��Us�^�yBo�4��ہ聉5�x�W��'�ēh�����I��)٦���(�� ĕrG�Ϗqp�RwJ��D�d��V"O�u�VoIȲ���*νn���g�h����Ԭ���?�f
�rs���'n�`��2w���ԯWN�n �'x�D0p�K w[��qP�g�xU�`�I Ю$27�Nʉ��I_>�p9"�7fr ��Ԭ�5I �󄖷gv*�äL�K��4|�T��sm�h��̛p��u��T�"���F.���
���+t�>��<�ȗ�v�4�j�K��h�:X3&��M=~����Hm�����"O^�!Sk��-����i�Y���{�U�3� ��"�>��f>�gyBk���f���L��MjTiD��y��B�j�h�E�J�ܑ��?a�&	 \f����b�P�"��W�^t8���Bg!��ǁ���BC��{\���&A1[!�DG���!`XeXR9�q��=!�DG.ѠD��I� ���9!
�4�!�$�(��`ǰ�,�H	F.N|!�d�4P�Q!I�>�r��(�Ao!�D�/8ͼ٘����p�8၈Z�#�!򤗳6�D�v�a��9IV�MR�!�71K�M��
�**8���#gʲ3!�dB;O�.U�4�� �b��F�l�!���)O����$H�3���Pr�Ҭi�!�$ÁR)(���MT:�\Ģ��4�!��0��@�go��,"0��/�!�X�\��`V6!X%�g X�!��<75$p�/V�N��"n�I !�DA�͒�Ӑ�]�K|���'�t*!���Dbj�Ñ@=P��j�`P�A!�dJ�})��(�MN�Bc�͋s�!��Y��f�H����0��B	C�!�D��N����B��9	���@�!�$ ��aR� �&�Z}3@(�!��Š:*�IPeҺ�
=�f�!�d�R�D�����+B��A0m�::�!���R��t�sS7k,|��L]H�!�Dۤ	���A�.�=-B��+	_�e�!�2�T�(&N�tG���0	Z�>����F�`�0a��*&D�ɑ����y����h�% nL(��Lш�y�!���Yb	�U�����&�yBN�5<g���ҦX�C����$��y�ND4S���J -�\�7�܆�y��ݱ��"n44������+�'�b ZcO�-\CΠ���w`؀�'c�!*Ղ
g#^ͩ�f���'"ʄ��.�8+��lBÈؽN:�y�' w��J��Xa�Q<9�F!��'�L���<UДs$�ũ2/�p�
�'/؜[H�A���SZ�����'��e��n[86h>��qI�x��D��'��I�@�~�x�tEU��#�'���%Dr� ����|>P�;�'��p*Db	�O�f��ƄG�hC���'YN���f�b�5H�ܩv����'
4�f�. �>�m���
�'7.���� Kw
q�	�u����'�>�RT�Y	1���Sq�S�k��$H	�'���Ҁ�3O���(���:lZ�j	�'��H�#%O*���_�lH4��'$�D`��Ru0-B�lK�fD��q�'h�C��*S2�dICƯOrF��'�*АA�Ğnv���BG�;�v��'cb�@�V�������<w�Z�'��l��[�KY��&f��g�F����� \���C��ک��������"O����UW� [%���Y�dyB*O0ip�Y� m�i)��I��E�'��zB�T��0��$��s�(H�'���٦d�T�F����mQ^�c�'�|I�����\�y�V�P�f����
�\�q�v�M�D�-8��I+�+�&m�X#�ծQE!�Ą�{�ы0G�W���Ao�=YM�'��9j�	z����)N;嘙�4���&4��MT''(!��
�?�����1�j}���7q�����c*?�&�m��>�O�-���NY���{!��M�NQ�QO�!�҈��|��ӢR=vi�1���')R֕"�'�9),݇�	�."x��(]O�����&�_ �?�1��!wy.i�C���;�x�'H��D�2�> !#������_
�`��	PmbF��>/ $�' TI4�ا{i�@�`W����h���̓���(��#RQS�"O�5�ޫ>e���A�C<1�H�^��C��*0,<1����U��3�
-�٠��>y��i��/[�?��9���6A|lSa�2���I@!C�l��!BG���#��l�0
t�@f8�����o��f%I�O����#�Y�6��il�$��J���؟�y{"�5xn �"���U�"O���*��q�)Y�� �L��cf���@B�NΥ�uK΢k�����9�ʡ�#.�(
��[�cF4@�v�S"Ov�0ܓx�� H�E)-�PX��3u�=�'hI J��bAg�$gܒ�(OF<�%V� =��O�q�
h��'��!W�A$JP�2EJ�@r���N�6�u��	�qM�p��h�X�p����kQJۋ8�~��Cn]�r,��?9C:I��5|:���8Q�4P�'@�eJ�qU�J�� 	L����J|X��L
�X1*W6lg�<`�$�74C�h��n��lY�Ʀ�Nx�?�a�w���M�=$|�Ò��,7�N�J�'+|��w�ߓ)��HFۥ`�$Jf�֙xw��B�Lsn�arV��"c+~��'�Q�'iޑAgS�H�][\lP���F���"e֙�$����8N
	��Xd1�uKj�� ��(@ �	-�p>iԮ��+��-�#�®p@
Bd�<,±� p�`�t���~h�8�ҡ�	�m!*���·ϒeYr��Z�!��� E2,C�A�c��-[��M��,S���6�  S&J�1s��4Ɉ���O�>Q�;}�\a!�!G.�J�ӯ
J&	�ȓ+,LC�������P��� ���.4HS4�ڐ'	��a%��5Bz��2AB�G���<Q�D70��9��MĘ%��Xb��[��t3Q�	�D,�,�"��=�.���%ϕ��������o#�X���9mT�|APj،�p>م��#+��Ӕ�69t��2'C{��P|�3��!e1	qg\'�����+Ŗ��iɡa���U�<r����V0y�!��\T�Y��1<I���/��Y �������wC�wO@��b�<§X\���l��D�EQ�&Ȫ� �)�C�ɘ
L���6�B��.A�ndK�팅&i�m#1k� k�D��oF�����Z�'�z�! *hU#v�Ϥh}X�z�c��X��G��d�b��X�m�T�j�H��(
I�V�n�M�fn�l���;�G\�y��d3�$b�07�[O.�|��I�!y�%�w�)�'VV�l+���Sg��0u� � <�ȓ����B?B���2iO:8
���Q(@�3��8���O��AF�4vl�	�E �^�E�W"O�D�V.[��̲aA�kҖܒe"O>l���j��+G@I&N���ke"O���i��;�ڱ[����v�^���"O&�Jé�*H%: ASO� ��p*�"OR�"UG��5�a�ɕn��=Y�"O���Ҕ^熕�� YL��I�"O�5C��
0ON��i�!9��@�"Ol��/��k�p��k��r�c"Oj���.�,�уL�
���"Oj 0 ,P�$�ґ3	#?jEs1"Oy.�������CӰ3�A!R"OV$�&��	u�X�'ǲ@V@�"OfȰ�W��M2$A�^�5�"O� �@p�o�)Rsν�C���8L�"O�m�Q���,(*�W:SQ�y��"On��$m)cSj��A�9@|,�#"ON�F���l#����0�"�"Op��U��XC啻w�0]�"O���C�K�L:T��4����$X�"OH{��L�jHJ$�"-��Ţs"O��%�f.�\�  	"3z2�7"O��+���)��ʃ��D8���"OL1�0	\�4x`�鑜���5"O�JR�M�i,8���4v_�4�"On�h Ɉ0��%�v���AHZ�i�"O��Z筒���r���8I�j�"Oh��6�)]�5� �.7]<)�7"O@�s$@C�C-�H�F��_%���"Oj�BE,�=e �pSRA	Ap.W"OPYql+7�T�gI�.UhP���"O�Y9��� t�dQJԽNG�c�"O��`�d�')�hlKP��P ���f"Od�0�M7A�dU����6h�f"ORh�� ǁd�A��N��8Ӈ"O�xvÃ���7"��A8�"O�Y*��ї<�,�I�'��z�"O8�B��������	o���+c"O�p���Zo�L�4*B�5���a�"O5h�]�F6<�ѫ�,,�����"O�e%e�D9�J]�K�R�"O�]J��Y��t}hQu�Jq�"O  C���?�Iy�S�6��@��"OpA#�D��r%$dG��0�ܤ8�"O�\ Q�՟tV��d ՜<���4"OI���`���e(\;l���&"Oꔃ�i�-kh��%@(3�> Y�"O@���!IX��i�Վ~Od��E"O���E�
�4rf!b5)K�b<���"O����8`K����'�@�"O���"�HbL���Ӱ�u�"O��e 9r0~�Aa�l���"d"O�ys��#ig�ո�a��A�
���"O\E8��g~hq�DO�w���h�"O�M���͑;Bp}Y�w�~�P�"Odx9��EB���A.د}.�#�"O@ ۰*7�)+��KP�	��"O��k�(�2w{|x�A�Y�(H"O��A��_밉{�T7<e�	b"O扩T՘>|B0ĤAh��sD"O�؀��ڭmc�X��
1dUƝ�"O���! �lGH��&^�C��"O`z��ͧ\���B�DK�\K����"O\51��Q
<Z�հ��8h=��3"O�Q��@�Y h�c94*0�"O�,�&��"mӐ�S�L�;�"7"O",Kc��]2��)BJ?>�!I�"O���%�L)A���1���)8 Dр"O��c.�|d�y���0k9�"O����-~��t�C&I����"Oĕ#� @�<�J`"�D��y�"O�mB�b�)N�x�ċ�"5��s"O�8�+��1��탵��+}���
"O"���kȔS殁�M�m�hY��"O�X�P��J��B����eEJ���"O��X���
B(yy"��7@\ɵ"O�`�`ő��$x�,F�3:�(�"O��h�"���b�L�#C��"O� �+���F9��Z&��G��4�6"OF�[@F�$b$(�dL�0��0�b"O�e��֧0���p�	�.���ж"O�����Ϫ`�t�Y2ʎ�H�H4@7"OZ\����5���B�u��5��"O�\�@ ́)���:F����`E�%"O��p�ΊI��!u�������b"O�ɸ�)��M�� � >��H�"O�UqԨJ/�|,�&흆�T�"O�$(Fˇ�$��x0�] !�v"O�x�#HB)\uP���0��0�F"OtU8�S/S���� L^l 1"O���΋5B��𹦉X�:�['"O�h� ȱ|�� ·	�!Kxp�:�"O>d������, C("���Q"O���B�ő"��p6�J'E�Dɂ�"O>� ��Ҩb�E(Ul�IǶ8�"O���������.NUl��d"O�My`ď�z]R  �'�>#�a��"O�ċ�żg�<��dF��\~�TS"O��Q&�Jc±R5��Z�%��"O  n#q�`Rf��DPbr�!򤔓8!��� B����E%�;�!��)/�z�Z���@����J�}�!�D�F�P$p7NتMSh�k���{a!�Y}�<�6%ɺ��pa�j�L?!�ǫ*�ab C�2S2hDȡ��Q!�%�!��"�7��Z'a��!���-�q�k:���PP��!��uc�\XÌ;S�Ū�L�!�ę,6��%�U��+"u��h3hU)%!�d
(�JVl�1��xQ��8"!����ǧu�t�c�ۡc*!��1
�^ysF��Ϙu���@�<*!�Č�T�� ��$�8r'Z�8s!�D�6Fx<Y�Pa� �\-���!S�!��&$*��^%�Yp�O��
!�D�$<�8���ÉA�~tsՎӥ!��T�<�����-D�,:�͏6�!��?Pa6p1���d����54#!�$�-jD��(�i?��ЦM��
!���|��T�}L�Ǧ���!���u����B-ڽt\���%Ǆ?,!��b��=@���}In�B�ٰ!�d�g�(���$m�)�u�W�l!�DP
e����`�wM�Ă�N�M�!�dĹt���yǬʩwHܓ����6^!�DJZdp �6Cئ	��[�<3�!�Ц*P�r2
	���hS��
�.�!�_MiNa�Т!8	�P03���~�!���6&���C��)�.\"��/��S�1*T�(C&��
�9�	L+�q*0��.�>:H�ճ�$�~��'��lX0E�.�ɧ�RyR�<(����Q*�(����M��^8Av�=B�bUE~����3O��:@f�2G�5(BJ@y�8�tjP)e�,�O���	K! ���4<
�m�I�Ab�u�"0�$Ӗ%����iS&����I?��H�M9O4�'�Ӂ�ۤs���iM
t�lqJ�BS m� y0 -P$TH�	*� l;�#�?㞨q�#@�P�F���$Y�I�( �De�t @�)�'�D!��i�-���o.�5�pm4�P�?a������l�у�E@(�����	y��1��>	i��pkr�;��E�s� �4���E\���u8��OB��'�@�h�����0|7B�v�����Ks�N��1H0q"��b�4T_�y�q�	t52>�N)%>	�O�慚 ���,�r��`Úr����O(	3��"�7�7�"V�a�T�_+�",�"�}��ȖBKT�A��
�� P6M���Rl�q�� �~� ���헯�ܩ��d��2lv�B�'�|�nڻU����B��N}���ߛY+T��6Έ�.-B��Ï~���m�
6��9ąhy
ç,�V�S,�W��Lx��C3tH��I�=İ%r��O��O�ͣ!�T�Z9�,�2��t�@L�
��3NA�>E��O�hD��$��q�
Y�CϏ26��I��&�;�a�D	��L�]2G>i�!/�(��'[ṽ��4�F��7#[��3�^a� E�7�F:�&ON��O"�)�e�F��՞Qy¼j�	��r�<��Fx����*s������2D���g�נ>�"'HK�����@��G��"�-ʇ�h�z���;D�܁Q&��d��! ���V�qd�8D�8P+����GBٽf6�A�,,D��i�gJ, *��Z�dإe�>�W+D�H�Ai� �v�[�U4m�^8�EE#D�� ��Rh�u�K_ Y�h��p�!D�8b���(�~���Ú$�6��@a-D�h��oҏn��I	�j��*�	.D��Q �[�/��h�
�d��K,D�����i��HJ�$uQT )b*D��@ҡ�w���)�苜I;L��o4D�<�7�PO�dL�¤˳v� $��1D�ta�؝ER�1�Qk
�&Υ ��.D��P��
)R��d�3M$
����2D���A阊X�|8��[&�m��0D�X��B�}�P����*<�R=���,D�`b������@=L�L���6D�T�0�Ʒl�6�yA�t��2�W(H�!�$�Ebz��)�W/��gg=u�!��$���9��]�A	��ϳN����E��b�h^j����lI�~|�ȓj���bs�T; jL �`�@�"J��ȓA�XH�k��i��=�ӣ�
W�i���,X�$�[��0��NCR<��A�"���X���Zai�v��I�	�,[�%��J�A� X~���x[��:�-�Y�̉��M5m��|��E���CFZx�:"�V=2�ȓ=$@be��= m\2'�Z�䵆ȓM�pr�+
�LE9ڦ��R��ن�?��2%��5-�A�1�Wn���b�Aj ��jc<K�I@JN$��O;�P�&�ݩ`W~���`�s*|��}�-�TL,c�y��.Z�	���ȓ^V�H3��N�lۅNK�<� �ȓ^$
�pb�_%���@C��¾-��:RH刟5ICؕ����0/RE���2�2RgG&~�~0�b��${\�ȓ|i҉k%�8w(���`x0�(��?W ٛ�#��o��I1��A�i�t8��v� �-���4�TcX�XH]�ȓw��\Ӏi�+qR�1#I"3�0�ȓoY����ya���'C�JmP��ȓu@�����&C#�) ��G$?�r���H𡂄
7*>t4��@]�&�~9��"�	2�n�I,��c� �bjt���ؚՂ����{n���(��ȓXb��a��ؿ=r�sP�_ Twnԇȓ,��� g��v=(E�9". ��h"VͱE��$�ް��mZ1^B����P�E�\�C��`� ύ�.�x�ȓ�V��d��(o�vY�1.٭�`��j����㡄�qI(�`ai�$i�هȓE����a� @U��D-�y��q�ȓsߐ�c')�y{��R(�]�T��S�? �� �Nm���z��ϮaGH�RF"O��j��N+��(�	S�b�H���"O|�(�S��.4�0���''܄�d"Oc��,�*���a�<�6�rv"O0Z�-5ΐ��'�X2&i�}Ru"O�<[ 	$O7n���՗Z|*���"OX({��N�0�(�!�+�6H���P"O�8�m�"��������Rȹ�P"OD��#�C�_v����M7ֺd;f"O
���ٟ4��<�F(oW, Q"O�E)�/6�x�ZD$�
A8��2"Ox��'LΚg��A�O>��YV"O l�I�P,�1��7���b"O�Fc�U��L!��@:ꐕ#�"O AP��4�f �q����<��"Oܹ��䌃h8*���H,� }��"O���%eB�+ZL�P悋CӰ���"O����ϐ�N��$�#�����"O!X��N�Z:!4$�q�Ȑ�"O̪���	�>|�d�щl��A"O�`궩�1Y(�Kd��[g�X�"ON����H?���ƅ9<:Lܳ�"O��ppGt�f�1��_����"O�H&�K�a{�W9jl�3�"O��Q�gP+3#:��'��yH�q�#"OZ8�5���	kn�ՈS4\(c"Ot�9�ʛqb�)[��OF*�d"O@d�3��7�J`�����8"OX0�)��,���KR+�������"O��8e�"]�ƈR-�;�J쒱"OH�z�&#���K`���S\$�"O2�Y�jI�%��	�B�%AI.���"O�U���h�4���c .F�2��"O�x�#E!S�����,{~�m�T"OR���@�og��2 I+x4QpT"O��K��O�JD�8�W	ߥ`�\�p"O<|����0"�s$ț�BAt�J3"O����F	<85����ŋHp!�"OHx�-� B<�Hr]� ��q"O���w$�Q�eY�6m]ڴ"O�Y fE�K�X�p2�2v�q+�"O½��E���d)T�Wn�r"O}�Po�u>h��-]�+_�m��"O��sMɔ��tZS.�0+9���"O؜��D�x�CCc�+fʊ��"ONё�m	�C�����S1k�H�IV"O d�Rg_4V����b�Z�~���"OP�� Y�����'P��	"O�9a7Ǚ�.<�0�lH:#�Y�V"OB�A�bݵe�p4ѕ�8Q1p(2"O�̃�aɥ'��z d��B�K�Ye!��91 ���+ߦFBА�P@[�!�(f�D3��@>$���`% �!�$,T�Q� �D��FMz`OQ<
!��=_�b���$v�&�"t��1L!�C�N���Fą9v�(�@d�Ŧ�!��Γ3B�p�SI9�|!�iM�h!�V�G�*uA�(�=.y�Z�.�>
�!�d9T�5��eԶ|`���h�!�ͭ;nJT#T^S��0+��P0!��Z�S�5�U��%9�����l!�+%�vt�B��(�� 	T�W�U�!�D�MJ i"���=8r��qk!��+���%�X�=��9ڦ���
��� zMs�"\�g����3�^��~"O�LB�(�	h��U�V�F6<���"O�i3�d�P��"��Z�m��`�@"ON�Q˘�/�6���F"n��y"O���e�ҟT��k��S�^r�X�"O(�Q��*�*�c�J��S\��s�"O�ro،]Œ� ��R�sE���"Of4�b�%�h�4�~:���d"Od���Y�T�S���d)��"O&i3����+�~����  Y�nݛ�"O����ם�0��Ծ7��p"OdH�B��H���cd��=Nʀ4��"O\�K u8��h��+�`�5"O�KE�.0i,��G?h�^́`"OB!�㚥H�p`�V��S��X�p"O�DB�o��JKXAP�n[��K��7D����`�v�d�B��ŏ6��9+��3D�!dY C�J9�'�	]��� L/D�@� ��m%�:��T6�2���-D����C�̅��D��*�b��7D�ppeH�/]��
��F�cE!D�pH7 �!��a �,,���He�#D�tr%#��.����K"G]f��!D�Y�˗,a�Q��(�0�u >D��8�L���A��?�jH�#�<D��rB��K%�x�v�0G�>��"�/D����sвj��¥%0�p� .D���G@֜
M<���*�q����"#1D�\Yu��
d���Z�t@8��:D� �b�V:1����"o��q8D�$�vO ����UoV�cU���q
6D�l�r?G�PI�!�"��<�"o3D��!&J }�rā��9��� �f<D�D�C)�^O��r�T*�84N-D�,���T/&�0Y �呬 ]zp��,D�d�F*-LP� �FH���-D��2��R��b���Mv���S�?D�P��ˆmd�s�l
�|�PeY��?D�4S&��5d�>A�$[�6���1D�,I�)w�pd�q�W.�ָ9g4D��JS�[�[��E3� �K��H��h<D����G�9�)�dM|1�''D�TbҬ�xŨL��혥5�f��)D�L�Ah^pU���0	�=n\Ve�RO<D�8���Έ!���S!�@�";Z���9D�2�@�# F�(W�S���#��<D��s�m%xX|!M�P#�i<D�T��I�xez�AK�/t�	���:D��I�ձ�BH#�S�W�xE@6�8D���b�ڗ�<֩�N	V�r�;D���Wo�7;���Q���Qƅ&D�Գ�L���⭊�zV��%D��j�-� w@y�2���d48y�/%D� �2kкleJ��3�YM���#)D���7@�< )��� �� �;D�;aHN�|O��bBJV.0�"yK�K&D�̢'K��A*��S6 ���JS�7D�&�B�y��S�*��	�>C�ɲkVҝ��c�HuX��ϋ�jC�I���	�(�?6X ����B䉍�r� C*� {\��*���B��+7vt۱�W-�(в%��NF�B�	�\Q� �ɋ�n�b5��
��C�	i���jFi��!�P,u�C�)� �ݳ��T�{j�]�P��)"�u"O�5�r!Է]�&�1�g�>*vP�"O�����7�������$�tzu"Ot)�� ��g������'�� �"O,�����7q� pC�9i�	�C"OĔ�c�����ԏ�"ML�r"O�ɚ!"`f���Gt>DE�"O6Q�<;�RYPg�) 
�3�"O���D��I.,�RE����	D"O�a�0�OEr��Y����T"O�XP�MH�L��m�)�%�)�"OV9çg�4+t�����C"�b�I�"Of%	�U+J1��1gNI��rD2�"Oj�30�\Z|4�	�ظA��<�"O�T���O�l�p�K_�JA�A"O��a��b 
�h��=~�x��"O��   ��   �  �  �#  .  C8   C  kN  �Y  �e  ^p  7y  ��  #�  Ԓ  S�  ݪ  U�  ��  ܽ  �  x�  ��  �  _�  ��  ��  '�  j�  ��  � 2	 r � � 9" �( �/ =6 �< �C J �Q �\ d �j u _| � b� �� �� �  `� u�	����ZviC�'ln\�0�Fz+��D��g�2T����OĴŦ��?Y����?�`�҅w+2���6R8�@ ���Hj2�2˜�E �b�U����d&˛\��.[�
���fW �	H>3'���bKݖ
�ش�TcėG'���Q��Q�m�QDQ�1��A�#Z,oR ��vJą9�'v�Vm5(n�Jb�ܔm�x���7?�~ �0�H�3���^8V�����v<rqmV$�U�I�X��⟘��-x*e�D�0:��ա��M�$�zpN�-9��شR��f�']�d�O�8��P�O�R�'��zGjD�W�3���6���'��'�r�'�R�'���\w(<T� b��y���G*�4:�@�c�8[��]"G�z���\�$ƿz�Q�@y�*�0Z�YVGI<� 	�S��!����'B�:�����4�B�FD��9��@�rφ�74�Z�ḷ
�R�`A�'��'�2�'z��'DX>�λ�Ҍ���uId����ZR��I�M#��i��7m�����	�2u�B�g3f�o)�PA�qi%N��ߌfj8ȩ�_O9�O�Ԩ4.H�����/���OA�$6�~�i�%��	��?��*F��,h- 9����8�Q�3d�REa� �o�?����:[w�Va�U
{��R�#Td�)�пi
�+aܡ_~�@�L4%��!�2�� 6�œ��g�X�mzimڅ	���E�ΞS��d�s�?6�%�q(ޝ_*��0�L,�M���ia~6퉯{��@&��d�Y�,M��=0�C6g^��be�HZ13T�(Y�e��E�QT��mZ��M{°i�u�����-g�ԃS��338�Ȁ=Ar`�i���$�GN�  -6-P��t̫A��`��-�� ��F��D+��$o�R�E�#H����7G;J�}��[���?q���?���i���$�F�S��%a똨��Μ97�D�<	���?I��^X�q�U�0yQ��a����R�W�4L6yh�㈼NǄ���*
A����P�\�'s"e��^�l�W,h�t%Y��O8]Ha�¡u)���ŹG�BMQ�\^�'U���+O�ĕ'�^l��H�� 8&k�#1.��j��?�����?���D�O��c(O&p��	F
�#d�X;&"�O��$@ ?���õ�(�����4�Ld��6G6�l"7�ׁ[J��,�h�Ī<�u�������'X�p��-p?A ��0�Q��B�"��$�O�!Y�S�2�n���(�6pt�Q�+�6Q!(�?���)Q&/R1#�̱	4Ɂ)t~b��P1��B,+xHС[ע7]�D���}�	Q�)pi!�.L�h��[ڇi��	K�V�$�����It>�[bD^��	xƪ������5���O����O�#~�g�[<#�F��s�� IX����s�'��k�TmZC�I�'J̣�I�1%�I� b۬1bD�R�4�?,O�q;&����D�Od���<�'��S���N�MJm7��]���6O3�8��G%x����,�����f�M���O:����B��<�BLDt1�$��w�C�*"�X�1`M~1�d��rG��~��[�\C!�ǸxZ �{B-^�n�FM�<�2!�П$�SG�L>! �Mq�8��A�-93i�`m��?���82�f� EhF-/���+͖#�
��	ϟ(�4S���|�Og��\����޺b ��Z��B��d�����DA�=���O��$�<y-�D��<�6!24��	U !����#������N�h 0��J*dj�O��	Z���7�	�O��|kA�D'=��U�Q�^�r��pF�4z���"L<	�$�D��|��B�	/-�D�%�J�BbD$�-��}����g��Oεn��HO�⟤�&���H�o�"F��`LOğ�	���E{r�JI�0�Q����R,�&�A�m��'Rd6mTҦ!�'��E��df�B�Dz�L��<����Lr*���sJ�O�˓�?Y����4$��ƩjG�T�M;��J���P��ߪ;KRav�Z!OPJ(�j@��(ˈ�$[)58��*u꒺tp��)eL��1�f%@���UD�	���G�}�5�c�\�`��Odr�OX�`��'��6�ЦI�	�%/��J�皤f�9�m�N}�'��VL�O��O�T�)^�:J�[�`�"h��*�!��y�O4�O�D�|ڣ�i��r!�*~�0{A�'���G�o�\�$�Ŧ�Xҩ�+e��)�'�oy�O��7�|����6sL�)��IU�\*!�O��$�'H��P������ �'�|��f�'r�������[ެH4,�w����O(4���@q��T��".ن `�e���X�2��J�JP��I_/B����ֵmjP�a� ����j������a J|ʋ�$E̖q�|�Y�j�'6�����
4���?qH>q���?Y)O���B���um <3��NT� ��b�~�'O�i����_٦q�	"T� fHW"_G�H��Q .���)�4�?.O<�pt"�d�O���<	)�l�"eI�C�.�1#�L6,��q2�@C�R5B@����?�l�)�J�ɐ2q�Q�O�|Qt.�zX$���N�$cL��c��E� ����]Jd(��@5=_z��Ȱ|*g��:�̻P1�8�,�5A$��S@@U�'���ݴY�I� �$ ��O\��O(I%kֲ�����v9� �!*�'�S�'^+�	�!��CB�2u�NGi���	�� �4��Ɩ|�O���R��14 �� ��T�����L�G�RmZ�Fh�7��O"���O˓��j>e!��ʰn�T��f�93���5��gnM�+ �u(��*6�d�BİF�Q�����x��r��ӵt`��8�R%7M��:Ǔ���
�KAa�U:��F�D��&�@"���kd�)6��u�^M�.צn7��D�ۦ���<%��QEH�� �4��+<Z�h�I_�	�$��Zy��|�BC�&x"�	�$�t�1-k���b���ڦQiڴ��)�(7LZ�mZ՟�I3h���Z�%ɅS�tl@�g�5Gp�	�L8���ş��	�|c��.�q�E��)�T��Nq�? ����U; �n�8���>�p��!h��	r���R8.��M9)ӎj"ȻfO?h�$����3�|��6ы"�F����E�4�J�O�1]�ޓO�	J��'�r���)�C��X�e ��!$��I��1��O�����=�9ǘ�o3���M���O��=�')�2K`��ٓIp&��!�[�?�,O(���#�ON���O��'.~���h�(��ԭ�5���8A�ͯ8��u��?���'�|�p�^c�����R��8X��@4�����2������6}:�Y�QB��	)Z��ș��`�1��N6��4���&1t$�C�oJ�k��4�ֲ_I��Z�}�f�P*��$Ǵl���'��>�Γhx�S�I�R^����B(����ȓX;0%+��U�8�2$If$�X�E{2�'64#=I&%E�Vkd�7M_�'���	s��$S��'�剪'DvE�S蟸��˟�'���0h� �����6��)�D�*����MF$ZN�ͪQҚe����?��5�J�|J�]].��@��?;È��j%k�ȡ��ƣ<��Y�0�F�'���[�E�j4��O�\,ӄO�yׂ�$k�r�1��žJ����$`]�.�fD�<En�����s�L>���?3�05OJ�xXD���A��?�����Op�?]�'���8�˗�WXX[��B8~����?15�i 6m�O��n�k���O���{i5�W��&��K�&Әid!bV�ja�I���	�0�_w�R�']�*@%���f��B�ީ&�R�c�F�NDQ��8@�4���_V�Dku	��
����҉6�8y�����a���!���=��2EW�0g$5
���#��K�ε�����G{b�I9(I�d���0I&�y"��L�Z�B�I�w�@H��ǲMJ�X��ݚ�O�o�ןP�'
�*��8�	ݮcjP���e=y �x�ʭp)�W�t�	ȟ$�ɚ}O
�8�I�3����G)���â۵U�U0?�M�T*d�����?o�*�<i�쌂a���5�Z0"�L��1���cfp;�J�|��i�D�'C�@xY5@
*'���k�.� ��$���ٟ��'��萑IKv���掇F�d4xK>9��0=ɱ�ݪA�j�q��8��I;E��Z��hO��$���̘b1̡�H�<W�����O|�D �����i2�O���̟����#`��ts�(��p���!�Ο��	3.�n�
W�T�t~"ܑd���R�0�Z�*DjH�'w7`M�ǋ^3�H�2��;!�l���O51��Eb CtmK6Y��E*�`VT���X��6Dՠ��M>H�㦞8bR����R�	�p
��$�Ϧ)���ii>a ���-�t��1���jb "S�+��O���S?h�p�� ��H����I?[D�=!��]	���tӦ�O��s%n���\�O�5@Y�����I�	� ��/��d����<��ʟ�Iͼ����.#/��6�A�J>!AeFH(/|x;1dY��l�DQWg8�|�Sb]�c�����\P���:7�0T:f��b(���`iIz�0r�(c���"f�4�S1T�l[��O�AUjɇw������-1 �J��'��	ZbF��OL�=)%풨������wC�m��$��y�%�8M��
��F�X99��Ԣ��ė`����'�7k�-ӵ�O@@���v�E(p�Ȕۧm�)������0�I��(�؟|�	�|ZU�Ш@誘q,��xJ��t+˪^~��:�nC"�"�bB�	!|�Xt��5w��<�. n�Bt��Ƅ%,^�! ��7_7ZmІ�<3%t�"#��a���ږ�ٛY�ȓ��ͼ��Z�H�3�C-A��PHW�VQgvA�c@���II�'&�t����k���&E�J`�aT@:|O^b�4 �%M!�`���ݵ5�̱��7�ʦ���iy"�5pR6��O
�䉥I@" h�!^�����'	h*��$�O��)�!�O��Dw>R'�:>H����_O4U3'C�0^\���D#|��fg�Ǧ�E��-!�(2�\�K��ǣ�.�(a���L'x�)�� �5p�����	�0�\���G�I�k��`���>|�7�U�8�B�ɫ'��Qc��ҬR��	EY*~d���ԟ���F�h��E�#�.gl;��%��LpUio�˟���c�dfO�?BBO�N@�(p�7�"��N0$�'�0����%�؀�gC'zN�Ѐ�E���T��?�B���k����C-d�	0"?�ևɘmV��"cOa��$�a��/q|���vE!��h�(xys��g.�ӖT�����.��'��>�ϓj�QZ�G,iI���(�40ߦ���v}8������)�vnU�}�(�E#ڧ(�f�@�
U�U�^|�8��ڴ�?���?yņ2�������?����?�w@r�5Kg.���h��~BH��f"�"i}��n�Pj�ll�g�h��Pu��!f{�a	�ҶN_�$�e�b��c��j�[��i̧X��ɒ/O����Q)32J�z�]�H��'���:(:���O:�=��4{1� {w��q�&��t!�&�y���-P.1��K� c�6ͻ����P���t�'n�ɿ-QT��u�0�%��&"DPڲ��5!��Ò������I����I:�u7�'��;�p�a���w���I5��$�z�����tD	��W�~<�àH�2��0A����(Ovt�� D}*�*>t�����f)���$��%Qę��C�H|p$���Ҟ}���+�":Q��O��+���:]r��(�7i	��d �|�R�'S���(�'Hs�-#�)�<)ip�`0�+O&p��IJ̓HN�eR�V.+��)QuN�'-�dD&�Ԫ�4�?Q,Oj��FզI�	�4��G�9XȒ倭HhB���F���Ƀh7��	蟘�	.T���5D�{H�����0'��Pa�,)=�0M���!- �E�A�щa��@���>�)���A�: t�R$�X�4@����F���V�KrѴ�12/��_��=iW�i����3�|��^1�?yv�ih�ɴ��Y�4��]���ށ 5 �O��?9�ϗr?��9u��U����!���C#d��hO��M�� ���g��-2c�Y�����O���5OV����X�����ӟd�O�Z`��'s��P��	l���*�NB�PUfQ	��'��nC�D�$4���d)JL�	։V�r0#�i��gT�S9|n�Y�!N�{��͒�%ȎKR�������)��.�4�"D�N�� i.m�ny�o�,�z�G�&yRhj�D��X3P5JF"�q~��6�?q��|��X]�0i��R*#��Y��nU�R�!�7}j@y�H�,`��Ի��Q��ў��	 �HO�LE�O*CJ�M)Em�~h��i������I����	�xH�#,Y۟X����������V"�&t4m�DB�W�$;U͏�]�h�a^�}D�����P�`T�|��(d���I".�(�Ba�!����kQ��
���+7}:P@DU{�,���MM?��h�O7&-',�,�yf�4O���G�f���7�@1�?!�O�]D�'^R퉅Mx`�S'J9mW�ђ�"�0G?���ȓO�2�(�
#�r@;s�Wܒ��IПPˍ�4���$�<���7~Ê᠗�N��Z%ʓm��	�#bU��?	��?Q�?���OX��}>�/B�m|h̻��-"I��a��hb\�&cK���S��ӓ)�j�m��6���<�A��	*��P��ѭeudĘEnĻcR�����f�ڶABn��8Zݴe�6�M2m�x�O�a'�]~E@,�R�aW��p����'��=�'3�xM�!`�J3�C�)-N ��	z�'ޚ��K�b��-�|&�\�ڴ�?!,O�mr��W���'"ly)�"�#��aPm�O��HҤ�'8"�ʄ ���'j�)X	r�	���
k���G �O�k��_8�(��AA�wӬ�H��'�\(��Y,?l���u+0a0��w��B����B�ZF����0<������I~~2�-D��Z !�r�.Xk�i����0>i��ڑk;�!���k6�)RǎV@�����O�es�"�&O�T�h� q�t��Ipy��2@������O�1���'����O�3!Ft9nѣjӐ����'�N���2T���$�|�Ο�-�)$�	q-��sѮl�㑟T��Tw�n�AaᎺ5�F)xFB9�' �m�� C�f!��X6L{o�x�'�@0k��?q��i�2�S.~
�\�æd��*����e��O���O��=�':u�(H� Y?vV�sg�"C��GR�w��o�~�	�N�D�Q�	��NH�d�V�t�	��4�?����?�!�!^Xf����?����?�w͔�2���d��h��#��L[�ybH��0=�ׇ�'�[�(�?}~B,�a�NO̓^����3P��h��ƈ `b���e���t'��8���OXb>c����G�&%��Y��'=D�b3�$D�����ud�֢�"70����<iF�i>1$���z�B��r��2�!���_T���ޟ�	՟h���u��'UB3�ޥ�g �"3d9#�Ј�)��Ս>���*ÅL��=��d�*o)�AE~£Z�P�m;4�(�MZD�&�:�����>tE� Q�Ҭ!$�q"K?���-��Ǒ8Z�)3�#?]��+4g��D��w�'��h9������e��_1���� D�xJ����<0`%/Z�>���Z��>�ą���ny�(��X�n�'�?1��E/SZ�!�lT��z�S����?q�P����?��O�HvF89�:��q��>�%��-Ю��S�>�LA��j�,�5ʁ�]��h8gD����d�?�p8�3��.T�y12����0<i���֟��	]~r������w�ܲ~�4�[!e�"���0>��@("-�����]����@�P���Z�c�|S�J���梁�o<|���qyb�
�8�'��_>Y��eȟ<sF��>qN���� �.mnX, ��PПl�I�cc�M��Aq*��x��J�BNB,�'&��Y�(�O <pQ�F^X\�K�h,(G�P��O+�&p�j@�B�Ya�� �@Hg>�4���7(3X��u�Ol剣(�"RDD���#��i�O���p�'t���<����f!b�{��UK<T2 �p�<aC�	��5M��y���i��U�'Q��8�����ŀQ=U��sn�e $�q�i���'/R���z�0�A�'�"�'u�3�8}��C�dX*5häD��8���-Z��0j�皘 8�Pـ(�U1�����H�~�._Q��&��_H91t/٠n�"�ccU|@��Ђ��K��-���a�q�L��S�? �b��d!��`���F���X��=�D�F����$� bC��c�CZ9H�L�p`퉛$_!��E�,����>uʺ����XP���HO�i9�d@�@�fL��%ĕS���@nZx"ĕ0��UX���O��D�ObH�;�?���d�� /�����L��y��!��ȏ����o�V)��J�4K��$P��'��ᛔ	��)��FH�L���ҕ�P�n�8�����n\@���3�0<�̌�_&��j1GW1�¤�Iğ��n�����U+��]������l�<U�A"O�{B��P.Eh֡H.�l�cӜ|"NwӀ�D�<yF��4s��so�(���4���MWoR+��O�����	Ԧ�$�O��Ӡ?���C�� G=���do�xjrQ:"!�-"�L�B��?l��Q4�Ѿ�����-82��AfU&|�@��WC]%$f�r�	I�$;ҙ�D�U	������L5�x 0Q�ɁU����ON�cE�v�O�G3(�g���_Ò�%�̅�ɂ\B�Qbd��,��B
A�<l���$��P�&)y�@h� ���s%��O@�qW�+G�i��'l�S�G��]�I�N����nƧhB����M,m����<�s�� \�|��Ȕx�X��苹 �	6q�ˎ$���)��W�^��
��;}R�T2T`�cvd_&?L���ӫ�Zc?=15�X2f�P�뵥�1k� #�& ?��k�ٟ���e�O���P��ͬo.llr�E�R�!��0H>��[���)z�"��أQ�џ��ɞw��t�
�j�<�H�( *�7�O��$�Ot;T��\���O���OV杌3,�c�.����0&g]���H(1�V�0���Y>Aۣ��|FybK�k�0];&�'��ѵ)�95Ӵ�E-�(_r��сI�w�>s����M��I,?��A��a��{��@���S��n*�M��� 6�0��������O�$-P:-W�|�����L�k�
�O�=E�HNA��kee�`9�
���nr�I*�MKյij�'B�� ��O���F��ʕ�#���v��M^� ��+.<�
���ڟ��	ğ��S�����|z"�K�����ta�19��D8@&�Y�<*�
�}7���ݦ�rf�N�}l�yEy�C�
�%��Ϟ
1�V���nݟ*�� ���ޡm�p9h�L��MS0R���`J�m����|bgS:~�X��Q����2�Ȳ-[*�����?��� Q�����ܲG���*��@�i���k̓BS�4�b���LO�)ɁkuyV@&��2޴�?I,O-��q���'J�E�D�ۜf����+Ah3Dx[0�'����!}�2�'s��\c��V�M�NB���'QJ �@ �V�@�
��ђ�j2�T$éP:��Y����bj�u�4��~d����.O�\3g�'�Ҝ���g(>��c��[�3q��c��!�d;�O��0�(~A��E�-Ҽ� ��d-�S�4�Oĭ���n�T%2��@�F` a@��'B��4��'����O�<�o�/�����ՁKҵЁb�O���ؼ�I��/P�a���z�#|���ܪ,#�)���'�����Ms~� 0�ԫG#�E*���i�OnL��L �L��j����O2P��'��7M�K�͟X���|Z���M�B}ɢ�\-3�.Exn�n��៌��I7N6�!�"��B�$�ҍ�yӔ�=Y�r���X̧{P�EKf�=�T�sIܲ$����O&ʓG�½(�'�?����?�,O��Hc�8!��`�V"һ$��P#2c�$r"\b���-TQ�AS1�.(b>�&��Q��7;�� Qj�t�-��Gֹ�R� �)��c�׉]]�c>�'�D�&D�{��]�c�O?}���kׄ�O�}�`e�	ɟ|��x�%DDD���̤$Ӳp�0�ky���'�0,����@s�Q��*Ēa�� ��?���)�,O�=)�A��GxZ�!��^LZՙ4j�.
��o�4�I����O�Э��&&3v����TIN�A��[1�0�cå�#�@TA�	�f�?Yr�������&�V��D9�`Т:��QmA��$ ���K A�!'�$"���z�a�m����'�'��'�O�"|"CK��9��C�#�td�`�]����<�hP4E��X���
J`�b�lT�I���d�<��٦h��O7�T�w#��03h�5c�5l�x�������O��D�O�Q���,$�U2�V7)��ai�<"�����C2t��@*6dם_BTpF2.׌9��Za��j ���3�"Np̫���8"tfxsq��*�^%� �	:����O:�W�db�̘.,�@qCGK�U�z)$�$�IO��P2%�.s��Q��E���HTb �	r����o�OKߨr���� Ѻrȇ��?a*Ot9($n�a}ʟ��'�?��Л]����\�~T��;2o��?��X�͒�c�6�II�dݓE�ш6��X�~��h��ݡ�
�#��~ �	/rix����(���zW�E+ ِ�� ��m�A�-e�e���x~�� ��?����h���d$� *�(��_���:@��i����t"O6A�&��k6��PL'u��I��I��tA��D�0݆�1�i��w�X]��@LH��m�X�'Ŭ,�B]>�<���L�z
~X;u+Bp��	"ņE̓a<p�鉯�� ���hHiB2�b�T��"LO�9��+�R��(��?X����G=�D�>^��󤟾���O]7y!�P+'�
�g�!�X	l>n���� T�!�!�&C�剼�HO>����/�*Y��a��M�Z��W�4GĎ �ڴ�?����?	.O1��1[�b�grؑ鳌˗FL�a��D[�ME��`���'Q��9լV�j���{�b��i@Eׄc���Ӡ1@���뉺l{F�[�b� #xPbVÞ�r�\�@�O��l��M��B�2�6
�h����+���Ac��+�LC�-,p����"/�^�S7�Mz(�O�`�'���
1Jش��I�v&!�dҙd�q!g�4u�axB���OB���*�i��Җ"��P���'���ҏ�ӬS'�M�
}D�x�)waxR�?�y2͂5��kb@���1D,H��y2��K�Rxг��{8�c� ��?y��'Ң�z�`[���X��^��bT�J>1���?A���R~�Y>���TQn���(�26�~Q��͜"&�L�Iҟl�anY?Z�pa��d=����S�OP�H��L����8��Ѐ6[�i��O|�s�D�zܓ�/Ɔ}zR�}�kY$i!�H�#IҘ`I�X16΍]~�'���?!��h���I8,���&M�Z���H�ԧ^��C�ɏ��l��L�S���3�LцC��?AD�S�H]%Q ΁��f�*�g��4������z,ʓjx�J�������?!.Oa1���j���#�Ƅ�y����&�sd5�uh��X�Ӏ��KO,c>c�����Ay��1�mC( $�����		J�0�{�ǟ�{吴Fb>c�$����Z�!낥��WF�O.�H4��	ꟘD{R��'C���ș:P,���H��!�$�:4��FąL���`'�1F�剥�HO�SZyb�ѫ��L
��	(���D���>L�F�ח6�%��SF�����&PX8ӑO��?�QT	̺���Z츈b�ǝ`�L�ٓiK�x6H�Y�������?���m�fX��_��PpO�>ͧW��2� M�|9T���j�teG|��KS� 3mZ�HG�ـj脵R��<ORiP�iO���U�7hU��9��\�T=��'g1�tu�6��;5�\ѹ��'B��u\����	&p�G�W�Om�Lz�F>p~�����Ay"�W���D��#ԓ.[�͈�A?��$F�Gb���OF�d�|ʢ)��?��1��X�ϑ!?�P""�w�8����-��ɛ%�D"�x����M�҂�sN��	��(g�����K�m6��y�mR���$��Zcbؗ�Aa�����i�������l|�`�}����J��%����[���ˇ��y�*[2�?Q�����d��d�b��2��Q積��f���$D�� $�V�a����cˌ"A �K��/�����4�j���*hŒq C,P������O����O�Ip�,!��$�OR��O���O���E[�v=R⇂,Q����g�_6![Q;��{}��ek�9P����̟�M���3��g�nDS0� 
=��(��K>F�r��-0v�t�	�2f<�!f^b���<2G����˂�yg�W1nH=�3�P"4��S��9���D�:c��'4ў��;�t02�O\��
A���	j@���Ep|ђs.F�~���b@T\���F���ǟ4�'�Dͱ74tȲD�s|Ҹ�t�!/��5!�'Y��'���c�E�Iҟ�̧�T؋�$�T'��')F4C��@6�f��rv B2F�a{�i��w���0eU)6��:$�\�=��IAu ��?P����7lO l���'��$�6Ŷ1�7����'�ў F|��N,�R�8g+J�ST�PG��8�0<y����'42��3�ÖJ�8{cn� H��ɱ�M[����$BC3�!�O��8���hb�B!e����6cʜ��}1F�'��;6�'>r�'�. ��+���J[d|��+ԗY�B4aaj(''�8�-ރ85R��qʇ���=��$+)Hv����ҋP�0��,�.�h�2EC%�1�a�M�;/4ВI.2���S�(/��O��S�'����ܸAK����%<��2��;��	ޟh��6:��;�`� lDu��͗f�ȓOH�=ͧH��	���Hbm�B����m��sn˓2;�غóiZB�'��S�n��]�I��x:�D��4>J�H�-�vA�!��BM����ڗr��$P&VoB���ʣ>�g�Y�'DMR�IR%¿[W�t�3��
N���6�@ڶ���c�<�]�wM�`(Yw�n�Pc@�2D��'x68A ���('zr`qE�[��͓A8����ڟ���'�?���� ���c,�:l�@4CA	c���!"O���ȠBl!��U#!��)�����O.}Dz�O���@���3=��r��S� @H1(��'�"�'*=�a��TU�'~"�'BJ�]֟tc�3��-r����Tg�Y�v,���s�T?\L����φB���O�D|���V���KɈ�B�eK��vX�Ƅ@�9��q�wj��6*�#1�GK#,,��h�|B`�ȹ+:��SnG����W	֖��Z�!զ��gt�)2����ǟ���\����J��a^�r���<o�lѐ���xҢJ�>��i�KO�=M�e��gAB�4��|�����=ёT��"OP�I���(Tb�J5xh����O����Opԭ��?!����Tlܲ(�	� )0��Scχ�0����6!�H����N�R��i�ʞ8C��Fy2�A���@��K\&��8R���PԔDS�)K�ل5�tdU�B
l��,_�l�Eyr�Ɲ�?I%/�F��q���g�p������?���7�w��8 LX�w�|l�`��)�hą�C�V��7��X����e+��c:�X�'��6��O4ʓA�I��i5�'�_�Qy���OD���娘�y ��q ��'�c�iL^h�D�k+"9�H�!CF���E|T�h��Ř?K
�
��e�&���}0UiSHɐ.� C�K��W�ꙩ���}�T��n�xň���h~z���͋
���Ot嫄�'���?ٰu�͙|�A�T1܅� �/D�����\?p�[�A �-�4�*��=��|:@[�t��H�M�Ҹ	�
�; I�5F�<A��?I����d�|�ϟ�Ur�\�>�<\����|���R����?�O��S�'0�jИ�@Z#�R��c��
R<��?yٴ��t)b�Ш7FJ�}�a�ï
�	o���Ҧ-�	2,u�P͓^���	ϟD��՟�'���k&kR�&R�����[;���$�P�M���t�t9y���y�$�$�����c�?ט�$>`$[i�Ex�I�s`�)�X(Hb�'�Zl,�0�'"�.�O��d��$|��(�L�0�ʑ��^7<�~�K�e�	0�>�D�O^u�3��O��ɉ3�4�s���Y?!AP2v��T�3jJ�y*��-���?A�,Nן���9�z��D�d�O~���O���bL�]�d�С'�C�v$��󟼛���O<�DL�e3��dk����Ǫ?7��;?�V�wUhЩ�#H�(R�rao��<��mȟ���.lt���?���J5��47�.�P��Ш��i���%��x�'��r���?������dm�(��a�?7��1oovE[����J�ZG
�v�L��&����^�N1�ݴ?]���!�~���	��M{�Hƨ.F�\�"��?�l����_���5�U�<�G� �I�?�I�<���|�J�t��f�<Q�|!��!�M��BQ�?�/O�$�SΦ������O-V����*����"���`)D��A���%���x7d��zS,l��,m�P�d0��ZZ��X��Oet�Q���'�P8�`AӁ;� ȹ��>N>)��$��` �/q����K\0{h|�4�=�	[�	\�'xɀT�^ )�tX��E�j�� ���$8O���N݌F)|a9��̃!vs2"O�Y��/H [�9!ė!^}�Z�"O�h���Kl�XLH�B>qbA�"O��aR�ƬI�`�]�>3�Y�"O`�+1�B=X��XD��	q� yG"OLM�!E�@��uH�I͕Tpq��"O��b�ɤ&�&E
�Ȕ 8:���"Op��T�U 07�t�ehT490.�Ig"O�D�1�ʺmb
=)$�����uأ��Οd���0����<ǣI�<�����0����eX��M[��?����?A��?1��?I��?ٕG+��(����R}I$DI�1����'��'���'}b�'S"�'l�B�T�S��M#q��ׂE��t�ie2�'|�'1r�'.��'"b�'n�u� �ΝH�d|�"�gndT �o�H�$�O����O��D�Od�D�O��D�O,�9�o�;il\�6�$Px�%�ڦ��I�����៰�	͟��Iٟ��I������)/ɶx+.��j���)��M���?A���?����?����?���?��%��~�fPC���{�<��o (��V�'C��'��'���'��'R�[�.���5���00<d�CB��C��6��O��$�O���O:�D�O����O����{���[�&�PD�FTt��n�ןP�I韜�	������	�T�	�~�K�p<�8�$��v�e0]Heo�ǟ�����0��Ο��Iҟ�������I	m����N�Of�=�T�~t�j�4�?��?���?����?���?���0e� (��
(�bՈǺi��'dR�'�R�'c��'.��'r�HQ�(H-1v9+Ȉ��%.0�������}y�S�*R�*�+Ցv�"�R��>q���nZ/]�tc����B�i��d�z��dcP�L�<��a!`dؐRO�6�HצA����1��O�7m���J1��y��+F��2@�Rk�m�Ot���G�g��1�%��|R�'6��1�!�k�i�H��0Ƥ�����D(�$Z˦�{�#�a�? ��c�J�7^Va�(߭A��9���TO}�fk�<�n�<�)��!#�'?x�rl�f�wB�(�W��˱K��iBbM:�g'?�'=ِ$�\w;��ɡ<SL\�A#��Y��A���a���$�O�}��n�3�Ζ+�i�5)˯o��I��M��Oq~��`�X��+H��p�'c��>���P��0�	�M�G�i��!N,ӛF���%Q�\(�D��̱p��.x�H�u�Z�$�� �7����'�1�&u�T*�),� �
#�H�`\���4M`l�<i����8��{e��nj�͐�#�x�#���vӔ�o�O����I��9����.	�h�4�k�']�8Mk�Oj�i�
X�w�H�=�	e}��W/A���C�Ĭ(�ޜ����yR�ۗe��0��\!��3bF�͘'x��+"��N�UF��$(��r���(~f0�XjJ ��b�*.L�G�R�̠�`!42��CsX�Ux�F�7j���`d�0+V�QĄ]�=u ��' ��YKӡJ�P���<m8)�s��O�uBd/?Z��c���<缈�T
ңO�T���>h,0ij3O��Z�,�Cs@�Q|6dIw�(r,u�%K=:�(���N�B�P���^�e���O�m�,�uj��T`�]𧯙�&��@FC�B�tD���"����%��D�  �xC"�w+ٵ0�(`p��Z�k��4u���k2�HL��bI�
�0%��/	 �% t��+,�<p˓�^��z��^xcr��N�6����a)4��E�����t�p�LX�k�&���H0'���X���t����	D�����n�)У��υX�(lZ���I�6M�J�V1w�H���.�������'��'�D�P�{�-[Bths��T�1��F�H5�?��?+O�̐&�[P�������x���YEǍ,���F�8*V2�&���'��XЊ�ԟ:��¯|�J�Y��G :笐��')剖i����4��	�O���Uyb�O�g����aˉ�B���q�j� �?q.Op)���)�ӻ5�,�j@@Z�5g�\�7�I/V&����Hm�ܟ8������S����?�UC|���D���.��=��ԙ�?y5��`�����dY�A�*u��<�\|rP-\.6�lZ럄��ʟ�t���ē�?����y��!8������W�W����$�8��'��Q�y��'?B�'qXy�ba��~r�0ҭ�G����'�̏(�b���IM��9B�
.`+�)
Eh���@SS���>�	ԟ���쟸�'R.U�c۫d)r�	���i�VDѪP�њ��x"�'!2�'(��ty"��-J<~�rH@�,�����`�yR�'$��'��);WP�C��F	t�BQ� �X6��q"I&	�2��'*��'��'+�	7X&��0[�l�!�7Tֱ�g蓅x��˓�?���?/Oz��`�[Ⓦ0)(�G̛U�
��'M�>(d����<%��'�t�ڌ{��Q&k�p#�!��5#��#�·$�?����?Q+O.��HZ�S��L�� �\���<)m��2�	[�:��e&�Ԗ'x�0��ԟvR
��m�#�ߵbF�1�'��	�Q(�m��4���O��i�\yI��S|{�#���%��E��?1-O�S��)��#}��M��h��^�`�iУ	2J���DP7��emZ��0��ߟ��ē�?1F@�+�b�+�.I�e8�(qr�C���?��1v0�S难O�d8����R��OZ�D�O��$I^@8���	�O�ɽ{�T�[2 .X
h�a��_�(!@���Z�������̟����¥0�"�6C��D����UH�ߟH�	 &���I̟�O��|b�J50�j	��^y	ڠbI$y�'���!�O����O��d�O��C*)��A.��T�d��|�ҙ9��O���O2��O�O0�$q�ԡ�2&���ff� �h4��O&ܘ��l�	ٟ$����(�	�
��|�'Z f�GO3+�\��ƿ~*¡��̟8�	埼'�<�Ieyrm�?&3��3FQ-R�Z1����W�����Q���IȟD�IGy/�5n�SƟ�q��A9��CvH�����4��蟐��q��蟔�I�=i�,�<tJ�n�ܻ��C�i�ɺs֟(�����'l<9"U>���ퟠ�S��LJŎ�)	�`� 󥏁>���$������X�a�e�S����ZQ�߄+�%�S�U͟��'O����'b�'G2�O���*ֈ�"�)�&��P��F�|��I�l���R���U�)�S�q"�����/�Fy��Pvt����%��$�O���O��i�<!��?6l�d��
�n�s�Q����?A�fN���������v��yhC��3ڐ�!f- :���O ���OJ0bp��<)���?!��y��J @n�ֆ��b�����H����'�r@�B�|R�'���'�� ��A�#%�!e��9V�\���'����Yu�Iҟh�	ҟT%�l둈��H�V�~M���)X�{F�"!�`=%�x���@��gy",R�1� 0@��L�z$�]B7(�|!J4�SY����ៀ�Im�ោ�	/2��i�E�8U���
�.��S��2�C�_�ş|��՟��'J&�cV8���"���%��8��ŨL�l��'��'�B�|�'�r���lЬ���fT,���C�P�3������Iğ(�'�(�Z>9��"kS@K0b^�W�˟A������O��$,���O��#k<<c�Cf��!	����t$$����O���OR�Iw�Er.�Z���O���=� 4X�"�w	��h$j��V�8���|2�'l�$�O���0>�Ԣҡ�9��I�ĮK�/VQ�8ˣ!�����Iş`���?�'�9�����LA
���P99�'zb�'��83�'�ɧ�O�Xk5�^:(�V큄��=�n���x�����?���?�����D�O���,����F:�6��F�YF �d�"n#b�"|
����	s�Шq�h0	uY����*��iv"�'�lհ\mO�	�O��䎒CN� ��o��)���A��O��D�O˓��9O�d�O��H2(�:X��H,M���g<mϾ���Ol�c���`�i>���ɟȖ'Ee��'4y�B�`��c��'��	ß`&�$��şd�'�PSΞY����q\m2�`r�`��n�Ol��O�D�<������CU�$��T�"�St�NM3�H��?9����?������7^t����>WBV50H���N/W֭2,O����OD��<y��?��V:�?q�?��\��C@  �� X��Ĳ���?A���Ċ
н&>ը�J�s�v��@U�Z�f��m����	꟰�'���'IHAq�'��SKf�2�P�a����wn�,�P�	㟼�'����ʟ��	�;"��CW��Q6j�C�v	BsJ_[�˟�I
y�L*0�?Q*�(����M�q��D������ODJ�'�O��d�O����0ʓ�,J�F./��d�'��c>P���?���2Q��r�	�z�Sܧed�hQ�"��+�c߶+X-��'<s�2ڴ�?���?��''E�����Z0c��hK j�"dB���k=Y?B�ߨ&���'���'��Z>�Iϟ/H��ZƆ�=�^�S 	�8�rI�ܴ�?����?�W��+������'8��j ��+��z|�Ԙ��Q���'���'���C�[>E�O��8ON��� 0��M�Vf��-�� ��'�)&dd��h����Ap?L��
��#8f��ц_����abDEd~r�'��'�� hh�$���$���J��x�Ve��a��ē�?���?Y*O��$�O�bs"�H* b��(#�0s�G�)Jn�$�<���?i,O|����rk���,ش�(�#@6A��X�IH�W����O$��%��ğ��	�R�H�`���aG�Mh�!O�V�ja���IR�j�'�0��]y"�'�N��Q>��I�)Rr`D�ܰN���ӧ��9�,���Q��?1��n0T)P��h�dܽKh�Pk4p��4�6�48���'��П�J�PZ���'L�=�d�KF�Al��teZ�<3Vԑ��|b�'2�O� O�)�y�OQ,���C���%j���d| )����&4�>�m�H���'�t�<q�b²b��qx�NїK�I���Ο(�Iǟ\yQ��ϟD$?u��D��LG;E�j0"7�8����_�T)�#\"n2�'�2�'[��V��'2�ğpMf� �Ã/K�V�Y�n�Nm� �Iu�S�O	"ȒFK�D��щ��{����6-�O��$�O�erc�P�i>Q�	ٟ ���Q>,LJ���2A�~����ӟ����,�	�y����y��'���'H��S�14��pjF/RY��Ii�'n"�"m$O�i�O<��<Y�"i�j��5
��(��*���?���)x��@���d�O �d�O>���O,\Y�N��e�$�BӁ�W�D��Ɖ-e���l��h���t�������<��=�X���G� ,%s$&U�K�}qu��c��?���?���?�Bo#��6���(|(԰�����StcY�t{��'���''��'u�IޟH��>��1��v B]`W.�e���0���\��˟��	l�O���0-y�z�d�O���񎐍d	J�$DI���kt��O����OV��<!��� �'�?��'�.�ZW�P���� #��!T��i����p�	ϟ�ɹj� A�4�?���?�'_+�J��®X�����K9�?A���d�O&Q�u.-�i>�Q#b\�Q�ޘ.}�0� �K�ڟ`��ɟ� ���M���?y���"�'�?1���S"�t�N�NC�#�����D�Oܑȁ��O��D�<ͧ��iX3GU^�2M��g�a{�d�1E}��I?*k�7M�O����O�i�V�d�O���M�$�̔�s�N�^�D�aW!�@ ���'����$�4�n��Zb쒓 ӚFGX�*#���|��lm�ΟD�	ɟ`ꆏU�?���ٟ��I��$��<�(�t�_ þ6�$:����џ\�'W�!#c����'M��'@�ͱ@#��A�p�h� ai:2"��?��%�`h�߈LF��'5��'��'�y"�);I�0��6S��h֯���$�-!��$�<y���?���?��Y�p̹@��I�r˅F������&�w'�&�'OB�'���~�-O��� �%�ܠ!�I�a���a�R?'��"�;O��?�����O�xx�馽1��V ��SBh�=t�ڜ10,������\��ݟ�	Syb�'Z°c�OE$]ȶ.ԄM౒Eڍ�8e��'��'�b�'��S�	�J��޴�?��ql6����C�L�ʠ�s [04��1��?I��?�,Of��ۍ?��2?YG�	���LȲk$�8��j��6�'%Y�XBR �ħ�?�'PE���Q��"�y#�9�40�O>���?i�I�5�?9J>�'i���l����1^3(��u�' �ɼ2,�̺ܴ���O�i	eyb��	v���V":eJ�Q�hų�?���?Y��W��?�I>���䦓�HԪ���3�!��.ד�?�
�(1ߛ��'��'����;���O*� ����J��(Pc���va�'�f!��'Sɧ�J���~:HBGiڞ4qsǚ":"n����	ӟ�HQ�E���?���y���K�f��P$ʇR7�������?�L>�Qh?��'�?)���?�Tb�4a��fY�h^Tq��
T�?q�ʴ�Iѕx��'w��|�fX�3ڴ}+d�X;R�;��\�T�	=Ks��Fy��'��'剓Is�0��&khܑ��%�6쐀!���ē�?)����?!�%��Q'��a%�I�w(�䯟����?���?�)OQ��!N�?ɒ�KѕK����b�Y�IN, 㗀�<���?1H>����?��<y���j�T��N�TE�
@�ۂ��d�O:���O�u��b��tM	�fh��.�= ��P���'0�'���'B$t���'�	�!?����6�88��uR���O����<��O

Z��O���OLȍ��CJ@	�w�Z�蜘r�|b�'����:p?��|b1�~�X��X�#������T��'��ɠf6|A�4��	�O>���Ry��߽Bpd���
�0VT`�d�?!���?�#jυ�?QJ>�}� lBO�$�%�W�;���D�E㟌�����M;���?q����x��'^T�J ㊏`����Ri�%_�T<�`�'k`���'�ɧ����Ns2fՙ��C2x�B����	��m�B���OD�����-��O��$l��Q-G�g&,S�K]?[]Zp2�+��>�Th%�����4�	�J��`�p�@t�C92��	͟�"&�F)�ē�?������2����5�d���`�1,�)OX-��j�O�ʓ�?���?1+OPX��%H}K���3�-�b��a�<)Jr9%�������&������,G��.p	����2k:�N�J���	py�'@2�'��ɎQ��t��'M9"�����R��-�H��ԕ'�r�'t�'�b�'�$Hs�'�L�u��w\HS�S�/uA6P���ȟ���@y�K�N�:�H�j��Rkdd��Є�t����e�O��D$�D�O����]n�b��	�邍�|0�'��!=������O
�$�Ozʓj@-�W��d�'��.�O�Ȱ&��|5b�#�p�Ob��G�K���=�'hf��wˍ�8(�p DJnvx ��~yb�"ľ7�|B��b�]���C��D�R�K�l�^�P��<-O��D"�6!�U��= �Zs ϜtqfEХ�'��i�n`�b��O�d�� $�擨���a")=&N����P!)di�'��Q�lD���'���3$	:y^"�4�6.>��xӨ���O �DAh�N'�H��ڟ��I20CPl֏4&0��X:,�E�?�SN���?i���y"N��=4���L~?lr#k՘�?���n^�x`.O˧�?��y�A�5E��`/\�T��e��(\���c|��sP)?a��?����?���,w�U��9{�|ف��P��l*�k���?����?��?�I>���?�"�^�����a���B��c��B��p~2�'���'��	?{7�� �'%$��c�Cߊ/����l
%5�\e�	����	ȟ��	f��?q�'' ��Ω��U� O�)MEnй)OT��O`���O���G�g�2�d�Of�$�
M�24�Q�(�إ�po�-;T���O0�O��$�OJ�+'m��s�M�4�����oE�8����`C�I��ٟ������ɳ*����ğ(�Iߟ��ӛdP���ǕL�N�����0Zb5'����^y�A���O�ͪ��$?t�5���ɶJ@�裠h�Or˓_w*]���i�����L����$�P��Պ��΁S�
��r
¿F(�'���ab�4��Y�|�I�B����B���	=۔���#;8�I쟌�Iϟ�ן���I�t↶0ʀ�dK C�H<�AG�J:��MN�ɋy��i�1���2s��%HD�1�h�*#��<���ͬ=�P"����U�H$���1��i֧LR����4�	�7�.�p���,�Αa��Y(Qt����Ɵ8i�#?Q���?Q���?i�O8Љ�B/]`i�(�
�d��2R���	�l��ϟ$��� Q��s��P@�'K�i5ş͟��I۟|&�P�O���/�O
��ˊ&qʝ+G�49Lr�+�d�)4"����O�OF�$S&@���"'x)�s�Ǐ�Exp��0Il���� �r	�Y��E�3`X��� �T6Y���'�Hbƭ�YXrDz�G�("
P����]3oFh���#��9�ta��P�HeCw��.����E�^^2�拀jK�XKclJ��r$I����e� � ����Nd��H�j6��e��V3H����J��
F�Z9)��{��A�Pz@�
��)e���"i�>#�,�%o��k�RXõFW����Q���f�(S�J�))W~�:�&��\� �9�!�4e�$!���'d�'���U��?5�%
� �,nЎ��&�U���bC(ܟ[��S�Y2ʌ鱇�E.�(O�h���фKsPm3���#�"m ��ŵ1�A(�eM�^���R٦F($����]><�'�DT�\��g��)�}:�ǮII�e�"�M�3��y��t?�����>���X�7F@�Bp� �/��Dz��k�$,��|�q�>�W"�5j֜�`A�`�^M��$�e?�����	G���'S>�9�Y���IѦu���Z�+ ��*0�=s6-�ÂLG�pu��DT�5��t��KȠ��.�IF#��\c�R�{��tb�y�R$)>9�Q�4^�Z�cH%<z0(ʧYBr}K9��SC�Ł���d��b�sZԁ�egnD����i=^L����?��O�Oc��� ��B�ֶB�,��͗�s�
y�"O�i	vK�wL��hm]�	¢�S���O�Ez�O[���)H$f��!�ȿYp`�e!xi���<a��[�?����?��O��Oh6�؊>4k-���Z�F Z��d�3^�*4u�'�"ri
�b٠d�SM�8���Ӳ�lHk���2-z�����	4� E>l� �AMW:�k�Иe����'x����'Q7��>��Y�l�	m}2n^;tLL=�@+�f$0���O%���~X���2�Ru�(����� !`��R�	AyR��i�<Qԅ�/�.�6�ۓ�n0p�����oT�?q���?���~ƚ�����Χ&��q��
(v�F�Ee��~t�����"����8�O�@YwH�.J;��3ht�to9���w�=QpP��k�D5�I�PL{Tm]	6�8��!�=aגlH"KQ��M�����O6��'qiĔy���>vӊ!�c
�T<żȓ{��tA�j}Zܫ��ħ���`}��ey"�g��7m�OV��~��oR�T h!&I�d���
F09``| %�'o��'ń��P FBl؀ ���d�6D����|�R̛�
�(�sK�2ga�b��Lm�'4�� �/F�m�f�i~��E%��|��(X��Ph�!��(]k�I� Qj�'�V�*��?1p����i��ٙ ���h��d�e9���Oj�"~��3C��)+�	�i JhZeY&V��<#����ݦ	!�OXՉqA�t�	2��]Nv��'��$A�ˬ>9����G������O�7��p �g��80����	Z <��-B��|�C�� +|>���S���i�P����a< ��JK ~v�(��4\��<���I9XP��h�·09�G��4k�"u�@�?,n�1X,���|� q��'�l7�����	v��M���U�|%��Ԇoz5�dg�x?�����>Q&T.z7� �4d�b�yȃNw�'�#=Y��8h�gپ~R�릈��,x�@��ҟ���H8�&$F����8�	 �uW�'o���ͧ-H�H2nޗ(��K���	|���DE"��i���ܧdf�������iF��lT!�W�j�&���d�Um4�����r�m!��B
M"�x+d�R����)}���;��D�$K�>��r��Ȭ%�v��"L���BM���W�����4��'<6�S�^�p2DC�F)��xS	V�1/�C����3$�Y/m�򽉑�A�2>�b�/W�<͑��ش�?�*O$E���ЌfBz�1 �V<��7�ˎFiB��$�O�$�O���T����'����2�k!�i`���ꝭ^Hر�FJ݌D���"�:�X�@֮�צ�q�`W�KR�EBJ��.N�,�w"0�O�dY�'����΄��}#e�1) ��r!76Z���O���?ٌ*��Ģ��؆Yx��ϑ'NT���"O�t�� 9@z�`Р�=T��q�O
��'��(c]�}��4�?������N�F.�3so�����ɀDV�� �GS���	蟸H�"b�*�:��;sk!;޴9X�ᨐ$)�f� !���NHN�@!c�?{M0H��$���M�B��*C�R$���j���ãK*mV�!E(L�h��5A���,$��yiR�"j�,�M>yB�Ɵ$�ݴGɛv�'R���_�"��aC	�o2\H�'�Q�iaR8;�������b
�qj���! bI�냎�)���A���$`'}���>��@����n1�u��$�~�J	7�f6m�O����|�G���?y��M�B�"&�ysǁ�%�$�Y1a�Z1Ґ!�TָK���!}�T>��|n��"��#�ӂUm���h	�Cs7헿m:��Q�-����`��M{w���x��	���M�3@�ڦ]�v��O�0m��M��舟�vh� ���pvb'_�V����O8�D7�O�cG��JL��8���!G)0ݒR�	��HO\I鐤xӞȒ��ףg4�途��,�B�I���i�n�{�����������	��u��'?���� r�д�Y�azr]�1 	���$M�,���ꐉ�1;ay��;�.����r����a�Bu��(�B	Ϗo_b$[�,M� g�dQ����<#f�C��3geT�w�*D�g�V0co]0si��b���
�����H�'r�a��F1u�� c���%d'� ��'�XY��A�c�j�
ю�Y�F�ApjJz�'��4�'��ɹ5\���`Mȿw�F�a��Oy��V�>P�����ߟ��şP��N�������|��jگI�H|�נhp��h�Ƌ�&q�<Kǋ#Vݨ�ӕV_Z��dմ!�ɒe�c�|]rR��':�@bJĩuD�R���?��٫Ǔ��)��n��1���9y�����44�D����M3�"�%��l�*޼�$b�	Ay˞��� 4D��H�I��=���3k�p��4�����O˓<��) �W���	u��7D�lh� ��N�,p!h!(�=��$�Oj���O�s��;/�`)��H8|��$	��~�s��ې��A�S�msܠ���Gh�'}�i�w���}I1��ޯ),��a�c�q~v��q�z�л���+�8ly��&�m4F��	��M���IU/8��P�g�7y$I����b)���O���� �%1&+�%VP"�rq�`�<�d�'�~�'����5$̨M�L1ą�I�+�'8Y�DgӾ���ON˧4��E���?�4%(����FW�"����P�o��S���y��a!�**�`��nW�ND��a���1�k,��7(݃��!�>@���ݪ#��ƂM�C�:Ef�Z���*"~	���-�%Z72��Q]>�"Jj���%�P�p�*�G
8=�7�<=2Dn���mZޟHF��4;��m�ѠA%T�xK�C�-���?	�Uj&\z �S�4�X竍�J���=���9�Tr�e�ڦ�� �;n eZQ�9v'�$�u���?�g��ic�1�?���?���v&��O27��N���ȄT�H����e��L�;���J�F�V�Ux��I+��3 3�3t�|B�I�:9^ �s�D ba:⩍t��(�åK?1~Z���� 0���l����/���ଟL���J����t�Ti6!�>��Ƈ����	u�	����	p}��"rx�A��$ÈOι�v��/�Px�iӲ�(&B�u{t�)���2\!�0̈́v���4�'�� &v�a#QLȟ1^D��b��
���󉏍0m���	������92@�ޟ���|���A#"HP��>\�8,�@۔*�(�G	��}��I�r:�i	��^4]����A[~5�ߜM�`��o]K�h�&`�O�7�M.E���5�R�}K�A�R�c�|r�']�T>EoH.y���m7m�P���<D����E3�0	)�k��2� ����k�O�ʓB��ưi@��'K��tBęv�g���	�$<r�i��?���?As�J� 쐼��c���T?i��C
�Q@
�+U�����?��Db�gԻ6`:��~0K�*I����#E#S$��H��F�'�2����?	K~��4
������;��i�l,(���� �'��O?�R�[� ����о_W޼
˓&&��|�?}�� /��	�E&P��.�~��'4�INy��+L����b��u,b�A��֖FC䉷n؊@a���/GE$����*{�V�ɠ+bR���8�H�G*��kJ��=��$>gt��ǣ]4|H�cKg�<"�& ��yC��{�Eh�!�`�<��! ma���ƪ����ŅW�<Y�nڮ� �W� K"��!��j�<�����B�I�kP�Y�n�huN}�<i�V�(�]ا�@pG�P01�t�<I�fS�~9�A��'9@MO�<�BE�%�љ��I�1Z�K���<Y���X<���e�8���ӅD��TZ��ڨ@�U�g� D(B�I�-�죕l9���:3�Q$��]�b�'ȴ8�3�(2�I��J�~Fz�(�1�t�)�ŉ*R��`��� �p>�:c��%j���-p�d�!���2_�E��� nƺ�"�+;*����>��s���{�1d+�#:���id'ҳ7 t�WF!?�@{$�X�䍅s�L:t,=?��ԋ���y҉���=lڌ��*N�nU��i�'/��HG��'{NIP�(�9�"�+JT�U�4�*�'�|.(������%*6D�k���M$�B��hO�>�%P�x�D�ݓVp�SD8\O"Yiǔ|�.>7Ĭ@%���`�^d��	����r�a|��\����S.F�w�0���i����'�T���ԟ`(��f"��Ve�N���!�o΢EBB�	9+����>�� ��H,��?�1ICź3�/ �ӺK�o57�E��¸�*ԉ1�z�<y�鈴T���p�^>IBvy�RI�w��Xc��A��(O�>�8��&,�X��쉰h�$�HѬ LOdy�>I�"�6^T�Q�#��2!���F�d�{2)-�W���R6���
�J��hO�Ӌ{��T(��1Eь����D�+�y��"0 �� ̟A%�8�˚��O� ��)P�!؋�Ɨ�ic�ϑ�!���.Ƅ�[���M����΂'��ɓ�Q�"}��a�'��|� ,�h���$�Ji�<�!I��0�@�����=_7��Q�@�o�	0z��{�#V�4��	U�Q�a^J`;�A�ְ?��
�O,�[�I��y$��+$�
{P%��"O��t���Fn X9"�L$-����'�	%:��>�p�D�.�8��a$Z�)S��!D�� ~�
g�Y?�b�.ϔ|���X�� ��)ҧl���궫Go�֨��m�/"�� ��o*@�+�Y��,�#O�]�A$�,I��'�
��%�ۄ~�@|�Db=����}R� 5?��G���Ot�J�i%����*A�\n��"OL)���!�D�Z�Ȝ�9y�m��cԃ�d�$�hˆ��l䋉��5�L4)�����M��$�a�8�y�nE*:�
�R$�=_�|h����R���N��FW���?)�ቅ2X���G?q�PG�\��䟹<x����~��l�jsβp��)u���ēd�a|	�j�n���@�&�NH���O���'�DT�TCN�4�
����O��t��c��U\B��D {�F���'�\�a��\<'�h�Ǐ��D@<++{�ͧO�l0���k�g?�]�m$�P H(�̽ ���C�	�Z��	��W�T.�y�w��[��Ƀ5+P�v1j�a��/�^�"��L�?7*嚠��15f��I��be�����d�+w�[��5��D*ŗ81���Z��\�U��+ �s.@(Ҽt#E�2�	)װh5d��Y��O��3lx3�L�������
�m����5�:�`b��Er9��ɭXQ�@y��� '�[�����Y���)
��Ѓ��vZ"���)D����'�B1����+`�-:q�g����ah���>�҉D6�����^����E�<q�L�d����2�O�	�;��G��$cၕ3��%���;�� ՝i��ir�"O�����M�0gԽI�eZ�E���K4�U�=&�M�����%{��l(�d؞{{�T����r�<a�ꍏR,p\����>P�d� ����8�����%�>E��c��P�A@j�Z�~�!�D��$�pl8wH��R�Z�`��үu��I!C�Z�:e��I�ay��RԴ�A1K;?�^XB�.վ��>Q��U�c�ؑ*�O�tM�q��2u6)�a��\�B��-��TH���aS����<���=٦�K�1�P�-8���CN�%qC�ET���!���zB�	� ���8��s��ޫb��D�˂���9��)��+�x�P�Ъ<��R�OB�a�� ǂ,q�
�����j��$�s"�;���ĩV�2��pP�!�<I˓�\R�X��O�h@��f�4M�u���~��$�^�#�oϗb>Z�*4	�� P��I�
�4`)�T?V.�!@L��u�	�b柚w|�MI��i��®0bX��k�NO�(�6b?��,ʪ�̰K5��)䱣R�)+�f�a#�;T���S�JY�Cg圦RT��O�yB��-q���3eTRR�l��@�%6"���8YR`EeK4�QC�p��+Ob�k��f�׉����&,b�dN?b�r�`�˯c�:�@�&§IV��BU�;�#����1 d֞iB��8'4�H�@
ۙFn�V1O
�["�H����M��'�� pu#��1&�)`��	|hŨ��W5
��@�R!x%���V�
(@�#A>"��Ӽ�ꃋISH`�nڙ|�:e����N��$�eⲵ�GO��J�]����*t*����jT&�z憉'fѾ��!�߸i&���%�.ao�@֭
�������:�	g���\6�T�)�=�N���!�S8J$##H�SM���ShD8�(OB����U4RsC�<Y�� ʙ���"uu|�В�	�P�p�[+� ���
.���`oXޱ�%��r{l���ɼ��gq|���E�ԅ���c~"���(�s�%ڈD�z�(��'�_
��iWݑ \�Pr��+}������5t+�1QP�D�!��B��iv��F�Dz���I�"��A�N!����	 �`'H�/��'�,@P �#CxP��W�P(Q
4)�7M���~��q�y�!��s"���8$���@�ئ�1��&v�ZjGⅵ���dBDiH�x��އi��a뛂:�\8��ĕ���]�Fk�#��!�C����ڬ��D��
$3��R��>�} ���*d@���'X�^�{��_�px�"<�0��V!Ɯ��E�0����q���O��ȃ�(��'�&�!�˦�ц�vHZ1uC�&@5�8c)��h����ڀ	��ק��UKg�>	3��.M&`y���2�'u��D��n� P<�C�����PT��Jî)��7M
�pM0�ш�Tq���O�lK<@��	����qp��.W¬*�ƞ&�:��!�|��&�>�],#q@���i`R�s3�ӊw��nҰ[��p�����D�~,��-|],��'��x������U>�<ٱ��mr���F��p�B�[�$�Fy�n�66�J��'�"����v�S�KHq�1��,	�5���θN�B�hp������� 2[����D��0g
�� �a�d-h����d7H�a����JTP�e,Y�Aè4�Q��]!0�`с��W�A���2�� �C�I�L���*�"$�ap��L�'�X7�W[����ı�:���T�<h�F���4��� ����KŅ/7��âI�7en��)��'Z>5�f,�8�8!�	=z�p9��R�s�"�a�cN)*�|�'�<Uȓ�SW����	�h�8��J�3R��:P(ɯ�$c�b��%O��;&����@'J��#v����U�vo1t���	U��݅�(�@��x ��x�eK�	�,(��	At��O�Ppt��ؒa�w�4�@��r��Ǌ]
,��TPȖ"OD9��DN*�u#CK��,v��X%�iÜ����D�kmx�z��>1eS�v����M~���bz,�s$ƣ4����AÞT��8ZsJ
0�M�r֐	�.V�J����KU���'?��3o�#�,ȅ㉠G&��zPHL��`B�D�?7H�#<��F	?@�N��[󄞣A*����dH&k���i���#d`N�8Q�Ƙ
I���NԴ4rE��2Q
�p��=O%�Ȱ���C�X�r��)D�>i`9��wWd�J�CT7v/!�ď?kB%I�A�$Za|D��.?r�\��l�DE�u&�5h�K�"~R'K�9@@��Rm�6&��i���Ui�'��&�	�t�1�T��Ʃ�dv��hv��9�+&�>��lq'8+˓fR��I �?��J-J*68}y��$��m�+7ר<�b�SW>���9ʚD�� ���d���Eoh<�VD9u��ƃ��W���)RlD`�{+��l=�H�o ��.�ю�dؒ��İ�F6��L:�CV�Maz�BۋXw(��qk�
$Ă���(ĊD�Er��@_���G�:�V� a�'B�x�B�,z�pՈ�	Y�}���(�y��ف���E"j�ye�׾R�dP�L~RѠ*�M�f��s�lp�LR�<��A�e�����;)��T!	K�o��hV���;�����J��!��L��T��31�H&KBi�ÎF8ȹ���>4�IDC�+���`�!�j��@#׆�1F>�U�RoZ�u�љ&̎6we4	s��dދq�B�a"�	{�t�0�7V��yb&ǋp�D����6W�� �o؇?���3i^ql\U��*R� �e���;�OX s�n��w�&��P*Q-+���3�|b�ѯ.���c�M3�b�QG̒?�1���']:jF �c+��"�"O���WƘk�X�j�*)�T��L��|#j����8A�b��`��z���,��qSvj�8��5�&�	���d�� ����'�ԏ<�X�0�dP%N*282�Z	}F����'sn��&�K2�q���HM6��qۓN1�y��<�Ӫ��h~rp���O�f��i��`�b�<��l�6>>�R3�*n�h�"���Y�<9�C�'#Y����.A�,�(r�<�I���Ψ�cի�.(��Ei�<	���,Y�R��7ĉ�<�\Es�O�c�<ف��Y�ФR���2� �@�Z�<���[6��+�M#>f��T�<a���(�>��K��z���"Ei�j�<��)'0��k+۴D�T�"��\�<97�p�9����37��B�i_�<���H��aw/��S�h�C��g�<���k�Q�KC&q�AKE�<�0λH<�H�$��@��Hˇ�Bn�<1��3.�@����ށd�D�7�n�<�f��5��e�?DD�� �d�<�Lخu�Z��WP�΁;��~�����9�ꌺM<�p�8fr�)!	�!��AE�b�<95ꉏ�q� b��`���i�&
Gy�mC	&��:G���哷s�2L��H`ؕ�ȹo�B䉺+;,uBw�Qה��d�$?򁃂��$å���'Oj�'?�����<i�$��7ŬiVf"�O.[r�] o�l-1gFk� �ɴn�	Nv-��,�pb�~�J�0��$�M�|)6Ua�n����O.ɒ@.S�3���d�~"��X$Ku���S.5Д�E�_R�<Af���t��4���H�A�"�aD �<��l�'GI� '�A~��)Z	]�"��f�4i�����#�47�!�d��3�2e��`T9���;�#ޖ��&�8��=.�c>c�HR��	7j7��p��'�:1w�9� ��D��UF��a�?ΔH{d"��G�҅z�!4�O���@F��A�����[J$��"O� 0<kD�Fi���ŭb�s�"O�$؂@��K:��_&b�i�G"O��PbLW�t��8�K��B�i�"O�9pe��/ ��Q:���	;q�q"O(�[1K�,8l�C�BK�d�("O4d#7n���`������
�����yB ��Ո�)͛*l�㫚��yB���Dj@'��O��0P�y"ε*�r��͟Q�$Y��F�yb$�)��Q�	ZM�T���ج�y�L�{Q��4oR�S	[SFH2�yB%.rA +��H$�5�Ҁ�yb��B�\b�cѩ\.Z�j��y�+9;�p��ុ��,!�@��y"���@5�Y�� D��OS��y"����%i#��06�ڶ3�!�U{�b�:�J��&��Mh��,�!�d,�	�
�v�@�0�^�!�	�-������㑋l�!��ڹK!���5k�g�$�bp��?>�!�d�/2˪�;��4� �3g ��!�$��i����U,Y%4`�{�?=�!򄃼%-l3�S/n^�����!�������Z9H���LP�[!�eZ-��nfC�ן�X�����4��MY�H��h�h�&kV��_ep�dBiu�]�Fں+�,��P)�	(�G��Fq�� �Ʈ"����S#����dO�Y@�fP�Z��m��zK�l	1�W�_����NT�C����#@�E�G*S�^�^���@Éi:���U���"�& Pp�QnQ�'ż�G{��<T`(�{0lCނu@�`Q��y��X
n!��C�H7n��s `I2�y"��d(�١΋�Z8�"���y���iP͒Flޓd�������5�y�&��F�RqPf�*['ҥ
w)��y�wG\)uO��Vq**�h2�y���dS��J�Ǒ"L�^@�����y��LNlD<��a&A������-�y�m/>�"}�d�>cS.hhW�F�<�ȏ��a���x����� l�<�0�e�t���L��uxr%�i�<�cʰ.dy�!�+	�x�g%^�<��P��%B�(|����X�<��O3�n�p��Ǡ?�]�gl�k�<�&!�xM2r�QK�[vUq�<yg]%@=�eCA �"}�3΋j�<i7gA��m8��L�y��0����<I7o �w���*����Y���B�j�}�<	ᯜ�X��\:��DK�����e�<A�W/%���C���`�x��֪�`�<��`���� ��@�pϊY�<	1Z�7Dx���`�p��{��P�<��M������>xT�Q+NO�<q��ߜxn��q1/ϙ Ǌ�,�f�<�LP�tyFų��7e�����e�<Q�n�/>���	�]�qf�V�<	�
 Z�a�L�B�.��&D�w�<�'�;Y�I[1�C�/u����v�<�Gh��E����Ui&Y��p	����:vZ��[��[f��禍� �����s�^��c�H��Pȓl��%��}�d��e��2���A&d�h�n�o���K
nV,0`J��vj���#��I����b�'����-��#HX��'ǜ)gh���DԦxp*u	&�2{���5o�9ZiDm�	(����`b˽Q�y��i��.��&")�� �q���ҳ&�T��1n�	K��rG�'�(<i�EE[c61����
7d�p����<%?�0���4T/\�A��Dgt� 	�l_x���xb*�z䐅�'��y8Ӣ_ 
QK��)X�=��&��c`0�D�O~ *@%��$``h��OJ@R��gQΙ���8 6pÜ|��?�6	rǤT�3}�P�qX�O�[�m����^�\4[W��h����z0����U�1�X">�p��*��٣3�� 8_.8�BLR1OJ�v�>q@�>�b�ވ[��}�L?�;�@��}G�%����^N��r�G�S�D��lM@X����N�d!ju`�ҘS�h��*�=��q'�LӒ�E���禽0�MJ�|b���+�z�
a&���X��N�"ZB���$�S�Y��F���d��Q9��(�N�=k:}[u�T����*#r-�U��R��u���
k����I)X�n1�я	����#nQnvO��'fA+.���O`e2I>r�ҊX��A	EBG�?��U���o?>W?*�B��U�_#Ux���˯�b����٠$�N[�BG�_:�h���MK�H��Q?��L�h�ɪV�b��=Q��L�!Q�A�Aɓ�����	e��%X����>I���1\}����
�1�.�"�圯��6��\R��;[u.�q��<��A+hg|����� ����/9��S��	2�ه�U���Q��)r!�$L0b⽲wm��@��� ��4�$s�&�)�vX�'t�)Đ�8/�\��)@�qC<���Oµ����"-�Y�I�Aݸ�+W�|�Y�]��)S*LK?i���j�|� �hĩx
��abG��,p�	+��-V��#��>b~T������0<Y�-C�m��-Ò`�/&u�)��_2U�"T�|3e�|f	��]s�BH����4h>L���r�n�����?����3�L[�,Q�J*ڀ"k˕J1&)����5MT���B1�DX�m�t�]�n���(rI�uk�썀Hݤ\��&��V��䝠]�]��.�UgV� ��J"w�\��4�h
X`[�a�,>l%r3/Sp�����E�&���FB����~#��PD�.{nlh�ɟ6%�'�nmj���A�	�3*N�ME@����42X�qcG X�u�Q	�%.��I%��8w�d�1Ju؞���	$h�,��n�F��U��~��A���R8	`��i��N�A� �=A��0�Ի�ĝ	m�b�rBF�}���!f�� ڡ�����ԥ�0�˒m�xMs�+�����CMzܓ O�0�p[���)n�@�f]?bե�('LݘǤW��9F�9<OܚìG7G���;B�I �j����Q&,"���1�*��ȥ>q�`#w�$��RAF �|d�a�S�p�{b)Ȣ�X���<e.��Ɂ��|�.����7|�-x5ɝ�
X���=��#X*sL	�]4�L�y�L�H��� 5�Ա0��dA��|��l��œs� HUC�+S�)H�gͦq�Z=;�F��D�D,�9c&�Uj�=/�e�&@P����@�+�v����,?�N��e#�+_,J�W(�Sj���/��L�"�j�q�ٚV�܄ �Lа�X�B9�|�gP&c��	)Q+V�E�џ��w%F��$�#�T��h!R�@�r��8 �Y�� �ĉ
�,��'����d�T	�`�]� 	�̌��'��å�HF�����Z�ݩFí<*>j�j�`p�
-wmp�����!����yEO�{����/`���s�$�&*��u�#��a�h�@�a_s@�y"�DK_�|Sa� \�j��e)�*d�H���m�U��¥��8��OFSǪ�'odX��_U9:I����X-�d��4o���+
ߓ,����R14p$��CjH��F�XS̞�k^(A���՟�ç?��嚰JŸ"v��*tm�a�$@Y��l\Y�Ƣ?���@2��aiN�1�dt�M�h!V蛥��)6<�%�'�p<�4=34qB2͖�";��c��c�2G7$�x�'g/p=ju��2��#hT(�2d�j2~Y��
�<���ڲU����a��
@,L��� 
5J���|B��<M����2F�P>����jא0��i9#DL ���,-/���R9"l!m��i �iǰ�yr+�;��L��Dy2-0�)�-7��1D`� ��pJ'� w�D�6��.݄ J���kѢW�p����.sR6E�vf,Y�F�W�̽rFiV�I�P�����R�E��A�kWV�p�N�kM�����W�X� �O7:��fU�|{6�@	�2-�f���4ѩ�$��	�25d����?����zDޤ��]*m�����F��8��'ČEIȤ��n�| �ɉ�>rR��Eqn�ە��f�oZ�]���b%���GR:A�&���G2	H�'�PM���ܭ �ɧ��ݯ$��)Ƥ��c�vi�����H����^��zl�$O��(��6nu�H�gi	�'@fH񒦔�Q�I����V��I&
�Ȣ��0�= �eJ)bu�L��!�I	&}�l���hb�!��k�!dܦ�b�'�
�*v/�S��y��4h�E�o��B���0�!����A��-B�%06�*r'�n�';t�Pu
\���YaIb�L�3KQ���Z�)��QTqP��ޔ|3d�I�Q���[eA%a�|M�5Gq���f��J�^x1i��43����J �Y�v(����)kn01�>y&��!m�-�"훁9�@g睩#���'ڮ9�G �u~N�{ ��?A-2-��钓]��`Z��˼;�FR� ٨a@�[�t�RPܓ)B�(���d��n��`H�b�h�*5� "�?6B\ �j�S��e�ҫS(j��a'�B��0��Q6(=:��*�!�B]"�b�1:�d��'�*<h@I��+��wk��Ft�4�ңF�H&���I�C�8hєiT�k~L@2*�h�d�F���ۆʑ�����6&U�>6��2;�8��H�uF�����7i��(�/�4=cvd�'�I'����Y3#R=-G��h�8xXl���9Ӓh�(X��� ���T��n��ఆ,P#I�8u�R�+�<�r�	.+H4���K�g�d��Y�h���F�%\��0&�gv��тf�l��Թ	k"`��f��9m����B�]��$�Z��.��W�@i�� 9n �c���%-�qO�0�A肶,�|e��{�AZ�|�"}�T�
=FZ(�+C+,�!�Q�OO��#ĥ�r���à��<�Љ�Z*�#Slj� �U�_�<R%��[N&�3�LL14؍/R�t����g��t��쇱`\Q�\'6cLʧ~%�K��PN��<�r ݋T��%ϓD�
��� ߳I�P�Ks�N�>�� E|�%ɪ���p�e�#�ڬ �����~��!(�x=Sn���N~R�n�?�`]�q��<y��U(QS�؞N;���ݳ�\�D}�PE���K޼ѿۥd�<J	�`A��E�n��Y[v)�1�"|OBWӢ����bψ:0�puBB0�H	�f+�Xܓ$H�j�'U�FՃe����'�d!"�&�Xu A$w��|i��D�,c��}����n!��f��o��dH+ɼ CeʝT�����=m���Д�TЦ�Ka����5Fy�<�Rh�.�(7&H�G��A�S�<�i@�2��{`b1>ԓV`q�'D�Q�!)�h��XI $�2�&��U�,ʓE�)�+(9��T�c��<��!��mP` @��A��(�'� �B<n���h4X��{�w]��q!DՉo{����.�NҊX�۴z���d_�����')�,�붿�p�2�ɍu����lD�[�`4�|dT�a0�`s��Z���?�O�()2�׍"��T��e�18�vس�d�xv�$��b3~�*vZ��iо�y��P>>o��SR��$mɔ����,~�
���.�e�8MВD-Nݰ"<��O|�"ng&�{�I.Gj�������)�vnR���p�N	!�ZɈ��">9��V#�����@�,�8�q�L�,Xn40��DL?i�+֮C}��o��}ж�Ǩ����H׮oe���dD&&�^�r�cǗr�\9Za��;����$��7�صȑ��3Eay�A/���i�+C?'
$�e��U ���k]�GEz�@B��:�L�?1&&�5��ED)m�91�g(c�v���cW��h!����^��ZL<�F̑+?=D *� �.|p���E`�^�jv�K�Z������4���'�j��S�ST ��ǒZ�����dB�M64{��
^E�t2B��i�&�`kQ�Gʞ��Q�^�p=Iݗ$d�zs�Y�jj����d��|KF.�w����ߏW��	�c]9D\1b�Kޠ
�a~"g@�!x~����=�"���X%?a��4�Y
�0=�C���pr�d�$����X��`��+�h��`hO.�H��{�'o�9���b0�׌[ e�R�A�'x(�Ȓj�8rH\��b�"%~Rp��y�j�e�Rq����l)f�'�ԕ��'�nut���2|�]�B�� �?VO�=. ����j�0��NE�'��	[�IG�P
b<1�A�Le�i�@���ut	�(�3�� ��t� 0�T=�2"�M�Y��\B�U`1q���&k��P{>�S�(����!�kd.1�CŒ,��4S��'�5Q㮏Y��-��#N�Xc � ]9Rχ�P��R#_�� S�ӗ'�l�J��?@��`����-)�XY��#OT�R����cGM&�=����3U¬�`��4zؐC��٥>��E��>6XڗĂ�X�P�84o
�8<�aiac��y�,��	E�s�a����V�&y�4��'�61�#�V<(���$�Z g E��Rnā&؝�p�@4:6���Gl������Kc(��4f�ƹ����0P��Ϥ�@F��q5O�! �ԝ	
�l����PH�>��� �'�;�>tÅ��M��a��,D����g�RPX����E�T�ϖ&lq�5 ^�rz 5P5	�0='_}�����2��5[s��w�U��"8`$�$���y�+��|��'
k�p�J�A�	�ε�C�Ӝ{#L	�7!^�7ʡfԐ��Z�ʠbİE48̻3ʄ >��4�=��W5U��������P��T~2ɉ;���*�-h��ਢ�	<��=y�j\�m�>s$CW�%��*Q�-�$�b���tt�,\O�j7*���X�(��~-�E��6#�lC�A�%	BH��ɨj:�t�IW�H���!�J��LѰ@���]Ѹ'ؠ#}�ӺS�$P��Q�G��7K���� IMQx�P�C�����A]1E��� ��	`����K���7c�Ʀ�;��>@��6l�v�0�Ϭy�<	�1F(���f�(ٲ����C���'�ذ񦙷A��a�ʜ,&���4Y>�i�!�fo�!�u��n.�,{RH�O����� ��(A���ܒg���D�>Pf2#��6��|�t�Q zR4�aN��a��i�@�O�#M���s�>I8˟:ـ���8t�KT� 9�><����-H�!��[��^�XDG��cl�9C�L]M��$�z:�7mhӚ�I�Ǘr�����#�1�BS�L�5�X�6�Œf��1�"O��#�"�ul=�T�������B�B�Z�.�>Y-����#U��JL�D�e���T�\q$#��(�
=un>�OF����1*uK�E;]����0�^(y�*tI�U�0?�"_)#�6)kQ��#����t"�w�'��0�`��V%�|2�#|��/�L��X��:	�L�����yb�-]�:=�v�»"��:�I^�~��ٕ��$���1r±��S�Qj
�q�fZ�`�J�u���4�:C�)�  �@J��.���Zs�\q&�AW/K$�dǺKG��7I���3�IH��gH��&9���PH���$�l�h!�3�_�N���$n��eCɂ�P��ęu���0?��ᅠ����(�5h�aa'��o�'�|  ����@	��~�H�Hc  :cbB� َ�R#�n�<ɔh[%r�0��G	��e�����[T�<�p�Ac��MA'`�4LqK�O�<�G��(��-�r���,s ��w$�O�<��
9C�V�+�G�> q'QC�<��!O>���H����!�B�~�<���;\���""��A�X�daDx�<2�!%XvAr�͆m?0	��P�<�s땬ń�E$G�)�Q;,FM�<�"��8�0��4u~,`A�<�S�ӜF�!�Q��vVu b�@w�<��o@2:b� �)_�<,`��Gt�<)�� "1����B�U)>�h���l�<�3���$�п2F�=�l�q�<�U�hzt,stœ:9zxq�i]j�<�GPQ[����fXy�xi�h�<��1~�(QQ�g�	Qbl9`��|�<	�J�Tnh��oڿ�� q£^w�<Q�`�<pP�0d��y�(D�K�<�e�PY�dX�.�D�r���(F�<qe��t��!��K��M�w�B}�<�s.ؾa���Q�(J.whKP�j��C�!��|3��7a�� �"���u��C�I��,��
�/�h��D�%t�C����\I('1<,�ǉ]�j:�B�I�'p��i��7V �3��Y��B�ɥ`f4��B���ʝ�R�9+�JC��_Nr��En�nz����ɛ�$�C�	�R�$��!@7�����4n]nC�I#- l�9�G��"v^���քA�DC��W��*��΅!�P������C�I.��HxTO�5�,�͙�Qw�B�	�z��Hy"	
!paj� �h��B䉠.�X!	X*`�B���V��B�I�a
&t�����yҠu"�.ʕY�C�	�� �pfP�|�&�� /� oxC��1^7��� ˗�T�ar��~��C��?]�<@a&(:A�!��4ؖC䉑[��q�Ѯe_H�c��P�KqzC䉋	�lxI�OŚ �"H�qj\?dK�C�	7	4 ����K'>�8<jfk�Uf�B�&4F~<J��D�Gެ�c(�UCrC�	�cԢpHĂ��k���I�&˛h. B�2Ngv��օ´w30-y�%ˋ`��C�I�,GF
�	����ԄH�%4�C䉟s~$k��=�^���A0�tC�	Q�P#��]b*�#_�?�bC�	�n7�зL�$~6��ek�O�6C�I�,���#��pn�U,��D�2D������onl	8�Ď @�b�%D�p���T�|�`�Г'�t�
���C&D�ĹC/�57c�QD��:o2Ta�,2D�LbOC�c�`U��F�Dr��Ad1D������(Wx*�"ϫO�5&�-D�|
�Ή#v��GN�׆��uc*D�H��'A�ab¼�q�X�Pm�q+ l2D���0�i��ʮ;�x�xAE3D�$ِ/��>��s3'I9Q�rAA��3D���`�?7�BQC�ƒ�I&i��!1D�8�Un\zܐ���QG�Y��0D�� :��dϲ'�,�[@ŗ�#�F!��"O��g g��r��w�~<b!"O��8�&�  ��iR@ĽO���0R"O��8׬ęL�ڥs��ǡ&&�]��"O�вea�4j��Uk�-V�*��{V"O6L�Do�<O|�Q��l�%'�p`��"O�X�b�/��dѤK K���H�"Op���-�bb��k�;�4=i�"O��ctE�&fVIpK��Ot���"O
��ġ�-Fhd<X���+��L�W"O`�P�E���<p2�E7?�P�"O��{!ቓa��E�A�i�D"O�D�I�x �`s梀:K *l��"O��@�DU�$B����,�f�@�"O�Y�-�8W
|P�¦�l!"O�e��(U#v����?�: �q"O���QM:zq��iW�G�p�"O&Q �0��Q4(;J�"�*�"ON����lJ�Q�Y��:q�"OP�`���!r�(]���
�6����"O��90f�-x�� �� �,u(��@"O�\2v`:,��� E�'F�
D*O� Q��ڱ(y�Ԩ�'�7g0���'�
��7,P�s̠HI��Ǧ��ua�'���_���]���J�|��"�'l���fK�$������#��(��'2ؔ5oF�" $XI�_�5���0�'�=ʴoP3KP��a��~f&<��'6���a�p=΁8�[�{�x�k�'#��Xg�D/w��h2�M
tt�b	�'���:%��n�*�؁�� mվ$��'x�}X��+&6J����2�`��ȓƔd)�-�.X^�j�F�0�h��B=|e ���]��D�C0V���ȓ6��-��w��$��/��U��Z�"И�K̔i�|�r���I��zc"���)|��@ #�i����q�^�
Q�NzmpA��a�^�ȓJ������=|0�yM�ȓ9�V�+XE��^�nK~e�ȓ(�FPKw�
��b�^:2j�}�ȓY�ZUy�*O>�tu��E��$Ih���2�p*��@{x{�'�2*�l�ȓs�t�!͈�^z��R(�7
���St|4���j.
��!#Ժ,�(x��=�ҍ�g�,wF�ԱC�и�p�ȓ�V�*���A�@d�֬�E8�Іȓh�V0�G%J)}pԘ�5��6=:l�ȓ���aP�Ts$�@Y�ϑZF"4���L)Pe]G}8�����~��B�ɱ}��U�gM�0L���;?�B�ɺIA��S5��D�Ba���C�ɇ�Y[��F<.ލpA�S���B�	"^�)8�@��@���B�#� B�ɇB���Bg�4G��M6��C�ɫB΁�K�^��Iɒl��4P�C�	0a<Xd9�O+-o�ەP�'��B��. n�Ĉ�1X$���� Q|B䉞J�Xcá�G�6�ÓeK�U"�C�8i;قcO��c�$��4�V:^�C�ə:�������%f 4{��R�?��B��&��"�V�"J&hc�9H��c�'�B��	�lQzF�L�X�y�'�&�և�AZ�8#w@4:����
��� ����ҚU�F��,I<;W<���"Or�2`(
 S��z�D)�LH��"OY���ԆY�PĥX�U��8@ "OL��ǜ?@L��V�g���"O�t{�<}H�� q$�败�%"O aj���!f���wa�^z�i�T"O�,��J)6*�sUn^#`F"O���qa^�1�)��.C"e\~]@�"OB�됍W�Dܻd�6wt�4J"OX	�gE�$ ������,QA"��r"O�4��Ä<��-:G?Z=�`�1"Oر��B3�Ѓ d	H4b��"OL	���//v���B��U�܋�"O~�b"b�-\:*����
2�����"O,��K9b�ta��J%	|�J�"O�ݲ1� �gR~���^�:��!"ON��6�wU ��4$�6{l��91"O�iP���j݁��6B4�<)�"O�E���4�(����6�#�"O�E�@!�?���q��-��D!"O�]I׬�C�,dkah@�(��B�"O��Ѕ��,$ȱ��(K&H�� �5"O��9Q���q�`{r���lή���"O�ph�A��7Ўe�' ģ.��æ"O
5Q�+ܙh"(��%�c�A��"O �(Bw���B၎�&�l�r"O<,;2i�߸q��aF��H}y2"O���宓�;�B�bjD�u��{"O��UOG
�p���^�N�0��"O<�B@�@ �`�hH'���j�"O&������Lr��#-Ο�h-��"O(8�bŚ3K���Ԍu`��"O���D��N�n,[��=;��`�"OШ"�C���`a��?V3�
�"O�����
��T��U�R�k�"O� {��۪f||� �o�^u\�Zu"O(\	%o�7N��=s �_�^��A�"OT�0W��1-шL`�+%eI�iF"O>!3�:.����2�T4l��YY2"O(���:z�4j@��0�\�r"O�M�\�"pB���P* ˦%��"O��
����Y�H(2GѮV��К�"O:���S�j��p -�0Z�*(a&"Ov�0l�+F3t�:-�#a����6"O��S!��!�� J_�&*U��"O�����B��cE��
O��-Rg"O�\�,-J�d`�MG͐�"O���=Gb��A���F��Q�0"OJ�I�#�:9H�� ��m@u"O\$�R�:.xH��aF%�Q;�"O�)��_=.��Ū@��LZS"O"1Ð��41�<���ʐ�QSq"OD$Pro���e���k.�Ӏ"O��sn�|5,}Jf��F�v}b�"O8�
���J�z`��.f�8�Ѕ"O����H�~���ۢ4��I"O����P�Q�������,(Ǌ�A`"O.���9a�����F�N�#�"O���-�@�9�7��*GF�˵"Oʈ��J�;hBy{g�O:%�p�F"O$`�ce
7x�G*�?o��!�"O(��d�O�00�iXaB�`f6�[P"O��Q.�?9�Ip�@߽�2���"O�uX���a�d��`W�Y�:��r"O� *���B�Sd��0@��,���"Oؘ�1Wc��/@���y"O�e�,L[.��!A`R K�T��"OjAb�,a��Kp��.�c"O��&b@t*���d��{*Y�"Oh8��H�ZL!"F�=�P��"OH9���"[����A�ޤL��!8t"OBq�O��9��Q�h[<�f �g"O�p 0��:|l��(H�}� �"OVQy�L[�'����3
�$�j�"O�9��)ƻZ�P�'Ɂ,���`�"O��H��'�bt�e�UWP���3"O�QK�A�$ݒ@�QR�
����"O��p!�H-#W�-�kS�w۲`��"O��C�tj<X�	S.�8 ��"O蹰��ǽ���B�怔����a"Ob<Z�$�@��z �
@LYr�"O�-�aѼCRt�$�?1I�e"O(1Q�c�7�6��C�!�Z�"O�I�BU�1o������%{���"O�1A��R,��JP���ڗ"O�[�IJ"k�H����x� �0"O�ܩV�Ɔm,�J�"�J�9qv"Or����S5b�A�g���3"O���FI۱<����d�ެJ8|���"O��i�Z�,@9��Հv��؈�"O,�R�eA9�:�C3"C8e���"O�u��j���q�@T�`,�A(�"O}IT�/z<J��n�5@H��6"O2(�AA
x�&y�v�Z	P0q�U"Oj��@��?��8��Ȍ}�`-��"O��B6d�O!�I '���.�VD8u"OȈ�4�..���T�W�|��,��"OP��썤c�ʰ� :r�H�"O���c�9�LX��\	�"Od��Ƈ_��J��T�͔_Pa:�"O�D�`.&Ff�;%h��m1�	"OR��!)�<t����Q��`�"O*���G�?C��E&�O��8�4"O��
� �=z�U���I?B�`-q�"O�,!��$5w��U�$s�"O��j%D�S����Zjz4��"O,Aň�"9k��I1�9wW����"O<���C�;0�����̓p(NX@"O-�0�/;�M��f�o0�"O���e�Y�A|�s��)�=�"O�0!ǬI�z4�E�Ǆ�#!�Q1�"OR�2"��	.޼�����%l�L�<9u�ː!{�9�H���D!�C�<�0Y�r�^e1��Gl=� ��E�<��#�9���R/TX��j��AC�<�EӧPmX�(���H���!�{�<A��
r�q�@j�adnd�ŀx�<�&�D�vjdU �n��xf�΋t�<Q�O[V��S�c �H�Z0  n�<A���\��Bאh��8���h�<1�@�O)���@	�8��b�<i�b" ��9  �m�H�)`l�]�<��-'Z� P�ޠ=���dT�<�%��*7�X� �I�#�2�$�Q�<9�L��d~��CGʷs�.����Vx�<I�lU�Blx�̗695`D9T�N�<i1)L�ey"�q�a�s� p�N�H�<Y4�Z�?H$hC�D�7^R�+�N�<� ��x��Y=Q�b���ˤs�N��"O�lK�ą�l]��!���Z|�$"O�<�j�(1]�)[�K
&�&"O�܁�#�-f���r�Z!�"O������H����' �g�e��"Or���*]�f*�2%���|�"9"O�] !�ZH>H�����A"O���e��yڑ�"�G8�6#�"O,���&��,����F�j�Y�"O�{���#�8��\�uǐ@��"O��xPV�'��b��H+e��$�`��6\O��O[)<
ŘqB^�lǨ�Q�'��T�~��T�[�b��D�¼Μ �g"O�$���..�����/�%T<���"O ���,�r��]��n+zLB�C�"O�����5�j��t甃4P>�+�"O�����_�Ű���T��\3"O����2)�\�AH�0P��R�d&LO^1N� O�P�y��V�>Č�"O�� @[+0��QIAFI^�Pe"O����Ŝ2 ̱�#�:H��ɐ�"O�i@�Mq`!�v X�l�ܬ �"O�@)U�9Y��ño�aA�0"v"O�|��̍):�^�J2�Q�f���"O�\��J�^D^��'ڗ��ňQ"OF51��X��t��L�)g� �p�"OР�@Ĵ1�jU���.m�M3�"Oa����*|T�@�Ν�'��]��"Of�*��}�hmqa�_���� "O±���J,�z)��	R!�$�Ie"On92`��&�����1{���c"Od���ȉcX�Ȗ(̊U@�"`"O�D8�I<~�T肕� 6)��"O$�+���;~G>䩅�+}#Z��"O8�;p!\.4��E��+<�l��"O*ɡqȉ<�,��秇1�T�""O�X�'Y}�t	3&]���Q�v"O�bu�\$;�nؒ��/� m�c"Oh�af�7P,衧)�Y��"OR5*Q��j5����<M�V�;�"O��1�%��5 į�<5��Y!���1lO@M�A�%B`KT�@�x��!���x�)��"����J�W�ި`%H5c�8B�ɲ� 	�vf��^�
0����B�I�H��P�'��#,��9)P�  {.B�I5I�S.	-:�A��
oDC䉿[J���W1E�H�v���2C� .�x 3<8�:�`�;j�6B�ɏf$8�jI�r��Ex�<C�ɐ���oL$M`��#Y-Q%lC䉊4q��(�D�V-���RaԘ#*.C�I?1����6�U?0�xb����*޶��d(�n 9�W2�DA��� �x]��=�J����_�.JpI���;w�p�ȓO �$Yw�ܪQ `�+$��7�&���x��d��e�9}Ne�M�_϶���X	ʉxsf��mx`���G�i�zt�ȓ\�R`ҹ!xȈ�Y;A�(u�ȓB0IrSf��f'����A^��X��s_�D�%-�*´�+�f�,�H�ȓV�ބ@A��%�&�S����_���ʓ��a9�G���		6��,u�C�In�l�:��҉�F���.�
� �<��Vӌ�ї.E~�d�"���$�T$��S�? *����7L �!d}���G"O��S��� @a7oҠZz��b�"O�!@��$�8ڶ+�6!a$���"O ��D:���$MA"J��"OTp�/�X�d��Q�i��q"O�!��kC<�D�Z0�Mn�1d�'a��'CB�-uY�8��˱Z��I��"O8�Ak�+p&����A���&�'�!�D�00̋�I��}��'�
+!�dY$0��<c��Pो;�!�ē�E�Pz��1V[8�A&ʬK�!��֭j7z@�+�ufؕ�0&^�f�!�|I����c�")ڲ�F�/y<Tq�'��E���;��2C,Z��ɫ�'��2킁R�Pd:�	�>����'��� `UήlC3�=�V���'��d�v&�-v�L���.F&+�2|��'�h���/K�`GБ8��Ǔ0d>e���d������T �%.�1��O6�!�$��B��P�J:���֣�)�!�$ƣ%��lZBӜ؞�b���P�!�$�k��b������3���o�!�$�n�:�z$��E���Ӷ�E�S�!�H�^�- � �25|�A�,�*j�!�Y~:5��*.Hl �ʄ�ZQ��x��I[ ��@���(�cM!o��C�	�!�\��gc�:
�p
��ׁoފC�"T|<id	�n��h���4%0.C�.l�~<`�1d�(�4C�^(C�w&^���J0x`��P�*ǓX�B�/g	:��N�|���@(�u���=�çNQ��2p��y0T�z��!ZBY��@=��QPkװM��	�j�N���Y��)J�#��m�3�ׂ/B���$uRuR嫝�e�6�q_�Ԏ��ȓgW��Æ'	R�*�(^GN��ȓbz����N��ٹ�m�N؄ȓ����#�X�M\��)�䛋\wTP��)��Y!̋p�\1�b瑀qӮX���l}r��$C��X�!��#M�	�Pnӄ�y�I
@iѓ�M����R�	3�y"�K��:sv)ŝ]\@$`�,�y"�X�9��C�+)���dĎ�hO����Љa!`b�\� ������&Ib!��6�v��f�C�e�������Ox��Ę-P5��i��&N�D�%��`?azr���Y�� ��H�*oj!�ݕr"!���ZHI�VC��a�=kAa�e!��
(~{�}y�i�%	P�2��G�!�&
�Bq�f@A�2�^5Fl�%:@!�$M�]+���'_�4A��B"O�lꂈU6=B��1���S�~-pW�>����i� |�8�rp�	y0���"i���!�䂑n��p�� �QgQ*]�!�4Z�L�2i��NZ�����!�œ)�ܘ4�N}:��p+\�t�!�$ׅ Ĕ��IX�?�9{��J�S!�$F{�"E	1f�}��7�C <�!���qh5�֡}�P��g"�!��ֺ<v"	��H�l_Pԫ��
bY!�$��;�I�R@L@!�WG_02�!��M�q�H b�e�;^��pj �
!!��	�X��� �a�*L����Q�!�E�"�n�y��U��Pł�SL!�� v�Y媏��Br�!;8=i�"O`Ya�D�a�:��dm�>ހJ"O�eq�&�V�F	QU\C�r4�C"OƁ
R�Ddz ��)J�F�ف"O��I�}-d�j���1����S"OB�!��K�Sv]�B�A����"O<[�G�@T�yvE�cр��"O�`�`@U>��X+�DBC��峦"O (�a"�4&`Ơӱ�Chc�p�"O����*��F"ʐzc"?H.�ѡ"Oֹ��K�-��Q�&g_0���"O,���(�� �4�k�S 6��5"O��ʤ�^v�v�j�g��`'"O��I0*��x ���H�A���$"O����J&�	�.��	|�m��"O��ywd�GN���B`8�"O<�0�+�S�9�O*[N�!�"Oj���΋u��`�`�jD��B�"O���4�9��͠L	�6Cv�ڢ"OL�[R/ֳ2��q4��VB���V"O���k�E��Z�d܃&X�R"O����X'аH���Z0>�z�"O"0��\�O��8�c��dX֘+"O��:!3s<xsIۢTQL+�"O&8�t�_ z�=Awȇf��#b"Oⴊ�����ڧ �:�.�b�"O8�c��Y������{$�h��"O��W
B9f��E-�$�>M��"O,�+f$1��h�� �.�[A"O�a�Β$H��h[q�EJ��K�"OZu��)�@��y2�荵J<)��"O0 .T�d�V�3GED�W�dq	"Oj���f(��Ѡ��bupq�b"O��k3�u����M� Tr9�U"OfM����e��� m��y�t�d"O�aC(��h�(Y�pF.J
"u	"O&l��A
�Ot~<0&UJ����"O���,D:e`QZ6n�"Z�Xt�u"O�T��,^�NR@�K�">�����"O�%X��X������tx�r#"O6-�c���0��5`E�ǀff�8�3"OH�C�Q.���a��|X|��"O�uY�&
��I���E�	J`��"O
�HbI�>�P��FE	��P"O^�� Ğo������dlD�"O�Q�VJ�EA���2�#\>��(�"OĈ��HA�v��%ٔ�\^4AD"O���Ì�/����i֭$! �"O����C^��8p��$Ρ�"O<L�aBڱ]ќ��$lO�C�z��"O:ɒǁ�dZ��
Y{���h&"O�� Ƒ;M�!�"�2}��Tf"O�=�`��=���AB>y� �*�"O�p���U�'(n�IS<6K�"O�����S^.�J�.�0|�a��"O�eJ�m�-9�y�n��!y,�Q"Ox����$	�T`�� D�* "O�q�	�jM0�E��,A<!{5"O�i;�
�<�ҘcAa���pQ��"Oj�Ⲍ�*�ڬ� ��Q���8e"O��%ǞT��� O��Kc���"O�ih�� c�pY���'Oĩ�5"OL���l�>BĒ rf��VCbe�`"O2����Q�b�L��B�ތ6���[�"O� �M�d2z�`�"��W��H�"O:�E�h�iJ`�-�Lթ"O����"4�*@#;t���"O���@�ݪzz)U@�V~|}�G"O��P�,-F̡��E�� g�Y��"O�A��A�#c���F��AR�E�"O� ��z��P�c⟦sR:��"O2���`�*fھ�c��2Q��Pr"O��&�$!H1����`pTM��"O�I�v�́w\B$j�b� u����"O!;�i/x�0�S��9FwjT��"O��6��%W,L�g���N���`"O�bs��hvn�t�۝���"O�I2��9S�0H��a2�,�"O�%�eh}~l��� W\0�P�"O�=P��E#:\���o� {0�@S�"O���`)�g�
�I&�n LQ��"O-�E��5&����Ǎ*xy$"O�@��ˌXn8�"ǉ�؞�Ȃ"OJ��CԴ`��Ȣ�Q�pX��d"O^�x��
��AK��9t?p, "Oҭ���	1l� ���@�.H�"O�A�ԇ
��2)�!��^�\3�"OhH���F�Ъ"oիg�r�r"O����=-, z���;Wct�"�"O��AF��xf.$�;�j�C;!��;�`�F@S!	&��$�A��!��S�Li�c�$X�r"��P�D �!�$֔p�L(R��S"��i�!q�!�$	�&4����ޠn�`å��7`�!�9ހ�Ul��+ِ��Pᇬj�!�� ��H$�\4�ZҶ�� \�!�f�L�d�l�\�ψ	�!򤙼��DB��(P&T��z}!�40�\X��D�"�m;w%�]x!��Q���2u�%�j`�doR8DT!��ʌ��ݶv�
5�p��*<!��%i�|�: ,�:b���҆ �3*!��"ǲtq!��d�t���!�D�) ��!^�V/z� eK5�!�D��,~��C�J�?=
|��!��k�!�$�8 ���R$��T�8�B�K�!�ԟ %����ȫ$��RN�/!���=��h�@�OR^ٳ�햟_�!�ě	�"�2"G�V�ER/ /�!�d�K8���uL�3~5�9�Vn^�I�!�d����d��.�o�����.U	N�!�:h��ME�hE���%!�ē�R��A�A�6f�� �K�E*!��,7 T���B��ً���g�!�B;^��paQ*s� *0��!�D�uw ��� �{tM�F@ͷK�!���w*����H�ĳ�n,#�!�d {�A������y!$���<D�XsB������ ?��T9�l�w!���G�<�s��l��;�+ٹ'�!���T,08(�
Dz��{�K�-�!򤙯;�UZr"׺7ͩ���n�!�$��@<L�l%骔MF�I�!����M8�3��		�D՚qm��Mv!�d�� @�%�-�&A"U#��8�!�A֚AU���-�`U�\3!��N�Y�x��@��O)>q��`F%#	!�$�%an,�AD@-i`4 ���w�!�� �� ��6c�ī�_��JP"�"Oh���D�k�pᙀ&*:�fUJ�"O���kɯ/�H�(����<C±)�"O���q'_�e��tS�&Q34����"Oyנ����DP��@�U �"O�@�g��!|zl� oä=��=2�"O�,Z�I�UX4�XÎ��E��"O��"�F
KJ�=�Q��*���R"O���DϘ0Zx���.@���(�"Od)��ƸaRv�3pd�@mP��"O8��G�F�Uہ��e�`�z�"OD:��2}
%�-̑_��Q�"O�d���3�xU�Z�!`J<;s"O�	���&_eqa��:E�iё"OD ��"�9�B�i�́:0�<��"O0)��ɜ�4����ö+zx��"O��)��)����Ćǰ8&�0�"OH-X ��1vd��@Fܶd�F4��"O���C� P:]�R$��;o.��"O<���k�:S��x�W#R�KU��j%"O\0c�J�l�c፠NP�=S�"O�i���4,���ݏZ-� ۱"O2�pP%�*le��s����"O~1BMM /\��p��>�e��"O�)"�2�A�@�-״l�3"O�#�0����Nlt�}��"O�L��-��@��ب���jl<���"O�ݹ��5\@�*��-_&-��"O��-9���E�N$Nn�{�"O8r�N���A��5D a��"Ox ��&�=k$��㍃a�N@�7"O�T*cH�Xa�[�"N�x0x�jA"O��áO�w�`$�ҡ��C-z���"OB��ʀ.){�$���	�x킹za"Od��F��a��HrЯ]�@�<���"O�T��4O-X�[��6��� "O�0��ꈻ|"�ׇ+#��]"�AF�<IT�C�fD8x�̙=.Db�����l�<	㭔�f�B����c8`�I�g�<)��Eq�r�36�3�h2�C^�<��	�li2"�k�)Y��|��Ib�<�7Ǥw`��a��R��`��[�<EW�q�Ωʕ��}�ep���m�<	 `2�Jm*"AӠ;uD��G�f�<��'�� �)���#F�F��(�a�<����hZ�)��E���@�uds�<�+D3Z���)'�W�v(`b��n�<QSo�#�<�	��Y�@A@���n�<)��))2-h�-� L�x�y��\Q�<yӈ;2����?������W�<9s�	�v=x���E���g Q�<)���2;�dD��/O">Ե�6k�N�<�&Iy���a�ʡ?hAC�^E�<��-_�JSBʉ �����%R�<��ӱIe��p0#���2T�T�<q�K�^T�S�E+�z�B��O�<�F,��T	m�'u0N<"@+�N�<�vB�$~�D�%���-�xŋ�Q�<QP�A<x/6a겤V�Sh��tAJ�<!��4fS����-�I97G
�<!�j�*�`�ʔ�z�� w
�V�<�ѩM8e4�)ggC�+��$R�<�qLF�7��H�W��6 9^`Ǌ�J�<��ho4��ӨB-
��C��C�<� J�J�)t���,[�b��m "O
�:��ۧ\��a�R�Ö5�Q�"O0UXt�,U@02lO�
��{"O,�9�i��R:=
U ��L(P�"O���I$�u�`L�8���y"O��TC���t�Bk�Y|��"Op�yU�	&LIބ�w��_̱�"O�];�E�E@��̞=��$2U"O(���F�
!�^#���'A� ��"O؈4%�e2@�aŜ[�~�1`"OT4��$A�y2�`i�?u��Uҗ"O"�����{�xD
ԨҹYV�1W"O��%%�<C�P�k��ۓkY����"O֑B�,݆c�f�Æ��d9|�5"O��HA��=f� �[�,R�?-�Ң"O��S!��$�FD i@q%�<�"O>�d� �&� )�@��a(b�R"O(�)&����@��M�=�u�"Ob���DG������L2*����"O���Ҧ8b`AS�6i5�H�%"OR��� %V�
����z~��r�"OD�:�-ӱc�:Drq�ű~l�<�"O�9�'�є A�Q IWNW�Lh "O�Ae� 	*F�i��J7EZE##"O�X����oYt��V�XW��HR"O����-�;�=�%A��PK8�!T"O�@�(V 
 ���؄)����u"Oz�"��ַd*�A��٩?�`3�"O\PD, ��n���$v�J9+"O�Yk�D#Z����E�Z�u����p"O��R1QG���Pp�<3�13"Of�StoS'/W��s�	�9k,P��"O���2mT)�,̐{r��C"O�� )�o �m����v� �"O��ST��Yu�h��I��K�*P`"O�uRF،]�2 a�"�*.�xrF"OIiŬR� a2u�̫eA4(�"O"TۢcIʅJ��>9��t"O"D�s��<��`���:S{0X�"O��j��Cn$��p&E�"O�<� [(F���?ڙ�"O��@���u���C�
�<:@}9�"O��)T+�8������N4����"O��!F]�WE�!�0H^*^�A6"O�؀hZ\�  ����K0�t"O����B +)�5�C�K�z
�p�"O2LA#H�BX�!w�D�pQ`��b"O��,�)�`)S��=):w"O$��T�Z6��[�@��q��S�"O@�+3,�..&�D _�@ϖE9"O��������	��9iB�`�"OF� �G0a 0х	V�4b@"O� A�69��@�pL����"O�0�Uo�oO:%��ƔQ����`"Or,�o;�D�x%O�}�X��"O�0���� [���"@P�D��"OB�:r�_ *�°�G�&KaƉ{�"O� BG k��0CNH�IJ\�xd"O���a���v��A��#1Z�zD"O*�9�.|2�1�Ԍ^�n��"O
J ��.^T7�v��.ܤ!�D�Ff�4�ק΢wn��w�O_�!�dѻ$B\" ll�V��g}!���0X^��ŇX�A_*`)m!�� �Dp.�
YF,��#�]����S"O0,�5���p����6yj��g"O29���ÿ[Q� �� �,qJ�"O��a*�'K�R�2��֗"�P<��"O����/2���Vk�nH�ˢ"O
�`̀/�1ydo� "�ڙ`�"O��ZQh.���)�CϞD�B�X6"O�0jv�D�j�2�!T�_�x�@��"O�$���H+{q]�f�ߔ-��QP"O�,�4�Q���Z�bX#$
XJ"O&L I*�
5�Uˤ�J�`"O��"�,�@)f���&��'<�9h�"O�P�`�v�2���G�c+։�0"O��30��6Il��f�&{~,� "Oƀ
#�ϨW"�3�F�0�"O~)*W� <cS��U�җ�����"O~$���MvlڄΣZ�$�"OB���䈌G�@�U�:{v s�"O(\B��CM�@Q0�,qlXa�&"O����-�[^2m����Ta��"Oz4	� �ą�%�v�a��ߟ:�!�H�
�r�-�\�豂(�/�!�O�Q� lz��9З�G��!��B�ƀ� ��O�(`�$�	�!�V"IW�؈1�N0'������Y 8�!��ҵCD�tY�ǚ6�*��e�M)!���5|�|=T�/iE��X��U{�!���;Q�$ �j�"IL<���Sc!�$ܜf[����+^�c��,1Ł*c!�$J�=�����dvS��3ef��/��B�I�W��y�A��|u#�Ʌ�O� B�	�S�Cӷ|�HQ��/��[�"B�	��iѷE\$3�����M�n`�C�ɣwEnp�g�.ڦ�Z�䆆0�rB�ɎO6��!����@��L]��'�����l؋]h��d�R��:�'ب�{ �I9~Ԧ颃�K]��;�'�Z�	�*�$y	n��M�%�Dq�'�B�+*��Uͺ�Z!��\��'R�YP�K�)'t��6쓚i���q�'��9��hQ7"��:�$-h����'dR���Y�9D�,���V1e:�-�'���!��:��Uh��E0Q<Ĥ��'�>e[ �u��8
��Il�}�'�~�*�L�p�-��c�v
��	�'��@ӇƧ^p��2�n�8l�x|��'0>��䆋5l��`��`�$�	�'ZPɱ�B�/�h�0���SZ�q2�'\�$o��+(�Jv"2����!"ONQ���FUİ2���o�~��"O�i�!���`���䃖�W��h @"O0�H5�W�V@8�J���;y�5ч"O(p��Nӥ9CT�+G�X�n���s�"O��IAeK]�	 �W-뒜��"O6�BUg��p�\!����~�Ku"O��a��\��P��
�s/��)�"O>�8��C](��#i?s4�U#"Ov�"��̷�BE�3.�8��"Oi0���~�iÌ��i�� �"O����/;�<��k͊$����V"O*�jڍ8'|+U�+-�5� "O���e
�/4*���ۤU�~�b7"Or��"ݮ"6�A�/�	�f�`"O�̰��Z�T\�a��ӱrJ�"W"O� Z�qrL�)kG��E��<-t�zu"O&�c� �4"�k��A	W����"O����!V	*����6X��@��"O4�$��$[2�/*�@�"O���B )y�D�P)�9	*�
�'��l:��!���7�X9���':����j2[V������'d0�iq�ܙM��BB��~����'���x�+ǩ@"��
�kͱ� h�'E�x��c�1��Xxek�.|u�l2�'����F�V
{?��ՃD�y���9�'����Ǽw5��%`՘;��xs
�'[T���R&>�LIuI "�l�)�'�HF��/��UgH)�11
�'�$�@�k�3	�l���� x�:	�'Kʄrj�>�Bl@�9v�T�	�'�Ҥ�@��~)bmy�#�w4
��'.���J/[,�Xc��<�����'f�q�$��5::\����	X����'�����^.�ꡲu"V/XNp�'���۱
�m P`�n�}A�!�	�'-^a;������q�l�8t�((��'fz��@�@� ��sba�}�t� 
�'s:����G1(�L&�^P*�'��S-��C����.M%H�
�'��<K�#B"*����<G�e�'-6�Y�Bɰ>d�ɸ&�əm�����'A09�5�D#? ix�+S3hVUZ	�'6��3��6��}�Ħ^0^ע�	�'��tS&��w[vIyčN$]�v���'3�����Z�a���K�����'¾
�f�D���)�G�x��'�(��ɗ �䬣r�0r����'=�yX5H�<kFZe� kF�h�YH�'_L	
��^�Zuɇ�Z>s�p�k�':���B�$�%c��<U�zvA�V�<��L#Q��hv�R>0��l)FO�P�<�_��P���3�t��Āx�<1��Ւ'�uv�O���)V*�i�<����@����A"F�1#�M�f�<!b���#Y���4��`�@hg J�<�׏/���C �� i��J�F�<i��@�E��A�%K؉rH%��dE�<�� ���+�A�1�����	��<��M�+
���#�EE0~�Cd��~�<�������fn-t����s�e�<ᑏ�Q=d*2�ަ>�^Lbզ�f�<�֏�-`�	�jX�5�rT�(�~�<Aऐ�ZoqQ����X5��|�< F�}7�����|� �n�<9 �D�^��d�f�:�l$�э@�<ٖ�1>�"�Y�5eL�#�c�|�<�ыBH�hԁ�S?0^z1�V`K|�<q�l�q<���u���4��0�g!q�<��KZ0o�����Q9-&�|�AE�i�<9�A f��)���g��!���{�<i��*e�� @��)��e�A�@S�<�d���2$`��|ep٩!A�C�<�"�M�R�a�/[)�y��}�<AlF�]�D���n��H!6�Ba�<IA���&XRi�BM
�0q`CW�<I���)hm~����P�"�����bV�<������D�1�k��@�H�`��U�<1�E��8�����4UҀ@i�[�<� �� tG�$�t���5�,�"Oذ�4�]����hǀ��z�^��c"OD$�36x�u�lʴz�d�"O�p��k�ˬ�	��`��ar�"O�l2'J'U�0b$K�>kz�-�"O���!O	b[6e��$��H$9�P"OrX��C�-l��򩍗C��d�"O�$x��Cg��!)�9hdY�"O�8[7�տm"�UB��к+Wx�k�"OؙH��!A���DV4,N:!p2"O��z��f��d��1}'�C�"O�h��KQ�#����Qy�F�x�"Oȵ���Z#C�� �eE%aM�aQ�"Obi�(��&&��e!ע>@ I �"O���S�ď#	^�)��^�^�r�"O����Hdy:T;%"O�dJ�n�/@����6Bϸ@��"OF�����9W��mA��R7@:  �"O�� ��\5JjmBV/G�MV2X��"ON)����?B!M+d-��(�"O��g$�L&�M1��z����"O$Æf��LZ����S1:[[�"O��Q��B�(�H�B�{V� @'"O��
fZ�0m�xx����$N�Y�"O�ё5���<� Q.">KҠI"Or���Îan&���,J��9w"O�Z�M(h����
�3G�i��"O>t�6dD+Ad\� �,h,x�"O�1�!�yJ
�+c���*t���"O���T�D�MbA�#F/"Z,}p�"O��Q�P�V�N�i���3o���"O�y���|t:�w��j�T�"O��ڀ�R��hh���K�t�$��"O�!V(	�4��41I�$_~!��"OB�H"�A�qH�����I�I�TyR"O�mC�S?]�<|V��@�ݰR"O��F�>�h|�KʜT0��"�"O�+�,��l9c�,.60���"O]!%��
!`Ԓ��88%���"OpbֆŒ�b҇OZ&%e"O�i��1����Ć�P�t
f"O�ْ5I�Crr)��(��P8�t %"O��y'�¶b�9p�F�rt�7"O�x0��S�%�\�u#Y��	{�"OV� �z��!D%ՏE�� H`"Ove��n
����xt��a���$"Obi"��luh*Q�Ʃ���"O�uI�&Rk�UP�!�2����"O��5,]�;������̊&�`y�"O�ڢ
I�X��3p�[�˰��6"O(��`�Z�`�L�3_�H�F"Ol�P��5m�b��J1���3"O����ǂ�43Vl ��"�¼�"O�-���!e����΁�w���U"O���*O�+Q3���@�*�"�"O���6C�8��)ʹ]��EXc"O`P�2-^!Q�M��̕xJ�)�V"O��cfB+?���٣X�'��s!"O tJ�$��q�B�6�6ű"Oz<@�/�F��I#Z�5�p)� "O`��Bi�-����w�1?�2��c"O �Zua�_pTari�_�M�F"O�H�֏�r�y ���m͸ؑW"O�Y26U-�$	�H�$iyQ"O� @�pU�� 4	�
� ؐ�"O� @+{m���K��!���#�"O^�P�ʡEO����ށ1Զ�Z�"O��x� �Sm����Y�*�"OHib\�z�y��@1��y�"O��Zg$�48$ۀ&��-����"O�i��g٧��aф��/r�`�"O����ǣ��<�䘟��@q�"OMzӇ��,�ې��$��}ڱ"O�ʲ�E���s��N���{q"OΑK�M�8V�Z sD=NW��Z�"OZ�P���r��4�UA@17dU��"O�<kdjA&�����@��(�^�K�"O2���R*|;r�rq�JϪ0"Oh8S-�Wu�=r7�X�S���2"OL� �a��m�����K:kA�:w"O^���띰W���(��R�
p,Rr"O�uҰ�H	7 �x�C�t����"O�遁�43 |�e�K�>�B�і"O��d��f�0�G���(�"O�ay`igp�@��S0@�̔9�"O,����[%P������.7�:��"O�Ȃ	͈"�x9�ŇS�ӶJU"O�=+�ɏ�Q����W�#��z�"Ol�C�c%,�$ȁ%bޙDP "O��v��U�u@'�53\\�K"O8����Q�y���~E.J�"O�a�&k�=hox�I�FA��4hd"O�4��@�6md��-ے4�����"O���Pb��;8�됶3�r�h"Oh�+��*^��9{e��/$q��!"ODm���2!lb��ő���z!�D��h3$!�*y*%xbAM�,!��3br5�dNJ4xF�!woDL!�d.h�:��SdXu���:`!�C�;������C]�a�e�9V!�DԹm�|��_!G4�����!򤈎|`�l�!��w�Sc�!�O��6Ti �B(��qb䉇_�!�\6u6%� �V�Ɣ�`���!��J�N��y�h[�� �8b!�ҶF�89�MD� �85J�h�-+!��g��iWMI8sj�%�ph�5b!�$��=/`�#��k[
�J$�Ɠ#u!� +��e��I���qKˏ c!�d�M'�����W31:A¦��G�!��P-Aל�-N�;;~ 1'���!�$�)ٸ$Pq��)10@b��,G�!�D�%.���4c�0l��k�!�D٫+{Ѝ+E�F;=��eh
�gi!�d�$�h�W Җ�����'�^�!�dT��h���ȍ{�R$�� ��K�!�d��<F��h��R������8n�!�dA#NB�{"�S�t�8���-H�!�A�!�"���R�`V��[�]�!��ج?+�	I؝@CN]{�J��>�!�D	��d`bíٚ[:޴{C�C,'�!��h�,2��A'uCB)���*PG!�$�~�*�)����\?��
��ܦZ)!���3��H���s�2��+�_�!��L(.�\�HwlR$xa=�1�ȵ �!���]8�C��&�u	k�XW!�D�;��A� H7	�T�q*ZW!�$̈́ZZ�ɳ%Ԕp���&Ɉ�[�!�� t��!gS>k�D�0�	�s�\�˕"OD�A�W�m(F�&V$��Q"O~m�E�/�,ݓ��T?�XA"O��b�H�5O�m"���*rY	�"O�ئ�ɋe�)�#O�%UHp��"OBd�F�� Z��N�G?��y�"O|�����5U"���d�C1)6��"OL)��%�P[l�����"~��Rr"O���M_�m��� ���*j�)i�"O��j�+��p܁raW2(oxu��"O��aQ픣HƂ�`baT=AȨ���"O��	�&r��|(%aΰ	���#"O��kգ'9Ny��e]�K:PI`"O�$QKc���ӡS�ZYA{G�f�<�`n
.X�~l�'�F�L�X[�`�<y���  !㔪�[,�bA[f�<�g�n�����(�58�|�FCBK�<$$*��P�nR�}9� �y2&� �� ��J�h'��*�����y� N�2|��*(�*$���y�oџz��!��Q$]R%��Y�yjڐB9PCi�;�A/1���ȓ��t�t��?`NJx ��r��������@���K��]�AG[<p�ȓNp:)����D-��
��;O�\݄�<^�RGnT5�t��#�.�����6~���*�V @Y�嚦>w֔�ȓx�P���
_0iZ6��� V<��H��<�w�n�\��&��B��Y�ȓ1`��a��]�؈H�aMt��,��I��	�8dŊ�k�`�P��ȓg��: �H�r��m�g�Q�#��A��+v�u1@�52��  ��m\( �ȓ-?R��鎔Z������t�H��F��� 7L�dr���`Y�/(�8�ȓQl`xۆNPۚ��uJ�0����ȓ.:DbPhX�4��
��r���P�F8�ҏ�!���ؔMӄq��|��~�nu�&�h2�(Y&�d��ȓH�~�X$�ՅT����KS�Jx�ȓ�$	 �g߹3�-;'�ӽbr��ȓ]�v���ř�i)D�ӄf�� �0���j๦(�4&�����˱|�
|�ȓ ��E���Ҟ1}:��9lsPp�ȓ6\V���/�����Ǎ!q&�ȓI(ڑ��l�!C�A9$X������TlR5��I���0'])a�����'z����A��8ـ��'�R�-O
pi�'N|�0HĨem||A�'":U��'<��N�0�`�j>�X8�'E����8B�h��r�q��'�t�v$Z<U��f�{�'6lhU�A5*�C.�@LJ�'�M(��1+�u;�L̝{��u�
�'�@\��.V2Xx�ÍK"v����'׈l��Yn�ҽYc8p�P��'�9�W�����y�k�`�tqC�'s�]y��8D�0���T@�\��'�n�z���.(/H�0��B0Q 4\��'W��0���%%,�ó�ڙMJ�A
�'��={P����̤y�ŧ@v�أ�'������]�(�,�¢ŁG�R���'�='�W�n$��I�1֠���'�lLqф�!�����k�`������� b�(�/׸h0�a
��xh�"O�!�Ξ-,�XЂoP�-��<�"O���֒ZP�����QΤ�y�"O�eJ�ʂe%>$Sg�O��M9c�9D�ib ^8k4V�h�T<Q)�k8D�԰��5g��J3Iǻ-UĐ�uL6D�$
�@���H�iH�7�4 �0D�8��=Ǻ-�K�Zu���,D�l��+�<-^�P�b�O�b@�
1,D�[�đ�X��b��0L0p�Ƅ*D�DwJ��Q�4y���7y�,ܱB)D��j�+Y��|;� �hl���ġ&D�\���[f�t�!a�18��]�&N0D�����$@k�$�CiG�@`�(�B$D��Cq+!�P
M�8�]S��$D�`��H�A� �B�R�9;�Ñ-D�(�b@�M4��@����$L*D�L0�$L�P����M��z0���-D���#_
%ʺ���,QD0jA�(D��p h�J쥩C�7�����J$D�0�i�8:����d��T�ԝ���7D�\�Ph�A�r}� �*?��9Q�5D�H8Oƶ�tA��LԐ����e�4D��q$Q�1x ��
ppz��) D�Lcᖅjw�A ��m�b|)�>D��c#O�=c���f�N�3ZfI�/D�̃cZ����&JG x���)*D��wC�F=��q�)U�~�ad�(D��JͼNƀy��j'-�\�2�O'D��i�`O�;�6Q3R�P$)���CM%D���5��-Jo�M�A�$O�mI�!D�hX��"������#|Q����, D����m��7_l� U���z5Ѝ�c�?D�4Z�`ݮG�U���׷'�LP31D�<k5���Rҝ����x�.Mq�.-D����A	-,���D��>2_�ǀ%D�d�ԧA�!Cj�r.ԤD���#D�(�bA�Xt@,S�pZ��@K?D��2��x�y�6]
|j�#=D�4
U���4�)
B0��9sC�5D��KA�E�6U ΄8=)��IQF?D��IToZ��QD%�p�-{PB?D���a��=�t����@P:|�z�!D�D�T���,�^E۴-��`�ǈ?D�İg���5��5[@
ܞs�"!D�D&�[?`�*Y ���tV6���>D���e�Pl��,��i��m�B8�4*OL
�	�f����÷dL(��"O*�뱈E�j-p�%C1%
,��"OF8A��B�t�L���$Z�/�p�Y�"Oּ��ݔ���3f�C�f)n�"O�I�fh�-�䅡�b��R(�l[&"O��Y�S+{�K��l$x��!"Od-X��^�0J�-d�т>>�r�"O`�x�#��q��
g�:OHh ������G�Z�>��W�#O�!�$�.m��m@�`�(#L$�`L��!�D�/BZ��G�P"1 a��-�!�䆷"��4W�!!�}��^�#�!�DFl����K�$[�Q06��%-�!�d�5J��D#=�Լ�K��}!�����\� �.���{��^�]!��2p�H�ݻ#�p�uIV�9�!�D/�jx)��L5i�02�H6F�!�� ��)��TEZR�Ŕ����"O�}S⚦��=9���|u>y҂"O���*�BR���*dl�Z�"O:���l�6g�� ^�T�1��"OH���b2�&��#O�b5J!"O�5�r�ԪJ��ɂ�M ��,P1�"O�A�҇J�7X���*[�0��*6"O�8��VU�2H�A�8$��B�"O�8�ӥ�����͈�
|J��f"O��x�/ۈC���P�M=)tH�"O2�q��	
PvL�s��vrp���"O��B��[+�2�BD�I�s��E�B"O�Aq�ܶE�R}0���)t&��{�"O���ҍ&7X\�0�#I�S7"O�L�րW>k�L$��� L�X��"O~u�P���I9��E5^1��0"O�����C�$��B��:V�eRA"O��Ӫ�+ �xh&.]2z�R�"O~�[� ـP�R1S���T"O�-���M�s-X��l�C�LH �"O\=Kv�[�0��	�B�a�`���"OĨB�`��_jT� 
K�J��uð"O*=H�đ1��T��I� ��A��"O�!����JB�S׈�'J���"O�����=u�� Ŝ-B�L(�u"O�\�&+�l�$�H�$��m8"O�h n�X�z#�g���$"O.�3�K�%g�e�Ҙ9���ZC"O�@�M�v6�-�1@��^x�5"O0��㕶\[``R��"Wu��"E"O����8���"@(E>����"O*�uk���J�BC�QB ���"O�a�Cʒ-9�����ܩ)7<Y3�"O& ��,WδTY��=��0�*O�2	�@F>�:w��=Z�F��
�'�x���� �t)�]�V�D�Yt<$�	�'���SAݸo��Ta! ܗ`��r	�'�������$����a�8W�}Q�'��j�[�g� �� E�TFA��'�H:�a��YR��Ɨ��$��'ń����G�3�l���ΖQ��'m$�C�EݓB-�Q���&>z̓�')��1�o�8�(�����h3�'+����.e���h���`�i�'�܉k�	�W�HdsU*�])��r	�'����b�J%Sd.u���@^�� 	�'��e���y~�2Dm�!Q�l��'��ّ�VX�器 ��q�'�asHF~Yt��+瞀��'��I1&��1�,��A��s��H��'=̱[F�3
%+3aI:hS%8�'�&�Ƒ.Qش�;3��]����'�H94I�C�(%��G�R�����'���ӆV/P 0a�v�]�=� s�'Y葰�a�%_J�#ɸ}yzD�'lʴ*�� @�`�4��(`Dy��'Gp=#�!�-����6v�)�'˚�R�
��<@x��nݵ[rz��'B4����.8��GB�#Ħ$��'7>XЗDJ
�Fh*!J$&�
!��'%Z�{i��~�X6bƬ��]#�'R�iY�ȃ�F6�e"���OJi�
�'�XTe2,�V$�b�#N���'v\{Y�d�,Bhӷ���
��� e9��&I��鱵☡y�n���"O��K�Y��-��A�9 �r���"OB�"�^���ST���G�>��"O
����-R�
����}aRi��"O�A���F�:����P?-:"$��"Op�@�"alч��K2���"O��Bqj ;'qr7���fC��"O��R7�`�'o�?=R�s"O�D��'2V�@��c(a"�u�"O�UiA��&�z���l�:0Pg"O0�(J"�A �ňM�1��"O�a�����w�`ȑ��)���"O�1jA$P�	�h �2*�=[�ށ��"O���J�:�$��I�1怩�6"O��:�a<e�ZQz��A����"O�#���&/A� �-؋]SLy(�"O�pxcB�-LP�0�i�"T��P��"Oqdۯ@���'�Ҋ�^�Zq"O@Q��F*
}���1Ps���r"O����C�Z��e��S�Qm� G"O4y��7Kd,k&�P�ed��*�"O�H ��H��a3a#QMl�(��"O~}C`̓�F�+�3��-PA"OpHBDЊ<�0%�N\J��|��"O��U��!K8�采K�[�� �"O@,�Ԧ�/ �K�&�0q�$Y3"O*�y��\?�Ե�E�0b�R��"O&mB�Ȱ�b��gB�i��g"O��ږ�2cԥ*e���-���"O�i��ʒ(��}��m�.Z+JX"O��k�����œf��W9lE�t"O�Y�R�4L�4)�RT�k�h�r"Ol`�V��	��/�IVp����^��y��?k}��[�jQ�E%�0�5���yB!�)F~�0�c#H�đbP<�y2ܕw� 	���xl��&W�y��L�'�`���]8\�\N��
�'�� ͜�*�ƝC�Ȟ��<��
�'̖,���\�v�&� _�3
�'�sw+��@h��j��O�s�B��	�'�\�RI�F�402я�qKpY��'��Ii5"݂?�d����T�
0��'^�Qp��=-�2a�G]�F�H��'ތR5%h{>�К���=T}"�'O�Iz���tsl��,McP���' �wͅ9?Δʇ��f|X�y
�' � ���+F ���)V�X�	�'A&��j�	>��(@�R$K�l	�'��AX���.ML���/��tK44��'��-���,�Ԋ��X�Z�<m��'(M� X�3���,U����'�n�rP��]yt%H��v.B�'|�ͻ'�i�b�L	i��Is�'�������R �@�q�[Tk\A�
�'>����FȊY�"2��]	#*���
�',�4B&��%�ԄJ��� ��[�<�KJ�ݚ���7<I� $��W�<�L	�c0Ҡ� �Ԝ3��L�aA�O�<I��U?Ԛ��`��J�6tZ�"�N�<y$�� Jb�q�P�W�t�%��F�<�c����ib%��^d����@�<���5��AZ��ȗ_�B�b�)�u�<�ݸ��xD K�01�0@��q�<��Ə�"��x���T�>/�T�S͖o�<� \4�$����@S�UN���e"O0����֫b��sO�-?Heh�"O>h)�o�:d��� �?o�z���"O:1�e!��^��w*,r�H)�"OMj��D��UC!j�$���B�"O�(�DN+`lr5��űVv�K3"O
d����ִ����Q�`8n��A"O,���2v��j��?(*���"O�� �̑�� �s��X!���'"OZ��TL�~0�QY���#J�^@�"O8�%�  ���ؠ�E<��L	�"ODT���Ã4�r-���\ �L{�"Onc1�2��X E�ٺ�d�:U"O��ƆS2Y�Z��v%Y��� "OR|�T$	^�����.J7JY�"O�����]��7��2t�s�"O�m��>	V5��+�G<ʰ��"O ��2�[!O@�4*�V̹7"OV���$�;,U��!IR���5"O�;���Dv�  �]�E�BHX""O4|@a���� �u��,�B��!"O$�{�!�6)
萒\1n��+5"O�	�w�
)��,Â#���B�1�"Ob�3��C�<�zĘU��+��<j�"O�DRrf��l�|!T�L6�P!Y�"O�]2��[-*��=-M�3u�$�"O~�YP�оQD���\:{U�dc6"O��E�Y�J�P�E�H�Hp��"O<|pa�ݯD6`jV!��^�"O�5
6��Z#���F�uߔ��"OY����H	��� M�)��d�U"O���E� 5��x �;7�biq!"O�(�bM�%���ɤ�	p�dK"O��c@)ڋ0<~�xBo؃�^�&"O�|1�G �����P��,�"O�	�lNxlTp�2a��O�H(A`"ODQZ�
���(��l����"O���!���CF� "�|Qj�"OA2U	��&DT���~1�[�"O�������((�fH,d�
c"O���%J�*%�Dt�q%�I4�I�G"O�*�݅Ri��S�\f<�8Pg"Or,cɔ�0���z�(�>b�7"O�EÅ$�(%��r��˙i<x��""OD�Sgo�?:N����	$8����"Oliz�cT�X'.P��B�B��#"O2��j:�p�`�)q�:���"O$�KedX�G�	�"pqJa1�"Ore��_��P3 ��f��"O����T4���!Kڮi&�Ʉ�q��E��ܽp>��A�KJ��ԅ�X�h=	6MB:T:ıkC� 
�,��a��Zg� t������;k�ȅȓ+Xd��ꈩt͚�!E#D��ȓL��Qã)X�r^t�� �G�_������\�0�E$\<b �g��e���9Ӑ��kN
�P�$\R�̈́ȓy�I�BԲdq
�9'���i��C�I9i��[PfǫH�\2$lN3i�hC�	D��1�q(p����z �C�	S����r��;ap3c�I�?�C�ɏs|��� ��3M  [քɛ~8�C�ɢOdf�(#i�'E<�ѫ	�<ۤC�I�nP���hDt�T�(W�0C�)� Di c5.Z�k5��v	�7"O��Kc�ճbt��!T�.�|�#�"O2e�R	)aN� ���nWD(b�"Oh�z�+(~`@��`��3.-��C�"O&�A�OƳH���2�������"O�h��A0'�(�j"��ml�#"OڤH�L�i���!�	�(��q"O��[����F\xh9�BǟM����"O�A"�IJn��wE!{\��2"O~�q%I�����$J&j])�"O�4�v'�����!�0�ޝ��"O�L�/�2x���B�:��p�U"O��DO]�	��88Cf�M�V|�"O��Ǆ_�J�)��ʐ)���B�"O�i�G�K$C��� n�+;�X!�"O�!��
�1\
��nY;F��5"O�M��S
V�(�;���p]�0"Ox�Q��·\l��r��z�"O�(�Ղ�P_��G��R�xG"OF`q�"��榙c$E��u
:99g"O����ߓv�r5��m�j�d �"O�����Y�Ap�c�.*e�z!"O0�Q���N�r���:uF�@�E"O��{ׂX�_�<���,��iB.ա�"OBy07�JR��u��MEpP����"OX�CpbC�/��a���Ԅ:1L`�"Od��Ҧ=4}L$ApM��8�"9P�"O�q	�g�X�jŹ��H�$D`���"O��S��KT~�y&%���D`1LO2"<y����d��%��mʹd�jp�`-D��!��`k�H0�e"""<��(&D�@w��&U�}o�G��˰*'4��r%�w�6A� N��%�-hb��L�<�p.� %t��{�Y8� t�qn�o��0�?��-
�'�ӅHY�y�2}�FPA�<�I�6.I.��`	�k�<T��cUs?a�'��$�<��OP��|��%�vQ�i0&�f�����s�<)�"@�
��S��V�W������l��M3�1�����b�)/p��b-U��j��ȓ�8�#���U^@�p7J=�ByΓ��?�FH�C8�AA��2�\�ّ�aX�4�O�A���	���s�h��]L���"O
 ��(��H,Y�d��Cĵ
g"Oj�#�N�MYE%�Bx@�"O���C�X���*1���31d�i��'�ў"~�DOתҮ��B�	�E8=X�BO��y��(&;f�!�ab�u0�����~R��`����%M�[Z�@�e���N �Cw�W�����F',o��q�f�.A��p$�A&I!��/2� ���C5[��p����( �d�[؟��e�ɍ���3�G�
���f+>D�<j��)K�p���ߒ5#d�d��OT�=E��_]`&�A뙃�^ܒsO�_�!���P qK��/UzYj�^ !�N [W��W�,\��C�+u��G��ħ�~"��x�vE�j܍"� ߂�yb�V&f�ҨB1���]�.�������Oldz��i�	�KJ�.�B-R`��~��	@	�'dt<���+k�aX-x~��R O����؎�B0�dZ�=Ȭ��p�I��~B�Z�'e������V�cBZ�@*LUT�]'����	�IH�aU,�u'r���� G��든y�/M����|"փUe��q*dB�+f�`����?X��C䉠����7�Y�I�ZSR���	�nO0�8�47j��W��u� ��3���rp��B�*Κ(rg�'-���im u� �煊W�qX�'�b��&��G�bm�߸�I��W��H�ᓰH"8@ˢ$�
2 cP�ēl� c�yb�'�R�;&-U�xP֍��`�Y��j�{r�'�v�I�Q�kS����[%=����'x01�U�
��;�,�8XN��'I��&�=<�5J�	�7
�VP��/רڰ>�O��r!��v ���M�6�zD�5D��
�'�!�L}���J7Z��Hg�5}�)�S	O�-����/u���+���R�C��?6p ��˜8�~�P���9Iz#?���S<��&#�i�����A7aNC��2Y��#4 �7Ά �FE�9��B1��<E��aX�%�x�$Ϛ�89���
�y�]�%�lԑF�ϰ��ap� ����'�a{��H"p*�r! �⠻�$_��y���+C��0e� 4/
� �	�y��R+_�y�/6L��[�ᙗ�yr�տG|(Q(4��-yJ�iA���yR�L�C��j�B��&ًC�ɇ�y"b�J�4�P�4"O2x@��8�y2� �&�H����0)�!�]��ē�hO���8C�
τo��7@�!*���B"ON��E�*Cr���	�' �%�"O�LӲ
��3�n%J�9'	t�SOn����(��$�Q�#d��3��E� 7!�$�JdV`JCO˥���#,<0��r�*"<�O��`bP	(P@p&�Ĥ`��Ls�'7@���3�FH�R�W.W�%������.�)�q�h�ѧn�	O�:-
r�S�L�"���'����r�7lHj�`�n�G�:@2�'��@+�c_<Rjd�#�fV�:*pz�4�hO?73���i��C�w\>�X`�"�!�nͤ��/�(i
M�g#K��Ɍ�0?i��7rwhQ ��O�DL9��eSi8� 2���S�Y�ǩ^(0�����2D��Jc�7��pk�/W�sE�(��"ړy�^"J�D��` H� ^.�\�{�B�f�<���2I��uJ�FC��8�M]|�<ɐc��	��dƢd;��j&_�<���o�����H�4�Ej@��B�'p�?	��KW�t^�}�HѴG��
c*%D�A��P3ͮŰ�����h�A6��<�e��c����b	N1M-�����}�<1d>sڠ��7ᜑE�h1e*T�����X\0�"���t�P-�>х�(�S�O�f�zhD
&��ꆀ�	+�!��'��=cbO��2$�v��?�^�Ѝy28lO��$/�7�t1Ȕ,Q�/�<�r"O�T�& �3G�HD�ĭ�>�ؗ��(OF�=�O��P����"X�&	սy��@��'Ox��)��2�T��U
־p�J����)��<�ghS�:d�������f�$�EW؞x�=qp�)3��bte�1vȰm��
�R�<їd��3
�*r{z��l�I؞�'C��GiT�$Mq�\`���!I~���>?�Z`���EZ� 87'� �x�'w�=�~�e�W�yõ!\�xt�vf}؞��=���.�|m�/Q�d���	@x�<�F��+�J���4!���(OܓsB66M8�)��S6�p�5cԷvaZѺ2�\�/�!�$� �Q%i.$T��{U��<I4�(�d�.
w$�\�d����$C�e�Ųdʚ�V�`�g�Q�:�!�� ���ID��R�F4}"��G�V?p�!�Tڴ���j(h����
�ax��	�3�Ĥ[��56����J�
�'��Aa!=X%��Méx�$!�'kB��'dY�<�e`�D/~=v���'fd�0+�Zƴ��,��n���z�'/���1�)|�L}C�DH�|�ii	��'���C5킍�ƛ4K����2!�!�6<(�-"�"=��4�b��vʑ��r����j�����#ʁT�n=ȑB!\&�O���$�4H�"�*BLv�z��!�#k!�$�{ ���ś�"���� a?!򄝺u6d�cv�:�T�rOYf:�ɰ:.1OTGzZwU�a b�G�QҊ���H�oN.M��'r�	����UC
�"J�v���')���c։MmF��p����d��'#��(�n�{�Tl+G%�,i��` �O�ܛ	�O�8H�-� $���A�X3`�x����@yB!
"j�F�i1�H�����9�y���#1`����U�Վ���'��hO4���N"~��B��% ����aB!�$�%V���&�R��E+u��k�!�dS�E2�g+I��2���OW�5Q!�Dʞ_$�H1�N� ��!��V9",!�[�sޔ
Ĭ�.OX�Xp�^��!�ğD��tj�"Q��háǻZ!�Ĉ�]u0����x�z�4@ L铃hO�\@��l�4B��%H��\�>��YW"O21
1(���H�s�յ9������.lO�	)����:�4(2��I�hJU"O")0���0������7X�x�"O��`��;-��C@�bҸYQ�"Om��A:��
�
�`���"One�����,���;'%���'R��0
�V��pL��'!��ǣ@K%�iB�����4��'�h�@թɚ>�2�ƦI0v�N��'m!����9�HP��*��`��H�'�H�	2i�2D���U��Px��'r�5AF�V���x�6��)�j�'~ ����^���#�d��
�'XJI�P�&oҚ�1��%:La��'��u�1�'6�necp��>p����''bP���@*8�
y���&i���'�� T���?=jI���8����'j����K((��DP��n xj�'��%2��J�% �d��6?���
�'xt!v���~����]*%ь,�
�'B��9��ӝ3gh�c��A7Ӭlx�'�.��is���q�*�g-���yR�T.�`1�䂝98��׬ε�y���b[VX��뒟C���B���y���&Ȭ��:[N)��E��y(P���K�g�8���6IG
�y�ɞ=Iu\iUcD��i�P�ن�y®�`�>����%;u�L"�N��y�^<���H$5������y��p�8��rn�-�z���◡�y�$�7z�aӢ��s��`�b���yRT�"� ��#��lQ.}V ��y2.����a���� 2��������y�,ъ�P�r5�@� �Z̢�ǁ��yb�C0Y��I
uȖ{l:9!���y�&��{����Ď��cН1�)��y
� "śDF�E�,L��e>�]"Oy�g��� ���%����		�"O���w(5D0��	4�����
�"O0�Yd��5qs�,����az�"O2�Qu�q��42�	c��P�"O�<��	��p�AÐn�
]�A"O��;`׫5n:��TA�&��	�"O�����Ȱ f�H��3r����"ODH��'´~ͬ��'��6.\n�s�"Ǫ0�سr#�hFJ��0Fz��E"O�R�cZ�{�
��R�ZS����"O����ԥW���	��H��yc3"O��������C�'T*z	#�"O���F�-Ɣ��p�8��9��"O�H��`��] �B �hy�(+�"O���M�=���1�S%wr~��"Ox�H�,+J N=��C��xq� ��"O0��6M�tǾ��QbK�UT<�"O�a�(k41K�Ô�fN-A�"O�`��v��)��"��yd�I{4"O��)��V��<�paE�;�īV"O�af@���Pu(c!#@��"O�l��ǰ0,�Z4�N�j"ODa%EʛP��Y���9�p"O:	�1 ̠d�4 ca�!��=��"O��M�@Bj[��?q") 1"O��R�R_���s!���p��"OZxzS�U$p�,��E�tL�IW"O�@�B�Q+��K�D�;srx�"O�(P�g�h�@��́�<_�$��"O�)��d��]暘r��!�Z��Q�'�Q� {�!�$iuR��(�<P����h<QV��FHt��sb�"f��".�w�<�� ��Zو]��BF�a��Ap��k�<�tÙ=�ƥY���
e%��Ӓ��k�<9¢�%BP�&ڽ,v	жe�<� #�4+H"`���.�c�<i�H  B�ܱVfn1��e�^�'ay��Z�qO<�v/D/(H�B
?�y�G�dK��K���\<�	js����(O.�Iky��G{�]�:��6,�BX��6-�$g��C�	�J>��JC&�=9
���A�k:�C�*ii�q���S��	�����UB�C�"� 8�P,T�Wm��8���HȖC�	�Sf�(B&P+u��9h��؝npv#>�{��~�g# ���`%�]��J����h�<yBj[g����z0F�zbA�<���R��d@'�Q�C�d�y��2>b�B�I3��h2���.�J4Ƃ�$��������O�m �H�1q � �MМ��	��"OV��w� �B�L�WG	�%��a�u"O0�p���"v!(0�b�	 �<�R�ixўb?�'֖� G��
��@��� e�����'�5���F��Q�����Zߒ���O���$��f��d�a���S�:���)�	!��ǆN�4���_�v(@聄6�!�ć�@�T���I�<������<%!�d��>o*tx��;/|�q��[�9!��w�beI��	i���#h!�D��\ij����14�В R�_	!�$X�� #�)�&��/ʨ^�Q��E�����a_
(j�n�=vy4U�f���y�,S��.xz a��h�J �&�y��¶�y�F^���|�!N��Px�� ��X&�"`p�9��	i2j�G"OJH#e�	<��@�3�Նw.J����'��'E|��1��M�D�sb��<��}��'�^�[F'�?B��ƚ8p��N<�����\�Eà�Ki|� Z�d��ax��O�b�4H�W��	��a@f�˷��4\O�%�7��GQ:X��FՖ6��5������s�O(�]R`�
&"z���G�r�R�'oPӕ��l��+J{W����O���1��D���hȕ怆Py����Ř�y�洅ȓqbhX�M��S�0���G2KhL`�ȓ3wB��ea��I �3g�1"��h�ȓ�`�ȐH��r��f�0d�J4��^�\�@"_�(�~�(Q�^�8�$��ȓ68F��� 1xHU��%D����9�Lʴ�G.5�؝�) ,T�l��	9���d�g"i����qE&�SJ�Y����'p%�$� (�R�r�Y�vPc"O$x��٥QL����Y!	r܄X��'��'-�ْ%��*����4����I<.O��	@�O����K�sw�H��(8T��{��_���'@>�D(�Ŋ��A��%��w�,PmZD�����`��7�h�馀U;o�*��T�����<Q��.�I3f�N�*�(�?��UXT��Mr�B�	���)ZQLWt�R�Jw"�;VA�O�=�O�f�'�l��ih�R�퐬�E 
�'�~��Bmޫ4���"�*	��@�y�"76��A��w�1O�� I���`V�
� �b���B�ɝC�nT��=d� �#kɷOC� ��'ў�}*P��\���c̓�j���"rO�hO���I�'��K`��@���a&a��[ѼU��yR�'<��r�*|^Ab�(��aI<9�'
�'�Q>�a���l��"�O@�Z���J2 7D�h��#J!��z��\�I��8˂-u�$�'�B[��g̓#tX)&T>4h,I�rA���P͇�g\�IS��`O���q!�r�FX���
��&�F(N��E�A��}��IP~���. �J�� ��L�>	X���yb�P������4C���s�N��y� �ONmz��:ɫiاh��X�ׁ�|��Pr�x��*�L���HU2�+s����� �O�T7-�4��9#C�4rY(I�A��~�����'�b8���B �;���[m�% �'�TD;gB2Ys�m��+U���Ó�hOdh��miQ����6�P��	#�'2a{b�b��r�L\q�LT�jН�?�'����iEfq4I���.J�"�'�n��E�s��}���A��bI���*�=�
����a��[�/�	���,��x�/]���x[D�؂J<p�ȓby�a�4i�=�J��$��|��t�V(kaA�X�� ��*L�QsFU�ȓ-ܰ��vh]4`.��A��Ip�9��D)
�b��,�Dڠ��Qf}����(KQ��K�6��\� W�H�ȓ	�l��"��/T`M�JP�MϚu��1��+�ǜ�v�)Q�kH�xnF9�O�p�N
�#�&acCéFz��Y�����F��J�O`dq���)/  
�״�y�&ߌ_oZ$���ݒ'w Y�"��hOt�	n�O���ˇ�D�D�(5��5����	�'|2� ?8�T@�%�((Xh��'��)��0n��!�#�(Hl�!bL<�,C�ɍ:Z ܓ�ĹG�>HR���9�C�)� �Q�&{���fNНAJ�K�'�qO��@�F�J/�E/c�VeR��54� 8�� �FOz�)G@8G�����"D�I��{L�u�cş)@�d��f� D���LKt�V���Aނ&Drl �1��hO��?]�T
Dm�8��a�Wˊ0�C�r:��� A,~ؠ@��1]6C�ɦ: qq��qjq�4K�,'�B��$9�4:AZ,UG\� �@y���u؟��
@���A����/Y0��0�O^O�ehB�Ě�� �JɐS�|)R0"O��е�C~�)ӧhE"��
A"O�Q�ĭ��P���[4�S�wLuZ�"OVU˓��29���2��4�P0�Ac�Q�������e�||4�/���XQ E$��xbb��L-0jB�����k=&qFp�T�O@��DZ�N_�P��Րy��Zv��'(!�$ψ:�ԜY)�h��!����!�d��N���:'8���ҥB:�!������P7Bx��i�+��i!�Ā;p��1�NV7IeB|�1�A*!�O�^��Qr��&xF�L��L=S�!�A�W^��nN/?p��צ!��P�t�"q�I�h5��3u�
1d�!�d�N���Z).�(�+LS�!�D�*�^�s��
b")B��-y!��-RE�ԯ��B��R�S�m!��I�J�\`�,�!؆i��G�=k�Q�	]<��J$d�X�����BPN-0R�Uwx��n{ܓs��(���X�5�p&قg��y�ȓ�ְ��Oc̰l�Ձ5�Y��k�rգ����8պ�ˀ��2=P�@��a@��WȈfQ������/b%�y�ȓ��83��ڠj�8Tz&�(�r�����m��T\PG��U5�u�4f5D��"�!.L%��%��b�|��2D� 	®��2���-V+p�UF,D��+�N�	1���Ӓ�ӓN�S�+D����I�2,����&e�i�5J+D���FCw��(qu+�+*LP�C+D��2JP #��(�j�=��E�q*D���&�Y"X�quؐ-��5�/)D����ޏ*�-auF��Uvu���%D�p��癣y��9���F�[�X� D���c!�V�r�œ}H`��?D�r��8C��S�U*xᶄ�U�:D����Z
�n�A� N�Ӗ�8D�Ȱg ��B�C�Q&������6D�h�)�91�*��0 Q�@��Y��@6D�����W3OV(��h�8r�vt��!5D��
��I1D٢��%��i���r`5D��W��C�P����S�2��0!3D�A���q�"X��z�Rp�/D�0x0,�;5V��I�왉9�"��u�,D� !o�8)H��B�	V�����m/D�HXu��2���k`O�zZ�г��+D���H��8X�bb21)|��*D����ѪR�8� 2M�&j�,�bA�&D�"Td#㰸�K�l��Х�)D�������1��]h`#ge�k��#D��3�Q�+�>�Ke�L���0�"D���q&GJ0�K��VGr���>D��9��K�:9�Α`�\	�W�=D��FM��WRE�$�=z��:D�� X�Ò�֧?H�<BcՔxUX*2"O����W�CWxT�\����"O�����M\X��暎g�+��~�ҔQ�z��V�%Z�l�fJǜ�hO:0I�A�}%�B����"O��2 ,�9��-�u�ÏcsF���"O �i5f�'E0 ��o��Oz�e�"O��{�e���ꖮ�Ts��0"O2i�խڽk}Lq����H�"O*Y@�EG�p�I���\��ͱ�"Ob9�6nԳR��lAdKh��"On�C�B�I�@��k�3v>�?O�̈����0;qǳ<E�D�B:0����W�(8�D���y2 ��S��b.ݠ0��j�E�.�<�I *��#k�!'_��������mɡ$<P�x2OѓS𞸲f#�OL�kª��i�y{b�E0��l����>E\D���1v�R��M6�0?���*����ТԢ]|�	sT�	M�'��4��;oP<���!E�G����X>E�|�|�j��R��*D�<� �Y�*�* �$���M.P��b�I#��<E��'P9U��620	аKF����	�'Zi��۽m�x3��G$�by��4"�q����ӂV%`"�J��C����M����8E��'P�� �l����9t���ՠM<!c�'y����ݾ
���p*������{���O�)��<�C��>���`�MS�}�*��%X}�<	��>�D��޴i�4�W����'��}�_w���EyZw7>cs+Ft2���BӮv�j�'�(�+1O�=O�Ŋ�-X�����¼�p���)�'h*�3 -Y8/�j���.�B��ɗ��'j 3��L�s�f8jbɜ��v�L<i��2|O&0�(7u��#���-�l�x�2�S��jLğ8Pl�o�XȘ��G�_ ��yG+D�P*��R� ��0���D�I(�):g�(�7���}RE�N�=�J,9�nC�`�-���@�<q�#��"\���^�xĪq&�t}R��E��H����F�0ajjh���ܰi[uY�"OJ�)�oK�7� ��Ơ��Zb�Ku�x���{�������	�� �!
�K��U���(�OY�D2ؠ�T?�h�0��5����9~���JJ�sf$��(L�LD~"�_�O���B��Ω=�r�a�R�I0���',Ε�0���P
֖u�@�®OԌ����Ӎ'���3g��e���M�{�!�䜢L�F1���*Ԕ����K�Jۉ'V�-��ɼ}FU��S�C��\�ug�%/9�c���F��s�Q>��LmD)3�h!x`� �?(:�1�ȓAH@y�nKz=6A��$��Z�X1t!�F��'�H�;Rc>�i�*)
37貸��(^�8��b*D���w'$\WV��P�.t�tH��D�|r�]�%��1Oq�O��Fx+G�_q:ahΑ�0�H��3�ϻ�0=��_g��������|��T�B1BEH�/��2�� ���@���`����xT��iN`�0�� 扏Lg��Pr�A�	���Ӯ��}[Qkќ&�䍛5J�S�.B��1\��A����,7�� �c��"X�-��Hمi� @�@;���Og,3/:��ek��<ݎ�[b���y�H_+�vDqf�)Bv��QTX����P�Fb!���=!��d���*��W�&Ig��{0㞀{�azҀ�7����@}?���G�h�`Npŀ丣E�ay��'<�`*���4P"�5q`��Aq�Q�yrDϬBv�MÓMf��m���5d�44ꦍ�D�8��RHN�!�$^�C��̳C(�Y���1��z��4��|��Q�4���|�'æ@�0NT�lkZ��lH��,+�'��h��M�I�t�B��s����۴M4F�9� )�O�q��?7�u�&�:�b�	�"O�I:��T�LsL���D/R����g�'k��z�? �I��
��P|�bX8'���1"O�d����,6�+�D!�p�bq�	�m�E��f�'i�Eɑ6�0ie���n�,8��Kg11��P�B-�[��	:�:��IB� ����Tj�S�OL���Ĵ%�,�ckL2n�k�"OPT �E�{��I��`��Za�&Z�tG���xn$K��'���Щ�W��B�(
�f�h�g�<�
Y��vE��+H0t�0���P:<�ڴ(7$�d���.[>N	( �y��:¨3ړO�j�tKPb?�wB6fPՂ�Lc��{AL$D��t����hst�L:�2L"5��O��ѱ��5AM�0�K��?�3�oP9+�^p9��ބbJ��"�g� O��į����I��	*g{"<i�g�)�%��j�ʓd�J�f�pa���Y�
J��i*?k����S"
�<�����4b�ҵ�`D�ux����66)�\����/l�I�5��&��d�S�3h����:
���R���osƤs�=�S�3�IkWDF{��	d#W�W�8\���U�}�m���ɠ���I��ǯV��y���1�tȅ�hFR	Q&�ѻU�v�d� <�L��F�'�u)�D��)�SH�;jCZI6�:��Dn�M�t�M-���`���D��|���O�|� �pR�c$̏&8�"|�����QC�ޅC��ݘ��ի�X�C�6~�ep�]T�B�,AM`�߆E��Ɉ��ܴ@(��(eNߑw*��E�4j��|1�b��?q�⋠TNU�&��A-��H��^�t"�4����?�;p��m�����,���3	F63���?Oly���Z�:�nx#ώQ�L>�G��8��	c��48H�'�J2M_|�2PGd;�cQC~��8�4E�.r~(�I�20@��.�b1�c�����Xf��	�����>�"!�C�f�X��D
��� ���&˓Q^���c�E�LN�1��B)O'�\He�K=�?٤��\ б���RT�����čHC�	�EB�O�t̻�Y���)$6�f��Z�м�'Jf r�-�D�8�Q���6�Hx�#$
�'��I��j�h��)&��v��P�����\�ц� f�<9�q�iH���A�h��M#`�J= ���Px��Y�(�7a��'k>��"�̠b�
����J"��fC��~�;2xL�ãӡF�ű���1���c���}�h��=|
�񦔕�������q�"�F���%�Q㪘�*ؔ}ITAP#[\�IB���D������2mN=Ӧ��A�-H�d��������U&�@�_6Kt"<a��	�'����O����$�*A߲,�D��UΖXӆ��#")�'����ئ�(ઐ�)�(%�U�T0#ܤy+��m�O�!6�T[D�@4s� ��>�� &m�a& #ҧ�A�c��M�j\+�,Ôe+XM�S-��\��6��h`�M��ĩLs�����O�Ѩf晆(�1����q��&,��Pp���8qE����)���'D����i}��
��K,?�f!ܹ!�LI�>�*m�%煥_�U��!O>J����ҧ�yb�P�~�����_��3� ���X� �C�/#y`}��[��1�R����S��X%��jƒ��G�z�P �uLX�<��Rp�@d�4�af�%����o
��p?a�оi�d��D�L�F�n\?U���v�A���I�|���W-����i�>�;FWLm�E��'6T����Y�L]��&6��15�_�j,v"E(ӒT�Fo�84��ȓ�mD.@� uB�*�<�/N6�
�&?�#�A�DrrI�ҋ(4t$-"7i:lO~�9%O�C�(Y;�R���82	K�Uۤ�y�V�����O�A�W�D2�A	ÓMʜE�g#��W�X�5�S�>R��>�DFO�".KFe?��O (85KvEȌ{��3B�Gc��z��-
�İ�'^*\��o�)b�z�AJ��2�[��C�]�����>9��K�(���a��Y��i�ِǬ֦>�ΐ��
A���)D�Ѐ�F|LbP���:mr {P�j�|�б �L�=��-}�Á���+���D&�d!���������X ��=a`��6q"�'Q��S�*Z�x�*,��֋ .(��O�A`�O��R@
�al �N;)\�,SL�}�^�Gx��Y{��D�=ɇ�?g`8=�ի�;>Є!��I��f<���_�>CቋY�TI`�KW�� UP6��WA�">aq˚(�h��Wb4��a�e�>!�t�&�ͪV{~B�ɼ���� 
�&K��S�>0�JT�sL�N��x�axD��'�0}���؎�8����1':�q�⒜�џ��4�Z*U��|Z�.L�s��5�g�FC �(�S`�N���jq(',OybG�:oO��CB�0:x̒�'wFZ��֤	�=#j�3�Ǭ	}a��"-o�\hSև��~� PE�41/��$H6��Ċ�I�}2]�!�B/Gl��p��-j(� �'�ӷ�8�B�&(��A�$�k4@��X-Q@�յt�����	��$���*;qvt�����=���M
&}Je�3V���Za���J�Ę^X�E��#Q<��ċ1�I#S,��d���VI��5g[�45&?!I�F�E� cr�MR1(Y1��=D����[.Cn����u�|��{@��DA��-BȩW*�{n��?�*O� T���+������!���6X3VOx��n͏>���Yd`(�$�x�؛d��̐��Gn�R�	�37��E���&{�d��W���e%&�I�Ś���<�'�A1`)>��e�.�q�7*N�Rݒ���B�7����(@:�� 9��'�RH�+ˎn?<I�"�2r�DͲO>�RA0w�P����A�����C��OR�- e�Y�`hҲ́�e2��'od��`f�J�±�_�V��c�E����!�Z��u�Ր����l��k1"�2��i��&�C�		�9�tdD�:�=��<�$�8�A�"HBN���S�l����ȌPT���!W�^0��ɪBUF�+�Z����)΢qy�E�(�(h4�%.-D�"6NϘGKm��'	r��"�(D�� �%� 2��
�!�ج��H2D�X������H�$�7o�ֵ��4D�0�Roқ;d��uBL8*BJ9��c>D��{�.зPUv!0�Wq�R�
:D������^fᚵnO�W�TŃ�f9D�`�H�T.IR�B��-"}k�(7D�<k$b_�d�^�#��2'�� Bo1D��!t�P��p��d˔���#G-D��0�$�5řBl	,֦Ԩ��,D����l��h�A�k�
'�F}m�W�<�'�	�5����ω'
�B`j�LL�<�AN�)Z� 	�ќyT���a�`�<i7��/\�� ˶n�w��a� [_�<��.݅/�j���jY�9D&i���n�ti�U�U�b�1J<)�
�j��؂��/l+����k�<��
ՈFq֤xw�I�X<ʉ��ky�B�%�h�W�K����y#!+�B��lF��T
��a�C�I�t'ZUJ6��=&� ���WZ�pG���9�cV-!�($?�,@r��rŢ��E`�l�U0�>�O�1���*y�0�r��c����u��jʅ�g��!,#�~b��|������*�`M*��"��O�����8j�L��~jc��:+nP�
eOiA�}	r*A�<���m���G(ʩB>$���D��L�!*������v6�S�O�$ݳs�L�H:
(�%�H�)Z�'D|��u陛q�1�t�D'�I�7�V9@����d��YR��adP��^ A�`@�����,+֞��jͳ��!�jE�#����T�Y)-����OB��;�`�9C�@�B���y�lZ$r�Vi�A�(�T��Һ�yB�O�	��s�h��0�sWό��y�*N��"T��� ٔƯM7�y�B�Vˌ���䘖x���E�'�y"&\�R^�Uɣ�!qf����Ǎ>�y`W�_��t�ĀH�w��t�d���y�d�#(媈�n�5kOز4JY%�y2��	\|�)H	&���C&�y�(=B0��R�s
�X���-�y���O>f-B3��bI��sc��yR	�pl��fO[6PЦ� �A!�y�A�:�@`pm�0\�t� Q*ю�y¬�0`�D;m߱B��}����y"��Z��B�*޹<�.e��#��y�*Y�]��T��,���(!�5�y�ĝ��#�M֜8�y�Ɍ��yB�΀h�ؕ��B�C�����@ҁ�y2@ʗdkn�@ѧA�? ��렃ß�y�.�;&J�H��c; ���Sp���y 1�R��-�?�]k5F��yB��I���2 爒Z�̨cڻ�y�k��(����o�4C�V�q��,�yO�:�^ܲF�R@��lg�§�y�L�<Qn<Q4�QG���I���y
� �eѪ[�7a��YFD�w�~�W"O\�i%^�i�H��ABҴ~���Z "O���F�	X�N 0���3����6"O(iŠ,>�N���`��q�҉��"OJu*�h�RP�GɄ6�H��"O ���^�Z�ȉ��h�2���1�"O��G�9 ����$��M��"O ��fU���Q�0�Y�dȪ#"O�"/��[��J⏛�nQj�;�"Oh�)7�N-8�M�@ψl&e��"O���4�U�J���AA/}_����"OFD�rf�|��媠��3jtu`�"O���APSg�Y UM��h���"OʈY��~{�M���/4"O�,8U��4i�}�ଌ:1���"O"I�T�H5�V�JQ$E�b�^�K�"OLq���D��! ���:��]��"O֌c���S��
�Oȯ[�@�#P"OV��,J�	�hB�KN��=:#"OYQP�ҭ��I�J�$�b�X"O(Xs�kCd,��C��D��D+"OxT:QkY�S�,�`�+_d���"O�$ƞ(�9���ϴ:=֠#�"Oh��S	с
,�	�E^�??�a��"O�a���FO&�s�%S<!L@[Q"O�����f� =��j�;m�P�"O�Q��[),�uS��I)�"O��ʑ�ݹ%(\��7�ڦ-��h�"OH)Y�ƨn�����D5Sav�"O
�����M���ҁOd4Ȫ�"O�4qug�mMt8��$��+P(%�"OH�'�B"���E�ˁH[~�g"O���hB�V��1kp�J�'BxX�B"ON�
&T�4������cD4"O���Q����Y�A��;l�)%"O�(��N� b��� � �L��-�e"OX��� +͎1CV��p9�x�"OZ�pgB��f�|Ha�I�(�a�"O
�i����jR�%k@M-8���"OJ]�uLޖP<���&a�
4.�A$"OHѓ(P�r�uAu�
�:��"O��Iف"���Z`�<Psl)t"O�-qSԗʜs' � ^}��"O���uƕ'q�
b�OݞzԜڃ"O�q6*D/O������TĘ �"O��@#���7ĢM���K�Q��L`�"O� ��!@�N.�hS���{���q"OB�ӑ`T�
V��#����z6��� �����)��$��NB�T���&T�!�dL9Y�� #M�M�ճ©I<[q̀�%�Jr�	<ZuQ>��
�8#��e��%`�/�#2��M�ȓ8�(H�ňXU4&��cҀ
�>��(�[��=xeC"�O6���B�	H�̢��������'n���K}yP��R�z�A�*!+�����o#�ȓ`.���W-^5��i4F�#�L��<yd���%�T�0��=�'}!� ���3N��eQ��J�.��|��Q�E�׃T�$��� a5hsա߶y8L�'�`4��𙟜�r�I�i�����R&��9�E5D��C@R�rl�*�i��SX�)wҎ80��( ��|�B��qڛ/���;��V��0=�@-͕V��=H2렟��F�S#�]
��Z$OT1�(/D����` H%�a׀V)��F+所W,��r���*Q?�:����J����.`�e�2K,D��(T�ڝD��5h�e];31�h2�D@���AL>9&$�gy
� �����
qN�F��:Jj��A�"OD{�C�Yn4)�`��i�i�fp��Cx���&J�J����_�k´D�â(D�X�&�Ʌ?z4��\1a�����&�O�9�A<&�hTP+\5�HI�c��{*�'�����F�A���bvc�=^5���$W��Ҝ��1�ӲazP���� .�N�1�*5�C��5sf��L�V(à}�'�'�^�AV�K�I
���O?ͪ��l�̄Dc#g�,;�˃]�<����%p��9�郟,��$�I\yRgH�tZ���@X���S�8?�b���a�2Z~�����/�O���k:�Ҽ�FI�ZwHl*1#��`�P��5d���x�a��1a̽)����D���hO�l`��ue�yы���%BD�E�2��!԰��'���y�)2@�Y� ��־8i/>�?����1�0�+}���K�a��	��5>K���E��~�IBfj�Qb<P��'�Z���S
2dYG��l�Y�+Oܨ��ܶ}��"��$}��B@�N�y;�ǻ���<gբ�Ie��_�N��Ъn��}",�k�0�#&��+� qѠ	ӓIȚ���0�R�mZ /8}BB�V�$2�
��O����B̕~��@9iA��Xq�0��-PP+����-?X�l
�gA0W^ ���~�3��5;�k�-<����V;{@�J��ٞ�� O��xi�sgT,7?�'�l̻�d�r��M��7Y�dT0���ON1a�F<q0�E��"|�0�]��|��T$nw2�b�͝� �|���a٦MO�Y��'C��ֱH�t���[.q��f��#2�}"u!J�W
�� �Ƽ;�fe)2�'�DS�P�wfЃC
֖&>�Mr!K�R��P��yg(N�+\��v��/K0j���-U���ص@ujq�ѣ�%�OP-!@�ι/�r 鍒Q=�4����':q�t8�k���,i5�H0?�zL�ӧ�q����S?��S;m"���#��~�Х��C��r��mT&Z����I�M��P�͎K�`�'|��W��c'���2�G��`1��|�R�گ*�.	1�o]�h�����4a'�&���<o�$q��AW>Y�1P1֪�	.{��`��P0>P���J�(����A�R(2�<Y�$�O
�� �U�"�"��L��p�H�L25��&
�q���P0eF��ğ.��bDU��{qV���S�"�24��j��F
s�����!�&m ���&�Gm|%	�P�`#��6l�p J���w�2h��ߩg�Jɀe�ڻ=���H���:Vk�Y䪹˃A˾:��	�P0�i�~q�����R7���GMY0P��lK�D�0�J�"��$��g�N���ٓgL�ʓz�\��L;f-g�cm�F{R(��%Δ���d�\��V�9 ��a�`GY �'8([�@��0��S�i3��a����(�b1�RLX�D������n��L	�{�ET��̛��2Lv�x�5�r��'(��S�P�*�%?e�E/R�.��s�hJ�h�*&MP���V�`%�х�n��x���6�*	K��Z�bTX��>��	��Ub��n�\�O���[��� ��*/��4E�(�
�'��L���O�1���q�O�S�r��u�N�)��\:�>���>Ʉ�Ul�NU�r�ˑZ^X�Ī�!�D�e���;Rş+J���$AC0�����J��35�Iܓ%Y�
�?�H n'm��	ЇW=
�ٳ�ٹ?ia{�
� 9wk���П|i�f��*v���脧=�-[S�6}��шMp�K��'B��I�hW
7��}�5���a�d�X�}��(8�8��Yb�)1����ٻ^SR�� jРF*)X�V<^���%
O`�J�e��:�h\`_�<�uʖ�Q2����#}k�,]�d�C�ކ �Ӽ��I�w��LJ3��>�2�А$�R�<��E \�^�c� �V�����ƛ����+�+w���
�y��3T�V=hR�5��ju$��D\�KC��ɢ�1��{"��.�� S;O��c��E��A����.��V��`�TBR�bQ�=��'b�� ^WDN8�s)�.p0�K��$��s+̚�{"���z�APi��9��0�%�Ͷ)��$����'���O�F���h5�	R�F|¤@9Bȉ��XZܧ�H!�D�R�rW� z���#Q����L);�J]v� !�4x�ܑ�晆B��%�p�W�#�Q��� }������tP���)�� Ir��0eџ`����f>���|J�"� k0�K,7^j!�s$E}�$�l��b��(,OT�K&��#�n�y&��6"��տeh<�QK�f��SA�,.�a�¿�
���$ٙ;�81񥀥X!���<V	�E!�F�� �Ǉ#��s� �@_t�1!Drh��!�H^�����9�k�="݆�Ix��EJ��d]���&� L$��&M�.4�`�DJH�	gJ� ,n�����ct��4��� )՘2AF�1O
Ũ�Ǹ6� `�H�2!2��0�i� a�D˥�Y�O�b񊤎Ǉ�!�d�.��D��B��v��){�lZ�7q^P���++
�W/0Ț@��Sty��@l.�$! Q&u�Hd�EG�8�y��F'"���$jN!nS�i�(��Zdhrb�ϩI���V%K�S�b�ۀ��@�n )�� �b?�#$�S$&���D0��!rU�Rh���R�*��WC�c��E�$ɑ1Xc&i��"�O,15o�"�x���7��A�Ĉ6�8��R��`",��1���Ic�5n�F]sl�-@��"O\�g�^MA�k�|�+ (�=2v\���UE����oH9 �>�!��YB��
\R���cK>YP>��ȓ
���z��ض`��`"$�'#�$���L/5n�}��'�>�;S�ŷ[1,����NI*!ۓ;�>Թi�<�Q	a��çR `i� [f�<�6��z �h���	)�F��SC�]�<)�D��4)���2\�CrDDv�<d �|#���a@>[��8cd�<Ӭ�/�y�G�[�X��Y��G�H�<��X�}�̸9�%��&�+����y�M^!z��'�]g�a�wg	5�y��ɲG�%�G�aD�2�m���y"o���H��@D��1�����yb���_�D�B� ]��(�@*P:�yR��W�P`�ee�9G���'#��yBMY;"\X�S#��"��@CK��y�*s&� £�/T��$�e�\<�y��_hDmp��W8N�.���CO�yRA�<����V.RDߺ� �l��yRiQ(4�����P(⤓D�>h �}���k!�Q�&��'���A�m�1�P�9�@�2=#��
�'�8��8J�詄 �y�F�{*Oh<i�GR���2���|���6'��k���%�:�zeSL�<9dŘT���g�G�D��0�'d܊FFP�k���1��H:��g�*ZN�{R��xJ9���^W^����)QP���C�ql�Y�֫V(t�Źb�O(6B�A��?�O��s��ܬzo�wf� ��̕z�'
���'��:�ʅ�K?��$�SI4)c��Єj�tS��=D��h��F�P�p\�G�P"di��<�!�ԝ4`4l���T~��	�)y� ���C���� M-�!����i�fpڑA:�	�� �\�t%�`;%���^c>c��P�-E#7�h}9��B�g�g3����"ƎFH0�KO����#�n��d�H�d!�O�U��!n4ҡi�ϓ�<�>݊T"OnYrEQ?��c���2�=�'"OVL�!LL�)�\T�R���'����"O�q�w阀7Kr��b��-6�Usp"O�c�G�@�mÑEН| ��"O8̋��3Z|��p�CH�v�z�"O�8H�Ɵ�IyQ`D�΁P�i�"O�Bmא't*���-%�O��y�o��${I�(Z(�	*�\��yBi��Z�J +#�	^����ʍ�ybfēL�PICC#_p0LU���y2)�k�ډ�Ц��S�	�/ �y��p���Ѵ���}4$P�Ai���yb����a ���u#�=�P����yBX-MP�X �՞>�N�Q����yrLL-2��0b�U�5�lE��%[��y��Õ}[�b�!��Eg�Q�����yҢ��S>�;��41��t��,�y��@>i��Y��%�1}��"w�Ԭ�yR*	��p3E
�3)I8�u��y��@��PGQ#(����y
� �jT`� q3�c"9Hג�z "O��q�J�>>@����X?Ȱ0)F"OB��v�X�udTى� �,�~�3"O8�"(���|Ӱ+A���CP"Ov�{d�I7}Nʽ�F!E%�C"OF���#h.���V[�>d�I�"O�a��DtUXB�Q�]A����"Oj��G/�%9�"�w'B�bN~���"O������5���S��%2�mZ�"Ol���7[�)�+X
	4)�2"ODD�� I'$V����� /�<!��O$�@�Q@Daɪ,��`d�%����<!���#
`��&ö�J���7�ZX�&�@vy�/S#�j�bq�;�4�A����ͨ#�&���]��l�:�z�	qB�X�a��M�7��sՠ���v�2��W�M�޴�^1`uED0]��)�'C��1��)4{?t�q������2d�X�9��D��c�<)��0ʧ��D��	H�5��r���*�^�*l��@Q~2HΦc>{Ж~�&�ûKH~�[NJ<'?,��fFM0kC<�pS�=�q	�3k�]��OyTh�.�?!;(��a	�^^&y��'x��QaN�CIj���O�>��U��p?�]0g��@�B�� ���Mk�G?�ne��O?�dڢ+�28��<;�|dz��߮JW�O|�=��B0�f-O`Q�0��;��u`���)w��N�A!�@+c8`�s���*�>PS�Ԛ�~�ޫu��S��S�'gD}��/��p�D"�Ȱb]-�'?�%�'\)��rߚ��\/324KԂ`�i��&z:˓Q
��<%?��㜄DѢ�@ԭ� E8��5}��;�S��U�L0P��ꉲ���(l�%�j-���ј'��Ū�I�Se�i��
Z�J9�ujl��蟾�sΗ�e�0L�Ј˘d��ӑ�K���1�8��1�j��	+;�:��]�4u1��>)6�;�l�r�x���Iܢ|?h��N@�^B&���B���~R`�vx�"	=�T?㞌{q.��n��	���T�k#j| ��8�@�&����P���JBA�)E>�
�Pa�_�v��:��O�3�����p��H"�2J<�@>F�i�O"���t�t$�b�^��X�dP��xq�N` �c����~�#�jp
(_�(���>v(X1���0g'�����'mR�Ii��{f�@Y�)�H�Q��TS{���`�?Wp���Q�N�9�LF�!��;U��֫֐?08�ȓ949�Z�i����[�2-��v�bi�!�o�|�+0��|](t��'��Ջ$����l��A\�:� @��FunMJA���8�AˆlL.?���"r<Pb`b�6S�ptb I�N#<��Z�e�p�۹e�1�F@�J>�}����Up��C/��}�2�y����N8!c�@L�^W@�u�@�jم�%�N�9�Ɉ�U"8`QG�>��ąȓ �x䣅!� N�N�CS���Xąȓq��)�$ߎ)����шw��P��uw����	�<�q��_� �ȓV!<���	D�(��M���L���ic��K�k,j�������;<����ȓO^��ģ'✹2; �"���Vu�QÖпqn�1����=r�DQ��_.� �A�> DT9J�W/�T���NV��a��] 7��Q�ˉ�{d,��ȓ!<�k��<H��(���	G�z���bRbH�A��1�1���>�rx���ą�B I)�SqcV����ȓvv�@;��L�B'���+�J~0�ȓ��{FG[�h�pE(� ��6R~�ȓo����&_/L-~<����x�ȓ��D��E?�1PR`�Y!ށ�ȓC��e���Qf��ۣ��>v��a��.���h����s���#%۱�ܑ��S�? $�G��B��8j�-�7]����`"O�tX$�Tq{ԕ��\	��qB�"O�-����v�4�c̎�8ئLg"Oʰ����C ̀�
�-��q @"O���#�"O�Z "&��bJ\�1�"OF����·=ȩ�@�E�D3�5�p"OF�A"�ɓ7�d�5� *'�V0��"O�(�@4�f�: ��w��y�"OĘ5e� 	5ؕ)�jW�l���"Ol1pr�X�xN8
2�]V̀�"Oh\de[;�\�#�*�7�c�"O\P3iM�[�^���@-��E*G"O�i�2LY>+�<A� �z ��iu"OU
+X+��p��'kO��C"Ox%Sb�I*S@��/��Z�"Oн��)������@�Ÿ�H'"On1��'7��k�*��1����"O�ɪ(�Z�Հ�
�5���ڠ"OeC�ݴ?����W!>�d�4"O���-��x;�Ó�̞:��${a"OJ����7�ƄS�H8��E+2"O���E"��?cb���K�"j "O����Ċu��e`��Ζ��t[�"O����5 z֩A&�B�W�����"O ��e�9T�t�ا :󲝱�"O6�ڠ�^�v㴘
�FČc��5��"O�p2a��
,��ť0;.��"�"O��2���{��Ձ'�U���r"Om��E5�h�UѳD�z�9�"O(�)�/JA ���d��1�P]�"OJ��@�;w�|�G�\���e"O(�W����|1�"T$=b>��D"O���K��.4�ڕ] 2 �"Oyش 6}J:L3S/GJ�H��A"OV���Njw�!sgnȕ
QT�a�"OhLx���:̞t�e-ïo=�aa�"Of�yƦ5������N5��d2 "O�D�!�6Heĵ���ш,	U"OU�"D�m����Ƒ r�p��"O��A�Fe�t���D}�N�Qt"O(�a��M�z�͘�#� Y�����"O��!7�d��sB9MND`T"O8� t��A������ۓFG2p��"OZ�*F�F,���9�I�>;LK�"O�	�6�G��,A9"�T�D>�i�"Oj@:�I@'�z��-vY�,t"O�=��ۚ#s"t:#��; I��b�"O`%( ��L��ӆe�07A�ڃ"O���#Gޡ����0⛿.��A�"Op��l�0ʆ��v`4Ip��X�"Oey���[q =�`*�_�-k&"O$M����O����tC��C�
P"ONU�$"�/En\��Ә8x��"O�c�*��<itu���ִXM&�R"O�=�Qo��6�U�[hJ�а"O�-��]x�Tur�+�	�LK5"Oj�
��:�%ǒ/^��Ȃ���y�W�����+A�G�Xɻq$�5�y�
׊~iZk�6�i�%�&�yB.ӬQ	��+��RQXt!\�y�hʈj	�jQ!�)&jV���F�2�yfQ�,�A��'v!#c��ybLU��6$��h��p�Q�bG�y⮜E;��v�fK�I����y
� ��s�R�Q��$�LJ3*��s�"Oaa��C5F�@ነj�=�)t"O�x�Jy��
6��	mʴ�"O��P厄�qBEj�,6����"Ova ��G�c���vN�f�@!�"Ou�&l��0Y4`���[4�� �"O��`V��cq��3L�
v�R��"Ol�{�d�\��!�IG�3�J��R"O�ڃF�|x@�UB��Pw"O��3w&��;}������Y�G"O��0т�(i���x��G�q~���"O$�&��%�V�T��<o��Rp"O��Q2$[>�0l��nA<vk��	 "OxDaC�)�`r��8N\���yb�M:[�J���15q�`��Е�y��lc`��U�3<t�xWD��y��;]rn)�d��Ԫ]�T���'�
���"q��D[�l�6P��}��'��5�`m_7�z���F:I�HI��'�"d�5�F6Lͨ�q�#ÏA�xq�'줸��Ɇ-�&�!�L]�B	�'�`�R�x�}[1��	7ΰpB�'Ռ%3g70Ҧ	����4ZdXZ�'?�Lpa��9�|8{Sʎ2]V$��'��|��	��P@�5pd�7V32���'V(�2%�ɰ)d�	G�L�@B�'ⰽiV
!�M[�mC$�q��"OҜȀ �&J~1 M��M�ʸ �"O�T(( $UP!�P��
8��<�0"Of�,�1�:d��֢a���"O����pN�H�iU�r�2"O���6���P0�'���Ń��yB��ې�O�Vi�买AUa��q�ȓ/y�̀��I��đa�[o[�`��9�HB��?��QUaJ.��T��d�I�"�� �F�3�Ŏ�~��$��P$��AG�����ʦC�$���uW�i��fVr}�EC�uxQ��r�V �0@�T��o�P�*��ȓ�ea����� h�V��e�ȓhz��3a�Ǜa��(�d�O&w>D��0:ptc��# Б�jM�%����ȓG,u
��ú*,�u�cJ�����\��mP0�n
�� 'ǉ=8� �ȓz8�{�*��?���5'Ɋh����ȓ0IH�a ��"�d��AE� �N���^A���!�e��0� ��, �ȓG^��ȴc�P`��$B;e���p�P=�#o�b�Pb߷,�Ԅ��z���UM�.`։3 t�4�ȓw�>�#�kԲ��YJa��Ml|���gu��&��5|���;��ʈFC؍�ȓ��k���T,L�C���8˕]�<9��)�rt���ӷz�����V�<	�3{~	��2o�Y�4��]�<!ƀ��S�.ĩ�Ѫ6�����~�<!���"(���S������y�<���{:�gI\�@j���x�<	�H62L�|�G 
�*Y�v'�s�<yg��&W�`I��&T[yV� ���q�<G\�X���k��ħV}uH�]q�<��H�*8 �,�0�ܥ>���Æ�W�<ɒ$��Ly���O�)[������V�<a��^�ʾ�Z�̛�yaR(�%�Y�<� �<�����"6�ä3좴��"O ���U9!���f��-nt{�"O��L�!*���.M=D�<�"O>����ʁ�p�`���_+fؠ�"Ov�1�͒Gk&�c����%���"O��U�S�X�Xq�
���l�"O~�Z�
�6y
�r�$~,��"O�5i���4r����L���ܘH�"O�1���9����!��8�ə�"Op{#��,
7�/�i�"O�$[g�[0�Mx&'�#���["O6IY34�тRء���5"O�D�v�\y�t���F��@^x\B�"OPhA��A(B�(i�Es+"k�"O�!�#�I�n��}��D��<��	v"O�A�cߧsv�a�V���Qh����"O 5Jee�J�J$�ɅSdp��"Ou���B�j�uqA�ZPbh-;�"O(9��mȂ,W� �ԆA0(Dj�j�"O��)៬#F��S�]���d"OJep��ר-C3�L���b�"O��h�JʁQ�x�Q��U��ĝ9"O���6�L) F}���u��	 A"O�̀��P�H�@���c��T#�"Oڴ���\m��+��ϢLDV�q"O�%@��A�PB4ig!ū#��(�a"O��� ˈ�3����nO�+��ʂ"OX���Y�vy�"
�yp�"O2�ʄe��2!2	Z��5{i���'"O��RnΗb
i����d�N)P1"O��V�ӊu	�ZAL�A|�y��"OTU�#D� d�x�0#�¦|�l��5"O�(CЬ?	�|T� i�r"�0��"On��@�FQ��L����#)B����"O�d�d���y�4Z`&O�:t\�!"O4���%�cKf�����)C�"O.h����g�(�
5�Զ��9�"O�k��Q�4к�A��(c�V��"Ot�����ci:3�A�n�r�1"O^���c�*>�D�s��ߴ Y�*����I8�`ٻհi>�?Kt���A��X��.�=Ft �����ɭU$FX�ȭ(W\�+T�Q�kQD|+t�U\�'~j�5e
O*:��=�C�
C�X�%��Q�ʓ/�R)���)7ƨH��:��!"ϵ~@�ԛra
\p��'��3�≌'1�����@���gݽC��4 �jyFE3�i#�n ʓ�hO�(����ϬR#�H�E�ځ)����$���kٴ�ēY�HEfN�J^r����0=�L�pDq�����<���?�Ez�kQ�Ҫ�K��֡*��Ze�A�����
�4B���b��Z*"��`�?���}�T�97�nˆD|[Z�z��=+���9RCJ8Jْ��Fc$>#tP��k�#*��Z��t�.
(���Ń�W6e����'��n��x1T�i�b��'r�	��S��T�Iݦ��I]4G#��{�"{Va��'��䓱�3�@�l����d��T#� ��fA�D�O
9mZ��Ms�Cx���'����O����r��W<a�9+�n�;�R�c�@'Xכf�'%f]�qfθ���Z�s\$���R�4��8����r,S�K�m���p�K
�,Y��D�t�B_�����J�2�+eD��ʡ����"ȴ;E�N�q��A�*@�'J^��t,��S�Nl�#���3�*+�?!�i�6M�Odʓ�?!.O<�l��Ȁ7Oh��z���!bU�̄ȓP���闇-E[�E���I�!�t<	�|�v��l�By2!ͳ@p7��O���f���Ϛ�B�>(�$����O:��˘f�f�*%��8|^@6M��(��fO]�<|�,I6n��u�0�C�G�\�ԅ�0%ʓ)a���%�(\��"�Aʐo�~����#AVH�6j�� ����e�HxD�Qqb��T�>��<YQb�͟��4
��ě$M&Jy6eW
�@Ċ�gZ!��$�O6�d0�)�S�>�23��G��q�!��4o�(�'�i��O���t��-�����.��4Y
<Ʉ��<g��m�̟�ٴiڦ kB�i��W����?9o�8>��h�P���V"��1,U�#v.�	ş��� �S�H���O�v|��QN�&�Qe�|� l��!$X'�����	��p��x B�V`���E��5 Y�0�r⛣ C"d��'^��	��y���N�0'u4�����V�'M�h"�S���-;�	%�P�"T�Zu�d�c�L�铳?������'E�*���'M��ٲ8��2B:Om�
�MN<�`���S���J��n�����7m�O�˓F�~AP�'�HO���DW�,q�M�E,z��Z�瀔hi��rg�NP�`c�')+5|�'��5DBh?�来A%�P�bǗ9z������rNؚą��=ڴH�@�8��C�~�'Q�0�4����c��[�L�Ɋ(�h��d�M��i�bFJ<��,O7��!Ѕ� ��4y�hV�vt$����4F{���Y+|:%��(i�����;6��/��h�ʓOx�G����eBL[�&+���(��Z�
�����?�!'Q   ��   -    �  �  w+   7  .B  K  W   c  �i  p  �v  �|  	�  M�  ��  ҕ  �  X�  ��  ݮ  �  b�  ��  ��  \�  Y�  ��  ��  ��  ��  ��  � ) � $ g" C&  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b��IV������—3Q��y��L��z��	!N)D��RM��wu^�ϓ�v5��r��4D�`S�ٮe(|��+E�?vu���/��hO���_�R���
�_�\��Ö(�B�	5W]�lS�	���@P��qxV��=�S�OO��J��K�R����6���H��'zў��G�$Lg(pTF:<��S���������<9��`}j�ҥk��A5���-S�a}b�i����	���c�%k��\�
C�I�H���.�.!5�P��R�g���?ш�i\0�� ��r�Q��gf�!�ׁ|{���FH�DY|%"!�Jb��hO�$�Jh 5q{D����P? f�R�"O�ਸ਼�?������IT~Y�"O�a顃��M�T��'��I;F��gOv�V)GT���.&+Dr�@�m�<!"��:(�1xg'K�+�2n�{�HB�ɀnL��+C�"��l����
-����~�Dq�ˏ �R�S�n�# ��0�1M5D���Sg8
K�!�P�	s���h�o-��w��>-,�|�f�[>6�xY �&Jut�B�I>���s�B34%�� �J�9�hC�� f!�N_ C3f$cv#ťS=�U��'��,�!A�8p ��ҩF�5I^���'�e��AȲW|<�p�::�b�'g�5Z>F��)2!!"�������R�����s&.OJ�= ��C�9�:�ȓ~��;v��"g:5೩�KFGxR��{8�H��eԖI��D���^��^h�G%<ړ�0|� iZ�`U6t_^�8���7���"OBr�&�^%�p!Dmת0��Uֺi�]'������;�I9e�N���0~�v��G6C䉞�fXք��e���j�*}��9��k��Q ��'�D�d�ыH�L(�N�{'V��Qʎ6mǽ��d7}�ѓÓ<�􉐶M���Q���	�F�-�R��2m���q�X)ex�㞴nP���'aQ�Î�0�~@i`��*E?F��ȓ#�Y��$ɖ�Cir"\N�<�'�j]'>=2���I�Q���ѷ�ާq!�2�C<}�~���#�D�24�$]�O޿6�~(�d�>4�!�Đ�T<d3�A��.�=�5�q/џ\F�ԋ^�W�~�q)
uG2�Ȅ$���yR�F�?J�SU��l�2���K�<���k���O�vMPbW����q��ҥ����'@�-è�6B�� PBÜ�Z4�'�����U�#R�^�HHЪ�5�y�"�+K�TP��P	h��|˰"Ǳ�(O���I�{��`�c� �q�,��`_�tB�	�1',)
�\8JX��I%c�K�D *w�>�0��Єf����&"9`~!z`
5�O֓O����h�:�t�&+�L��Õ"O�L2�o�y�\9��/���(u��"O�� �@�>�K���=-�0�Ҥ"O�1h��`.F�9�#�/�x���"O��\e�����P�_��]Z��\j�<�q�K�P��`TK��R�l;��Mr�<�bX�k���+6�"V��;�f�l�<��G����"/H�
����h�h?��ͮ�P���b�[�����}9��dn_6,�m�E�9q��,��l�&��T�ĖVT��;� L,D�Ƥ�?����~�� ���1C
����H:��J�'|�?)*%���,�w B�=q±�b!���%�牫h��+��s����X-y��C�(y8�}ؑ �U��"�ρ_4.���'�a�	�"Qgv�r5�ϼc)x��p�C��y�lŞ>�Z�p�O>Ug���L��Px�i-�����]�1y`F[�?wvP��'��A���-J��l��FX�.��M�Ǔq�Q�pY�#��M��Y�c`:!���3�o5D��i��Q%ml8�&@�&Gk`�YK3?Q� �S�O���ЂK�.�֤��[j����'X�I�� K� \�A�KՄ���0�}r/px�Tã��;k��i�e�J�#D��#J-D��4��b��6A"�x��+D�\q� �#�b�p���
vl<�R�<D� ;�a�!T��ḁ	�%6̪2�9��]���C��B�,=B`�.ʘ���6�O�4�`)�R
J����"�Z�x�ȓj-(�	�a�Ҭ�	v%�?d�X��ON t�R,Y�%O]�&HW=��`�ȓp�LT)	�~�2�����:��t	���l<�V��&�����f/$�3��LQ���RL>���4�Vq�"^�(�tءM�N�<�������GDR�	6�ZE�<i&	��Z�z3C�P����B�[̓��=P&G�F̠�h���t�@]!��Y����`�HUj�$#���Q�\G���ȓ_,�d�FB�V�L�A� ׌Zt����hO�>!��"�X�i+�$�< �i*D���(�>N��dh�#�#�&L�ŧ���'���h��`�w��yX\(@C%'>���0����=��]Fy:GiۤR4�`�I�5����`؟� ���$�N%d�T���b��Α	a�O��=E��B��X�!����$�Q�S��y��ܴ��"OT�{t45K%�������M�	ۓz|yǋٛF5��J��p�4L����<��� �~2 $L>�Y�aa�l��<��ƞ��y�	�O����I�[Ɍ�
afŀ"�x4���1f_ўdR�l.�'6�r���$�G�B����IP�ȓN6���J�d�T��J�.Z��E{�'��$Yg/�P��Jrhܱ	��r�'(��D�J�gr��R��)kt���'� ���ʢL��9ȷ(ڲ`�Z:
�'h��`�N�.��TY�B.O���q
�'v�pu���N)������
�1�y�G'�Ş-b��EaSX�H��׾+4|��8��0� �L8�*q2��E7&΀Dy.8�	C��#�<1¥ ��xTyp,�j��B�I�yh�asǤ#����rf���C�	x����	+P$`���-����D��'����+��\<x�x@b<\B�Ј�D�r8���E��0,�������eʺ ��%D��طjX4@s
U#Eߒ$��a��%D���`Ǆ84A�Q�W}��%�Q�9O�����C�x�tZ `�mS>9��A{�!���+wĘє�S5!� �:�
2 |�'2ў�>Ӧ��HO~�Ӓc�x,�����/D�d��j�T,�Rc��n��{)�	W���tdƣ����\)מ	�2,���y���dD�I�"O3nFr���Ѹ�y�aT)-���c�(X�_��9�A)O��y���}����T{l�ч%Ӧ�yҠ��u�~Ȫc%�	XL�HW�N"�y"ٌi
B ٲK;<�Ȑ��@��y���?����>5N���4,���yB�'�@��+@8v�X)��Nľ�9���E~2e�l�|�1�7>q4��'Nl�0��i"�BP	���X�'
5���)����[�M�%��'�x3�f�m��:G�T���{�'�.�Z�T܂�F��v�6]B�'Vڰ`�D�Q�r)���@m�쉇ʓg� zѪ�;��� �E�<W`⨅ȓZ\�9 ���Tp�`��LA�|���nP�wM�<?tQ����H����N�P�R��`m�IZt��46I�ȓ|����#��.� �'E]�+!P���[@ʴXԨ1	�B��c'56간���pzDQ>X~��C/�$o\�͆ȓ� <��	<i��{Ѭ�!v����qh���&������4�F�D��5&�����|>5s�Nƌg�����\���oȑ:D��S�� <Ě��Um&�1/Ì55P��S&b܅�$� ��&

K�,������r��-!3�K�p�
�
7��lf�ԅȓc �0�C/H ��N��wZI�ȓ��Ҥ�τ$ �
��2����ȓ^�p���!�3LW7MƔ��7��ia*�d��!r�o��u:<����t���ێ.���Yj]�9�����5M�����7r`~P8tL� T����ȓs�u�&i:��40#��;�j�ȓ2��`�O�q��{`�W:B����|Db� �MA�x�t�wkE�tI�ȓ3l��+�	��Q��H�y\��S�? N�I�jĿT	��9��� 0����4"O�D	 �0VހTc+��~���ir"O������ %c�� �#�yB`Y�|��D�b�.X��]A����yRc�6&4�#6a��a�h���B#�?!��?���?��?����?���?���W�8�9����4c~�1QȊ#�?����?9��?)���?���?����?�t�E5p���	ZX��- 5_�hq���?q��?A���?!���?����?a��Rx��S�!Q$m*<�щ�,Yb�h���?���?y��?����?����?��eИE(e�Y���1L��$m:��?����?����?����?���?���b]�9��i]0	�&g�� ӚI���?���?!��?I���?Q���?��l�R�q���@�.I�!��"�������?���?����?!��?����?Y�Sˋ"C�,�R
8+,0���ß�Iß��	����	�	ݟ��͟��d�ϻ'��m�!��ZA>��c!ӟ����$��Ο�	ܟ����t�	��FD��)���u���1~`s�������Ο��I��|�	����	�H������1fQ�m"��������g�����������������ʟ��	�����N�*����d�}�0B��_ߟ���ȟ|�I���	ܟ�������ݟ�Y�ӅU�Ę�B�;>H�������ƟP�I��L�I۟`�	��M#���?Q�!X���b�>kU��a�{�IȟP������I��Y��]?M�p�t��#v
Q��Á�JJ��oЛV�4����m�����x��%��h
����9�ߦ�M;��}�KU��'��x'��ȧ�2��$�O�C�9�`$�.XFl�#��ODʓ�h�d0A�����u�w���qM̌I2�ߦYC��1��L�'_��w��Y�d���j4�5c�FH�*�
�pC�|�lZ�<�O1����#�mӴ�	�nr$p@p��5!�H���Fu�p��t�B!�*hjpE{�O�2M�O�@�H5"�����)Q�.�y�Y�(&�,�ܴ	��<Q�1��`�vEɃ*��}0�ү��'6�Q��f�jӀ�C}�+��錩�G@�{/��Y��@��d��F������ 4�1�>��S
|���}��k5O�2Bp�; �.C5Z]�/O
˓�?E��'+����L�O�8��Ԣ*Ctك�'��7�Z��ɞ�Mӌ�O�����
��jW�a*w�% RtЛ'm"6�R��	�ɇ{� m�i~�➧"XB\ �M*	Qp�v��{��u�&��pX�Z`��TT�9$o�_	��q��2���'[�U�~YT��X���H���(�HT���+�▨+C�p�ϒ�����B*��t}Z�'N	]�@�i��3���*�y�����C�����wFM�8,uYQ�<LȬM�`��s{�$��BP��Bpc�O�	�� ��DH� \��� &{ȱ'Oɦ[nx<��
� v������M�L���&Aw�P�"&<*#��p�J°OF(��5��<N�qr���â��>�D@U�N#l�\�R�  G�Q�����M����?	������k�G�z����./D��U�l�v˓"�X�Dx��G�KW��,h���G�D��X��4uy���W�i���'U��O=�O���ǥ2a②��W�H�4킧(Ǥ
�P4m�k��#<E���'�ȜY�G�@�"ų�%�#�	vC�v�'�Z��f��$�Oz���O�	�\@�<�����`,��0mJ�5Hb��3�"�	̟d��ΟYre��"��`)!c�1B�p�IӇ_��M���rP{p�x2�'��|Zc!uS�Y?Te���Ӏ��*���ɮOT����O2���O>ʓ$	��L2A����$� �J��dNQ5?�'"�'^�'�I)	"H9K�@89!��:Ң ��~���9�I���	����'Ȯ�B��f>Q��+��ĞYx��		v�qUA#��O��O��1	 ��'��P� -�0H�I�(��$���үO��d�Ol�$�<�b V
�O6l���D�/�XaJ�(S�+\ҹs�~Ӕ���O˓��� 1��>i ʖ1  4��e�ʥ0��*D����I�P�'L���8��O��ɒ1�>x�����&ڒ%"��ͭr���%� �'��ʏ�T?���C�()��=�`��@/x	CG�`�|�=��\���i���?1����I1Z� �)��ψw`ı�wI�F��6�<6�@{���O02��.���m�
JC�б�@�Ϧ�� ����Mc��?��������0����"-�{1 �r�1_0Hoڷm�l#<E�T�'c���^: 2�負��Zn��"Rr���d�O��D��&RM&�,��ʟ��������q�.@`����{.�>B��R��?���?I�	���s5�ܘ4�7��=D�^�MS��r߉'��'�ɧ5��9��L�����j��{5),��O`���O����Ob�d߿uZmȤM�2!�H���n
*8�y�!�<)O$��5�D�O&�I�Ue�Div��>�@
d��R6MS+W2�IП��������(��aVşlj5ƀ�iZDqA��k`��6���M���?I��䓯?A.O:-���i���)Ѧ[3~[ 	��hٴO-�X�O4���O�$�O��$�'���D�Ox��N�;H�ʗ�M
,���*���%�D�nZ���%���	`y�`�.�ēp
ʅIw΃:�<�����:���n������t�	5�:��O��	�?��k L�f�S�ƚ>��Q��0�ē�?�*O��Q��i��  x�lF�|���AI OH ���iQ�	?VB,E��֟T�	��@��|yZc~�(S�a�B9J�h�Hw�Ĳ�4�?���:��������N�#L��X�Bç#R��C���M�0�Ƚ�?��?Q����(O����O�y�ː*<h���CeA�$ܮ��ĉܦ���N	^�S�O~RJ�=��={�!5Qo8\ƣ��z�6-�O6�D�O�� �<���?����~"WA4�G�;fn �ҡO��MCH>Y�ώ2U�O�r�'6�G�P:�$��U�5�:�c��\*��6��Oq����<Y���?�������f`��qo()�rl3�MHJ}2� �J��'�"�'��S���u �U�"X`,�K ��	";�0�'�B�'	|R�'r�NHڌR�M��^��L�f��e���H��|�'�2�'��	�;��	��6
f��U�\�^��TЮw��8m�ퟄ��럀&�����LH�FX?	��!�u�v#�<vh4�*�%�u}r�'LR�'��ɺ4�@H�O���W9m(���J`��aqR�̟4��7-�O6�Ot��O�!��8�	h`�!SM�/V��QR ƎehZ7-�O���<���N���i�O �����('+T%h*�-v��L �%Qe�	ȟ���6S܅�	v�~�ѨG�&a
����$�iJP�G���'�d�0�'��'�B�O��i������1F92����a���g�s�����OBys«<�)�S�[�� ��>G�Lgi�,�7���3����O$�D�OR�i�<���?A!���N�4�v�L@?\X�s�VTӛ&��5?��O>a�	*Z�6����l0�Ɇ�iz@���4�?Q��?wF΍����O��$�Ov�I%;�񩜗wn�y"�LE�x^7�-��ݼQ�<�&>y������	�a�8�r��"���y��	Ғ�ܴ�?Y�Ӕ����O�D�OڒOk�X%N��]��
�-�u�beM�F+���(�q%�t�	��,��Uy��[�$�8���F�.������E� �����*��O��D�O2��?y�O�~`ʔ�o~�2�5:���4�?�(O��$�OF�ģ<��$����FTP�p�iK`��9Bm��ğL��ԟ�'"Y>���)*�fP2��WQ��)	��<.`K<����?�*Ofݳ�O�h�$S��`g ��.< ���&b�J)�4�?����D�O��'�?�-�ְ{�Դ�0����0!("�zU͈�a��۟8�'��:�:��O���l�f�W�B�J���*���(�D�i��ǟ��I�'k���	j���?�X�a���A��F�2%밬ќ.�^6ͼ<��웂1����~����ZԘ�TQS��=^n�3�S�Mbʩ[�d�����OP�����O��O]��Oc�sӖ4���@;!���P�K+�	y�i�0�w�'=��' ��Ov�)��;,z؀J1Ȣ���R����w����N�8���y��I��DBBt�ЁB1�C2�Bd�o�ß8�I���ǣ�lyʟ
�'��-#��xy�l����
��U�E&�	C�z�SN|���?)�e�P�r�4mqEE���|�T���i��'#HNO���O���<y�eH(�5Z#�P4N&�D���RH��'�����'��ԟ8�	���'��L20�ЍW;.|�Dj�#���r��G��
O����OR�D�<���?���]5A�>�+t� L?<(��kC Dú�b���d�O����<���4 XJ�O�,�BF[D<�L��d�h�^�޴�?	���' 2�'������McD HfGv��'L&�j���#�F}��'@"�'@�ɇ��L�fⓐ8�^ܒ5�P8,Il���B9BX��4�?�����O����X���=�CQ#w��I�p�I�C�Vl�ש]2�M����D�O���щ�|z���?I����5�1��`�T�+([�ǟ���$d1�U�<�~���?seH��nC%<C�5Ht��`}R�'?>̡�'���'(��O��iݥ�BHIf�0S��2~X�|#$�l�
��O�Ȼ�({1O����!��(N�d(���!9)0�ق�i��X���'#��'KB�O��)*���4M~l�c0Gɺ4�L���� �q/��&{�բ�y��I�OH�qsl�&J�Xّ+6�M��Eɦq�I���� J83I<�'�?)��n�b�W�9=��\����	,TBXHr�i���'s"��9e�ꧽ���OZ��+xj5s��״l�����H�7K�6��O��欲<�bU?!�?�SU�.Z�8/D<�����Jb�	;O�.��.*?����?Y���$��'�T9+�,M��BiI��]/r�B �"IHs�I����	П��'��'��p���+$�<�2�^�B���m�rZ�8�Iڟ(��iy���%�&�B����TdA*|��(7�ȎK�ꓠ?����?)/O����O�|B�J�OeKe�^�T ���2�07��YR}��'�"�'�b�'��e!�gx�����O�����S3<<ݠW�+I�6�vD�Ѧ����T�	Yy��'&�P3F���5G�P5�YȰ!d�ܺv}�)R��i�R�'���'�V5fFs�`���O��d�<ezDa��Z��Y�W�ayE�ZҦ���\y��'�(
�Oq�P��s��QsV��1- �X`����Ċ	��M{���?�W�	N�V�'�2�'R���OT��TeXE��7�Bɪ��i\@��?��L˗�?����4���O�XQ�す2H�BI����4�4�cشT�>l�3�i&��'���O��t�'���'l��9�"L8**Љ
�IiH�@r�OaӠy�R`%�i>c������ �1�*��莜�5jD�.Ł@�i��'���%3��7-�O����O���O�N߻jFT�����'���P��?؛�'�I����)J���?i�jF6���
g!� Ѫ���HD�i7�Fؐ�\7��O����O���k��O�DZ" x���_��(f[��87m�ܔ'b�'�b�'�rnԤy�&�:@n%(�h�c���7�I"�b�����O���O�@�O��I��l�5k�(Kֺ���NK��$���R�:���ޟ��	�,��������4��hP>�Mei��E�2���i�@�ϡO���'JR�'	B�'�	՟�Z�v>Y(��ڑw�%0�%ߘ}a�d�#����O��D�O����O����n��a�I��8y�b�v�(@� w��܂�	��M+��?	����O���Q9���'@*��q&F)/�x�s�ݡB�6a�O��D�O���� �m�ٟ��	֟l��- )��ۤ�U�	�F8cb�
	Z٨��ݴ�?�,OJ��@5���O��$�|nZ\.�	Q��ald���KT�aL7��Ox�$R42���n�ӟ��	͟���?=�I�m��P�ê@�ZEaE�b~�1U̬>!�!��,K����|JH?�G��-W�T�#SlB�n(��g�*2��M���Iʟ��I�?QRM<Q�@$�e���R
T����Dt�I��i��lR�'ɧ����+)�vP�}��eڰ	Ͽ��hl��x�	��0�B����'��O�r����Iw	 6�@�źi��'�:�� �5��O���O�}Q�K���X}��Ü:�|�gl��Q�	>�PxHO<����?qH>�1� �:r�Q`��Y�R�#�h�'��@k�'��Iş(���Ж'�.T�ĩ ����-��>��1Fd�O,�d�O�O.�D�Op,�V�D]*!ZP�0S��[��V�{H���<Y���?	����DSm��(ΧB�\��@�b["AN
-u�A�'�'B�'�'`�Q��'�fY�T�-^�%X�FU�d����>����?�����Dy��q(5��ίKGf�A�+ �]
�f�Z���l���(&� ���� �C�B~ܓm�X�{��['^Gh�"G���l��lZڟ��Imy�ΐ�A���V��x��dG�!m���F�֤<2���7�k�����I�ZUZ�Is�~ڥ�_�mRIat�R�5&"�p�¦��'|��$d��!�O�2�O�D�/B�!�[ ��ر��gt=m�t�	A�px�In�)��U&	
'�0'��j�:6�I�"�n�ğ �	ǟ��S�ē�?�0��48��+�'�1�Ι7(>V@lZg����c��F���?��ѣ_r���A<P�Хo�}���'��'&��84 !�D�O��d��hA`˂0�rUP�hG�5�\j�|�h�O��:��y�⟼�I�ܲ`'�$�0ɪ� �7f��<;���M����2�x"�'Ob�|Zcƍa4��(e����H�K�\�@�O��SN�O�ʓ�?y��?�+O>��FΊ�yR �)LƖ�
��l�\�'�$��˟�&� ��˟�Ib�
C�.K�V��I�K�(mT�$�T������`y�.��6J��SX�<��#OX�<���8A����?����䓳?���O�E��tFm�� '*>�
[6���\�,���@��^y�AT	d�|��F�w/|rB^�G��B+L����K�	؟��	3/u$���`��S�r��h��A�iO@�1�
Md��'�"]�� ��V���'�?���z�� Ì�"�T��Ec�/N�􅈤�x��'�R�O b�|��P�2,U�<u�9ɢL�$t���iC�8wh���4b���ޟ���2���ψF�(!�Ԇ����2J�"���'���H�B�O��a���\a �}�"J�g�4()�iK���c`�����O������$�擹e���7���3�8�#��P�\~� ߴ�~-#���y�Ob/G��㤍��f������7M�O����Ozɪ�.�r�i>�OT�Y�n�:�~Ä�T<N��s�i��IfyB�"���O�D�OT���/�/�^�B �S�u��d����O��d�G�%��@�'9��M=t}���B�*j�z c`�Rʓ�?i+O���OP���<aӈ�6i��Ze��53����L�'�p����xb�'.R�'�������I�k��#ň��1I�q�lϔ�A��.�	���wy��'7�H���E	F�M�H(����V� w�i�2�'�ҙ|"Y�p@A��,+\7mʼl<@(�􊊨L����F�(��	�(�I͟@�	�����p�IU?aPiނc��%�� ��,�D�����I�	q��˟L�	62k�x�a�/�DV���JE�M�4Xc��B!+����'i�Y�䚖����	�OZ����	Ӗ��C��UK�J�L��E榙�?Y��hOk��YJġAX%WN��ݑ ��&�'i�K�,Hb��'���'���'kZc� ��<Az���I���eCܴ�?��_�X�9Y"1O��$��?�(l�0�'.|HhŶi=>�xB�',��'��Ov��']�(Դ�r���#>t�7��~�¨I�OF0��)�S՟�r��vcb ;�B�$f���/M/�MK���?9����)2�x�OhR�'h���k� ��Y)qM 	�|$ː�1��,cb�X�I�`�	�-�;�Gԍ-6=��-D���5J�4�?YB��?A��D���ʟ4'�;�,�yM�����;�x�+�`J����D�T?�!"0���a�"��NʺK��� lDc�j�� ����� R� MP%ީ,	�Z��ǥ;�:�&,ޓ$T���h�V���8'[��G���>a�-�!\��3"%��v8UA��b�z)���̮;��Cbd>\m�4#ł��i�<ڒ�2.R�#�L4X8��ZR�Ǹ����b$h"��F���/V���� �k.��rpDHpT�J���)Gd��
.
B���waD�wd�0���H�FZD,sc��En�ț�a@�1�4¶�'/�xhRƁ%�p@x�bX"��M��ğ��	 Jb����]?<t�a������yrDT�(�F��B��~��k`� l��h0�4ʓ*Ҫ���«M؞xb�k�G�f�1�͘���,�%���
�IbU-ɶ<1�- ��0��n2�)���M[��	�88K����bS"=��Y�F,z���O(�����'լ́�'\�7~r���-Y���y���dD;��O�>e-(�h�A/��1�T>O�=�VȂ�m��០�Ox,����'���'�V!��r,�/TԼ0�H�Z��H��܁=��}��Z�
<V�\nU��a��w��ʲ�IN�|�
�*=8����Ƶ�@���	�E���`�ЭZlX��˄y��iR��|�]�k���ФT?������WMU�� 柄�IG~J~bI>	��խRq��۔�ϱK�
� j�^�<Q��O-kd�(�*WX���g�Y��?QA�i>��	���8�`�.'�z1�F�Fb��	^y���sER�'.�:�`�]ҟ��	"V�z-C��Q�ͪ	��� '�p�I�EF��K��4�OV���A�Sנ	���¸��(���^���x&��,��ʔ?��(�9�|9�"ŅA�x4��>6�����/.P\H��'��g��Y����_y�	�
Zx�좇�W�:^�C�����D:�O�E��B�-��D� �r���qtg�k}�T���)b*O��HdԦYa��$J8B�a��KfYHAG��֟��ʟ��	�k�r�S�,�'G+�՛�N���E��*V%�h�/�:�JY���&�Ox9Sv�¦2��Y���
�d�<0��!$}������p>�C/W����44�D���(����q ChJ\P0t�iG�U�x�	m�S����9l�R��6�N(k��2EE�8�yB��Eh�)Z���>�����#��y�˧>i.O���el����	��d�OP�0�˷G4,�b��AR9�)J�h��u���'��bS�U��X���?aX�ic�/
h@L��'E�9X�oT.*׾�v��(vO�TGy���w%6�YI�7��F+/k�@�'Up@�ǖ8z�qЀ�0g��Fy��P��?I��z�O�҉M�z�`5��1@�YiPLZ�)����s�T��%8T�J��z�+В|J��=�|"&�i���'�v���+�$���C8w��(�����Q���	L�4�����'v⫄R<`l��V8 ��(�[%P��(V��1<`U*�	V�r�T>e�|��n2�iZ1G��A����HU/on�����8# <��;�T9;c`�D��?y�gĲ�j$�t�U�O�ؼQ��'xD,��*f��%~��d(���z�-VI?ҵ��#��/n��4H�x�IBx���ƣ����� sǥ;�j� ?�葞��OV�e���D(��AčԢ^{���w�'�怄iڊ��e�'.��'�t����ȟ s�P,Z�4�������"�K�G�
�A��:;R�˂���t�ӹ;Dq�r�J'Y�P�9�D�o�D�$%�)'�z��L[�0Y�Da�� h|��۟v��ǘ'�����>���$_�P��փ��r� �j?!���֟d��4W����C�t�G�qe^�i�V~��4Ҳ�x�'�U9w$� #R��`3P{�ѹB.�o��f�'E�I�l�t|cܴ�����<�Z�8t�Я9��H��?	���?�����|
������4J�0Q�EGj5$�ô��%,�.I��IC�v�ׇ�OV�hD�i�b��r�\M���XE�'L69����?i�ň�M����V�?����ak��?������O���8^�(�h�ڎ��`�QS�:C�I5Q��� ��]��k�`�&,���ɶ���<Y��؝`����'�rZ>hbއ%��U��iم~aNS�'PC�M�	����I�%(7���>-�E��2�M�v�HX����鉗$+L��)�[�4�Y䂞��(Oj���4i� {�F߃
�<7��Hh|�3�Ħ�:0KV�F9�][GPm�B��(��FP-�	��M;�i�bU>-�4�(!����"��<T����-�ԟ �?E��'T֘����!2ɑ�E2��%x�O(�=�'xӉ'�@���U!:�4��F
�"�����'9nM�Skc���d�O�˧I�F�8���?���$l��!j@.�Ɉb��w�<����ݥ$��@{ө��$����i#��O4�1����b�Gl8c�&	�UIS�DC@iҫX�`��]2��_��"~��g����- *p!���2>�`&A�۟��4HC���'9?�dR�sEjD��H��M��B�/��D�O0��Ę }IR@,�_����s���k��H(�􄞖���<��SuBb��2���X�V���O\PA�]����OP���O漬��?��
(Vi�1�� ^�l��d� g�6��`�H�%گ����	�t��"k�&֪Y��XE2bV�
'Q�tKG�.Y6ހ�v#è��$�)� ��ƧM����©�,���z�j�Ozx�T��O�5m�9�M�gyB�'��ɘ���p�F���@�f<C�	�U9�Aa���.���I��ɼ �.̣���⟢�ħ<��@���F� 8:�(���Ŗ(q��a��́{)��'"�'���W�'��6�T���g�N���W'@�Be �  X��J'�A�?$��s_pf���;Cy\��@@P$AB����8LyN��@
�\_�9xs"ŗ7(F-ZǓ*7r%��8�M�,�;+�8 ��L,s}d��1�H1ɛ��DOr��y�A@�([�k��*U8�r��\��y�eݮ��	㤎�Hٶ�F&D$�y���>�-O����b}��'H��X�$��PON?z������X��%�C؟���ǟP���A�� ��i��I�$��RX�4m��y�6J�H�p��S��)I���W	C���4��p��)s�ϔe��� tJk�!@�#I	b߈ى���3T��8�O;�@��A�I��M�$���t�v@����N:y��X�h��d�O���$ܾ#�����-t-�s@��Z�a|R�>��8��4�M$�쳃��Z�$��`��`m�ܟ �Il���
|��'��*S�J���:%�P�l�FUz��R�%����g/�6gG�%٤�Z%3`����*z�.K6��wi���r!5#̱��!�g4��f�!gܝzQg�Iw�h)���)\0�1�.$	�eǩ|���!ھD�@ώ�[�%�d���OKF��ş��ݴH��V�'�?�G�h���k�eK�	�N�i ;k�D�O����K�/�C�dW�2a(@��/[�1O>�P�'�~y���'+�)#B���M-��9�iC�~�`�0"�'t��A4<���'�B�'��Ic�A����)kU>F�ؕK���[q)��a��=�_?F��u9֡&@$�ӷO��K���ܤ6Q��R�O��d}1F�D�(���kC��%�4EBRl�T,N<��؟�a�߉U�^+��>���O�A����}~H�� �c?ٗ�ȟ���C�	ȟ���FyU�P�ا��)H�pMnѻ�xb�'� �G�Ȣb<��)�����&>��|*����đ�n =l�<�qr��Ek����&RS���	՟����8�CΟd�I�|��EM�sbD��I��1��ô���?d��w��ajFX��I/;�ƘRǟ�bk����*ދ-] �p���}�,���&�O��W�'���мS���hs���`7��1�㕐<��'?b�'��O�Ӟ��`BE抗*�PY��O�:��B�ɳfz����(�"�Ba���k��I-��$�<m�-N/�f�'r2U>1�v�@���0�S,Ta0M�4�
����۟D�ɰ`^j���;�)���J^����*����ɟGSQ��'cGN�Լ��"�ӱ
�dm�c��j�
T�`ܪ"l�<!r����	t�S�� ׫S�Uj��S��Xi�T��C̟$�?E��'0�	#��Or�0�->�L4*	�V �'>����H�U�����:�4�O(���<1GA�L��$�-��T�2��F�V�<��Eՠ��-��U�Du��Hn�O�<a�AZ�
"�5�E�̛3��8'�Xs�<9t��M��&m�8�Z��sO�I�<9���d�D\�"#���D�؇*�G�<	��%��=q6�E� ��H��K\�<�fϑ}���&�1&Y���Vb�V�<��
Ș'VBX"G�0czZZu�NV�<�!���Vi8���N�D�h�fR�<�s�	8	-@)���_�s�y���T�<�`O��d H�fJ�v��e���PR�<	fJO�,v�%aG��Р��J�<q!#�2Q[A�!f�O�&3%�k�<a����<e�V�I�w��]@�Ff�<����^i ��	,��!����H�<���+���v@�9w��袄�E�<�$���5`WaR�K�n邖�JA�<���Q���a�1t������q�<�A�-�(s7�E�|v�`�E�<�#`L3������*5�Џ�V�<�Æ�@u��)��#ZshY��O�<q@lY?1.���Bl\V G��E�<���U�-� �欗�;ZX]K���h�<��H\.�1�4BD�[/��&{�<i ���(��V�`Gr�ڒ�M�<�D�a��
�MяfF�-х��I�<� ����Y'a�^DN�)�8i;"O��I�J�1n�$s@ɯ��l��"Of��U�P9�,�c��= !
YYGj��
��1Ģ� U����iA���p�x�ɑ=T�2K
d����fQ���>��܂�48p�ϙ; P��1���L+�fOj���� h~���f�.&���j��N8�t��H��k������F��h���<�$f�}z��ӕ)n`�ys+D� �VCb>O���b��P6�$�gB�*,,�Q,K��Px���-`L��eĉ�Ȅ��ǖ2�MCШ�Iܰ�:���;��P��)��Ơ�(��,c܈Y�cA�.[�Zi)T�'\�X�gI�<�	x�Z��d��9�4<`�e�5N��1�#��x�/b�ɂ�b�Y��Q�	V8�>��R�J�#hg�RE�Z� ~Xa%�"��N�����֟�L�X���E�J������n�D4��Z,yeLT��,O�j88��GT�?m�Đ��U�ܨOX�8𩊇C5�Q��v�Tb�ըC��'l��'��
�CT5"��O��`��	�V�t�����>cx������!(�l��-�A�z�A`p �"@&�I 0�>���P( L-�Dh8��Q*\��E2a #h�9Q�t#�
p�첤e*,O�M�2N U��۩Ov\�F ,�*�!Ef�4"�b5��d6�I�"��6Ɲ ��T:G��>)�f�hv���<	��%%8�볦; j��"#ˀL�I	6��=�AN�!Y����~��'Y�Q¥��4W���i��@v`�`��)X��mq��&<<q`�,&A������T�'�Z軅��;4�p���Kh3Ţ�����[p��'lޠ30�����^�Ч�΀�	gLF~ �iu�.yRa}��ހ@�yq"&
o����F$tK>�'^@1EO�L��\Z���ByR�q� �Y�aP�?n�@� �-M��q�$�*|������'�(��A�-x\��Ӫ�v�pa�EV~�����]��j�(	ty��µ3)��A�Mظi�������/hx"$"�C����u�T	$nOZX;��ȉR��!��'��A:H>��Q.i8�d�zY���g��>\��в(��M����:&
��!�'Vq�6�Bl㈅p�_�<��LP�i')����@}�'��a�$��Du
ű�d��?���z>�҆�F�9�fY�5g�!���!�|I!U�K�G5Ą�aj ��F�#Tć4��%{�'�0l�1��"6�O�O?Ҝ�dO[�F��9h�L�:A��]�	˓\qԪ��5�����W�sj(�8q0�p�iȰ	K ����F�r@`���+W����I��g�W���eTA����W�3�Xy'�k3��=&�J���B��WB���%P>�g�be�S�L)Y-��8�iɃO�0�z�'F�~%ȕ�Q*����=�!��>\r}�c�ёK\�P�hE;�ҙ��-�7zF���E*%VE�=Y��A#2��Xc�l�ڵ��`��U�\G��h&+$���1��F%��[�E�d@cV��"$���c�{�`�N�j!�"l�p��$
����A�NW^�Y��N-�D�!ӊ.ay�nٽ���2�S�U�89J���;S6�L2��.b�P���P:"���K,np�]��D��	[�&��@�w�#8)�u�X��q�I��dy�$���&�9I�]3t7����%�I?gj���f �:w��mҳ/܌t��q�).��1�f�ys�z"bP�7���,�S�<���ê,��yGc[�H���C�'FEQ���.��)A����eDS�x�ƥ��ɘ0���Qv�i�*�ЀN+zzdУ4��OlH�6�S�J�赠өW�@�
@�wʗ�)�$`�!��s �Ȳk��:�5Ҏ�$Ji$�hW��|��᠁�2��r����6� p��4&�R��Q��Q?)4��?��0ÒJL�z�;��Q�\�wg*�	�	�~l2�\�J�r�8�
E/�� l�t��ԡ/�P)x%��$�6�@&L���'���s�隡Qi����H"�z��ÏW�����p	�/k��h� %���J��$+y�5�n��.RF��p��#?�ì��q[p<p%j�,ߨm�?^�I�k~�T-�:|O|�9dB�H��� �/7��{���	`?���	Lܓ_��%�n�듈͹XN�O�~qS℘k7�3�i�`���ҋ���0cL$Y�E����6�SO�>(?�(�q�4�4l�5�.%��x�$&�IA%I��H��T�ٍsAb7��!	�i�fo9|X���&Y�ǎO�uGX9i���{�|q�I�0���Y�z�E�W��8b�/Úc,�5��g̓X��S�J-hs�^�jfٹ E������ܲVWj��d"��O���W�-L�J�Ss��[r���"A�?I�x|��G]�w��t#å^`����t�ֵL��и�1�:�]8;�(�[Ч@u1�-����,
����ቃ�A��eR�Ĳ>`����'@{^�O�%J���w24X��털6X58�ʐ+�jħOl�hts�:Ԋ����+OLY�R/�+=R��za�@;d~��Z�.�D��W�s6��E�	�>X�8�KӕN��t�Ob�#Ʀ:�\��a�2[�ZDr .@�y��D�.��5�D&#��� ���ܔ���0Je0�w�6�2�#�M;�"QzD���OVD���T�T��O��U�P��B�Ȥn��ɓ��vL\4․Q�ݨlC��\�8�.ak��M1* ���Ӊ�&tI���
�6�\5���A�\]�mA�'����f��Nx�9F�ho�U#;�	�,g��[U#�~�F�����'��0ʞ'=�ષS��U�����8s��1��Y=c���ecA�*ȾȊ5K)'
�0�Ca�'bP@�$t����`ӽ{�0��P�1MBc��u�&��GR=L����&0~���hÝ;����'"�� X��b(;��u"�'ދhҰJҌ�������$I�
l��;I<!/��&�T�
]�Y���%�["p2	̓T��U�ؚ\:�� #��՜TIT�,��ˡ�J���\/9y��Dë��@V�AN̓��� ��$U�;���1K945V��	u�&Qho�<����k�<(���Q�n�v�F̢Ӭ��26J4PH�a1�R8���j��U?yנǘb(`��ת���=��)D�7�z�+��x��'g
�Z�.{yJ��e(��G]�#>�RY�&
�O�� �pj�V?<8oZ
|�E�a�-`��,X��7���>Q�듪v`�Hʑ�ˬʤ�&�D�<)�Ɖ�q��H%D#,�H5%?��D�<Q�0�jm@EB�D���:e��<&T�e��&� �>I⌌֞�afH��4�����63t���V�jj�@d�T��Z��|��&f�E�X�I�9z����a�xa�wfñ&�m���da�׮!��2]d`�Ӧ�Y�qO �)SҮE�lѢ'��8�n
UdT(2�����/~j�O����G]	&���؈� !K��O��r�o�wm��質�v������xf0x�{�l�8;�)�.V����iȟ�*�&��3&K4�D�7�'`��B�#�E�G�<c�(��d�-&j|�Vɗ�1� ���F�;M��5i�l�[��"Xl�ל�$� \��$/��A�˒?*֚�9�LM���L�v�0d;Q���f�	�N����d}�]�P�܀~di�OF|��)��%HU���$�2Q��]�%��ш��$��0bT��y"��p�T��U)ld@5`����&�š3O��������0k*ў�2E�!'���Q�f%�ġ�!Ī��H�<3��a�W.0zn@	�ž��1G�?e��o�m�'���O4����ⓤM4���B^�hH�"�|�>H�@�o���i���
R���D{Zc�NQ1�+��tf�4�RbF���(b��Ě�?1�#����'&(eA�K���|3kY W���"��B64=Hٍ�d�C_��X��0)q̻ ���qA$c�G��2t�8%�e�Ȫ s���I<:h(�?�O�l�*�"��X��钷E30ip���B~
!J��x�bI�g�@��5ks:\�`�?c�(���]��U5@ZL�*R�d[�OL �"�O(���M�ui�U�ݟ"%��'����G�f׆D���tK<x٣␱ih|�ireX�9@�hB��	�|�?� �g�Ή>5J��%m܌Pˤh�	8��W��R��
�D� G|Zc����#.#L4\`�X03Ǿ����'_����X8�1�L�PR�c�6����\4�A�K3U1�܇��8�4�C�[���12c?���ȁ��0��I��M�3⹅�	�J��	A3,M/w��]���i�|i[{�>���I�6�@���8hX��9�I������)�/>47mB-mv���o�`�y���4n��E������)\�L���ݎ���?�V
Q.�k#e��E�@-���Gg�Ibb���-���@�×e�'>�0�� Z�$�8y��o���l0�#:���K���K~���у��5��B�-Vflܸa�D<�BI�݄�	�1��=�կKPf	���U9r� ���I2 �ׂ� ��H���Q�	��GC!r�N0��I�Ip�OS2N1�b��'T1`�;8jL��w%(S%�UDz2��3A*�2f�<u&|̹�����d�}7�Ҥ�	*%�c7r��'��a3	 /2$� �s�I �l���{2f,@hj�6h�=�~��sb��M� ]� ^������N-zj�v�'a���.M5WvWc�*�Zp�B�~�b�I�Mݵ�����p=)��_�0�T��Gr6�r3�äR[�q�a% �I��9�g�*3�*L�'^Q>qp�͓�n���qF F<.F � w��kX� 8E�ȳN�x0�!�,m�l!��[-+VXP�B�Yb�Ɔ1BJ���Ba�Q�0��-�)����Q�D���k�2�`���V(K�2�`* eh�,!���<Ȁ�[ݠ-K��)( ���߁���a�DҐB�L�8e��Y�����
�!+ JD�Q�F��,Ј�i� �± �Ϙ'A�a#�2#|���K�\gri��4,Ģ�[�k��>x����\-z����,�!�Vيa������4�u'E�=Xy�t"\�B�y�
ɻ�d����7���+ �z��  ��0�:�"���gj)��� @ѐ9
��f���]w�x�Z�?	��	�H�]�H� y������7����D�2@���
����w(���g��2�v���o�� ���A7Z7��u���ӞI��1���'6P�j��|ݑKc��D��ײ*]�2� ?�N�%պa�2�L��犓�h7�O^���� ?ں���r�v�y�[�h�Rb�*��t�%��,�4;&����Ov��cF]�n�v����Q�?̘��`G*~���bc)9��I�d�����,yo`�2U�+���H2*������H���غ]0|)� ȁ]9f��w��=3ń��13"BQ>��~�4��h)���7i����I��'QR�ۗg�r�l��&ǯ?�ݱR!�i�΄`�Õ�lxj'�k�����<��|
� �k����F���{��X�\���K��%A�������x�I?����C�1�I�CO59�峟��Ap�8 ɒ=_��FXΛF;'�d![��3b։��'�k��� ���kv�R�W&n���(P�Vjz�	�A��?ya���~��M�w!*��H�����.̱S�,�8A���I�:�\�٢�[/sB��ѧG�-$�̓m���0۴�M�u�)+��q�O�	�}��x�S�+I�B˼����SA�<� �U*����I�"L)�-s�)K�BO�Ѫ�Y�`Hd�3��ə�t��&��he�	�<i�� �U�sMP! �=�O�ꂆT�N�*+͜W�ĳP�!7��Q��Ԍ"1��{	�k� 8�1LR�nO,�r��"$,HD|b�$G��Hh��%b�.��d�Յ�w���iEc������"O"���cL�-�0E��_���5O�EۖC�����	.Pa����-�JC�3�H��Î9�y�P�M�yG��j	�Lz���2w_ D�"��UIDn�#G甸��Oz�� ��J�P�BN�\�x�7�'�<�ף�4E��a!��ˌ}���r7 ��'8�i� 	6r9�͆��,���C��4l�$:Ç	jDܣ>e�To�@��CQ��ħov��E�+2�f�[KÆ8�b9�ȓ]�}I穓��r�C:`�:���?JF,҃�܀.b]�გ�%
�4�ȓ$Y�E�N��U+��\@�e��d�n�ᦂ�%0
 ��oZ�I&�؅ȓ�}hp�ɡ(�q� g�4WB���J��h��e�K�/]cR}�ȓ�|�k!ꐘ�
P�gI�
E���ȓRG��`%�O����p/PH��$��7AH�c�Z)d���a���`��1H�&��%�n�[�$&A�L��mxب�QB���G�Ҟw漆��Al	8!��+S���r��j�<��.�%T��᫡G�����&c�<	󯘿����.�驢@J�<���J\��`Y+E�@'��G�<Q�\!j�<08�n���A�0A�<�r�2��쉀��9&@��9��Z}�<�Be�4�d0RH��[��C�c�<�V�˭[��fI ,�zhhph�h�<�rk�_���j�M[<dd�qbOa�<Qd&��� vm�f���wE�d�<u�I�7�ny��N>KFDl��Xb�<�@�J�j�} ��rA�0���SF�<!$;r_�)�7M�h`���g'�v�<a�✃^ȡ2��.�j= &�
u�<qwo�y\�k  �/G���Y�t�<Au��Z+Fq)d���}cR�B�K	z�<�T,k�4� �._����b]�<Q�٢%6�I�M�9w�����r�<Q�������%���C��X�r*�z�<i���.E�(q@��=^ &X�Q!a�< +Hv�`��U�0IT� ``Nw�<�W�rO�8�s!�h{,=���W�<�g'	-�$�#o�~���[��V�<'���.,�d��}��`;tOQQ�<��jZ�Z��<�J��BȂ=�>T���l�
��Ċ�	�wU&P�� D�4{֪��q�Ɲ��B�7640�e2D�H�Wꚣ)�R���KE#^�Q��/0D�����b)H�M*nv�q��Ox!�N�.�(H���#t���+�,��!�$7>�څ�f��5�&�PeF�!�[�� 0��2tlq����4Xz!��,�0��WƆ;_X��.�*!��%�llSŀ�n{J)aC�Ӏ�!�D&A
�S���`a2E��l�:7�!�%tl�G�,[�}�c��&)�!��5��s�NY ������N�!�Z
9> ��%���@bް|�!�d׼l���)W�E�=�r����S�!�ĉ�:�b-��ǋAn����W+�!��$-���ֽ]�� T�٨;j!�� �@�sn!D�ku%S�_��qb�"Oj�VDں]`���႓$#�pV"OV\�E Z�S����X,���"OС��"�&` ���?�t��7"O,I���C�̔E��>&@}�V"O�(Y��`<8��]�JJ�u��"O��[Ŏ ��|�윣y�޵*�'����9>6I2��V��2�'�쑐��ܼcи�@�,=q�I��'L2-����53��H�j�	9
l8��'�z�v�̃�,����۴8�J��'0�IS%��"n�P1b�GI���K�'2�0�� �� ԩ�{��a�'�~��rA�+5`!���� ���{2�'��u{��L�mm\p���#����ē��re�]�Y�b���p\T�ȓ7�c&#(L88��R3Шa�ȓ}Z\�V�I�Y a�Bn��dq��UH$� CO�p�P��^�y�j��ȓ&���W�U/|N� 
S��	z�ȓ5-��CQ��ܔ4�toFA�>9�\����*��v�Z��S�H�XP�ȓ���ks�;a����)��Q�F��+O\f�ܬ�d��R/�_����>��-S�͒�?�F �2� \����ȓCH��5���F�V9�C�W!Pt�ȓ{;�a�Y&6Ζ��E�^�m����;�L`&�ӤZŠpA�E�l���ȓ?k���kJF�<�Z@��1�B�ȓ08�9�1�I�;��Zf�յ��؅ȓ~�:����;+�1��!Q�vP���ȓ�I+ɛZ�v�Y���]��Ņȓc���z�@X���1&�ZfS�=�ȓ=�r�ApAQS>>��O�`'2������ۃ�Y�i���pm�.;����;T"��p��7���$)R�h]ɇȓ.����MW��$�V�d�����S!���Q�Ȕ��xZ�N]7E�v�ȓ ��!dL�!��A�OD1U�`�����,�&A#*]z����*1�T��eBI�0
X	dt5�.¡\h̆ȓ|:�.:�8���� ��yQ(]n�<P�9a���Q2g�l�4YuG�R�<�=jd��[ḧu�Q���=Y!C��ay�E�.�=C��w��&�S�'YF���*K�?�R�@�MQ�]��B���@^6�0DP5%��A�ȓ"z��s���C��yЫ�:�5�ȓo�@��χ�3_40aG!��pLz��ȓ?���L�b�� �3@�
s�����u�bX���7`Ĳ@�d��d�:�ȓG��h���p\�J������M�ib�%^�4�f��<a�����I$VAď��w�<ᱦ���>�e��<E��kahޠF�x5�VOR��tE2�S�p��6�4_�t��1�V,S˨B�I�;%����� dFQ�0��_�|B�� p�@ŃG
�vrl���P�kӜC��'3g��*&C��:�<�  �n��C�I(�Ta��ѥS�M�ֵPbzC�	�p���7'����"	Z�BC�	�)�Z�P���=q7XcNЄDB�B䉦�Z� �
��ڭ��ʊ
VUnC�%=,݁%W�V#�$��퉜,g�C�)� �08ԅ�H�~���FƲ|h�h��"O�l��H�	}
���+\�x^,���Qx�����sDP�I�,��W�y�v�.D����닁hh5"p@�N\�u� �(D�|���V6��jrL��3�b��v�'D�X�KZ�<��`����4S2D��p ��8JT�'�dhƤJ�"D��-��(x��e��3d �{c�$D������=-���CPH
�a}�>�GeM#�Ƚ낯��\(�8�"�]g�<!�,M�����R'>l�i��I�ل�Q�=!&�E����5��]�:���'W����@*.��y#�
Ud�E�ȓX� Y�����*����E�$�ȓF� ��%�L�kI�5�QC
��]����x�s���XIT�@��t��A�&�Q��(G������X>>#� ��)f@�!�K� ����&6_P��ȓ��؅ SOPU�q.��T��ȓ9x��{�/�$_�͙p`�!� ��ȓT[.�gh�!?���iPG�@T���	b~��@�oM�Iy�'S6��a�C����y+��UA���pJ�;Y��ٗ�ψ�y�"��Ns��*A�V���c ����y��@
>2�]!B��b�>Ҙ��ȓd��H3`	ߕ}�`�"�>V,����q�I���:��Hz��O=�썆��8h�G��M� �+F⑹T�$��Iz�'MN��k�i1� Y.�|�x�''��y"+D�(I��s�jV�Zd�	�'���Ǥ����,���\�L��	�'��+ׄ�O�>��C��dd���'&8Ij�f�$`�*Q9.D�A	�'���J�*�q�Ā�$@�SU�����$1�S�Ā��]� @S�'�LF(���Ǎ&�y����\q-�r��)K� ؊�X��yb�Q%uƂp �F�p�Q.���yR���d49��& ��A�L��y���! x�T���ΩpFp]�7��&�yk��J��JZ�9<.ш����yB)� �4H�`�:9,�*q�[(�y�U;��t9c�B�)��1Rm	��0?�-O����+J�|�ȧ�45���"O�AZ��I@?�}�d���[���s"O����-L'i{��[G(*{q0�2�"O�-A	ä�0ҁF�Hm����K8��$�J�lD��l�y�=�!D��j8� �3ɝ����w! ��~��HI/�8/d
��&#����d;<O�"<�PJ�b����A��` �QC[�<��o\�3FrX0DL�`�$9E��S�<Qb��X�����5�$�WL�<9����v���i�nP�Ĉ��G�<!�Ɔ�+*=i�&��jE�a�E�<��-|����
S�����~~r�)§i��)(	6p(���\�:�|Y�ȓ.��hi��K
��""��XZ�d��s��a��,��ݡU�A V�$ن�����'�X�3.)Q�-Z�ȓ�@L
Ǌ��갠e��HT���.�~X	sMĉG4�Ы��,�N8�ȓ\�Z�r�@]#N�� d("ׂ����F�WȜ��D���&_p��oF���#�(vD�k��U�Pvz%��S�? ������Cd�[E�Z��QK�"Od�:����]�T�b `�.@}ܵ2�"OV�C�E0&� ��nR�z�y� "O�����?`����k���&"O��sHؖY�F��2k��5� L�"O��[�ȑW�Ry���.l��kS"Ov��%��T��iJ�ĆFp0� "O��I�6=2J�r!*W����"O �%I�ݕ�Ĩ$2Ђ��A�<���BC�(a�"/	^ur�~�<��:;GJ}���F�)���h&��a�<�WbA�M����,S�&���M_�<!R��%L�S0O�'K�*�� \�<Q�eM+�H ���8:f�����Vp�<�e�$,WL|�5�K�{�q�Ƙr�<��-�1ݠ4
T� �NP��X�ɛo�<yե�a`���DA8a2����XW�<i�
8B�.�4�)�$(b�Q�<�`�P�O�2ذ�(��i"0�d�WK�<��	H:6p�A8�"W�FX��ۃ�}�<1�朆>&���N-Y��٫��Na�<�@�H����W�H�I%l�Sd+Pb�<ATjN��E���{����.�[�<٠jH+z*ە�&%o�Av�[M�<�B+�>O���`o��'��0�'��I�<Y ��H1����j��"ǖE�<!�g߅b\9W��D���32/�{�<�e(�F����"�/s&��@P�<�U�B�$��QIQJ�)p�Hm�3��N�<���Ax����M�5!���T�<���N3*���yc���:�~�Y�B�w�<��ʷ_��R�ކOߞ�j���p�<��b&�BQ���G�az�8Bӂ�k�<���za���+i�pLߔ=��1��|8�AF�1���D�L$`Ʉȓ2ov��R���h���{�`8͐�ȓ��a�N>h\��d�	|f �ȓ/��E[��">1�KeM	hYp��ȓ!��X����0Yu3GA$	~}��(�l �G+��ٱ����d��5x�̒p`	�0y�0��d'�P��}rDY�(�*"��C��6-{�ɇ�s��tB����}ctMԻ�(��^դ)2a�0���Q�+�HV���v^ �h"���8�f
JG|����}s�aIflX,�
C��H��U���2��G�	�4�*6�����$�9�'�'*hl*G�G<N�Di�ȓ_Wq����ꁂcI�����ȓsFx��Ũ�/)?r:�
E,�:نȓfA�-+�f�Tg(��c*(0����1�0��S�������&��R�ȓ0�6�pf�=�mC�ŏ�EL֩�ȓ#$���X'B�+(F�LE��h.�1����E�f}@C�H�����ȓ��R�e�;Y��Ի�&[�bdp��\~�b!�2)b�wCӸ�����"�<�6�R�%�lT�1B�<�����.�rX��*Zht\9��4��݅�a��yj�拐G�V�� �&�(��ȓ\��`J�-�.d��\���X�J��̆�<k����%l����) 	�腆ȓ|��YSC�7�f�I�[>W ��./�� w��fi��h`�߳�����S�? ���G�
CZH!��:�Ҡ��"Oh�gM
�S֠�g���7�R�r"O丠C&Ī)�<�6L^
h�Ec"O�Y��"P�;z�Bj\�%�uaC"O�y�:E(�)�Ȉ�V�X�F"O��iWہP�ּ$gM5�P9�"O�����1w[TY����Z��E@�"ON:�@�9���11���@AR'"O�q���,	{�����E�E�>��S"O�9��:l�dub"��4<�d%!T"Oj%XV���Ȗ��SÀ�J�T��"O�JCB� � "(��)� "O�0h�˗�yv�U�"~�4�7"O4��r�/z"
�ꤼ�5"O>����T�q���b&�8#�(�D"O@e����(�H����ޠ��"O�	�� �/��Cr$Ċa��Mɵ"ON��֧�Z�VŘu��l�NШ"Oh݃�&L�G��1W��W�$��"O(�ä��4J9
`�"7[ڑR"ON!a�7v{��A0V�L;���1"O��oԻnB�8u�S�(*8�&"O�PK�N��P�ʝ�e�~dl:"O8%#�	�i
�ka�S�i���C"O�8�-�}���@�^ h3��4"Oޙ�`�f���R��ϐ)&�H�"O؁�� ��fD�婕�\�����"O�Y+���qH8��e�3E���"Oa�A�6:U�ə�%3qR�`p"O��k���Xf��7E��["O�Y���O"�P�`c�7��YP�"OJ�B����v}�:WH���Y�"O��B�ֿI�j"���/|.��"O��� �f]�]�v�I�J���"Oj�[�f܁FH�5��fHM`����"O��ǀцjN��
g�ʞ9zf��0"O��h�d�<+*l�(BC?J����w"Ott@qχ����SD��8�"OȨ�%�P���Ã]�^�hm��"O@T�D	�'LP�$�dI�i�Tpw"ON���o[�H.�uQ�h�8,L���@"O^�Zq��23$h����I-�}c"O�Db��2b���B�2��C"O�Y��ɐw�� ����<�\ s@"O�I# E����"M�B�&d��"O�4�b����U�ЋUe�BI��"O(�a��
-tʜ�5
�8��BU"O�ʲ(K�A<"qW(�s�|l��"O�DI����0��W�̍4{DP3�"OĹ�e��0pt)y��ѝ]��0�"O��  ���ӎh#��u���"�"O������ i� �S%O��!"O,8���$JxP�by".up�"O�P`��T̺���j$��m[r"O�0�Slގ]%L|pTI�����*"O�	%�.v#�  I�2N�`��p"O�u1���n�x��k��2�"O��\(��e
�$�����"O�`�Á�
�a��b��iT�;�"O�\��� ߐ�;�]�+�� ��"OY��$��'R�@�ھ��ͫ2"OX�01C[�W�ܐ�e�go�@��"O�q1K$Z*�]���ա,��z�"Ov��f�
�n�޽��.G��7"O� b��������=aGdܶ҉pq"O6tI��Y�Ƙ�d��JF"O��2D��\��փ;<*�D�"Oމ���~x��#ԝ��	"O��*v��;����C�Vj�z6"Oй���A&Wʦ=(��S�fZH9�"O}13b�-b��D��%��=��8�#"O�l��T�a&���#�S�$�1"On4�B#�Q�I�C�12�p���"O�I1c�<9��=I�IJ~)y�"O�\�g�ՐJ�0�Q��5=�lCg"Ol���̟�P���Ħ@=-PqK�"OB`���X�(�
yR��	^v��A"O�hG� !��㤡� 㶑Q�"ON(`��у}�bi*c��+r%�p"OBh
ϔ/ª�9!i^�j�0"O���sH=[ot���F?´�s"O�q���%`�ҹ -ÝGK�|��"O������Z�}����.HAj5"OH$��G�5��1��ǔ&0����"O��(���77Z��`�٣^"��S�"O�l�&�B�'���Ш�N�8�"O<}�5�ܢf��q!�����yb� -����<�ف��yr+�`N��ˀ4��� F� ��y��މ�2DC���:'��h�(��y2ȏ��2m��(�
�y�a\��y�j�Cgu"q!X�0��@�Þ�yBbU-'"T`�'V���"ƃ�y��E>}��Y��?�R� � Ǳ�y򊌎2��T8����m[���fg��y2.E�jl��i ��:f��9F-@��y��V�5�FB�v��� ¯�yҨ�.|/�(��ԃN�!�V��y�K� �>�*���TQRRoY��y"� �H(&Q����lE7��=�y�ڍvGb����y���)��y�`�r9<��uEE���7��"�y�E�pt�$�ӫP=C�Z�2���y�"�!#	��bw�35=U�W��1�y�k*��s��B0���(�ڳ�y�n�9F@�N�oZ��h�-�y2�4>]r��㡋��4���B�y� �Dܜ���mn��H�D�_:�y"n���.m��B^s~���N>�y"��"(N�tPs�ؘ"�$ؙƊD�y�Ā<ve������9c���yנq���k�3!�l���:�y� <�2���`���f��0���y��B�p�p!�a�Ǳ#�����y"�@%-*�a� %�V� 0�E�yb��\�$�Cn�'[xX�����yB��,J
�i�sIh���Z$�O��yBo5Z�v�c���"s�y�E��yR+U
���U��Y&ȭ:`�
��yh�%*��K$J�&O�8LP��(�y2�B�JT0)���A����L0�y�Q�d��d`�-@@��Y�fc	��y*��:���4�;^�9�5%�9�yR͐xa��CX388�m�7nE�y�+Q�^~�!�@ӇF��*����yB��
Xs��q�;S��p	'�\��y�>�yQ�[J���ȕ���y�뛅{E��'MQ�I�����B�y
� �P���Uw��t�ޅsk�1�b"O,��Td�@��\�Z+_T�=*V"O�A�`��3PN���&Au:@�;V"O��*'�^�Y�F2�~��-k7"O�홁�V&wNz��D֞T�  `"O`�x� �>�
��tnګ1~j�9�"O�Apׯ�w�V
�M��WZ�ɥ"O�%jR�D*Ih2<qgǝ�Q!^i�G"O��T��
�\��%����U"O�	��N�[We�+%�8�"O���E�ڑu�����@�<�8P"O\�$G�N�d�)s�Wkݒm�'"O�UN8x��u�2d�&1t��"OL��4��1z�"�ɓx�Jٶ"O�x�B�ܧZŎ�����C`Q�E"O8�í��o�-1V�ֹ�V�� "O.8#�P9���R��~%��"Oh�"��Rb�f��#�=��<y"ON R$R%�P�Cۆ!��(�"O�J���b�|�Շ
�W�D�R�"OI�!L*8�y��Ȁ|�l�;'"Oa�a�Փ,p���ۉ���6"O�!���9b�� 	�&�,jR8�"OB�X�g܌|����%���L(�"O��o�#z+����B��"OzY�Ш7=�[!�EV��"O�-�殈�V�3���&�t�"O���mU�3��a�E���y2� *>����\���3�-�y"�1zR����~Ȫ�B^��y"I$u h��y�Ru[WO��yrJD��u�R��&z�p*�H=�y�a�bQ4<��)��w4b$��B��y��	�<0�L��X���Q�č�y�	[�bs�p�q�����p�Ǔ0�y�#�!^�
��N�n{�u{eDσ�yR�P�
qi�H)r���t�[�y�e��O0~T"���.nX�U��ɦ�y2��n5h庰L�[6Z\�UG�*�y�K_>r&�T(ӍR��H���*�y��B+C�$=�7n�4C��)���+�y��i휸2�C�@5�!Sd���y"c��։�U�T�3���(��U��y�K!P>��LW�+�h�����4�y"��w�&T�C����m��oG��y���[�8m)�o���,mk�^5�y�#�h�����y0�#!�Я�y�N�(�<q�:�^�:3��:�y"��Q���C�9�
�3G���y��8�R�yäړ@xzݠ�jP��y�
�- �ے�W�%�8�� U0�yR�	�=�\�2��[,*�d �m��yh�!�͈�* $\��,��iۖ�y�cP�Z�ց��A�U�ⅉf�J��y�.�(����"2�����D��y���.d	�-���Y�r�~I�5�ާ�ybfW<8O�����<Tvx��y�+�bVD#W��2`z>Y��c��y���x�:�j��/���k�����y�&_@Aڀ��O��"�`�ZՈÁ�yb�Đq�(+�'��>�Д���y��)������\.�.Th��Ҷ�ybHq������8;d}��cK,�y�M�ygZ�`r� }�e�_�y
� ��Ef�:4OJe rj���+""O���u��r��苐��� >(ER'"O�E�bԚEK�|��i�'/t�&"O �����M�z��,�P"O04�1���]����Agʉ [!�C70B޸{�"8j���[��?i7!򄌹do^q
t@%�$B���V@!����Q��!��{c��H�!�DBW}�����3c���@��
�%>!�dʴD�Ta3Cg6	��P�'Bo1!�DE.,��p$@%:�0ٖ�݈K!���ll�Q�׭�2&��@0�K#!�dמde�0�������sjO��!򄄎/=��U�fnn�H�h��!�� �T��)�YB}�ag�q!�$W�C����䍊0vD��1 恝1g!�$ "�0��4��=*���0*Z�sf!�
�|H|��T�'4�@��!�d�<��	���	+DżIʒ-Q-J�!�Ğ	s����W{�*t��m�.M�!��Ξ^O�q�a��B�lbE�H�d�!��3���*`�ޖ\:x���]�!�D�<-ɪ}22�F�i�`�\�X�!�	8��Ό��8�����8[�!�DY���=�a� 	��&a�Q�!�Q-
���q�^�Vd�Y���!�䝽h�֬���M�1i�У&�!�dK<��@��R0#
�p�T�g�!�̝
	(}i��t�� :�	�R�!�DZ&n`��I ���� i��!�$Ƕc�����B{� ��St!��ƿr�č �@� �^=Y�Ɠ� i!�-K�`�NQ�'���Y�F'j!��Z@��+I}���s@�]�!�ӿndRC��ڭxf����� d!����A�d�Ā�qa�_��T�ȓv��I"�ƎP~r�����!�$������Ug�!c�d;�ɟ���P��C&�]⡍C�a�*|r��,)���ȓ/��!�U̤H����]�9���ȓ4�z%94�϶f�@$��CY"I�l���Vo<�XbbI�	��T#Q��$��Ą�Q�Xp�ҫJ�u=��tD�}���6~PxK��Ӫ,��� ���87Nl���K�d��#Ł�0& ����<��a�ȓg^إ�PΊ)R����b�ۿO�X���� ��+��o���HԠ�`oޅ�ȓ3S��sGJH<!ޅ�֭�m�(Մ�*��X��E�9@��KNلȓ*�H1!FB �9�p�Xv�M�ȓN���̈^o~�gτ;7Ax�ȓH�D�ڀ�D�x~�Q�@��\�\��%��	w���)&��	�P����N���˱,5$��e(i ����R�6���Шb�� ת��?�0q�ȓZTK%��;[�j4Y%"U� BK:D�TH�*p����T-�+͕���y�!�4�d�q�J�=dֆp���E��y��
&n
�9`�Ah�r-�S��yBꐲs ƅ���5V�\���P��ybn�$p1�!���1Id ��eF�y�I�
+�e����6A�Hv�y�cѐ�p&K��X�R}�6���y�aX��!�t�"��C�>�y
� �Q�7
�
>G���qc��<��"O2�p�������AAԮ~�fK�"OtY�U�R�pj�I�.=zڹ�7"OZ�{��=~z�@@7��6|h����"O蛕o�	�a�d �*niZ�P"O�͎wǾ�
�$$t}�}I�"O�*�(��
��9�A��Qf�(�*O� F
^�F̀Y��DG�%�J���'F���q�2C�|�ER'k:�*�'��Y�^��A�$k5�'k�)Cd��v٣��f����'�@q�k����(�X��pR�'z�}���9�vtz7�U�fR�k�'�ݳ�e��T�)b�ƛZ��x��'0`�4	:~�Z2T�G�ZM�� �'a>�D�]vj�[4�E3ID��i�'�f�iC�M�n�Ղs�V:Q��s	�'6�8hL�1|�4x�!�	G#�E8	�'�ݚ�E�[�L�`�V6t}`�'������žy���y#ME�B�q�	�'CN�)1F�a� ��ʃf`TxA	�'#�l G��G7N}p�+��I#F�h	�'�zA�7@�0r�VD�򌎵?�I	�'ش�#���x�
���9�aG�<�1k�#ǲPc��x���%�G�<)�jL5�e����3u��ci�<)'&9���+Ģ-��f�<��L^y
��Q��$X�*��t�V]�<Y�I9dL
� ��`Er�`E�V�<��AK�|i�U�"ΞI���� �Q�<��ȴ �L�a@]�P�"0�N�<�6�&-� ]�⭚03��Mc1�K�<�W�"�\�b��&Ԃ��II�<�2v�b�� �\��`�H�<Q�˜d�����>� ���D�<1�l����jwȝ��� I�KV�<�ҁ�d�Ny"�
9q$�Y�@fSF�<q�`�Sg�8!p� p�d�E�<Q	26R�aW��6g������e�<�E�$�H2$��]�{"Kd�<�#�=UI���1'�
h�5�Uk�<�$�0	�l�I���\�����JFe�<�1Í�{W4ݺ�| ��b���h�<٢O�:{� 9a1��p,a�E!�o�<�vJ̈́k|�l��h׻/1���1G[l�<���[��� p�:T�xS��O�<1B@�C��s��9.,�Tʅt�<�W��r�(�DH�x��d��h�<��-2bh��bƬf3Zm�BF�d�<Y6H�;[��Q��T�7�i �,Xa�<A�"�u�!C(l�mR�W�<��!��b�>�����M�'HV�<�U� "o�I���	Ì��'�N�<��D@����P�fR�*�#�I�<�g͋4l�h՚Q%��4����u�M�<Y��.?dp��,^M�Z�@k�K�<!f�ōXq����su�a���R�<�ʝ1SfX���F?Oc�����O�<i�ϝ=O��Їd�9; �QC�D�<�Ď��5ɂ���H2��`BajTC�<�L���tY�u�_�B*�	�Ci�<��l����Ƭ:�	P+Nh�<���>��[0���V<H$�d��a�<�!���B��u�J�e���ka�<� *}8 @��>�`0�ͺ2o(Z�"O����ʕ'=L�� ̹WY�l��"O�ӣ%u^�R���h��ɷ"O�P�7�۞K��Jbn�03-2�"O
��J *�T�@ W%,:h�"O���q,62�jd�u�!v(jP�1"O��*2�G*�A��+���yg"OvTk3BW�U��I� Hū2E�d"O�,���,b��S�DF04
�:�"O8�z��0e0�pv�_�^�k�'�ʔ�c"�;K@��`H]�����'��4�3�1[}�MPЌ��z0ָ�'L-S���t�D�CCXq�'�����-BF��Y�n�S�8���'��d(���
hp�1�;;�V�S�'o�(@hT�$�2���*
�]�(Q��'&h��4x0Q@��J�\r���'`:��p�?8�AЂN�)\`�'[�Q����fᤨS��HUf���'���kS�������>?�
q��'�Ȩ��L�WN ��6B	/<46���'p}Pr	�ݲsu�E������'� S%At���DX�
 `8�'Ô9@��
�G!6L9tO��| 9�'�qa�WG�@��Ҋ�n����
�'|�xT��;��u8Bmݗ_��k
�'�6	�`C'V���Ѥ�X����	�'�����Gד6�l}��̈�[��	�'��ѵh��7m�m� o) �l	�'����@� &HP'�=2�"���'�^�²�QH����@(
j0J�'M��)u��*D�UZ�K�P ��{�'S�x j�?U��{ED���:�'dR;F���$8��pJ�aw��r�'W��;�����0*��ZF.�h�'��ش��d9JeٮYL����'��3��R({�䄌N40p0�'�VD#�"G�sZ��s��N��@��'����T�%~z�aKV��Hl��'�j-rl[0�$�h���;쁠�'a6�i.o��;V�œF�vd��'~�ܒd�G@�L���(f��'N ��A��k��P�G�:��1	�'S*��f�+�d����1+�����'�L�۱e��,h!�A��s2����'��CN�>'�Q�M�<ɲX��' ���-�¹B�Ią7��9��'��AX1�Z�![��B'"1�*T��'��)P Y�-'Є	Q�� 1۠�J	�'��8I��J���\���)Ẩ+	�'��$"�v�zAaM���p��'��!�%j;�E9���#����'��i	a�Gq~X)��hY�\2	�'�JL�!lF�P���1oƨ� E��'<$���NW�Y!B�q�6^��P�'#Х[ӧM�c. ��ᅇ���!�
�'\�=��-�ri���Tl�?x�ʸB
�'�Iav�,j}�ԇ�t'���	�'q��EMͦE�Ԙ	��Z�}��h	�'�J�PtF-vF$�S��|.J���'>+s��r���k#�x����'��6�V�7^��*���u{j��'�y�6�W�3�	 "f�d�c�'1�8z@�G�9�Љӑ�>1�& I��� @�S)�eU�a���7�Z0
�"O�Y���T"i�� b�8o8Y�u"O���D�o#�dS���Z:@�{2"O���"a[�yH�A��#H2^UBe"O�qd��< ���Q�f1��Kq"OJ<H���6�x@� ��L7b�8"O�������<�@����怒r"O��y���d�౳vFŭ)n�T"ON8��\�8��r���h��!�"O�qХ$�>XR�@$�
�`�h�"O�}��§%�6R�b"�4,C�"O�ܑ��#
iVE[� ���z�"OZ�[�e�5yu�l���Hn�j�"O��R6)��=`
9AA۾4r
���"O>@�W�Ɔ`�أ�4rl:�"O(���5��l���<iV���"O�,{qH!?D������0͊�"O�̅Y�Xt�\P��໖"O�|エߌH��oC6~ז�H�"O��1n�+j����.�.d��;�"O�!S�A�܈��-��}4^4
"OT�@�/״z�JprClzXB��:�y��t�%)�FޠF�4�cqƟ�yrL �;�r�� *�9;庤� �T:�y�ŸR�"1�ʪI`Z}�����y2��X�`��!3�px$m�y2��y#M1wY{��p����:�y�%��=�m�瑔��h�#,���y�I�{XM�B�@'�(���?�y2�ڈa�����a
;	�\iӨ��y�)Tm?8��$��� �#n���y�m��ȣL��e[�i���Y�yr!Rp�,��gӮd��� a����y�KM&9*�B�)B�^߆� ��(�y���=��:��'����2�yb��]qP�X��U�+��`XA �y+̠]��7m�7rU�d�S%F/�y���]NԘ��Ř~-��
�#U:�y��Q�U4�3͜�"�ec�i�)�y�#
���VL�-p�8Z@i!�yRB�/5��Z5��\��qb͆>�y�m�	�jD�q��Pe���yl�9I�@1F�#%R$�2�#�:�y��?I�����I�0e֊�y�bN/�6IQ�mH'?6x��ֈ��y���.DY�<�lN�2�Y�A��y� ʐtK��T�Y���؀ ��y���)J��A��G�D>|z�Om�<9�n�*��(���"}(x �Q��k�<���3h:4�,@%�x�S�,�L�<�qj	{�b����KA$�F�<�鏉-��y��G�9�0���<1C���H�@� N�v�XU c��{�<1J�#p�8�BD9|�p�[�t�<���Kq�qi�L2a��-�G̏[�<�ff_$Xv��E�%� ͓o�<1����-p ���$��n�<��&ݖ UP��{O����k�<�"��f�* ��D�l<^��I�d�<�/�@Jua���q�H�a�a�<���Z��2���O��I�a`�<)�O���(�NId%�(��̙]�<YN�;��9�ѥW [S�a����Q�<YC�ǼԚ�#�:Uɾe�mQ�<� �!���ɼB:B=�M��lhq��"O�4`̑���G��0$��"O	Uc$!��t!ۣY�LгD"O8]YC�K?(5K�@��  Hb"Ov��h�k	\��RoJ�u�č� "O���сE$'z,�֮��	�q��"O�x��E�~H ���l��]`"O֭���X�^4�E�]-
H(d"O��R#�Ze�����X:�ѱ"O^�ZuOZ�G+�,0@�(]P�tp�"O*t84��
Q�X�g�M*� �"O>��A�&KZ,��ޅD��Qv"O`����&A��E�>:� {"Oΐ�HȏQRЀ6Iҗ>*~�aq"Ov��D�2'��b��i%65s&"Ofl؆�C'yZ��Y IƧ(��"Ot�`�!ފJ6T��_�D�0�"O ��K�(�nU���^�ܑ�"O~��#)L)D�)�I"F�Pyx�"OD�xo��b��DgD9z�%��"O�Z���*���c��c����t"O�����U�������g(��b�"O�1���T�4����W�V�<{�و4"O���D�{���U/(Y=z��%"O���ĕ.1Yh�)��h �U�"O���rc��j Sc�L�X�&ܳ�"O�Ţ��T�6WZ�`'�"��is7"O
��1�C�(��2DN7(u��ä"O
!���	Ҷ��4�T'|VJ�0u"O�3�d)U,�,f�<2�x�"O�M[�(��w�e�Q����ZQ"OX+�ϊ;u@�r�&D;mAz���"O�0�� ��:��H�Z�".l$[�"Oୡ��c�6�Y���)+>h��"O���Lҗ$�������$}����"O*t�S�Osx��zvi�6Ama9v"O�$!��M��a�-_ڠb1"O��۵mF�kd}�V�P�8�d@�"O��8a,wߢ5����tN���"OH�2%�Z��SoC�.1R�pC"OV��&F ����H߽*n�a�"O�S��V%1�ʰZ��̎!�F�AG"O�d1��ռQk*����Z�:0�"O�I� ����'�>F�x1��"O6\P�a�9���J �9�<�S�"Op�фΟE	5듋H;��p"O��CU��/ܼ��b��?Z�N8�"Oj4{f�_/��R��6�<Yr�A�`�<����)'8B��� �|����mC�<9�m^�B\���Q�V�D}I�EZ�<��A�)����oД�:�m�T�<��i��e�d˖���A4��H�Z�<�V)�g�4T�g��/[v��`EV�<����=���e��,��-�\�<Y��ڢ(��m�({h��gH�_�<��
�LSv��C���kH�Y�<� L��:I�J��ǣo�����Pj�<)pj��[?D�w�ۺ!F�� ��_c�<�aW�o�]R�Y8RaØS�NC剷C�̀�7H�!���9��3w�!�ma��mI�^�"����!���.�����#�%����v+5"!�d��|:�J�i 1*L�A"
/!��B�����/[Z83'�0H�!�� ��{W��;�~=�U�=v�$�"V"Ot�M��v~tD��V�X���Ç"OP%��l�?5>v�U��w��p��"OT��A��?V�i#ŚTt�C�"O~q3��)�"��!d�7��T"OJq��S�p�N��EI�x��P"O81�eF���A���s��8��"O�����/q) �T������Y�"O���L�O�Z�"$��P|.ب�"O4I+ï��M�<$�A�; A�"O���S�-#��	����?�h �"ODɈ�hH HY�5x��{�6|	�"Od�&�Gj�@�OG=����"Or�sqЭ�D�+���.���q�"Ov�.����C#��^+(�Vb�;�yr'M8{�,sp���S�H��%�[��y"eϊX�Vi��$![�`0�R�y��#�)B ��"W��`��ݖ�yB�֛} *]�u�����Y���4�y�d����pp3�
0hz̛&.���y����el  ��_��0:����y��)F���Cw��VH��+���y"�Me4q������eb���y��Y�g9���Sb{�Az� ��y�`���y`�
�CaN1DL��yRg�1d��c4��$B�����]��y"+�3�ݳf
L�2�؄�C�3�y�$�1J�t鲄�Q�a%�d���`�<�W<<�L+ �4D�戨��EC�<ɡR	�����E,Y���0�h�<q��=[ʚ��/G�K�F���v�<!���l���r`���>H��w�f�<�C�ә.Ƣ���N�z���a�Xn�<�G�N�5�0�q�5]��Pi "j�<Q��I!R ʶ�Ԯ)�z��q�<�&/�9&m�a�mŮ{�B�p�AIj�<��fΧXך�A��4+�0���p�<��挗^�Ұy"�@�v�&�J�*Hk�<�Ӫ�.3|�)��\�.��1(	s�<�FaN�$�T��������J�<	@,D �$QC���]J{`dD�<)�lޝ��HB슺(\@�BqC�G�<�S�2\!�e��:�p���O�<i��-O�=�A�ߍQ��+�WK�<�$HQ��̹p�ǜ��<�����J�<)P�E�RE�󪒎N�|��b�H�<I$l�)`:��c�n�^z��l�L�<�¥ �TϮɹ��Ѽp U�p�<At&
: L`iH�o�7{���S�t�<aI�EH���"�1zr�s�	Cs�<UG6���&i�� H2�3�-J�<q "T}f�p�Z��0$��&_�<�A,>�N=2�O��N >Ě2j�F�<�����|�nY�CW�ZWd`����F�<iRM�$ԤS�o��s�rg%�]�<�V��`0p���K&�J�!��RC�<q�鈀S���w������`]}�<�PN�({�j 0��G�Rer6�y�<�P��E�9I #ǚ�,�h$�]a�<����%%����j�������H�<�ޚ_)��S���f!!O�\�<QC�Ֆd^v�(G����	���Z�<�a�!��}Zb��g��IP�ȃN�<�L��Lr�#G�t�P�!$�D�<� H�@`a�nq�p���н��"O|��2�B,9�0cFh�̆��@"Oڔ�a�T�|�R@��$�h�mk�"O��{�d'l���7�]�z�&u"O��0"�$�8HuET�v��"O
9Q���2����U�]-9c��e"O��[��>�ڰ�t�^�L����"O"Ԙ@l��^FNԉ�B�#���"Oν�`S�@�����G!|����"O��0@^=n{�YG���*���Z"O�Tpg�ƫh����F&I��� �"OTЁ��֞�"�p6Ŕ7,b@�"O�e��0u�\�����-/�+�"O�5�2��T��%���զ;f���v"Oh\�Sd$�n�u���i�~�Rs"O|�(�9����#Cz�~�p2"O��s�	[�`|����Is�9R�"O�yr�Q�A�09�CD�8s�hQt"OJ�4�@��IX���O�� #V"O4q��KZ����3���z���i"OF�3�Mۗb� x(!��!����"O�!3d��! ��PA���u�1�u"O>�mҏj+��[�ꚫ:r�e	S"O��W3r@^�:F��/LR��t"O���įA;� P��XN����"O�)��D��)f��)�c�!XZX��"O�8��N4qB  )�;'?.<R�"Oԉ��F�0`G����	[�i2��b""O,U�@�ѳ��J�).17b\h�"O��+�qfΤ���Y�H�A	"O2�;si�c�\
��J�anBDU"O^@Q`_�$R�q��Պ	n�q��"O0QQ�NR��<Q$�	l[~�C&"O�`@���?��P�	�HB֠� "O�;�� =S�Փ1��
)�"O��䨙�C�${ �w�&!��"O�4�Aoڮ|\0x�u� �l�"O,����ւ.���T���@��8�"O؍�vM�C�N�����5ެ	ڐ"O�9�k�%��`��� ��"O�`f���-��Aa�ΐ�Z��a	�'8���3 ���
 N�����'BX!�e�� X����S�§g�$���'��*�I`~Aa���/I��	�'<�wM>[juJ��4R����'�xћӄ��VT���&�TA��'�b�@��j`�dH�m�>�&���'�x����*!ed�W&�-�!Z	�'bi�#D�+�z�����Љ��'���i����C�*<�r��	�'S�A�Ej�>�@���O�9>@b	�' 4 ��@ʳ=���P�U/[��!��'됐uAM*{�q�p#%U��9�'��UX5�U>8P�S���->����'�� Hs���J�(i�K	�3�R�+�'�� ���̨A4ȁ�2�`��	�'e"=��$H�GC: ���P�YD}y	�'20ݡ�Ɍ
Y��pP�V����	�'1��J�ڹ-��X%�mU��S	�'�4t��X�G��eC,^Q�4�'�~�e��⠤�5 ��W��[�'�F-� ���0pB�`��M�^lj
�'b�10��Y�8�����@�(P
�'��M��m�.(j��&�I(?	���	��� \Qa�Y�2(�����ƶ[Ǵ�xv"O��Cc�U�pof!�I�Q�.�Yg"O�K0n��)�4���j���"O����+��H�'��ew�}�"Ob����}�bDA!mEk\�\ �"OP9�4��){0� ��QxLU�"O Y�@��>	ثK^�LwPk�"O�幁�x�����Pl-2�"O�3�Ĉ�PL�0�B��&]^�$"OJ�{���� �5��Y<�!�W"O����OC�}�d�����-�rF"O�Lv	�U�!�FN��t&���"OHȀdLX=���&�Uc|�E"O$|�����~ ��ʯx�m�"O��@ƤZ�'l4���]1F�L��"O:�)eӜ"t	1�K3D�ET"OH��Q#I�b�P�@H)�>�"O>��1�/d�(�c�ĉ!Wv�k�"O�uk�Ԯ�p��"�P�U��"O� a�_�+�:�ʡb́8�"O�k6 �	',���B?`�z=��"Ol�C�P0#V2Mɠ�T�'�Ҍ�"ORpٳ`��m8X�pEЍ~�,�� "OR�`�CP�ݱƤMq�6���"OR�����Sj�����I�w�Iz�"O����� �`D��KشV����!"OE�����L���7NZŚ�"O̼����Wg������#5V�8S"Op�c+?DNaq�+� _T��6"OB�E��35���=^�����"O:]
`���~u�d�MƧ3��H�"O�90SF��|�&,�f��/v���B"O�AdA�oRƼ�F�A>8���"O��׊��p�򽓒k�':�p�B"O4� �`��qL���ܵC�0t��"O��Jm�+��x�����V����"OT�� ��9_�\�����ev��Pv"O����5'6��Sb'ܷz~���"O8��Ul��]�dc�EK7M��"OP����O{�ԥ�	�����5"O|���60�����gQ/#�z8�"Oܐ(��;�*��-C�%���+�"O�x�L�2@����W����A�"O��$ꕸ{N�Qc5�{l�%0&"O@�ւ[:?m���A�5]/`=+�"O<�@B7x|:x��2x&L���"Or�R�̙{̰�8�OJqz�c"O����̈�s4������,@��1��"O��r��&�ST�ј���b�"Ol��5d�2.z^yX��=]v�2C"O64J0�șn)5	�
�%L` 6"O�dD"DӚ$�2HK�e�0}��"OV����M3�����ln}@�"O{�m<vD\��!E tr���"O11��*,.��PČ3O��P�"O��)4,єYH ���!�L�޴(1"O�B�E��8���`�k��0�5"O���Y�M|$��a��V,�$� "O�h$!�D���m����U"O����c�IZ��@�"�ȇ"O�k�ƚ�~l��&��y��4q�"O�,��߄gq��QvC #7& d"Oꝑí��E�Y0���5w	At"OF-`���[Q���%�+Vl��"O�  �R`�>w,�ذ�	*�S�"O�1��Δ�N`��NI'E�Zt�"O�5�S�\�<��BC`�6�"B"O>	3 �T�|���h���m��G"O���P��x��u��E�,��D&"O ��Ah3)����m�:{%6Lrd"O�|�e��)Bh�sbЅ`�58�"O6�a�ܱ�� 頇�&4@�"O��i�L��K�,��R턊|��"OBuS �x6�Ȼ�����Z'"O��{t��`��Հ�M]�V���X "O�q8��L�|�+��P>�4[&"Ob�#�,u)��aJ�>���"O��H�	"�Bp��?}�|5"O�8�0��9B��	�b��k���"Ov}j4�X jMq��>�:�"�"O���$v(�DV�ڋ ��<�"O��xӋ�']�>���j܎;�0 �"O��P1 E=J��Yw��t\@"O�UX4���aU$i��f3"�Uc�"O΅��g>���ޢ!^�(D"O
���	�^��i�mJ�.d{6"O�az�.��xt9�P��tk"O�ՠ��ʿhU�����D'v�۶"O �c�'�7w|(5�C�QT�0q"O�A�0	Q+]����,�&p�;�"O�Mi6$�T�Gj\c���"O�	�W�4���Ô���"�"O8�j�/�g�6l���$U�Jx`P"O��33�Y�e���"��K� ȑ"OP�#��~) �Y�^;Xߐ�y�"ON)pVnƊ[ʖ�ʶ�ɿB�HmK"O�hZ��ae�Z�r��&X4Z�!�D�c��4*��r/nͺ��:y�!�$�y��4�2�J�@�	�$� w�!�
������'|�8��/�!�$Z�p�Ȩ��H��]�܉`�D�!�DX9 ���l���){#`S�-2!�٨zE�$���0|$��u%��(!�* �80�Mǁ���B2$�
+!�P/Do*��Ξ��(�h�b<p,!� u�ѹ�	��d�R����.`!�$̬(��0�m�$q�����&,�!�bn�4�PW"VB�
s���~�!��V�^<�-:D�A�b?"d��R++�!�[�Bf@Kk�T��cD���!�T>8(y��]�
���Yvm�04!���&R��	qE��/�RIрk�$V:!�٠�
�B5��c�<	W�_����ęv�.�`ի��F!�ms"�Q6�y�c[��<���F�M�򤃐��y�+G�}�r�cq�v���H5
�:�ygö5�����ܬE�6�z���yr��7=��ACf���:���G�yR�U�'l�D�qn�~Q\	r.�%�y��U�$���k��ye=�L��y�̗&\�JT*�
�o.�UK���y�偫>��H ���`N|��E ��yBY4J�Ɯ!wJ�Y�BI�DK���y��E�)l]p��; �� Bd��y"�TΎ��)�<��p�؞�yr�N�pO����ĩ�,
@K��y���S�F�+�A�#|�Z�0�� �y��T�;5L�'���E�Z��y
� Zc�Сj%� N��S}Z��"O�غ��P��xx��V�^�v���"OX��C����*1�oX�,]N��"O�ڒ'%3�xJ�J3J.�+�"O:IX�� ag�:UK,4Pd��0"O${B�.v�a8@, �3����"O�d�5��N{Fib�� j��U�!"O2���)�2G�Q�@���@h^�
"Od�D�@U_���m�*[.�*7"O��S�MC�3��Cb	83z���"On���k50U������i^}"OT��Ѐ�Y�"��������"OV��fHA��*ê�q �9�b"Oi8��@�;|�aK�	��V�B�!6"O�98�-&5�����d�|��c"O�y��iU�l�� ��;gpx��"O���(�;P+^�kƕ[E�I
0"O����fWo��M��T&W�ex"OP�Z� �� ��(�A�܉B9ڼ��"O���N"� <�DE�o+䘘�"O�c�1T1v�+�%��>7�| v"OH\��X^U^r��ܗo�(��g"ON͈Ԏ�?cHD�R�)<eia�"OZ��B�p֦��F͟\�]�a"O�/�O�����LU)<V sc"O��A��>g�>8bw���8Be� "O��J���(m�q���U���H&"Oސ����*MD�HeJh���+�"O@ "!�G(`9��ڇl��X���"O،	s�3+?4����j�d�'�Q�,G!�p�P&(H�|��`��]�<��)�^�
��!a�D���#H~�<!��J|۾���	��C����!��{�<��!� � xjwǓ�5+�q8�/�u�<�+r��Kg�H�d�^��7�BG�<Is�}%��{D�.5�Ĵ7�MA�<�2��L
 ꧨ�� � I3q��u�'d�yҁ�M����`��,i�p�C�	�y"��]u�Q�6�
�N���`Y�Of��Ry�DFz��q�%(�M��T�vCV$4B䉫bBB�CL��<;�#UXB�X1�D{��(!�ZYK3N�M�C�I�?�v���k�6\�2��%AN�L�C�əS�ܩ�"A3ٲ���*@�
@�=��{����)���X%i�lxh�A�j���y��ω`��5�rBԳ7WJM6(\�?1���S0	A�@�� @�g_�h��+'Nv�ȓ����="�D�3�GѨnSlLЈ��s�ԺaV�m����#]�G�X��Ql!D�xP�̷h�@�q�ZW*����F+D�| �J�!ܨ�W�&!�Tl�q���hO����J� d�'΄+p��Q3�4f�H�ȓ̖�S�d�&7��Q�)�1����?ф�B�=aV�3v;�*qjNf�<��i�i�&h�#CƳ���3��`�<YU��݊2�*R�p-����0�!�U8̘�k1S���C�.&�!�D �v����T�;+����fJ��!��!uzb�B ���g�ظ��L�!���	$f<���z�D�qT%� ��D�TA�?���asl��r�ܠ#I�"�yҏ�)n>�Ȉ  �7iFb�s�"�y[?�i��.V�f��%�%b�'�x�'K��9��[�Ty�9�ł�#z�P��� Tewc��J{��4�A�j�Q+��'�1On�9�/��i�zT���ּ/H4,��"O�9C�O�2$f�Br�X�7C��*@�>q���	���nL�I8cŐIhEa_�l�џH����O�H�p��[�N�y�չ�< ��N1�	q؞hQlH�_�m�Fl�<h���P/�<��'��舟����ַG)^u�Qg]>Z�|�"O���̺$�$�y���uժ)� \��	O��O�4��P�>�5"��E���cA"Op�Q��Lˊ��`ܺQ�X�"O$�Tj��Q��)�A@�(�����"O�l�7�@�q�~�˂��1���9E"O`a(�)Lw�~�8Eiz���{�"O���"(��BD��{�'	"���0�"O�U�rhD�;�-�c&�	mh-��'|j��	H�
+�I�3��5 � ���&��	E�Ȇ��џȒ2(���>��d-��<�0�'�޷�y򧔚J� 52���91L�dj���=�y�	�a8�j����%8 ��5�#��	Zy�5O.�~�/ɐAd��֨��I��}2�YV�^���<�|ғ�_"?/���Ư	F���A!Q=�ў"~�	�}6Р��gta�,N�2����C�O�ڠ�Q �&59��F�9Zey�"O��C�G2T�1�4�	E_(M�OZ�=�OǛ0O�� ���%??`��gQH���"O@���2�NY0�'�_B�A�w�|�'��_}�Y���0٘����;��8�K�'2؃�+�9%+bC�ɞ[�Z� pH�_���0n�=D�(��'�ў"~�g Զ4 �p�b�~���!¢�m�'�RJ"ғmτl# 	�!w������	 ĒN>���b\��B)�b�CRNƥ^��U�O��	Z��J�Oo8���ŕH"h�� ��B�D�	�'M6]P`a�+a��h�̘�z<ϓ��$�O��S��{ҎY�]� ��n��S�IR"���y"�[��D�CXx�æ��yl�i}����K B���%B��>!O�����!zp�"ǬQ�6�	��.D�Ѓw� �(d�p�R�l� ���OX$���V�����/ug^���M�������/��+b4ã�	g���!iܱW�J��'��~���V)a���i�!v����'�ў��<�@C5@}K�Ϥ)O�<��s�<A'D�L���E��\�R!2���u�'w?	�eN��v�"�2�É�n��#��6�Q������E�b	z5�	�F�,��5�O��0Q����ڷm�Ĩ�#=@e�ȓC�*�A�N�{o�@�gO7�F}��S�0S0S��^�^Dݑ��K)n�.B����h#�B�w%鳠3JVB�/gq�D:��E"~q#'�;pg�C�ɼ]����1��%Ϭɢ3�H�eL�C�	kw�`���pϜy�G�Sɡ�d˂iy�M�"��T� t���N�!�T9:��ݐe/�l��E�:i�!�D�W89G/����ED^�L-!�$�$I�� 2��#? ��$C�0MTB��<n��s�F�*�����PY"?��(�"�!rB��S-mi0+��Q�"Oz�)w�_;u���j�& �-��IX?I���S]�( �ͣ/�
���ƧZ�!��5)c"�y�,ܑ+r��*�F���O�=E���Bkl=�d�H�y�D�	5f��y��Q�
1re�ۻ:N��Ht�G��yN�,z��xuă
9]�< ��S�p=Q�{�� Xy"�GG�c8����ױ�dii�"O8��b�+,j$�yD䔌U��!�"O��g)S�rk4��b(O�(��A�W"O�e�s�U9EN� SH�d�&�9b�M���	P�> �QQ�^�zod1�W��[n!�D�i*xr��b���#R!򄁱h���g��A��!`���!򤅰�2�iu/��5�D��aUU�$1�O�}�5 !w�����HZg�'�'j���p���u��aW�NZ�P��':�0x�V� ���z��%o���B�'�$�C#�!s�<�b��3~p�8�'���%����K9hJR�RsN�\�����d�2p>�@k�ʖ�`jQ�u����~ӂ��t��>n`���O����ٓ8O���D��5��C	�p�~��'V.U!�DUa[�,���ҋJ�^�ٲՖp"!�\x�Դ���b�<9HP�%Z!�Ĉ3#
����\9*� ����i=!�ܩU5j�u ��<^x��6��w!�$	W�E:���.Sh�(	�m��!���eC=#�Q�nU��P�L��>i!�ć[�dQ� �KNC���	K�w�!�D]SEDhHB��	w����3U�!�D�Ρ8�T�)�Jk!�.�6 !��~�:���M�Y�d*7΍�X���|�|a����J�r�GkD	G���Q�i����<�F��CA�,�t�S���2f�ayb�i±O^a2��E�XL��K�e�r��""O)�s#ʎIO8���*g��Գc"O8E��'&Ht �䪋�F@���%"O�@��"e*@ȢU��#���"O(�J@�*Edt[u�6s�[�"O�����F5e�0k@��48�"O��0ņ�/��I���+.΀s"O����-yj|�'�ɨD���C"OR���͓=3���S-�%u�"O��a��G}|��$&��k� ��"Ox�ؗ`�f�P`Ar�Q
F� �"O���t�RqBz���#�p���S#"O|aC�G�7/�P��O/��PB"O�|�⠚6S�Yr�R�P�a�u"O���tD4ΦU�r�\�?�����"O��iۙ0+�|��*-۪u��"O< ��E�!�]Xs��;6Ւ�(�"O��B�@��mY�����>��!�&"O�)V�0�~\R�-Ѽ#�(��@"O�)"�D�I�벮���X�D"O�3΄=(R�ju Z��Y�"O�L�d�F
�$���(��"O��*w��5�4�)�F�!��p�"O�}( ��O��-���J����`5"O�b�+�oI栁'���C���"OTQ!�0:��mP��O�w0�Xb�"Op�G P�. ΕJ���O��ٗ"O$q�d:h��T��B|("O:X:�(�.{�����צ~��LX"O� 0�a
;B�9ڥ��)&jt�C"O�h���˳<��`�N�0�%B�"Oz��#�޲6R�j���5�|��"O����Z�Zk�Az���UrV*"O ,u!E���L@�����H� "O�H�6m�"zq�uh�fZ�H�Ȱ9�"Op���+UD>A�
S�X�l��W"O� <��v���T����*�?�Bī$"O��`�E���m�.J<Tɠ1c0O:d��n���;e�۰Q��Q�	?�2Q�� �&]�Q����4\A�C�	R��Q ��bޔ�I2�N�t#�C�IN��ST��8��]�� �/@&�C�p7T!$hkOKȢY�)�	�y¦�8���AЏ>֤��E��yB�R�#2�@+�#�+1]J��H��y���}�L���I5��=�����y�E�6��-C6�B2ZZ4��O�?as�X2e*,�E����S�qZ�;�љgn�jS��#�~y��AL*�*��Z-NiluY�L6z����'���򴦖D��l�wN�PF{]4@�$�p���!q |�.*��X��I^��)[gF5v�IIg-�J���D�Z}yl�eG�u������'�j�"�A��(2��2J��I�t�;�"i�p�Š�Ý?2Xt@5��3o��с|�ڨم)N�xyC�	*Y佐#Ɂ�H�� ٓ���^�����VK����R8C(��S�á,~�RP�Y�(!�>1�S!Ƽ��,�C�=��Q��h����s BE�(;���~#�8"t�'��ڌy��1E�0���i��BϾ�`(����I��p>�D�c�p�j�T*:G��K��u̓:E��Gx�O��	?#��h��X�8M�u�*��B�ɇ��鈫��ꇅߩR����+u���9�Fy��0��t��/��b�e���2A� ��.���J@���lt�x�I�SG��M.<`���퓫B�~�c��ݺL�4bs̞)0f����]z��x�j՚5_�aD��H*��LU
ĤO�D�	� �I��HҒV*�4��n53�<�$�<F{��0u��'.�I�B33�x�$&0����	�'bl�"��9�B�$'�($`}���D�/�����FZ;���� �ŭ",|�"OX!�+���B<@`e#�����O,�p��퓨 r�%[��!b�����@�C�	�f�>������°��%m���'( 8��	-j�1�cʊA=z�qlN�{e���d��y�ڹ7ֽYf%	z���C��y⏝�¼:`��h.ȁ���['��Oе���	�k�*��`��\�Ā�Q��YH!�D�7O¶̳vGN�O�
��0�N�}��^��(O�>mQ ���d�f��	ZD��/#D����e���I��fXXq�� }�a�@� �g��R]6PA �C�u���!�:@q��Z��So}b�mȶy���0�j)Ԭ���y��H.�]rt'H�1�^Y!��M�����|��M����짿���l���IA��"o�j��MXKh<)Гe�dx�`���@��y�.�*2
%aV�F�	������dL�g��dC�O ����"�>�y�.����ע�V}B�(=�Ȱ3�°n�u��ϒ�����p>��nJ Z��GX�?��Y)�DTx��=��iIW�����l�02�d_"�4�P�T�m���ȓl�|�����6�3�k�1K^���F]�b'�����O��H`�U!������4v��dêS\d��K��Ƙ$#'�C&}����eDL����{"�X-��Y�K~��� �R��KvŃbI!��D*Q�@+��NH[�y2B/��m��	a�����L��7�8x �%ac���M3����ce���t�S����ħ[z(ܨb�'l�����=pGl��x�N�I�Zi� 0QD43u�ͩ�j���ɾhg�D��𙟜H��F�Y�\�eHo&���-D��p�\�>ѥhE�dJ�r�bE� 5���5�3�O�`��Ц ��]h ��aF�@ �"O�<j�ԧn�&h�v��`8�I��'��,hӤ;Gc"����Izp
5:pk�`�*
��� ��3-y���Ѐꂸ[l�����j�X#F�~�O�	���Kl�B4��T��L	�'�бZ�%��t�tqc��ڇR��pܴV�\��N�l��ҧ���fH18b*m�� @�9�Z��M�yrN�bJL�"��j�D5����8sfd}S������<��΄�n��m��a�x��H�SFPSX�ܹ4獣 �ʅ����?+��TH�jD��ȗa�ˡ�$�p����M-�	'���4`e�;M��\[��i�X���S��^�4��	
T�[��ax�"V��=��%[1Ur�=�'�G�D�v�*�ʦm�
ϼ!��ᠵ�>�R'L�/ۈ�aV��99nH(��ٗM~K%�g�����"y�q!�p��';�����G4]Z@(S3)�T��>�����J�4��@�����`Z�)*�����TA�Y�f9�����J�y�M�)f�z���G�5����~��ݔ0��d��� LN(4�F��I+$	��Z�@	nZ�'������?j�*݀�^(��O1hܲGꐧ$Ҭ�7ÖT��P�6L6}��=�q�M;z7jQIM>�1M9=~qyՉ��m��e'>	����N�����L�$�����;�>�d]�@�bKP����iùJ����q�T� ���o�jakM�]&0�h�5�	��h~�n�a�+ħ+�,�cX#��Rt`B��B�b����d᷎��QF��q%���4�	�ɖ|�qJ��N�Tw�p�m���p����=��#�*N���'�$)�v���j�����\ t�Q�ҍ�;?��=j�c[+J��5�1G�埴ϻI�p���Fp@����$MV���mׁ�( !�GU���x���r&�@�BL�%o��Sъ�>
�2�r���;���=���A`�#5���@G��< Ɉ���<����^t�- ���
UӢ�0�ϝ9W=HA��D�v��v���ҍk���;r�f��v�W����'}���[Ba͒����Fț/N���W.N��$�i�)m���aD�
x��������궨�.D��̻6�5�C/��BĞb���#��<!hXE���$l����O��E�@�x�b�nA?,\�eЃ �(e`)���V�P�г%��;u�����3:�n�"e�>-]q��)��0 ܕ��g��l"�ɍm��<+O�i�	�%1V�iZ��̉t�0��#��?��4�
Ͳs��qxA��ɦ/��Qm��:f(�1��1��D�� �����[�Z~�\��Ԩ4Y��K���k�a�W�T�U%X�b���a�<�f������M��t��6�Ĉ�&��R���]:p�yS�6w�|�;�o�%�]����X")�x���F�=o��W�H����Ŋ<���a�-K�r��X�O���3����M+CmՠP�&�(1"�<;�X��?��ł!V����2��cB1��7?���\�
��Bh1}J?jd�W��`�B�L�%b��a��=S�F��U�O.����:3[⍲j�<Y�0
���>-k��;+nR�`���ȹ�圃g��'�̱�2��f�d�����ɦ���a^�uV��c�wp��a̪3��+ҷ&���ʛ���$:#y���3$����3��:F��!
TB�{8nL
a���d�n���4db��q	W�D��c?u���Q�h[��Q���;0��Q�C�-�N�ӆE	4����9��C�؁;C ZchI"!�e��<��I�F:�)� z�3�{2d�C�0�x�o�?7���\��y�ŉ .¾��D -|�:�&b�Z�ڂL�LB�ڏ{2-�& b��<���P00h[���ӕ��kL� ��*b�`U7�� �F"-I�i�NJ��b@�\�0�ɝ1��Q��Byx� �e�5�Έ�I���Bӌ=�ɎBB�	N@/*A�O
R�Y��A�+F���я��N銥bsj�_�=���JjH<�7ǐ-_74��ğ�2}x�S᧕�{y��p��O*A��8�E��b���'���11��q�<�&t���_r!��S���˅�4p���6�'�>q8�>ZS�eC��m�d����ī&�6�i �/m��S�LΡ�p	��(<a-����.#3�����h�2+��,	���	�i"���'w���
�B�>��ɺ<^����C {���e*��d� (b@�txqO �׹:T��:��gx>�ia��#���f����xB.�1�4p�w��?y���%F��hOƁ��+���)�����Z�$fT�)$��[�"���?q�Ⓡ&"l��o_b5�X1b��!FH�$ l���߆a2�@B�#}���J{� Q�� <�K�$�-�#?�E@	6���dܮ^.��J6�X�Bb����I:��DT�P�� �U0<O���{�y�rG�0ᄽC_a�P�E�	
?ز`��#�p�ܩ�
ç1�|�įR.z���`F:r/���[�ԡ�#M��}Z�!cC��Q�P���]�:׼A҇e�32j)�p��E�����B"`%r����
j�ʌ�R�!<Op�ۀB�i������2t��Y	�ܼ��d��1�9�N�oT�C�	 c@�hzB��4���!f�5��O����0� V�
�![ �p�<��CG��jG��8�Сks�O�ʆC�\�&�	g�A�1��Ia��K�k��Y��ҞqcL{�j�����&/;��?���O
� �Kv�2Yqb�C�D�!��C�? И�@-ȭk�xj�L�	z�C�LL�؜�ꆇ
�δɰ��96�ax��#z��2t��&S���j��ϏӰ<I�̀H���˥�M��V�[4o�?M�(Q
�	N�4��f��)���ÄO4�y"�:"Èhy�Z�����0�x���7w?��s���3N��z�,�q��\(7��(9|>���KL�cH�"O��p�U���`:3/�n�(q{�b�(T!i�΍�2�VE��o�6T/���'����5�Ɠ1$4�� kI����'�Px�-�1p)j,ַ��Q!���	c 7�Oh�S1��0���dJ��eɒL��'�(���&r~2��Sot�:���	10�m��^��y��cAcٌ�N�c5�,�y���-q���zD�W���mB��	��y�M�-M�� c�iJ�"�C1���y�����5$k��}�5엟�y®�N��t� ���Z��u�U��ybn'��ɢ+�%\!<�#(���y�a�*nV��a�6.wT��̷�y�A� ,�P��h�X("����y�
�3MV5���'�h4"	6�yM� M'I]�F,��R�)�=�y�ɡ*e�X�E��<��M@�!�;�y�@F�:%ZH2��?��5k��y� �)8Xi����86�jL��
�y�Nَ8�t�qǅ1q\eڥ�Ŧ�y�Kۮz��]��B�i�6iX���O�M�G�K�ܠ�&?���n��wT�0��_!\�ٲ0�-D�x�0�A�s�����m\�"n��2N�>Q�n��(��V~���߇v��t��+��J%ʲ$F��!�ē�5�Dժ�U//�4��D�8�2��']�y1�ŉ'z���O6l�Í� �
�|�V����'��A�ǚ
���-Y�v� Ve�yC�ˇM@ȼ��	.N���`��t��PvD�
l�"?�7��˰eGr�+"���cfa0�<�p<�%D�S�E��g�&l�����aȚͣ��>�f���a/�!�̞u~���Z��\A�U�÷k)$1�¤ =9�!�DT�Z�p��4��K��hӡӗ?�@O��֣�',x���qO���D(M� ��1aJ� �h�PO���6!߫/�ҔY���1X�b������O�}�@���lXAI�`�,3���Ô"Ob�C���]�N��s��
S�T)R"O���q��g�.�!�KR�	&d"OP\��FT�<I���	h�; "O�1R�.��hu�3	��2pz��"O�*u�F�̪$Y&�my�0!�'�����S�/Ҕ�� cI/Oh��q�'J��@�g
k���C�oX4:��S�'�R<j&��	T��a��7�(x�'eQ�#
�� u�A�$��$�|�`�'�N��N��4R$Ü*,����'�P�I��\��F�����rB9J�':Z- fk�������&�=!����'���j��^ud�;$��%0�'jB��� Șe�����K����'���դ��.�<����WY����F��������&�s�
HPX��ȓdFV|�ጰk����Q=p�ȓ;��+� �-W������e�̽�ȓ8�N�:e�̯6�8LE2h쥄�qI�񨳪IŊ X���?��M�ȓc�r�rC@�R�HE��W
!΢!��m�^!x�j�gA�܈���x�E�ȓ2)HB����.	��d׃p�2��,V�k���#}{���F��?58��|��P�F��V��\��J�V��%��S�? ��%]-x"��	�뇓T!0T�r"O��@��GY��l1WdY�P����"O�I�)�R�a(DbC�	��X�R"Op%9e�d@��B�$�0�Hq�"OV�(���9~�C,-&t	��"O �v��HMr��D��8}��#�"O(8Q���=/`��P�(q.�9b"OL����ڜ˂�����v�=�"O>Pzr\�Mx����(�5w�&�!�$�!?��:&��-+	 ��AƄT�!�d�@=!hp-g��y'�<O�!�$׻Uh��SaTc8��e�6a�!�ٟ������] b��0��6@ !�DA�{�� ���/U���	Œ.��D�~�����H0��������y���tp����x��,G �y�ʕJ�����@�;��x�ឆ�y2�֫ 4&�H�@�/bt�z���y�#��H�#���#$��b�M��y�f���e3�?ǌ,��K�;�y�V�8L����ئ{�<����yB���X1du��e� i%�|y@��yª�!Jl��V�W2\�Ҵ(�G��y�eѲu��@��g�@\j�ۧ�*�yr�Y�S��l[��H�@��EX ?�y�
�?�j�b�Eg������y��3"���id�9fy�QI4�y��e��:���)ytȑcC��y�۵5p��9��_�	I���W �7�yR�]l�(��P���`�aS��y2i@b�5Y��A%	.��������y���`aB�C&�E(>�0ء��y�� Z�E��C7��qѭ
2�yrF��(�T3Fˉ�;l�8�I(�y� �6�p9��M�(�0�W��y�g2M �a�`X�p��٪W��y�LG8xݠ�ɖ�c�H����#�y��CS:$	���n��)���=�y��R�N��C�VҒ��ǬY.�y�%>%��E)!�E���3N�y�l�0v���T�ާ���M6�yb),���L��R7t��3���yb��yp�k�M�_ft|;�(��yb�:e��I;�I��x��2)�'�yb���͉pi�<���a/D��y�a�"8�L-���H`@ɘ���,�y�D���e2�.ǉCz-�0g��'�M��A�F>ͫ#�I�M�\�P�L.j0�	f�!D��:5�0}n�+@�Q X��,Q�'�\���?�g~�.�I�2�#��(#��Mx0D���x"���`�H�y�J���� 5@<=�;�oę� L������C�� �h=��B� v@��Ć#�|�v�����@'��L V��:Lr�Q��&!��"5T!�%��b0L;���'`:PkPN
	F�č�7L�)�%�Sv����yR��"���ю� ��W�> ��i� G6��7G���O6	s��
����HA���g�Ĝr4O�%�A��P&!����R�ɴ,�8k���>��ǈ)G=�
�+��"�8p�'�\x��*�+�'�(h�]���G�Ph�EcН6�a�!9D��z�/�'d<�h�/ѺN�)��N4�Q:H�5���T.�ȟQ��H�+,���8!G���{e"O�ق�~���B'�ǬP�d�ې/**�O�84�3?ᴅ[/h> �E�6�H�7�`�<� �d������E�	>UL���� 8��'��$�J��{�^�R�kM*'��h��'�
���D=>��6�A'$u�
���qau�z�H'���!���!O^��ȓ^B�!f��&p J�
(a���D{�b�z�	��� �eyF
p�v��DGU=�B��.d��x��_�&�[��&�6�ܛ�R���kP��)���ڗ�=s��x�- (~�J�"%�>D�X�E̕�i��d:����6���)�>����8���x�i$<O�� 5�p�DI_$��ْ��`~a}��;1��Ѓ1�P6gZ����J\����N�0R��m�ƓkK��y��2������;���Y��I�OЂ	3�Hd���z�L˪[ƹ��/I��xt��"O:``S%��6��4Icm]/:uz���in��b��#n���O�Xl��A�*�vU��� _����	1�(��*� ���D��mN�!
D=e��dk`��g��	�S'��e��1��޷���(5B߰B]�-��|R镐NJ�ŭ&p�����eX���W��
M�4�:r���'vQ�3�\�p("��C�C��f��/	zH�;@΅%#[�u�a�>�Sv�ǿi^r ��ϑ�����/\A��D�,1(�f'H�a	�@Ò����V15[t�R#f�Szl���fC�4f: j�
R���q��7_p�&��a�w�@��.�q�]�'�:80ߴ([��h���?i�.�[�#��t@�@@ݥZ��a�֖3����Q
ۍn�x�ש��p�r]9C�=���'���f�y���Pr�߂a�"�X�Gֆ-k ��i�'���B�xny���z���h�K�g�.�qg�,h
��k��:�f)��E���3�8� ���8�/S*8^(�Q��pt�
 &�&{|�d���/�D��i�>b�@D�g�5P�њ�i����H�O�D۠E�?q��&2C,6��GI�/H��HC=����cN)uџt�!y�0��O��-����AR<B$�	���Fڃ#.���=H0�Ip��;m�`�Rc�r��]�!F[���Y��0��Sт�ZhmXFBY�qBQ���èkF4�8a"͸t���n����C�:Jޘ[�!��J�b}c�>!���0a���>�d��`,���a�d0SrS$�R4	�Y�����>J�h���N�5�7�ؾɂ�i�aH�$�t"�����w���A�����3A��UL��s���!3�Z�b-��X�z��z16�=h�bʊT\԰!����Ɋ()�iB�X)��أ\7����p�Ҳ!����A�&ռ�����C5I͈d�#���}�f�2|4��A�#?��拳�Z�Fz�BՍ;��0�S�"�u#o5�ܝ��ITz���:h�u�ө4�tӧ�N`"U�O�2\Q ��O\�|�:��	�?�n�`U��P;,�sIx�Hi�"����]%�l���	��O�ځ�6��0�$�$j�@�Ӑ�=t�PaF��]�!�$�	X�J�IE��1P�-��|�qO���l��e�F�r���λW��P��!:�l�+�`�2X�!��Z8������*H�����NHξ���������|�'[Ω���=PJ��t�Q%H��'�yԣ�Δ���lX~p�0E�D7��a쉹��'��� ք�\̓m���Y��؁D~�17��&b]��	&Aؽ�$�HB���2,}ؔ;f�2e &��@>:��Ie�
XPGd^Ax�p�0�oA�e�'��9+��@S	-�	�P��Dƒ#�O�@���f��"�"�*�y`�r�*�͠��#�`H<��	x�Tma�Ǒ8jY���+������G�UV�W)G2����.H��'��|��B⍕8�&P�B+vՅ�9{���v�)��H����1��'�k'��2�-�Y��0�@��ڞ��'0���� ��
����B�+xa#�5zM@!����~2	����J�Oڣ*�`S�2��d��j��H"�E!װ<���ף+�4MA�F��#E���![��|<Lp3e9�	�=6��b�"&y��)���8�3!n^�*
YI�Oz��ǃ&��z���P�<A���	�B����Q��6���n�� ͖}x�$��G���p��'_j���֞m|P��� *%����J�DYh���GE9W"�b�]���
�J�b�չ"46�P�c۹�D�F~B*"%������O�U�X���+�@|3��Țz�	0%��&�GQx�@I��:!�B���	`|�h����e�X���)C�� �GF���)_�PrQ���#b�����؆\I!�^g���5	2AԠ�;�����Pv��X1�(3$����h��'V,��6�|>H��@�ȝ�ϓ|<P��B�̉��E8l�j�3�*ӎr��,dk�5`�f�o��t�!�� ޠj�U�L1����`i(���|" �dc<��pm�*�*(#E��2]1��p��	0���;���6V��җ"O���T%�4U�z5C����xM�}�L�HR�D{�V0�d��D6e���W0�m	�E��D�	
HB5��?�<uBu*�Y� ȹ� �޽r6-�%҅�Z�؉�B���ҭbÓ[s�dQ"G�7��H��9E�8D��I�5��(B�G�<P�E�$YJu�ɓ�-7�� �N���9p��W<1r]�;1�� *�^~~��b�J{�I\xn���:!%�ݙC#�����>�Cq ǒ!L�q�f���xs�=D��H��11�<ٴ�֧��9��K��3�O�L�nu�q�����?�'�j\��O�C������
#o1@��'cv�	%��	F;RcD�PZ�Թ"&WR�d݁��'�XQj���"B���ѱO�:@b�uY
דtxp��.0?qr�S� a�Y�Ǘ)z:�W�M�<��\�X@��Q���d�<�� ��O�<��ʹ���2�I	C̸(÷��I�<VO�JH��fku���Ǝh�<"�;bDtX*'��R8�1��DSn�<���	*�b�Pw�<F]ܠ�Fa�<Q�� )�J̈@@&5
�xլJ�<�Bε}j긠ql�6c�-/�L�<��,	��ā�FܢMp�{PI�O�<q@��� �S��ݚ#��D+� I�<yr�Ү$0H�g�UjH퓑��J�<	���%���i�'T�0#u
�K�<9���S�.PpW$
\��CVE�<�GC\Md��+P,"3�@����LC�<	bj�k�t0���1�<	��c�<iDJ� #`�	S��4I�LRZ�'����`�9ES����u�Ɗ�y>� ���ŃJ~���"O�m�R�J>8V��p�kN�o:���\�șrnE]v�a�!/$?E���A~<�t�1�����O7�yR-��Bl�$��
	�4 �.T�RҤ��9pf�*����'�(X�M�;[�09M��{�q�,d�m����A��l#��^�T����S�B?8�aį�w؟x��@� %
Uz0G�z��T
��%�5P�� <О�'>rU��>.�6� o�=h�B��#D����I��$��԰�˗iZ�ke�>��F�XR�`����k~��)�{I��ɀ���n�<�k���4[w!�dS	by�o�
��	��c�4WP2O��+tE�j����qOP,ae�^�s���LS��9�%OT AUjN?��Q��%]J xL�d��e�仑OV-�R�{�n�rt��	$!��YC"Oҡ�G�X����2��=�h�"O~ʂ,Ǫ	=�LQ�	T2(�=K"O:ˀ�[=��Ko�ԙP"O�=�@�Šmuz�I'��~�䴰�"Oȥ�'�Ĥa�dX ������L�"O�1�U��?�J�V�һ�v�{�"OK��8��B�
ts��@[�y�R�ι:sń4H�|�3)�"�yҮN&}�����K�-���2DV�y"M$c�B�k�.ٜ�������yr��/S���+vOQJ�Qp�Hə�y�U�R�@��d�Ϋ�t-J�_(�y�a^�F�
Q[D��{���X��E��yr��:��4d��a)p�g� �y��7���iԯN!\
��[��\��yRO5U��$1��̩!�ެ�e�y�ٱ�*��e͍ Uߜ�ʤ	��y"�ܓmmd="!ᝩ�5y%�T�y2H}Ȁ���F�ecr����y�S�����f��	�Ơ�N�:�y�NO*0t��b�?u�L���J���y
� ��Rqc��z��9kGN�=F���c"O��Z���L��{��V�;�j�Q�"Ov��5GQ�F h�wB�[�ڈ�a"O��h��\H �aԐ\�XH�5"O��뗋ݵ.u��+�`�Hᢑ1w"O&�R�N��{�\�ЮՓY�|��"O�����
�z���l��cg6�S�"OY�%�ˉ~U>dq�,0&���"O��`$��'!
n� 6I��U����D"Oњ�G3���	�=�r���2O�������;���K�̖
 ��Q��x=ذc��<�b�.t����O"4A��yI��R�!��AZy��I$1�B���~>�0��O�t�N�
$'�9	\�j���o*@s��k��������3�|S`��|�Z�J��'R�!��4o�0�o+S��)�'b�,T�)>g�T:w�����+&��0��$�cV��V�Sa�$+ӑv����QS~�(��]p�0qG(?Y��}��N��K|*`o]�&@�y�d��ar^�x��6��	�k	n��℻\���S�OR�<!�ƺ �`EY�����'�ޕyp�K"W����O?����W��>x�r�54����v��˦�'C��oT��䧈����4�� &X�B�z��� E��O��=%>��Ubȱ��L`�$�ځh$�$�IX�B"<%?�J6�%G@�å9��5C�+�~��.D��S��S�4'^����˦Bl�8d�R�$���']4��'H�Hç-�V���EX#w��q�o�\I4n�*2��	 ZQ�b>�R�l	~**��cFA�5� �8�.?���)§5�A�bŏ�Yc@Er�&?(�h\͓/W���и'D&x�n@1wd��6�M/v�l��QD2�S>���J�]-�!
0�2IjΩA)��ēe�֘[�N>mۢc��/d����� }��ڤ�#?Y!�Y�c@�l;��x��)^Y�z� V�G�<g���s�
s���`|��cFKL�~�>1#��c���X$e �GѢ�R����3c��1v��On��y��EB5��p�O©B�r���,�	!Q8XY�}�`�~ZAh����玗$%&����w��]�'IHHp#�5?q�K|��ӹn*
I��C��0��\�4.�&a�!��c<���$q`4���(K�AM,G��ONik���w7���'�W8Z6�ee�'���rg�9|Cɧ��VEu���:)�`��4%>��J4QF�̡��'S�]Y�KF_��eɱN�'{��ܻ�''��v�6��у���xȌ\k�'a����n����⑷�X���'F�3���~-�
C�$�h���'�����ƶ�|] m���b�'d����˄L��yD],M�d
�'%�x��S	O|*�kA�8R8#
�'X`�ɂk`��3�=d���
�'#0�C�͏k���r�S�+��1	�'�6�#�(G �cn���BU��'9F����	v������f�!�'���e�K2$c��a`�Qs:h��'zv��cd�����CP!˄xA@�'°�����TYb��&�+s�^M�	�'QHL�R�k6�S�nG�
	�'�z��'^�ĭ��D�VC(mP�'@����Q�GP(E��g��U7V���'�j�x��(w��BX�G�����'޲A)��$[�t+`�NN,ҩ8�'?"�xp �r��5�ȕ�=�V��
�'e�Y�Ӄ,&�� 2�i�3���	�'5n�a7ω&z���%�ޓ9.5K�'\�zP��* �42�,=-�L���'��h�g�ȤNFP��rv�A�'�@L6F �,��<q�J��b	��' �(r�$K4k��I�3 X\�H���'����F��޲��ҢL�0Y�'GD��  <Dl0"��E��z�'��0�gg��:�8�f���8����� h�0�I
L���lO)]LаT"O�KA��-�Xٓ�e�*)�}��"O��z�����:Eq��߶uAb�0"O.� 5ޞ%�>��˯$Ԣ� "O�2I-<3z�2�aD�wo�լk�<q�m �pbZ��vˀqa���f��`�<	B"�xϪ�!u��<Kg֬�a%�A�<Ia�Z\	9�턎ym��p��{�<qJ$@���ө	c`8�`a�w�<��͓>$�!�%қI1��Ĉx�<�W��?�fh	�N�Xi~�e�u�<I�jI�h�Ԍ`���,e��"���F�<1��;���ʀ�~��  T�\g��k(��
��w�F�a�8D�B&Vk����ǈY�Y�0U*��9D�����D�;k���R)E%�8�b'#D�lSŅ�3/��TC$�=b��j��?D�lb3)U�L�lTbQ)�-dU��#0J=D�$P��;B����F�_�\��,=D�\jd�`����ݲ+�4�I�<D�hh�` ?V�<㗋[�s%$���$D� (0����N��3��	[#�� s�"D�h�t��2y�Pl���h�I�y��%7$�!����ԕCp#V��y�ە��T�'�
?`�Q(A��yr%U+A�ɛ�f��&*��u
F��y���t�T��ҭ :WL ���'�y�E�^;�hY��+9V�Ӫ ?�y��� (��VN�4�nT���8�y�"%���EF�	,���!���yb�ǔv�aS��7Y8.���)�y2mU�(0ÎUP_�y�# �y�m�I�N����\?�zv�]��y�o�@��
bdU^�.���"�y'V� �<��gK�OC�dx�m��yJ��w�l,Q�K�-M)+#�I��y"F��B�)d��Y����c��yRkW�WH��`���WC̀����y"�x�2��c�"�f%�⤆��yb��?_�PMC����%��-ٮ�ybe9&3�ؠU�ӵ�$kA�E��yO��]c%*�"�ə��y��_�M�r��G�	��� A>�yb()<�(-�E%�D���+̞�y���!��Ĩ��5?�l���y��7uQ�Q���!t>)��H��yR���Z�x}r�Xz(�B�� ��yB	ɎN�����@ 
Z�XQ��y���%@��٥+�0,��R�D�yR�ުUԼ���I*v(4PhK"�yR��"�L��-])1�<�3#Ӫ�y���!G�X"q�ʍB�X:C�گ�yR�Ŵ�����ɩE�� #�e	�y�Ɇ 	�$)��@�,�r��y�\>��%a�="����*���y�aAH�n�S�cM;~,���%۩�y�(CG��=ط�Т/\���a ��yBkDlB���T��.�R���ց�y"bYv�R�YW�9,¼5�D�y�"jƜ����O����2��-�y�$D�D��"�MC�H��EZGA���y� �1�&��Ri�:b�$�Wc!�y�	}8�Qp��-;��8W�]��yҤ�; ���R�O/QH˶I�9�y
� )�ȕ0gO�t)Gj�+y  J�"Oh�ѓ�^8M6�Y1�(ގor(��""O�u3tBU�*��,A���7`5����"O�l�p�:)Gx �/�3xD�b"O*x�!�_
!
��i���zt��3�"O���"�>��5{�M�1?����"O%:DOI,g�u��+��F�( �"O�T��Q*b���r�)I>O��$z�"OdU�Ga�7S��x��o�?-���"OI��J [&�,R �A��� �"O��b'ȍ"���6��D��"O�H�EK�~p���D�+?b���"O�[�&�*?W��ː�z"��z�"O�-8��E���27��}�q��"O�!�&'�	�
`�&^�y@"O����Pc^)���S��Ѕ#�"O��B�$*Bw�Z7��d�!$*OR`ɀe3&rlyr!�*Y����'��Rw�+
V��(g(3dfX8��'l�d˵���t-��D^�2��T2
�'�:��u�S�2.}3����Z�p�	�'�ZUC����n~,�7h¥QI��	�'�R�Pc�=.���"E�5��D��'�ڡ@�bKd,��[�E	簽�	�'�� �1i�/�XM!�-͐pN�Ȼ�'٠1����M�)K�*>k3�d��'(4���LE�<r]iN�X�F��
�'���rW�n޴��	Z\�Eq�'F�l�2��+}B��co�gE�آ�'8�1Í4p�$Q&Q�� ��
�'P����,G�(@c�H |��l9
�'!��Itl�+��"-�>Kp�'ļ�����k��qqLI�H��t	�'����Ѐ6:,�h �1��,��'j0�����r�� !�.$��@��'���eB�!3��|�a���+� ��'.�D@v���&� 0ɤ��8~P�'-�J�@�B��j���AV�
�'uش�6#��8��|���ڭ7E��!�'cЌ��w��;2��-�l�
�'�db�EK5ѳ�@��d�h
�'gf�Y�
�6q��O����z	�'�����)�^�t��ū�LW�4�	�'�6e��k�"��o�/H��$��'�,T�2*H:Js�8B�G?:ǰ�	�'�h�pANH�xpc�!2S����'�p��S�c���́#M�T��';�	�K�(SZqS7�N<e~��(�'�z�Qe	�_����q��o���';���qB]	(r���IԬiNd���'К�p���&�A�ं�����	�'K�=�!�����$� �ԩ;�t2�'j�<���ٱe<��2��R&<�B���'�v����R�EV��2�"� 5�X���'M�0S�ɶh|
4B��B�愹�'0t�Y�Em�!��	�6Iԍ�'Q�ٖ!^1L�@��A/�3z�$�'
��:�E@>z��9{�럯dk��R
�'~�И���+f�H����_uN�	
�'Tz�1P.Åi�%ۆ���X��4�'���ǣ�o����(W��5C�'Q�����Ñ7Cڃ�`C�'9t�z�����(�a@ϙK`���'�1�� fH�ѠVIxPr��� L�q�	CӠ��7�ʉ�R��"On��0��l"���	U�,ޭ��"O��{���L��A�p�ۊJ�h�"Ò�E��?�p�av��<�ث"O��2���:%�4Heh�	~~L[s"O~1��E��B{���M͍w|iku"OйQ�.��0�"���N�%/��81�"O�%(7�\Z������^P�"O�`�r.#wL���'˛���V"O�1���{ ^d%�Z)�� 1%"O
Ը��ųGK>�2����X��"O�*e�Ֆ(�"�ײir`W"O&ře�ܭ%nAh��)� �"O����(H���R(�vg���"ORLs�Ńj�Xe@ug��7T���A"Or�+$�� 	T`��O��:�"O��2%�4^����凣1�X��"O��vNH�E��9�T?+�v"O�e:B�8BPd����ʎf\>�z�"O�-�C &L��B��_x��r�"O~�h�˛/[KN�J�"I9bWDD�p"O\��e�l[�]�Y#]f0���"O*�´�A��R2`��P��]�"O��1��i��+�n� �\Py "Op��vȌ�s�N� �hJ�.�ؘ��"Ohԩ��O�pD@1��V:䁰&"O$hr��/Dμ�
e ������"O�m�uJ��?���"/ïQ����"O�4�W���E�`-������R"O�
v��Q��0��	��a��=��"OD+ ���Ț���S�ਙ�"OXq�	ԛw�Fu����(�-�u"O�uJ��_�Z��Kd
�t��t"OL9��&J<�X����8o�[ "O�J�LI�Y��敗V��Ys�"O�mi��e��3I\+y@[c=�yr��A�\��DY8}�k��&�y�a4M#N� �U'aؚ)�)A4�ybN�u!,[W��Z}�q22i�+�yBJ� 0  ��   �  �  X     I+  �3  �>  )J  �P  W  _]  �c  �i  0p  qv  �|  ��  9�  }�  ��  �  D�  ��  Ů  "�  ��  ��  ]�  2�  ��  +�  ��  �  � 	 V �  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\����IG��FA����,Yeh���S"�� ��W-� s�C�> �̙�!��^\�%�E{������/���a¡W�R� Sm��y�
���(�oE�cp�eaGL@"��'[�zB`>Tp��%O�
��q���%�y"���!���r�fU�- 6��B�̻�y�N yǨ1{��P-��E�0C�y��M�`��i��l��jmBG����?�'�f���_4&#M�a�Y�w�t���'e ������#� ð,K�xkt<8
�'�x�ㅊ:@^X����(Mn��	�'@^��c	�sB pŎL!oV 
�'��(�E�����
�Ƙh!���yυ2;n<H49������y� ]�:U��h�-ӥS@��f��y2��>R��-���/LfL�zB͆��&�S�O�z,C��j��ψ3^Z�q��'���ȔT�����'*�2���`^1q,B��,���1�Ͻn������.k�C�ɑ1�0z'	&
gFtr��J߈C�	�k#����ĕ�"�6���,p��B�I**��#W�6ܵ�g$݌>��B�I"z�b@��@U�ұ��EZu'�B� V���Pr�&0��Y:����B�)� ��IE
Hz(��T.Քw��0��"OV�YB@�� ���1��ҰE�b�s��|��'I\�	4�U'*��g�XAH%��'j6m�y�B؀��Ry�~��� �O��=%>��K�
�,���H�u�3n?O��=YR���dbD!�-̓j2�O�<Y�{�=�g}"&T`�>�S�źE���3��8�y���*~�`�DC!�����A٧�y��'��}"�!hʬ���DF����KΘ'e�y�'��x��:|װhP�'M,�JI���y��{f�4�S{�&�ڡ��O����?�Pǥ�J iI�gvt�( D��1�	0���RUm[-j�N���;}��'�z��ː�*�ccB����)�'�X�q���QS�)��� 	���,O�ą�ɵH�bT�E홾Lz����%{��O���Z}b,���<���I��\f� ���y�
�8�ڼ�VF
 P���0,0�M���1��|�%��*h���.��/��x��h�u�<�'�U�-��i�!-L�Ir��F�|�<S���9�f�9���9oC��[b'^�'�ўʧ+���I]�cA�����}!�مȓjOR#r�X,V���9��Z�o&���<!���	U���H3��J�)J1_ �!�$�6w�B�X7�S7>Br4;��ߦn��O��	~y�|�'Ҟ�
���2)�1��GW��F~�Z��~Zv�r���qa��Or��X�m�'�l��D�N{L4A�B6�n=�����Z|�z��D�c�)U犠rx}A��,y�а>Q��:`��!�f�A�^z@���i�T�I�<��}��Of˓	p�e��t�̽�3�O��t���z?	�s����J;>@���Q�^8�d(��g�T�I�4�C	@�u\t�Ð#H�y��^!^�%냈�8���H§��듵����	i�\U�@�I�� h�&E�:/4C�		>7D1�Ѣ]�1��ٵ���vX������ �w4�[�"�RL����?|�'f��'�*DC��2'��ST�[��J�'>"�
�^���OB4r� Ŏ��y2�J	!���40�4h����hOF��R�O�`\h��[�t�2❧p0�'T�᲌�-{5�}�6�ؓe����M�����Iؕko@2)��m�)�69�␇����IV!+�R��'eD�HU�'�a~r*�!]D��E�S���P�$Ȋ�yb,V�D*���0F�ME& X��ē�p>�"��6�r	-5��� ��L�<9�_zd�	!�-8�<D5*�q�<���J:��hGK��	@� 	�lYC�<��$�=����D�c�>IS����<	�4&6ŻQ�	2dh�B��{�<c�1)}(�ye
�b`�R I�z�<锥��944 �h[>z�SQeAk�<��,�[�Ј�"cA�NbfZ��o�<AbaK(+>
!rs/�8.LmK��W�<i��#�*,�3&5Bp���k�<yRJ	��а�jϥ:�	�G��]�<A@I�r�-�6У0tP�c!�Q�<#�'�� ��ڟq��m&�I�<����"�Qc��2<��Q ����x2E!4t�b�*Sc���
H�y��F�8HH8��]�*�޽��iY��yg�6����!اV�9�aI���<	�4��'	����h�\����s#�#7�E��S�? ��2��'^<xk�\�bAPUX�� \O�XZL�y�n�;�ϵG&0qv�'��d�uj�BP'�	'u�r� W����RhQ?Yj��G�!��)
w��a<�=b��3��~2�i4q�|qjԍ��
<v�3�Μb���T"Oe��L1YA��ۄDK����Ҷ�I�a��5@��+p��]�l�+��C j�B��\N�%`N�97텆 	�6�%}�>%>��=?ydh�� Ɩ�t*
��}�⦗i����U6O&���W���܊���BX0�d"O���pUw��xa`5��X�"O0���#�	V0�X��"G~�"Oθ���^(PDd���).�њa"O�����9b����*!hY�"O*�
���8+-^�1�#��J��|"�'>�0SkU�W�!�S�? xJ
�'А�i4a�Ƃ�Fs�`	�'�48��3Z�P�`o:Jpz�A
�'pT�j�炱^�M80�Ar�k�'��=#�γ[��}�����7 �����'��V-Ǹb@a�E�l�!�Ċ�_��N�29�-��fI�X�!�DշUN`����6��`�Ɔ,�!�A.SL�Lʠ��~~VتD���)�!��Zp2���!lNqKv$�D\!�;"�(�X��?;j���bQ8P!��U�<CZ�h�i�S6��[6�;|9�IΟ�"�}��	�f�}�
��BC���H,!�^@��m�S���pD�xy�KB�!�Ėy`x����M�G�^�����)�!�.8A�Ȧe{ !��M�U=!�/s)tj�!�@b�X�q�%!��Â/�@0���_Tm�i[�5!�$H�u_B�ѷh�yF���D��aR!��pL�	�ɲx6d��sHQ2jB!�DY�4���!�MR�/�؈'� �Q[!�Ĉ�7�r�:�ѽU֐�u&�"�!��>.�$���&Md�Vi��!?!�$�]����BM/7� �Fo4/�!���1���Ą8=c*9B��:�!��qs��2��D�0�2�R���"Oҽ���Y�Y&�r�Mں��dG"O@ `��4w�8 b�-���+C"O�M{�b#���1ց�G�"ɀt"O�D�DG@d�\���`L4���`B"O^q9�_��<�D�'>� -��"O�Q�cC����PFN��r��T�v"OH�t�]:4�̍��N�ר��"O�}���n��P�S�]��슃"O�q�ϛ9(!j�)���g�����"O�e��h��P�^C�
^� �S�"O,%��H
v�0� ��6)nlzC"O�鈣�S�h|y&��*9�^U�u"O�@��AC>��ٛ
C@s�U�"O(ɪ��k�څX��*qn~�{&"Oh���kO���%�<�����0�yR���&���3�h�$4ߤ�ƃ�>�yr�[5	$��B�j2��,Q�o��y��@�	�6��f%Ȯy��4h׀�"�yBb�1�&Q�a�!vf$������y�ɎkG�����=~0�xf��8�yE�(ud��K'{��0��GN�y�	��#��	YV̰�$2�yB�A�G��%I�d� ��Z��y
� <$zqn_�&a"���:a��yK�"O����-٤M�t�j�L�K�~ܑV"O�ܹ`��9��m���Ҁ�x� "Om��	:�p�!��A�4��1H�"Of�@ϕIHju�Fj*?��(t�'"�'���'�R�'2�'���'hF�kB!�<t ��ˎJ�\X���'���'�r�'���'�"�'���'�Z`�)�(P�g$T���BD�'�r�'/2�'���'��'�B�'�p0`a�S;'(\9���\�W����'1��'��'���'&��'���'^�$̓9(tfIx0�K��B,���'�"�'��'{�'o2�'�b�'ٔ���oM/cT\�y���*���t�'���'���'h��'_�'���'��Bm�*b�(�C���:�D!!�'���'���'�"�'���'�B�'����]�~%t���[���D�'0��'���'�R�'3��'��'>`ŸjԢRI�<ש��7�Fܩ��'^Z��f�'���'[��'k��'#%�U
�����1>m��2�)N���'Db�'�R�'��'{2�'2�ɟr\89A�W�h�# ���hH��'���'W��'H"�'���'B2��?���j��=>��§NM6��'�R�'y�'�b�'(b�'<b�9;��4��c�6%R@�i��'C��'��'��'�7�O��dǐ	����#�4yG�	R�	�'	�T�b>�Ӣ۴.ƹ���C����Х�Q�4c!�z~��~�f��-�4��Ħ�:�Q�!��a!a鐩v�XL��$��M��"6�._�`�%C�����?P��O�����E�m�&)�s��$�t�i�yb�'��	V�O�>Y�H��c�0��,�K��]��K��'����oz޹�)	PZ`���Mw�܁a �;�M#�i���>�|Z�A\�Mk�'� ���o��.�1p��N�1;���'Ԧ�gE�+��p��i>Q�I�_3r�j��R�$��e���3<���	iy��|�	|�*%����ULKf]p��-`�؉�gD~y!���JG}2�b��nZ�<��Oz�@�I�n5@�lϡ}2�Ԟ�(�s��IǤH�U,>��L�TP��x�b �+z5� ��יF���r�恈Z�Ijy������ć
z��p��Q:&���iV �:���æ�Jg`0?$�i��O�	�6}�A�ff�ik,][t�G0T��F����ڴ�?�ѫˬ�M{�OR][��H2Q��t[5[28Pp�1��Wrΐhw�{�^�*@bY�k�u��|�P�iת0��'-�֐q�h���G�v�9�$W��r���=D��kƋ�=9 �BI�&}��r�A��c��(�cR)� 8r�&�,i�ɛ6��	,HEr`��,	U�2gC����d��^R5DP�nV�1$��	w�E�F���$Lc�NE��~�v��U~m�$�wkS�%�I��B�Z�x�5T�%8�Ubè]�8���j��Q�1D:	rx�3��c�:���O����p�'hh�S�
(��J�1mf ��4�?I��F8��+O�i�O�I.}�l�p�,tR�D��k��QY'�Y��M��K-����'U��'G�$K5�4��6�|�KFc�J��CEȄ妝2�g�Ay��''��Ϙ'l�<Y`��bRd+\s�!��n��%I�6m�O��D�O:F$�^�i>u��h?�֍F@�,�H�%+B��UzqLr}rY��@�7�i57M�O���Fs�*��d	݋�Aҳ���+Äml�şp��j�����|���?�-O(�K�I8�N��C�z@�b�Hæ9�ɡ�
b������IHy�F�[>X����R!eH��SS$_�b���e�5���OF���O�ʓ�?������*�/�`�����\|T-Q�o�k��?��?�)O��ADX�|2�H�� �TG��Ri�g�b}��'y��'��	ߟ��I
��'|/�	B2ɀ@��*��ӛ
N��'R�'�bR����AR��'s��E�GmS�[%�,+�l��zX�`x�i�R�'�����	�A�c?IJ�iT>"j��d�à1��*�&~�@�d�O����O<�a.覍�	ןp���?%u��0*�|�#��9�ʐJq _3�M����O\���=�H���<��!J�$%>����	�D��k~�@�D�O 	�v�CȦY�	��	�?����xy�K�N_>��!����aS�׸��d�O�����O��D�<�'��ӥX��]��� 1�fe�whL)0�7͒�]l�<��ݟH�S�?E�Iޟ���,g��8b�9/���z$�W��T�޴�0:���D�
q���<�����đGM1�,�s/^��,Sڦ�������:V��Q�4�?���?Q���?��\���0Ɯ�\�.�y��@�n��'���ŝ���8����Z5K�'z��4h�7�@;�����Mc�b�>P8��i��'R�'7v꧷~�B�>V[z�j�왭i���c����ދ,����O�d�Oh�d�O�'o����gJ���ՌЅ_X4i	��"z���'Bb�'��A�~�-O�����Gg䝻�`Fq��J�&��2E5Ob���O ���OH��<�tCցO��IW�Xwڤ��Ǹ#�(=�p�F ���[���	Ay��'Ur�'�f��'��БT-v��y{u+n�0��GdӨ�$�O��$�O��Ow���Eq�`�$�O���Ć%!qB�k�*A"k��p�#�Ǧ]�I� �IByb�'�l�y�O�L.�)TmL2Kl�Qw�G�
��lZ��0�	����������4�?!��?���Cw���$��Y��D�cͪlPX�nh�	~yr�'���ҙO�S��s�� Z��G(~��8�w�7�|�־i���'�v(���t����O��d����I�O���!)[�M��@���*�lY�%�\}�';���t�'��]���m��2��!a[1'�84F�DM�&i҉2�"6��O�D�O|�)ퟘ�$�O���O�x��#�{R��q!�Z��)m�����k�i>�%?�	y 2�8�7tt�x��?i��9�4�?���?��eɁFD��'"��'3���u��
�p�<��m�){3�5(��L�Ms���dY�3�?��I��$�I�p�p�03�GP��c��cV୫�4�?��*P��')B�'ɧ5v,�hJ�
�m�;y�����e4����r��$�<q��?�����ԋ3��TJу@�F"�ԯ�/1_x��G��e���t�Ii��p��6	aB�c&J�)!d�YbN�Y_��9uf����'���'�Z�@�E��$��D��.$'�x+�HR�Id ��&��$�O��$!��O��dL�<�4���]M�i�D��5��4s���!/
��'o"�'BP���-�ħ@b���g]�K-ڹ�ѡ{ ��в�i�r�|��'���X�|6r�>�� A L���G��-���q����I�I��L�'f�	 � �)�O��	C�yY29`у��QV�Y�W�D'�4�	�萠��%��'8M�H�f̧R&$�Cw��il�Uy�'�|!f6��F�t�'���&?abްOѪ�XPa�?�l�'�Ʀ��	՟(#q��ݟD�<�}z��-�y�f
�F�T����e�,���M���?9���R����rƠ�ț[��xª�Kho��G�}��[�X�'�?���Hbۄ�
e��K�V����[� Û��'��'�ё8���O��$��X �_Q`�i GJ�:x�Z��C�vӶ�OLi�4��m��l����|����kn��YfK	E����!-W#�M#��<n�Q閘x�'|ZcI:�*"�3|����YA����O�Պ��O���?���?�+O��G1�t����fg.�2�H~$�$�T���&�P���<j���^�Ը��=�.]J��ò_��My�'�b�'7��9�"� �Oc��ɒD��;s/T.@����O����OP�O����O�<* 6O|B� |�p�f)`2�����_� �I����	uy��������ёMߚC�R4�#a*�=X�E�զm�IN���h�I%I{ډ�	t��zZ�0T�қ?�͊�գH����'��W�(1��I���'�?���rZy�/Ƕ0�BuH���:=�-	�x��'uR/�/+m"�|��bQ�Aذ䖹q���=�
(�i�b�'�Mò�'��'/��O���5�C_�/�b<��ŴhU�#R˄�M#��?i0n�R�'�q���T͒=X�^�[�e� d�89b¼i�V�S�l�BPh��y�b���(�(��/V\��ȓ�p����0�����$
�0����R�9AA��*CqV�c	>� �$	�tRU��*$���!����� �U큯<���I�6DLĨ�J�U�&�j��;E��qGB�0������������3H+��$A�G�!��Q3)�(��䲠&ۛ7Q�B���?i��?������O��S�Z ���2ό�f�S�F ~�\�!0)W)(^�% «� ���$<O&��E�[� 7����mB�l��M�QU]n�	��U:�䤂�O1<Oh�	�Gɋk���c� J۪-�@a��S�2�'�'���'�ONЈŦP��>��$g�#D4�̊"O8#�	(�8L�seړZ�0��w�l}BZ��h��	��d�O��z���9!.�ar�A�`�t��OX�Dĵ`t<���O�ӭZ��zEβp���#1�^�5�U
A���B�ܘ����k6����C�o����2
r,�Y�ȉ�+:��%�+�S�)N�|���t��>Fx%
�$/�<lGy�ö�?1���0n�����(I��nQ�$o1O���@.��[�a͡1.���הC6��F{�O��6�Tds$��#H�Jp�)b��1"H�D�<)�e��	���'	�Z>�� �ꟼuɓ���j5�сx=���F��H��*�ޅ��!U�x�<0v��.f =k�۟Vʧ)*�y�� ��  �q��dܥA�f5�O�L�g�0|���c�cɲ&^̴�SDbܧhT���N,A]rIk"NH����O����'Wx7�O��D2��x>u�b_�(4
d���_�t�G�O��d�O^�d <Of�:b�*O�r\[ǩ�5B	.�ش�'�"=yƫN �$T"��ŗ`R
L���S�c���㟤��"Qў4��� |�I�l�I��u�N�6�L]���#<��HǞ��J�¢��.}�>�Q��	s#��iDR�$��	����3�Q.���ѨѕA���	ɴ�,l�T�������T�D�h\���J3u3���ԣ��[���O@���H=:��Y���	�HNz\��l w�B�صő�-m�хƓM��q�T�sz^�´���;.��'
#=����?�*O�0c�@�m1�͛k�f�HdnK�=�ĠT#�O<��O���]��k���?A�O
$���A4���y��� [������|(��	 �F8����x]�8K�Z�K���$��c�:�U�ƪ��|T���b�H��\R8Y{ak�%Ѧ��^���b*�$�OL�$ �	ZI�`���T�~���I]�<�C�)� �$*���b��T��4l�� ��@K}RR�D���	�MC��?Yc/��s�:�vo������$!Sr�'iqq��'�23��ɡ�`�$iȐ/M1a&�Y� ϓZp)���&
1��jHx:���&Z	�(O,)�G�4���F�/
܄�d�=7�pS&�K���G���?\@�0d��(Oh�`�'n�' N��LF�P��S�dˀw`���'�4	4��Z�-K��Ҷu�8I���2��|jQ�i׬Ј�,��ޭ�d #hdҜbb�|��Lr�6��O����|����?�����F�[��J�[�2�s`M��?���Mt����]1!��]�c���h�uj�f�a��-z(��H��Kχp.�+3'̻.�e�Ŕ>y��C�wR��'��o��Y��h˽F$T0$�6��!�XbA��E*0!K��ZP��+������9zOh�0��/��wIW�<�B�ɢvI��s��2H�xx��V�k�4F{�OR#=i5�A32Ԣ���E�)��
�G�]қf�'"b�'�����V�dh�'3B��y�׾b/*ɢ�(�gF���,JG�1ON���*΂p�џ$R�n�"�r��/��)-�%Q���̓B�P�B?�3�D�u��x��K�y� 9Qg�A����O����u���Y�X�I^��(SS�AP�ܝZb�+���Ɠ$�Fp�F�4����a�U�l�&i�'Ǩ"=	�*��T�'%4�
�	�q��,�g�;X�x�
2%x���b�9�?���?�DY�n�Ot�s>*�D�"$�e9$�hZp�i�L$_t��(��yw�q��G̓c�&ЃV�BQ�L(���-H�xKT�Q�lJV�"J�+M� ��O�~�eʦ&�9׸,����.Q�$��b�%!�a�բQt��0%�G�c���dQV؟P(� �~�Z,��ш[�X��,.�OJ�O��X��јj|q� ��{o^l��㦹$��_0mh�Oh��6	<<s��L�uffH�qEӭpd����Op� %��O.��d>m�D�R�b���r�0G�`���I7�:h@jҭ;�t0Zdˎ7^r�@+͜�Q�����?ڼ�{g�D� ,�6-� D|`Q���Ԗ_XA��B�M��NB40un,Gyr�Ʋ�?���i=�6��OʕH���Y�K��Nz�ܨ���<q��������r&FŌt�Z��+������Iv�����h��T��H B�>\���%?�Hذb�O�˓3$^<�2Q���	M����o��׬*��M@P�� ���2��� ��'uF�h�MԷ�1O�ry2Ί�j�Jp�S��fpn��mG���	�4�&|�0�7�)��3T��AA�
�Q���xq��'0,S��?a���?I���k¿3�����P9e?�(���M��'8��'�v�tl׺.�P�JU둑Z0}��D��\#@�(l�9�&A�
lH�3b�UBy"�'�z	�Fl�#�b=��O�\��'��aU�V�+�>XW�N�j�
�'�D�Z��̯&7hXF@�쥸�'� �"F.
�L噵�T��R�'��wj O�>��!�J�]T����'y�pap⁓^���ӠiG>\}x�'��ĺ��ݐ�
����\_vT��'�@����V	��dh�b��n�d��'�N	)�E�����O_ o�UQ�'�\��H$�.TKK�,�Ѐ��'��I B�ɧyh�a�$^%*��tk�'uL�	��3�����*Q�^�I�'b�h$FܗA�䀅Ȅ `yHdq�'S����jEM������Y�H���'q����
\h!�S" =�\Y��'O���ŭ]�dx&d� �x����'��`�IC��6ʂ�T�s����
�'>h�)L6I��p3��4�\�	�'��m��a�$���B
�-�r���'p*���$�ف�6�����'{���j	��l��e��<��;�"O��{�	�k�f=�e두Z�ʍCV"O��:$�
�v���z
�K���S"OV�Y��̨^[����C&d�B��"O�9PAP�Z��@� �'�� �"Ot ��2��xx".�pw>�S"O�1��Ꙕz�� 	
t�cg"O54�U&y��a�X�F�Zp8"O� �� *�>=< ��Ѝڢ,/�d��"O��e�"YD.ԓ7�qM^5�"O��p���*��� �Na."R�"O�$��
\$�x<!���"��U
ROXHb��Ժ���� �2z��2�N�Dh<i@�7\�h= ���l�*�Y�&�aX��x(��1}!��Y�L�u��d�2%!�B䉈�6|.	���h@�����1�O\Ij�W#*�,�O�>��O�,ϊ�	Z6���p��(D�$`��@�e2���C�I��4�`a(?qa�ĳl��4j��'��-��3����n�K��]�	�y�Ărf8:�䘋#�X�4Rtf۹j*6ɠ�O\(R.��Vb�kd�Ɇ�:�cc�@��D��"S,��O�t�b�EE -�=�*\x��{�((p�o�0�V0($�K�^�9��P'�h]Y��بB���'����um�<��䅺#<�3}��'�Μ1s-"MF�ISq�W�On�(�%Dϲ�;g�J8�ё�:O�i&����<G(� 3N�Q*�mQcj�<���F�R˓mvY�g�)B���6��!��$x�nױ�Ɲ ��*!�ʉ \b���I��?����$�U��I�"��9P��8X!�K�D�EU�̮TKP(7=X5���MNV"��$E$s�֋E��y��'3n�����Ա:�~(�a��p>��LV�}�xh���/��,���ÁA����o(�	#�f���[G��%2�G':�O�c�#��4ZX�tF�<Ra����ɟ���;�lW<s�����(9$��1�n8�@ʔ�n_���~��-��N$L���-/�Z���'�Z	� �2Z����*yy�-X�
���*�����qpkIN�+����Ó���P��Be��:V�:���O�8K�% Q}�Q:���<�
y�˚�T�ayr�ѝC�2��g��C�eH�\���:& �= ���!�#Or�F∠w �i*w���6R�!�m r���c�bu��ǌ8}�0%YR �D}���y���q!ذFh6�d��9�O��phZ ����@�t�1��X3��|i�$b��ӟL�̮��]��?!"�* �Ӱ��#�P|iA/�	d�
MI��A{�շVtBAi��':�Z�L�L���P��A��HH0�O*@ѥ6Oʐ�dDW ��H��Yb.�Ӣ˺�c��x�Ep0K"U"�)0���5�`W $�T��"�DQbe�BX���  2!*TU�%a�>E�%��j���<�@�O�`����?E���^�ALpijŃ��>K��C�$4��:�0á�/��O�.��N�ܭ�I�7[�5���	tf� �L����4�~��k��U�0H$��HQ�ãA:�/�tz�ł7��`�< S�ów�����i�ޥYD+T�Kh��3�)j$Q����
����~��@�&N5+�����*,O�-
�咬?��	C�.�bTE�Ʃق�y�c�0thR8#�HEĦ5mڷ:��آ�PF��Y������+a����O���X
pB���0?9%�����M� -�,��U�W��n�0B�V\Z$��;:�h%����-g�|�!]?�(�#إ��� ��(�$=��T��B�#���?A�P3'$� �U,Z�hث��.P�1F
h�%b��q�L\��L��r�zu��@V9�P�0O4	*��G��'SW�4� �|ղ!��!8��ݍN1  [Q"϶8�@[�
�O����U��m�Œ�M��y�!4��ń����;�%Ƈ'���wO_.�H	������b}z&����<��ӱ|�Py��_!mx<�ª��.:<<�g��W��֎�h,��ˣX��(D��
ǀ+,D!��.�jE.ĳU/p��/@x>LdB=Y��]��T�W��8�� @�L��PC$�J`aZ�{-hq�A. D�d(1LĘOKd�j�]��nζ!1���']x��	��D�1�R�r�ߛm�9ق̔�7t�[/��K��)e;xY٧�#��e�1���\�P����yR<�S
W6y���O��̑�艿8��M�t`�� <�T�YG��~t\��Ԭ\'F�
���GE�E��C�x��,���\<n�Ju2@C1n���qS�B����i"C�T��H?w�(��%�@�^ ��ɍ]hd�����<����S�g���I>���C�'����B8M� Hx���.�NQ�u��b.��H��bi�����"q�h�MD�NW�JN\��	�v��`��MD���K؋o�"9 �j9�y�h#�io�:qգ�&�j)�@�^��ؙ�Q@�r�DI��^cܓ��%�S��$ju��r��L�Brޑ%��� ʵ)����cN���#@�>��S�řEI1@�DP��4M�T�3�I���ɒY2.�K��?k7�ܺ!kޥ6�,�!�B�tN���rK܍[2�\h�O�� ��h���Ji�OQ1-Z�y���z�^L�'��op�F��ZJH�����0<	�%�=
Iԅ��Bހ"`$kՄ\�`�Q�آ�@5�'9q*�K���g��r���4~ݓ�B]x�p���t�~�ͻP�p4+CI�lhԉQ�b#8PNu	��OpeBI�t�|R�jx�Nt�WJA�� ϙ,BTy�CN�A+���?�0`՗]��7H��!�r��h��R�7�4�z��*9���U�f�(�x�4�ē/Ԙ��شh���N�\���(�O� ��;4EG3+����
Z(0Ѭ��o���t5��i*�� �JK�'`�P(�8��_��S��{��	�*���:�MK�7m_t8���'�;v�����\�>Z�iI��
�OP�=�%x1F�j���#Q����M	Ff�`R�'.ڕb`�^(f�F�h��Ă�vA!')h'<�!-�1O<㞐����S��ْ���}j� �V��بP	�t�̠�B%C �O�e
��2-��U�qh��C5���҄�g	@��L�1H�D@�W'+�4#�nZ�l14��6�I"P�c�h2��Ĝ$4r�%\�Y_�L�C&�L�KF+י���m݄y��h�=��OL�1�~�xL���Z��	�w�¼#�G�i�ucP�'%� ����e�qy��ֽhMڤSQ�R�'�f��y�,^�stz���e�xic�@�'.���-�	���߅2g��`����S��P�V	T��1��K��� R(��Ob���O�0��C�&�l(�s,�-{�вT#!F�ٰp%__�.�,]��/ޑL6�kF�B�0<&�D���(���ZGf� p��dg??����~boO$MΈ ��)v��1ST;����r+ZEkS�����8Y�8#��%�����ΣA��<����0X�v٘mU�<�`�3>_���\�8Y��W4s�0�;��ɡ�#�p?���d0?�]%2�����zrdI#�C�J1n��Q�l�$u�U!֍
�d�f�F)o*��A��)m��� ��K��	-r�$�L��(b?�$��++�l�8�e�	1|tqA4�N/l��\Q�OP�i�DU��ķ������ z=�$$����&˟>�,�3υds`#E+3�d�+{H���w��e���͡%��OF�h4,X:fV��)E�t��I�`ԬC��Qen�!REJ#��tX��Yu�DS�p�a�?|�b�3$����6 �M������%s7"$��g@>%�.dk�� ��\0˓<ʜ\�Ґ�܊�fJ�m�\k��� {�RUh$	����=��'E����nZ�Ov���eE���+so龴�K>)wg.Di��J�Ɛ+*O����8c�"4(�`��v�[�U$b�G|bDJ�F���І �#ˢ����P�yR��#"0�c��q�ȅ	�K�m��Ac��	�g��qL�7�@��>ٲ-�
7Ƹ%S�l�:r�@!!�o?1�%�g;Ԑ!�LxlےL��<qJ<���RF踓t��$�AQS�50k��*�	�HId�4u�a{�K_g��4+�FT<NNu�v	(<�dr��_��D����韉�5F	�/l���C�t�J�"3�K��xB�,4�`��S Q|�E�b�͖c��xA�yb�ݶ�ē@"�݉6=O<�VWL�%AR
J7dȢU���PF�`�I	h]� �Re�
B�@[�A� ɐ��!���,Lx5f�K�8{��Q�	���9y�^�L J5�Ҥ��➌a��G#EBh�(DkO/&������>F�T�z0�ìT ^�ƱXЫ�B�'�F��A�}�ε��J_Lf��d�OP�#�L;.���	�6�}�p�/ plPb2�ۆ �t�d�gX�آ�l�W�D�#Dd�ia� 6��|+G�9Va|"�K
G�ɳ�ρ&b�f�Q'�^�$�PR�$���[�}�Ԏ���r)+s5O�,2kW,~(`��儰D�e�^����Z�'�\�B��"L������l_�Zo~���
U�P�J���-¤)�����-�'B�(����O~�Ra�Tj:Qڎy��@H������d$ �L�z�僠bZ!P���IV"RL�L��[�,���L�'H�ƉR���]Tio������ a�j�z�ņRtr��L~� Cr�A6=�liF}"�Pǟ��H>�TkU�`�5�0'Xy�� �efM,�=)$GE4 >̭�!�Ɗ>A���a��F@@�� ��	p�:O66-�(H��5��@y��yb8O�X��>O��yg��(Ѵ�Q%+P� ��}��t�z��nt�E��O����tH6��j%q��y���X��-?��؟<��Wa��mZ0(�P�_p̓o���+1�E�Z���eI���ҁ�R�\5ۥ͏�ۖ��e���lz>7�'?a��[�t����|gB,�0�.f����aGG��p�s.4\Ou@��A�È���b��x�n�9�L@g~��բGq,�w�|���
�Lvx�E��h�y[2n@�>tF���/���ԏ�X���@Ű��|@�օ`�@PH6�S�.�1O@QJ2�CI�4�`4.yʟT�A��B�̀p��S�:��Y+��d�1V�A�1P'E
�1ʍ�����uw֝$1.��zS����C��}G`��Ib��۴y�v)z�W?	5&4�� !}���!�76l��Ӎ֩`!.	�oI?�birg�F}]h��O��>��	�iV�w��y�#Ó;�(� Q���*f$t�J�w�2=�ۓ8�X��$��08���&�<E�&劇��,��EV8
qO���*q� ��'��;zT�T �D�xv���I% �DL�co�118 �9��B ,��u�L�$r�Qgj_SܓE}�7mOs~ ��	d�Ӂ\�q4i�o�n{qO�6�48Є�4�G0�(�`°W^X� ��8O�\h��|JcOH�6.DFK�?a�����&��tv���'B><�']:����ХhCh(��y� :T�QUꕎ1���;�N��� ��K�8%^��DL�3kthZ���gy�π �E[�M��=��x��@�Z��@�L�Z�yٗ&���p��'� ��Nޞ4��9�iH6��B�!l��K�&��p����l����Oy�O� �F"ٺ ��P,� YJ-2C���p>)��ɦQ ݴ``6j�cP�e{�Ա�!ǁ�@`��i��dX���:Ԫ(�l(���(�*(�O�2w�:�c�O%���"OF���8 D�ZE�3��e�e"Od�lF;X��آ�ћ\&�c!�5D����Q��p(ۖ�ܧB��a�I3D���U+G)|@���_�dLxP!L>D� ��I��`2� ۞
�z�bE�:D��ICh��*���T&W3�@yas9D�$���!`걒�m�*��+�G3D�HQ HԜ&-�H���U�D&�  �<D�����W�$�|�P�*�4%� ��I0D�|q���L��:t�X
�.D�|����?��2��P�uC(�P�m-D��	fH<|1q�bN1p����2n)D��P�n�B<��y�)e�n��m;D��R�E�
��`�O(�b���,D�l�Ď��t��E�;�T�Y�)D����ÅRV�Ж
2oQ(P�-%D����[�h��6n�4)>���(D�xC��Z|x��A(���I;�e'D�T���L|h!�V]�H��.!D�����(56��f-��	�`5D��J���RĎ�h�OF���c�4D��b�nI��ʰIe��/c����K2D�D��,�-=�q�%�;>r�b�/=D�h`������c�� IH$�:Q'>D���4h�w���cC�s�,DȵC=D���6EЪ��ۣC������?D�l�V��ST4���Ňz}���"f=D�h����LL#�D�����@:D�L���)7.�=��O��]�PiХ7D�Hs�!RV(A����xh�m��(D����(�.�Ԍsǫ�$D�- �%D� �t�@>)��@� �
IIzy��"D��Ѣ뜄F��=I3��$^�D�#D�4��d�>�����-� %��k!D�����5}U�4�ROV�kv¡�Ԯ D�����9%�N�C���1��I3E<D�xEذV���S)İ�t�(W�=D�q%��Yf�T����)�b�#�,.D�X�BV�}���{� �2 � D��B�(�:C6`����B�	�@B��n�NԣC�.La��p�	��=&B�ɋR�	�th*����5�B�I�<���Å$��>�f��I���B�INS @`Vd�?<aR�;�+<�B�	�>�cW�J8}*�悒�xXHB�	�R�t���Q���3�ʃ�o"4B�=GA�L���RDt����A�h�0B�z�]���0D�P r�҂c�8C䉉t��QU�E"+pj�@��4o4:C�O��K������� �E�Q�$C��~�m{'��c2�-(F��4'�B�I�&_��iIE ր��mh|C�I�/�[���JҺ�z��2׆B�I<	4�9D¶�⡫�O�C�I*	�f��f��W����p䊘r�C�I�Z���� c6�
yp�
9K��B��
�<y�$J�J;���I%0�B�k
e�B�,L�zg H�K�&C�I�<�Ƅ����4=`�ǁf�4C�)� |D3�Q,����HE<p��p"Ob����i�rPK@����y �"O��8���(H��x3M��4(2�"O6	�t@˞o���j�Vy&�r�"O�m��ȇ�%�VĀ�)ͪ�֘X�"O�9i'AC�?������Y:X�j�W"O��R̃4,�Z1
�%c��25"O�ݛ�@ n�,�q�a�vaQp"O&�a�DJR����6��$[��R�"ON�g�J�Ϥ<����j���١"O$<�v&\�J�����<�V@��"O�!���?Sv,��
#\6�@$"OЉ3@y4H%۵�O4Z���"O>��w�Yo�ґ5!��{(����"OȬ��%J�!o�mc@���j#��#"O���́�lCZ��6����sq"O]:5!��7+,�2�h�Bw"O���S�,�x%ڷl��~�����"Op("�tx��ρH> ���"O~h�n۷G\T�)%�W�[4�`zQ"O�g@\��G�9*�X��"OP8!��
J��ɒ�@�����"O����ۊ=�Z8f��'�2�"Oni�O/J�zY�:��i�"O����;F�jD��!%ಹ�F"OT�R��
�Z� �աK���
�"O��u��>�$�"H3���r"O{w�I) ��j!�C���a�"O�1��'̹py
�{u�:Rp���E"OVA07��gF�H�<m�Ih"O&�2�G�
Z<���J��:O�qs�"O���3�F'r��$��/�%sZ*���"O�0J��}vh�����$O0�Db�"O`u�b���C���kpD:F!8|��"O�q#�ҕc|zE�AC�/RJ٠�"O��&�,/*m�w��=���D"O�iQn�*3T�)�C�x�����"O��Q.�蒱�۳1:H���"O �*��¿o�1�/
�7�ف"O yx¢D�'� kRK9��z"O�=I�fY�^��*:��9R"O��e�T�?Xx�N�2����"O���jK��(�ß3_��p�"O����	2=�@�ƚGs���"O��&���	 X�/;�И8"O� ��*=�d}�0-�� �bѹ4�	�/ב>�R��7)�q+���7B�Pi�+�O��=E�Ԫ_�V�`y���:&)�H��"!�$�c�t����CH�d����g�!���W�����g
��y�/P_�!��8<#~�3ЏE�ׅ��l�0Y �"OΈ�
�!5L���F�ϕ/<�vY�@D{��IL�:�hG�NJ/���Ł@�2�!�R6y5:l���P�`$��� 8�!�@�f������`*U�v/փa�!�о-�n@�� W�n���!����!�d	/U.壁ɐ"q����Э�+\;!�D]����Qm(=�J$k��u�	�'�$e�P��(� 9"�gb�d��'�%X�f̡�uHam�`�z�)
�'�>����X�|e9A�E5Y���	�'�faIGz�|��@̋,D�z$��'قac��L� HZ�"�:�<�3�'�6�����83��x�L� 5�xd���� �e���Þ�xD��cȓe�>t��"O.Q(�A(|�Jc�
/,pl���d�O�2��Ҍy��q�F��=�x0��'�NȂ�HK'g|���mÞ;� c�'�,0s"�Ї.C0ų��5�^���'\�qMY�?=�IA"	��" m��'�������Ȱ�݇C	8}��'\)�7��cOJ�X@�2&C�=;�'�TUf���T����I�)�ά��'l�����>�tQ����(�$�
�'{x��e��!�)AG,p��	�'�c �˓5��@	�oF�}���	�'�P��Ӆ���:;��1�(�"�y��Tu�����4�01�⁦�y��^�9u��.?~Xmۇ�y��9R� ���;fM�v���y�
��'p>��v�U8����^��HO��=�O���%^
��s�[bj�[�'G��A��_}��c䣇�r/ख़�'�d��3�/H�l��#Ϗp8T�j
�'� q�t�@1(xnQQ��{S��
�'�\���o���yçJ l�"|1
�'|�prF��iK��
�IU�2���
�'��z�
Gs��İւ�	[����'>P��a�
�3��	����$��@�'VTLIA�A
�`{�,�"vL���'�ɀP�!�"�ڠDB�+D���'W���1n�ne>�b��L)G���'3�`�'i���j�B���EB�q��'�]�/��b�<� IҤD~Px�'3R\Ҳ�
�	�4��gN74ʈ2�'��J���`�P0�i�}o���	�'�=h�#����ջ��6c&t��'�<X;���M��s.�x&���'7(<I%i�h�9�BK�[��A
�'d���Z $��`2�S�O�� ��'���Ӯ=4�<"���
]!*#	�'i�:��
�n��A��,EA�0�' �,`1��;;�p���85���		�'}��x��?(�����^��c�'E`l���W%�NUÕş�j!���'���(C�נ��u�Վc���'n9Y���?Q("�	��5V/B���'2pHhv�;*s�5����+D pj	�'�������*Ġ�E��}����D�<�&��)�4��A�זc�a�AR�<�-C�||��L�����w�<T*��"	|�jd��?\��kql�|�<!v��5���C%�\��JDK 
Fv�<�R(����19�b�7a2 <;��{�<�dW<T\D���.8f*�JajOw�<� ��z���A��ȨT�ƵB"�^�<��)�/"glMPѮ�U<r�	��T�<��#�.���*�+ꂴ1��US�<�v�U�v-�d`�� �ɂB-EN�<���E`@H�Gy�Hi�QVG�<���JWe�t���G"I߶����@�<�Q/x�|-���D�W�+�%V�B�ɽ\�{� @�B�6ԓ��^OJC�	3b�јF�$LLqW��DC�ɓ���&�R�
&z�R�H��C�	�D�Ks�����h�ч��ryB�'������T�~	���T�����'� #LC�(y`,���T=M�j�J��� �D"ݠ]�;��� ����"O4%8r��A�0q�%
�^|�[��'4�OF|�vؾo�  Z��_�<�T�Q"OҜ8��V "E( '�}�N�:6�|��)�Ӕ����A�g���	Z�pB�ɚ`�0#4�G�=Tx��ܔ�B�-m��֌]�r��-��B�	A����ˏ�U��pV�qٞC��p.A��AGv�N�ؠ�S#%}|C�	&O0�@�bj/yW��4�P�O�vC�w*^xa7N
	nip��fۃRS8C�	3]�3�o�=&!
1D�׶d�C�	�T����w�Y�jS��3"W��vB�I"�p��CB�DR�	�s*�C)PB��ZƦ�� Kr�����52NB�	F(�Q���Q3LlN�(�HH-]�C�I��	R'.3���B���,S�C䉭j�>���MI*y!´;�@�G��B�	�Jp��cG�Q��b&"ߤ0klB��)8S��T�� t\�+��K�2B�ɗ]xZP3'U3j\8��r��i��C�I;0b�"!�Q�% PH1�ĪyA�C�I��"���/�>~Z��%M�22�C�	2H��@����dY��K�C�	 T��(2���/D��a 	�xC�	;|<�6	�"$X��DT(!HC��7.�l�٤��fĖ�C%/�A"C�I��V�)�.�f9��@��r6�B�I2p!V�XvF�\D��*��B�Ɂ��ipc���*r4���OB�	��fX��-�aԪaÃ L'�C�	�%��4���w�0��1'��C�I�{|�՚�D͕]�M�K��Z BB�I�2����!��*z^�y�`i�U?�C�	�3-"�bӄM5���Bl�4;�nC�I�\�x�Чl�=E3��ba��i�0C��I�\�)�D�0�4TY��<xV�C䉮1��tQתW�mdjqz� �+��B��G����M�(t��]�B�I�p����a�".�,�(4���8"XB�	69�����HF�2&н��-��}�B�I�G[����ѱ{L�x��k`B䉓l �hF�p��DI�E��6��C��v�V� ��J1Z���k�yپC�I��x@ r	�!_\6Y��͝bG@C䉳 x2��&ѥ��5{��/i.,C�	�OBZ����W;�ٲ��
���B�	7 ����S+x��CfʢD.C��)9���e�ChB��EJ.8�C�Ƀ��4R���i{��r#�H�UG�B�ə	*@�E�҂+�pR�%ǎ^��B��JIȠ�)�X��Q�6��B�r�="
�[b�m�5�,g2ZB�D���(�OX(�`��A¼}mhB�	�qMxaص�K1<��J���2RNB�ɱ��9�QU(>�s�g2q"B䉁UP�5�q�V�fM�q��$�1l��C䉩=ӲU�ΐ:K�d�@B�̣+�C�	�H��1��7����JX#p��C�6^�>Ȓ$.H�2�̬��-ɷl~�C�I hqbSbY�5�d�����B�I�n�hLŹ5z��5/E�H�$B䉵/ϒA�
�"mQd��!�JB�IT���j�dP�/�&����_�,B�)� ���$d�#Vf��f�֫Q����"OJ��C�5 � �Q탓+��L�"O6�ٷ�� [&-ˀ�Q�D��hV"O�=8�l�m�N�2��ś����v"O "3K�>���R�
<Qz���"O�`"���
0��u)�/Ъ�p"O�{!ϒ��ۢ��#;��@s��i�<9���:+D�ZP�'kݚ`�s	�a�<Aq�$, fC�b�ۀc�x�<Q�a�"0qn��F�L��Z^�<)ǌڳ�f�X�cN968T;jUQ�<��oN�YA�ْbM[�)�E�<1�C�	h`�3RC�[l����w�<sP('T��4'Wo� Q��m�<!�#ڡA��}ʒg[� ��J1a�g�<�2g��2ER&�8R����X�<)d�'b�4#�I˵c�t���J�R�<�c�$�HzfKX49�r1ن�ZV�<a��FyZ��J..w���&��S�<��o[�Q��})�/~nҁ8q@AQ�<i�7t���`�K�$�[0��P�<�cR�kb`X�VA�0�
�E�<���Su�:e v�[��T��>�B��4������HՇ�0��P����C(&��	�P���IWz+���,|��ċԍV]����K5�$sD��U�4��eH��X�ȓz����[E��Q蟎q�z�ȓoO�q�oĮN�PL颩b/�M�ȓӂX`lK,JG�$i2@��=<� ��X^Y��Z��btJ�Eсx����c"��f
Ð!n����G?*:)��Iʩ���KK����K;Y��<��$�:�bv�,-���u�ܠ2�ɇ�S�N�Y���*�cR�XW�)�ȓq���	d����|��A�ed�ȓ�,@V��8XL�#.�D��ȓaOΥr��D�O8�-&�ZD�}�ȓ;Y�1Q�o�)@�h5�~Ȇȓ2�Ա�d>ZI�H�tD�=E�̅ȓ�Xq��EbB٨���<}�|��m<	Ò��/a��EKQ*�3}(�I�ȓTA��h��V�l�+�(G7p9��[:L�z�j�-��)1Ɓ��xz\�ȓ\M�\���!��@����a�@Ѕȓ3+j) pb��[�a��a�x�m��5������:l �a����ȓ �XÄ��?�@�C���]=��ȓs����!�~�.嚦��^�̈́ȓ{��A�O�( &�8���aV���ȓ%��<����&Сj�"���ȓ}>|�b�_T�LAr�'�<N�Ĭ�ȓP�����R��@�S�ލ8����s�|I1Q�- �~L��l�>
 ���6���f�V�
��s4F��{����ȓ&�ְI���L�D\�G�K8WA�ȓQ��5�2FT�yh��9a��0,�8�ȓw�T��N޳e$&�)��N����#Ӕ�Bw/�2�x�"t@DVy����K1���Q�,�65)WO�톀�ȓr�� �@�gxة�r��.HՌ��ȓ
.d�bgʊ���[4��g�\�ȓn	�h��I'���{�%�=����ȓ4�1!R�ځn�ifN�<{ �l��S�? ��ʃ	���|CWJ9H� 9G"O�D�ft:�2�)&a:�9CS"O"ɘ��¡/�&�[fH
 W .s�"ON�c£KY�l����G�y
�Ek�"Ob�:G�P�e�ࠀ��T�1��S�"O&i�E�$(���v|�)P"OL8sЁNZ����@?v��Y"O���c�uxv	�y]2��0"O:͘�i�+����c.�-[�8f"O Ě7��9 ��tP�ʐ�YM>���"O��2w%\����w�,.�}X�"O��+�*Y#x�zl*A�T "��i{ "Or�����j��I#T/J03~�� �"O�AA��α0�b(%�E�	i��;�"O�\�U��ȥ��>A�I�"O�D��AV�=�4E1�L_�N)��"OR��C�*���r6S�VH�pR�"O�P�`��[��D�Z@¦"O�xcXVt��6��e����"O���ë	�a
�a`B��;�`��"O�=�g#�73_\iC�(�x�%@�"OZ��1䕮lU6���[4l��9f"O�Q�P	��BzM�a�'�����"O�\���
viB<i�o"�е"O~9di��NHK��S�+��0��"ORL@�z�����)��3�����"O"ɰ��U�X|\r�H�g��5�B"O�H(����,�
�
�'�r�r�"O:!oȂC`�g�5S+R]:t"O��eH��**6�"P�H�B^���"O�
��+(B��GG�"�`S"O>I��+�.%\F�*���Ti %�"O��I��W���Xu'-UY�l6"O���O��,��07L�r�8��"O�d�VN�E�KĒ-_�+6"O��ia���i)~���W�qnVȺ"O��J"���O���9 ��1nXNĪ�"OX��U]�Υᄁ�����c�"OF��E�L J� b���M�ف"O�u
b&8�8�� /�(�E"O6�;�"�8�X!�C g��jwg�d�<!䍂�Dڸ`w&��_��0zr-�d�<iw_.^��rc�E�N�N}+��z�<9�Z	W�lP���;H4<�����s�<Y��S�����-�6N,���l�x�<y%-�'{�����9U��9�s�<�င ��xz�K@�+j�m���]g�<�'':ϸ�1! )�B͑�)7T�lJ���R�(9g�0G�ʐ�©,D�� �atڍp`T6i��D�'&D�h�cm�����.Ph�b��>D���&	�pܑ�%��v�h`�(<D��e MH��l��:�yZ��;D�<I�-�
EF&8��5��(b��.D����A�p����&��R*|��F�.D�0��=+P �f� 4"��f�!D�\�!�E�
���H�1MW��j"?D��A�ȟf4H�7���i�,Dx�C<D��B,ʼ^��$�#�GO��Mk�<D���"Q2i��j�KE�dD�yЖ�8D��k� ���u��(���N6D��a��.N��QLB�`�ၣ3D���3JQ#�B|i��׵H����f1D�<¡=G�"�;��к����e�<D�� � �g�yn �@N+&�F�S"O&tЄ_�t��ը��Wl����c"O�"3��)  a𷄜��"Ou#����|�'$^��bp"O,ʣN�y�&��S�̔+�`Q�"O@ zuƀ�L+�����F�~��}��"O��Yc�,�ִ�ڤ���F%D�L���@��θ8&�<&�x$D�xӤNR1 aĜ�ӣT&���Q 6D�@��Ļ0k0�{⬑M���xq*O�s4DŉRQn({d�ݿC���v"O�Scm�
��Q���\n��v"O>�0��E�7רhðř�&a���#"O�Xү�d��-�`�SY̩@T"O�H�Q�24&*�ه�P�y����"O` ��%e�zT�0B�	�8�"O�<�F�@��k�n'x5~�"O�AQ�A�[�Z�0�^�$��"O���F����[A ��<�u"O ���G�#c>��
���֑��"O0Aٗ��G����H	d�X4aB"O�RЇ��<I�ɣKo m1"O��AE��~�` �	�q�B�@�"O~}[dJ�.�Qc�G�81�"OB��Mm����ҵ	�t1P"OY�,ٽn�tM���I�L���"Or�17��'qt����]�#p"ORuط��:t�$I GҌ��\�G"O26H޿j�$�@�
;^pp�z"OniɅ!
�5��J4*g���3"OD+�#(c�mJDHB,�`�
�'��|Sb-#2�Z��C*zr���'�]��
#d.�t`�͉? ���'�"\����i�z��B�<�p)!�'Zh03߶;�\9yq�_o���'�����Ey��0yQ�K��U`
�'�b=1�_6h�y %Gk��	�'��Q���$m�&9q�@C�>��Y��'��i��!�N@y����4�x�Q�'��a��'1���*7Ɨ�,�&5��':N%���[X��:�!�� &��'k�c���P��U����:	�'��lɑ�N2�"؉ �]�h�	��'U(��F��9���������'��ŀ%�5!����� ��'I�!(%J�"]ZM1a�v����'l�y���S鸌���Qp:jLH
�'o(p�-�JWXq8v�H�q
J	��'��i�;<#f<)�ꒇ���c�'ඬ{���,��ٵ��,��'���U'X+$�Re��s�X���'�|x��K�&:����.��;���B�'�TI�֪,�<���\�Δ�
�'�ph�� \24��K�Vu֕J	�'䉒��Z���d�Z�U��y*	�'�^�:��ٻm�b5�ۻ����'t�RS��"����֎���R�'�jR�=ݺmxćd���'n.�A��
Hz.�I��A�y�$@�'�µ�G��	 ����Y�&���'�EQS䘡i�:�XT��7e�^e��'@n4h�ڳS�h�hr)%F�N��'������X��oD�q�"�c�'*�F��$VY@PlY9pNPI!��� r��R���k�]hC
K3Ԋ�:�"O���o��#'���Sh��*���V"O�xCa�Cz��)��P�rL��"O�u��lՎdB��� �M��U�"O�5�P&��ZI���W,~�9�e"O��@/ݭd���ۖ���~nB��"O�q�PWh���*�cP�o��(0!"O����U#)K�(s���5�PRv"OH���- �� �_ ~�1+"O��s���O!����)ں#�<{T"O~`B�GR�̫��_Z�l�"Ot�ɖP�( �	ڡZ?����"O�@c�Q�O�<���c��5,~���"OV��W�\�	�T�X�KQG[#�!�O<��ᙁ�
5v~[�fW�$�!�d��ah&�x���2T�|s��$N�!�$�2��NO4V��h�&R(o�!�Y����Q�X�f
.��1L�:o�!�D�uH�C�	*���F�5�!�d+W�pس���r�j5s�v�!�]5|��]�Bψ9�L�C�l�P�!�䑏!.��2�K�Y�ld�L�'5!򤓣 ��t:���_�ta�k�R!�$L�v8=	#k�70�<��i͈&*!��[��e:�NϾ5�1�A�K�}!���*/=x%�ʓ�ų2E.3�!��d�ԜSkͯ:8�맪�D!��&j��AEOS�t��9�b�GZB!�X�R�,�R �
oպ��6��`!�'Y�=҇)E4F�(��)Cs!�VNI��Տ^.Y����W!�ܴgÞ\�JN54��0��/F�};!��=Qb��c������pHB,i,!�ėh�� f�η���k�a��
C!�䕓%wPHS�E��r��v ٸN3!�$�	]��F݌v�Xi���4!��CwJ�v*�hZN�pP*IN2!���2% b�ͭ?jt�qbٌJC!�$�#D
D!�� l-n��G>T�!򴲰��.��%���U(RY��9�����~�С�U�X�W.���n>�;�ʐ�Q.�¦E�{�8�ȓk�	IpeL<�4)�f���*��	�ȓQ�<榚NٚR��:���ȓ��%���',֐�����#�NM��}ކMJT>k�L����_^J��ȓH�>�C�.s�D�1�^c����/�^����3 dt�Ҡ��:+Ņ�*�� �2 D�L*�1x��-A4���ȓ;��]��Č2�P8� �,>*�I��(̺���A1���P��Z:,ć�JJ"h�����sF�YS^��C^���[f�`��/��.�%��qAR����8%�<;L%8����Wd0�BO�1��9�F�)����oe����@� F�L۔�/��Q��k/��@4�^��Ė�Q� ��pZ@@�-J�3�[ GW�(�m�ȓU*d��A�	d-���rj�<�u��u��xz��SF�mb�$H A����+�"r�=.�~L
��ΰ^���ȓh�k�!�1VP�w������ȓ
txש��mhD���Y�)�U�ȓHۼkҭ�O�0ty��'2Bp��S�? 4���Ɔ�s��YS���d�H���"Oܜ�piP�|Dc�� �4�6"OB�0�(��:�,���&ި%O�pz@"O����
�[cL�aO�qM�!i�"Oz<��D�3�$��Y�|�= s"Oȥ�F$��M��Xa �*t�9�"O�<�1�R�=_�RԯL�tn�ѓ"Oĥ(p�ҭq�����ōD^�'"O��q*L?�����'�Z�R�6"O<UjaEB�\A�=��f�$�P��E"OD�"�a��*`�(C��.CQ���e"O�9@a���qXD�;6�N-�5�0"O���mF�?�����w��tS�"O()��݁S�%�B�L:���"OLU�ᐣM%��UM�-2�v-�$"OtzcM$Q��a(4L	9'a�d��"O65PУ�gG^ЧD9&�֥�"O�L�B��<;m�#�(,�4%�5"O�=��,V[�F�9@�Z�"O����#$�TJ2$�Zl,��p"O���e�W>.r�p��H�O0�uȅ"O�i�Zn��I ���t'@��"O�!r����T: ��Rf�+H�Y"O����f�y���9)�R�"O��r�J�]���iVo_�{)��"O���p$�-�>P[�N>9�Ey�"O���v���`y�e.�;u�N���"Oި`��G�M��0v'+[�P���"O��9ѡ�
c)l�Q���4��"Oh���勳PP�AQ�Q�DUSf"O�AҢ�$K����o< l��` "O��+��  �\���6f�ٓ�"O����Ɵ^ئa���	� uHv"O
�""�ޤw�Ązq�u�5�R"OLy2E�o��r��R���xV"Oj,�E���$h)q�L�b^5؂"O�@�J�w킨�1���J^l%S�"Ou���4^�hx:Ej��ZXf�� "O�mQR�]��P!q�V�Rf��5"O�`��l�`Q��(N�$+<�"O� w������U�D:,�$34"O0�Q(˹f�N����*��2"OTQF3?A�-�`	��p�22"Ol����Af�p�`(��R��d�T"O�U)£�\�&��u`���`p�"OYi#ƙ�JȐ�A8U⚙d@l�<I1�ñ0<
雑'Q�D�~�Q�j�d�<���78X�1!I�`�X��GJa�< oā#�~��e�`U0�cp'�Y�<�r�<a���@,�*q(���N�L�<)�o�^�,a�%�҇27�3@��H�<	q&תR����e�˺4�P�5i�H�<�K|5@����? �0��D�<a�M�a�f�c��!��1�"ZB�<�P�؟)��ys�"�[��`�T��c�<Qw�I
�Z̀`BK�
邤�V�<��኱O��h�eI���ܐ���B�	41tr�#O�YZ���+ f�B䉭k� }bd	4ϮM���ʇaxB�I��n��Q�@�O6�8",].�hB�	 "�e���|y��26nZ�fpB�&#T"�3"L�*LyP7	[ܦC�I$U�x(���?�!��d� ��C�IKsXc�&�,C���.~��C�)� �`����l$x�j`����b�"O@���ԫP�(�s��ӳ:���*�"Ob����ȝF��<�WDþl���"O���;����S�$Wqi)5"OXRAȐ�%�hy�FV"=�L4��"O� �6�@�0E�(>�5
�"O�x�E�~�X��'���5�Ez�"O�����A���v��}��"O�u�S��{3��)�@�}��"O�@��G]�2���������!"O��a�`�/&�*���H�:)tX���"Ot�s�@��X������ٝ:��D��"O�HS� �q��m�lԫps�P��"O�IwDZ:~f�� �ä:�x�Yp"O�<K���73t�Y5�]�l l���"O��p�l	�ms�}�$EX�+�Θ�"O��g�bԲ�(	�n D�#T�(N�(W��$SBH�U�L��"O�Pa��4N�ʌ`��D�\�l c"O�f�]�)V�)C&�L*FH���"O���&�P>
`Գ�a��8�C"O��Z1�˂ �0|�ˊ\���"OJe����5"�@�� �ZK�"Obq��.*Q=��� �0K��Dia"O,�C�Ŷ� HY3T'�a6"OJ�h׳ �t��3��d��"O�uK� FY��ԫ>D\UQg"Of��v���m�����F^r)0"O����J��rVH�(Y޸��"O�h�Aޥ5R���UI�Y/��(�"O��R�O��[�P�d|�ZW"O�0�AI�dG��3�hQ"O�c�K�:E�����m6`Yg"O��p�A1���Lބk>%��"O:����4RV|0
��A?��@`"O�)�S���{�6D�F�ĸA	�yR-�2|����.�.]��B@����y2%H�y�<�qf_�A�H	(0�P��yr�:�R�,�c��b��д�y⎔�k>�k�D��i͠������y��Ce^��c�7�H�i$K��y�%�M8t���1 R�9 ����y�KW�L>�H�`�X�M�t�&K/�y���=a�T(p�� H��0�H٤�y���l�a�P�լD_6�����yr��6irm"#�I66,���.���y&ًt����Ӥ$Z�{D����yҠ
����RAҶ,���`^�y"Jy�B]x�a�����#K��y���?�~�A)�8��)��y�+D6 ��x"Ɇ*�)���]��y�(���_�j
d!ؑ��4�yR�k���6�
�^g֕��e	�y� �(a�J'���1��yҏ�5����ʅ/�VTh��B2�yB���
� T�Fnǆ%dBL�Q�G��y���!z�D�c%��!�(��eF�y�a:�0!��D�cz����ɼ�ye�}rfH!&˅%Tamb�h�-�y�Ht���(��?LT��KEf��y��ƕ�$���*�?zv��T�΃�yBJ׎f��yAS	�@� ��ŏ�yrƟ%|��	SD*}	�I�<�y� �@ɼ`�q�S��,x�A���y
� ��Bq,�I6<�`�H�(8d8��"O�J҄u�x!� 8FJd;C"O4Y��`˻E�x��=����"OFhhƶ8�h�3��h�
sQ"O��)��F8�Rb$�N��	�"O�����ܺ80�z��O�F� b"O��k�OκrU�t���0|�DQ�1"O:��s� )]�G���P/�PE"O
Y@;4~20qG/�@U�g"O�-b�EZ�Fe8�P�3���"OT���۸L������1}ۺ�9R"O6�sm��F��P��&Q	~�>`�"O��(��"e��t��$%�x=��"Otػ�l��:�E��YJ� A2"O��#��i��pB��$;h�"O�T
�	�%t�2)�u`F8��b"O�x�����4]�Kt���	4l��"OBQ�)�@x<� �aR=;�d(��"O��0$� �g��� �K���&"OT���$Q�?Md�� W�Y����f"OpA0j�Jj��cr�!�dHA�"Op���BD��i)���8&�6�(4"O�4�2�G�t��Lc�X�2�"O�`��5*���V�2/�bm��"O@���H�l���5�>0�`4Ґ"O����⑁P�,prS��*�&�"O��J��߁)=r�����!g�(lB"O^(��>%#�� 2*7��h�A"O}����fr5�������p
�S�<ٰ�(�L�ٰ.U3s挂��P�<���0t�����lP�i�@[q�<q��6�-�%��\-���Ek�p�<Y�
Z�ܑ�J˂*���co�t�<��A��?��C5&�:n����-[r�<��ͩ5{(\���Vg�X���t�<�s���_�H3�&��7�4ݲ�&�m�<�4�"�^�H����V1^�1��Gk�<�s`P�S@���rBF�H��8js�X]�<���'0F�X��6�4��`IZ�<1ѩO Sd����J�$�n9��c�T�<�d]ɰ���<$�t!+Jv�<Q���8�&|H'珷y�ZD�3�Np�<Y�g��#NT�[�C���V�"#�d�<���ƴG��=P橒?Yk�mr�%�Y�<����� �P�K�;(�0�s�fM]�<!ũ�y.DA�P�jl�(��Gs�<�c��2"<P}��+�jS�����f�<���L����8DLX�gV�,����J�<Q�͕�O�m��!���V���F�<��J�8������²@�$��ĆRA�<a��������kM�{ta�p��b�<IuC�s��p)E�)/!�H�6(u�<	�!�)N7r��r 	iF,/�V�<Y�i�|�t�/�]�j�Z�&�T�<Q�+�"N��
=fP��J�<Qm��6ʨ�̏�W��h��C�<��ł%~%�,P,	�e�����%�V�<���D��*������Z쑄˔\�<��	�4)�s�Κut�)�HN�<�Q�9-6��l���'#I�<���%v�LH �N9J����D�<�� �0�psS�ڎa=����	�<�g� C&��o
���E�R�<ٱI͍E#(i"�Fː<�v5q���N�<� �a�m�+_Td9c��h,�t"O�!pk��O������=Jv���"O�,#�c�br@�����	��1�"O�������Ps�m�=S��"O:Ȉ��3OH��׍P���"O�
DD��n�U1*A
~��*#"O0�E:^!��Jr��o*<(�"OƝ!�+�s?j�J���x�Ux�"O���N�hliG���Fl�,��"O���##m^���FԺsVBt��"OT�[B�_�S|0�7�P ;v�+p"O�0+@I��G��tsa+ڸSR:h�"O��`�N�X�C�JR�t�E"O�@� 措c i��2]��)d"Oxa�f���e���)�b׆4�QYQ"O:]� �4"%bʈGn8I�U"O`M����p9���`@�W2!v"O�� ��Ϩ9����}�D���"O�)��Rd�|�#�Q�?���q"O2����B8}��˒�]6t{��ȓ�f�2�ɟ�Vw�U���*@��ȓ!��U($��u�����䒙/����jl��BF��I���OQ�B[D��ȓX�xy�e�)e��1L�Ѕ H�<�!�^/� Z1�ռpε��JB�<�!*�H׸��K��U�%�B�<��H�6���t��`~���7��{�<!P��!r�1j���sRڤj�HOz�<'N�*2��Q����e���7NNr�<����z�ʔ��GЌ6Tq����p�<!)C�̸�g�҈\�"��d�Q�<%f�l@x�IS�AIv�@I�e�<9%n��FȔ��@�HS�]�O�x�<!Q �$u�2�9�!�`nL35o�u�<a� lN�	#u+ш k
�J �q�<��L�T����q�%>�D�q�<F��v>���b�ɿB�^iBG��s�<A�5s�h�U�44����Fo�<�eOV)
��r��U�Jx�$�Ng�<	e�ܴU�
 Z�F�l��c�m�h�<��g��mj�`ʶd�����Ǌb�<A#J�u�P��E��N��]�Ga�<A�� ��4J��)Cp|�!�E�W�<1�р>�hq7Β�H�2���T�<���J52���ZL!De��C,�G�<�b^>�qbU��胖��j�<�!���0��}�cތ���ŭ�f�<qv�(�~%S�bD�(5�1(f�<)�W*{8h�XC�]�T0�f�H�<Q`��$?�MQ�b�@	���BH~�<����
6T0
fo�&m$���ȝb�<)6HU�a�t	��$U�Y�>P�3DJ�<�/�/8�L�P�.!a�r�Qq�Z�<i�*�X�|e)�nH$<�i'�ZT�<�MX�?�2���`څp"Ta�@T�<y4����0�׌^�@�P�)R�<A�^�\$q�JdH0��qb�E�<1�2/�����0���6  B�<YR�G{fp�j��-ij��@"�}�<��mB2�r0��.Y�FW�p	Kv�<)SI��X��
��!	3�u�
�l�<� -	9K)�)��ͣ� ��H�h�<�3�˗��, W�G�s�0+��y�<q�C �����Z�lt3���x�<� �D�t��5u�1sGfQ��*��"O�@RĎ����#��@�Z�x#"O���Vb_0}��-�F�+z�`@	e"OB�s�C�����d�߃,� �0"O�Hن���K������	�n���"O(5�ŧC6#_��Ciл>Q2ِ�"O49-TL��c&i� [�`�"Ov0y���DAL!j���H��Lh�"OH���:��D��FO�M����"Oz��ևۑ,{�kD0�L@"OVa(�	����3BkE!�<`@�"O��2H�6Z,:q��ɦM�r�4"O��
3,-YI��e�$u�d �f"OHJǢR=;�څ�եT�<�v�;�"O�t���+}��qrE�$`xx��"O*t�p���d[�b�:t��"OZx lI�'� x���*|�P0��"O�d���Zs�U��
�f�܀`�"OP<sHD�3*^X��O��.��(˧"O,�Rh�Bq�G�D��	I4"O���p_�#�x�)��@�K��8�"O`�t_�;��x���ʮ=��ĉp*Ox��D�,j����n�;k��]J
�'"\�vės��R�A�W�N�
�'��%A����dYy���HO&��	�'c~EB!��eI�љ B��A�(�	�'�b���ټ
�Dh�M�8ҹ[�'`R���B�o�� ��.��+t<dj�'� ��@;������x����'蚙���K-20�y��I|�`�'+��7B�'{�.� �h�>u�&�Z�'���F^`���qgNq���Y�'I�t�B�۴X<2pk7��8Y��[�'�z�GÆ;DV\��5��.�l�'B�� s��$�)�"��fs�ɹ�'����ȋ�m5"�C�B�`���'`��GK�'ҰuA�':eH�'��5aA�����aB�-���c�'�q��dD�{�"���P�)ݰ�'����=���\yDII�'���l��DLXMs�K'��1
�'���$��M�i���,1P�
�'@���H[(d���
1�M�+R���	�'�Bc��F8���$)ovA��'�΀�F
�8ٸhy�n�!�88y�'�H�G�?JR��6$���'(�p o�x�����|)~���'�����]^Iry�5.W�x�-��'~N���!� Zh��c�m++�H��'� ���	ߖw&�=S$N��c���x�'� l�P�������M�0U$�\P
�'��Ò.2D�>�H@��@� x�'�jy�AE	�75n��2��$9�*�)�'%�ؠ�J$|� ��"�'?�3�'���!�%¬iJ ��<!�4�'f�����[�^�R�PhO�(�Ɓ1�'�6��a��/G��|b3�%kؘZ
�'�p��N�Mją�b�@k�"��	�'U�1��ts�T��c�
z8ix
�'�tA ]/��x�֍F�mΰ� �'۶��k�v?�}�$/��k�d�
�'�4)��Q�IF�9�R�i�H9c
�'��9Q���>t���.il|�r�'�H5��91���갌�d;��Y��� ~��%��;R���U#/�)[p"O�iXÄY&��B�fֈ,/xaz�"O,b�^����s��5o $���*O&-�ƀ��d��2<��'	r����N�x,Bb�*wظ�j�'g�La�OC�O]�\b��ϒ^_�$a�'�4��T�M�zt &� �#�jԡ�'��k'��E��A�6�ƈ<)�'��4
��=4�D���("�8�'d���G�m�h��D�ϱt����'3\�Jv��p��R� �!n�Hc�'�ܸ����&�q�GO��m��S�'�h=�#��f��Ƀ	\'ag�i)�'N�%�7Ȗ�r����֬��(*R���'��aH$�ȳr'�U����v0����'�6lpq%�8T�sBf��i�F��'ј0�@�ta�y����y��|��'MT�5�[���G��U�*>D�()NT(}�ny�m��Ay��*3=D�8w��+M�!
��@��Ke<D���X)ö��W8ʎ8�#�;D����;16�bU+��)P��ᑌ:D�X���ŰD[d�"G ������#i7D��K�����Zu��3\�%��l4D�$+R��
I��l9��^>{�\5��!/D����Y)4��UhP�&nXi㔈0D�ز��J�S�n���*?��E�+D�j���zd���;2J�h"M$D���6�E������ATYvZ ! �"D�@�Ԡc~�8���| b�z5H D���F+X�bNq���s,!�&j>D�d ��:d��CˌB}��J�:D��6�ɂ4�1j�˞'3BAɁ�<D�TY4hQ�x�
	#�el)�L(D���# ��Nt˒�W�yf<Q%	&D�lK�lY"��D��{0�	JP�>D�(Z�!܎g�l$y��®f(*m<D�T�t�̳b\�p��?v��x'�-D��KQ�nJ<�t�[N��!��7D��SⳔ�;dͅ���1�S/ޟv�!�� ,zиzB+�;f�j�	Cd�U�!��/)�ܙPt.F�g.r��db@
J�!�$K 4���Cŀ�R:�Zk/k!�d�z89*�"�2�i�鐀1b!���#8'"|1�g�4Y(8K7h]�]^!��Q�A��Y�ʐ;&܀9R���>�!�5=J��P�J�8O^�y�`%I�9K!�$ǵ<��AD�^\X��DEII�!�F�Ȁ����:|�j��!�dZ	+uD`0f�-����ɟ7;�!�$��t|�pMw�\@�WiԢ�!�xY�\YI�|�+�i�!�ʑ.�*8 Ѭ͙,�f�`�G$�!�4L�AF�ۣ�>qp����@�!���7�`e��O�)��Pr���*�!�C�~4�?���@!��B&Sh��"I��o��@��%.!��ׅv<�#�'��}b�Z��Ӂ*�!�D�(��4X2�1��u��!�!���u5H\���J�z����TQ
�!�dQ������Tuf]E&�!k!�D�e� `P�Okx�kV��9�!�d��p.�8���Z*z�N�r�̅R�!��Y�!t[!��X��U��N2LY!�� �ݳ҆��F�J��QGZ�1�����"O�\Y�G؜���ږx����$"O�T0�R��-��k"��(!"O����	�|��c͇ ��e@�"O
�E�+B	��ΨlxE"O�l�7kZ�U���P��ZgĆ4B2"Oj��$J�6����-�0s"O$�@w�	�'1�)��^�$�Z�"O`�B���5�+ы��iXv"O��A�hԤO�a� ���]��EhQ"O,T�4GǹL&��萭>���)A"O|ij7����X�� �*^�T�"O*��J޿H�ՋR�B:~< 4"O.ha��[8-��X�E!�?	��:F"Ov�p��A)�z��"!?s ����"O�)sw��	a� h �@	K�]Y"O�����kD�TÀjD� FT�p�"Ova���$�2��3��&"OĹ"�`��
��Zu�b�pإ"O"}pq��j�=#�T[`s"O�iD�3Ťxr��ΟJ�H��"O���#!!s�$��CɈ�;���"OP(�q钑B����"P�9 e"O�p�,L3�8i$H�A�$�1�"Ol��4Hda�hޟMk��xP��!�ĕ8��٨�%ӾB����Ƌߐ;�!��-��jrL �dT����,ؼY�!�K�uV05
U�&���X�5�!�$�b�L@�a�zt�xRҦ6q!򄍘9S�L�1�A(h�};A�Go!���;P��ᆇ�9:���D�n!��Q�$� ����*���	4���.k!���`x,��u��=�:��"W'2T!���<YX�H@�ג���*Ìۉ1t!��:	Pٲ�Mݠ=����эN;V]!�Zbl�-X���h`ٲf����n�`Ti�3$�&/G�M}���&�����8Dl�����1*����?=p�3�
�*u�<U�5g��S��D�ȓX�V�!�e #�-��K�))(�C�	F���G�����Q��4x.B�	)b`ex���+�Bשм��B�?<�2���B�,N�܁R��!>GjC䉡>�Up��M 0��
��ڒ�0C�	|v���������1� N`C�I�7)�p�IvT�l��!;G�C䉠x�@(i�G]�oP��vP#D B�	/�>m���Un8ApJ�?�6B�	��p`$i_O!�`��͜h����86��i� �4�����~!��>6N�Qu�')N-�TK�(L�!�$ɔDn����E�F��(�L�=A!���B���ݣK�6i��e��E
!���YHQ�ү��Nj�<��/Mf!�J,������4zv�r��5m!�E,`�pMHu��p[�e1�%S*~W!�d�K��a�$A�g]�ܡC�P,"!�$�k0U�"@�6`<��hڵ: !�/}*�,���]/Сڥ��9|!���q�� �N�)�1`45!��=|��vFH�wN�!�$�$+�^u2c���E[�a��!�DC��&�zЂK[���a�D?I�!��1E&��;�W1��0��.�nv!�� ���cǡ�t��VЮ#Ĉ���"O��kPc��{Ծ)S�I��}��"Ox�8Da�]�f�1X�&�@{u"O.���N��Ρ�Ԣɠ=�-z�"O%�r��l^X�� �K�P��"O�ui��P�n4=(wbٜi�����"O�-h�DD5-�q�0o�N��"O>�cN�4i�����ǫ{䌴r�"O�D��JJ�G����@Ao�1�"Oz٩���C��;�-ӿm�H��"O�<q��2q�&�Q���5|a�@�7"O䑚'k�OD5���>yZ<{C"O�2��b�]��aǪ~w���"O��ŧÇ)�4R3�T�+@�+�"OZ��eݪ �J9( ���A��!D��#QN�7nyS�*�
�x��+D�� ����RU���=	�V@�ǡ#D�ʱ�JLR�-��	����� !򤐐J���`�HA
e��L�7�B�a�!�BG����R�N���Q��$j�!�B8%��G'8� ��E��$�!�Ė�K�zxa��O N�jP�iL� �!򤞻1T��Q�oɌ�0�ao�7�!�DҖ+�8��,��H���%���Q�!���*�@څ�ɇi�pDh2�D�X�!�H���|�E@�D����6虯7�!��D�1�R��$Ct�B� �=a!��K.�	8e�!�P�Ss�%N!�D�-�$�1p!�������A"O,���o�#����C܏*��Q��"Od�pU�7&�}Zƌ�x�^�R�"O�a����:���{F��%$���"O������_��년
D����"O<��B�P�K��eA��.NȰW"O�)8Dm<hz�����-/��XD"O:d35�(��9JBD�$�Ш�P"O�����ѝ&�|��烝V��E�"Ox����I��	:T�<�6!�e"O�����f��YslN�*[�I&"O�d�mȁNo��#�o%�0R"O�qX�퇕Y�ʘ�J��%���cP"O ���G�mBU�DDK���"O��@4�Y+e�1�6,�)t7�A��"O�u�oT�clڱq�*� =%8T��"OѰV�2m��H-��[�)E!��E�$�`E���ͤnzL	2*Q+1!���?�L�h��ħ"�4�q�ڌYA!�¯>�eR@�:h��CŇ	�e;!��M�'Ja!D�&W�Rrd�9,2!��򒁎
��I�� [�	뜕��'�
8y�fU�!V=Ihҫ7i��'�L�01h�I�P�� ����
�'��|�-��v������#
�'��� 
,�,��wc�z\z���'zJu�%| ���ƞ#v9>���'׸�� �Gƴ��kL'mܚq��'��iV�F��Fd��I�����'.&p�u��D��HOZ���'@ 4!1� �>�Ǝ3 <Dy[	�'&�D`�'���`:�ڤW
[	�'��PzDi��6�,tS�2f�<p�'i�0�'�])LF�JJ�#�F�	�'���v�Nb;~�	��0�Nń��Z	�����*��p�߆�ɇ�S�? Ɖr�%g�����ڲ(w��{�"OR�X�K"��l@�H�hfI�r"O�=h�/T/,����`f\T F"O�Q���V�]@�jR�pk���"O�� ��{�\����-`@;F"Ov�juk�D(tB�׈DPV�"O��8��%Z�,M	2%!�<4��"O���(I	x/��r&�\
��Q"O������ :�����%�*M�8�B�"O.]�T��w�����#*z0�&"O��˕��hp���Vi�W"O<9����2b# ��GI�Y�*�u"O x���<ko�٘��H�h��ei�"OLe)B�+��];e����@ks"O�p[�$k������� ��"O,c�iT2�-�W$	�C�H�Y�"O4�@$A-9�7R�7�HQxS"O�%б�קD�vb�)���W"O���� �"hW�I�c�["O��A3�=���3GX=@�f,Y7"O��h� /ml ���h��"תE7"Om���&I��PS�Dr�X��f"O0L!䡎�)�*R�8\�XQa"OJM�V�ٔF�Af��b�D��"O�x���S��L��i�� hZ-� "O�Z��,?�tQ�FP�HP`��"O�lc��Q�[N@Ӗ�L�0Ed���"Ol]�Շ/B�h��A��?��̩"O�и�H�m0d�A4��7Ԓ��w"O���f��% �CQO�c�| �"O�5�HΚi�b�ؗ@7]��m`�"O̕t��qun����W��j�"O�q��	�G�:�1���f�c"O��yu�����2T��"O�A�p�@�|ۆ&P�WƩs&"O�Y���7jU��K:�5:S"O�ݒu�(  &���0L�����'AQ��r�摬k�X ��$��N��p���<D�Dk��ۘax�����_&%���.:D�p�$L�@T�M�&
��ڤ��,D���L��fM�1���O�t��4D���"	Մ�2�9��:Kj>��C�2D��аU�F�J��s�2R^�l+�
6D��p%dGd�00p��� 9�i`�4D�<!�$T><�!0g�f��`�Š1D��T�E?'�0�8M�= ��d�������&��Х��Q@貁��=bjC��w�85+��R3|X@Y�k�=C��B�I<:��v�؛Tڑ`"�>ub�?Q���� 3i \slN,f��P���6 �!���Q�^��Ó�a�l���!�ă-� ���JV�|I`�)])$��$�/a��dAq�K��$���$]���C�ɦ	���rRE�ZjĔ-d��ё�;D�$p�L��@�P��+W#�l�f,5�	T؞py�,D#cɶ�k��� �Ic�5D��A��� 9������N�܀�@0D��;�DF�k#$Q���^�TS��c�Q���p��$/�PɁ.�?B�R�p"ORݳ����r��Dq��ݡD��H��I��p<�R�P����S.�2
�Ru�?D���R��Lgd����Ծj��a��B!D�p�1�X#��y(4�Qz����#A?D�$bE�n�`D�&Z��BQ�/���)� \�x�
�����/�-(����v"O��C�b�)f�1�F̗*�zდ"O<��-udDq�16��l�>1	�L����I�q��}Z�� �I�q���:��d� G�mp�M� ��+Q+�m��D4�Ox��&�|���{Q�D8@P� b"O�h+L�*��i��ۛta�)�"O=a���]���(vl&x)x�ʤ"O������#"����*K18(҈���Io�OZF�g�Ae9�Q�P��]�	�'j�Փ�DN�xё��E)[gPX{	�'Tȁ3��Wq'�����:r���'I�Qs��u����Y�� ��&�昦$ր�PC�@ ���y�Ͻa��l����G��ܻ�!L"��O�����.s�0��	O~@��al��AD!�6P�ڵ�E��(B>�k��ϵ
��	s��H����Q3<O��� 	,b���K@"O�)��Sòԛ�*E*B,��"O�P��N�o�vi��iC�1�q�1�'#��$	3@��l���O(j���a�&$�؃��;Z�l�FУ2�.��� ��ybǕ�Sd`��PLL�(Ĩ����y���zJ�jЋ��'�Fe�lV���p>ƈ!���)�e�Lk����i�<q��&�����U�)ڎ8[#FGi�<���+����u���*�!l�<r���Lβ*���4���4��c�<��bۏ�\�M5�.����`�<i�MA9%]b|I��
&X�cN_�<adႷ(�&���� -�� �����xW�6�&��Op!���y2+԰,��iu-��L�t����_+�y��@��']':E�ת�B�0���'8�
��
�&)���5A�qc�'Ѩ��>)9�,�P�T�,Z�l,D�X3U��C*�JŌ�&j�`,Y��(D�����5{�����Ӄ�V<J��'D�|Qw��U��K���pl���$D�DPD��-߬ht��3v
�j3�!D���2��I����瞉O��*�>D���SZ�nGz0B�[fP�E�G�8D������t�~U�t*��-���C0i7D� �j�)C/�-���8Ξm�3!)D����:�nI8�%�(QeV�"�&D��1$'�N��1r1�Z�	��4!��&��oZ$*L(��"��0d��J��4mNB�	�mN��$*C>:j�u���TC�I�A��y)i�)�I�  ��B䉍#�N��mX ���w �sG$B�	4Ei؅;%��]t��O�� �$C�ɲ^��q���.1@�j'�L�W�B䉸
�,t	�+!2�dE�c�� �B��#	�Ad�B/�^�h�%�'b	LB���f�z�aՋ,���/$��C�ID�=�0>o�����M�)zB�Ɍcz�a�Ė;9�b�Y�dMfc�#>A��)�a�j���&�=l� 8�cS'b�!��H)"pEC�-%z�����
�!��xk�0j2c(y~ �D�õM�!��9{�<���˯TZ��)���
�'���2�p�vc��Z����	�'�@ѹF́#�<)�=� ;�'>>� ����� �E�� Q��)��hO� 4Yq��7^��d/*�8b�"ON��0`��$�3o�#m�PM��"O� r�-_�2 \� �m$9�\���"O����D�C(D����r7���&"O�`�
ċS5�@p��&W?��b�"ONP�c��>k<�X�-�10����"O:9�i_PW܀c�+�n��R�"Oʕ!f�X�=���F�۬� �"O�$�w�?� ���΄K���0"O:㦌+^@��s����f���"OB�㒠O2d�	��MK>� i��"O��gr��p����3�r$c"O�X1�䋛uS�\[6�Ęr��x���'��D�7|�<d���S�]+s�\O!�n�d1��l�%��;gĂ\*	�'�FT��)�|��aP$�� �b�'e�a��*D7) ����Sf�pa��d6�d�ta��R���i�6V\	E�	1bB�8m�	
�.M.R�ba�uҼF� ��2�I�t�|@�(�MD85r��KB��C�	:x�4�P��+ ^B���(1�C�	�s~fP0�]�d�p���hӏ(N�B�`(�AWe��@���B�I�N�\j���S&��Q�aI�T��C��)Ҭ���aZUh�03녏	
�C��>v?(�Bw(ĽL�,dq0#�[i�C�I�"�`z#E�	?�8Ł� >�~C�I	T]�J�Nӛ+\P
�f\9gC䉊T����Q)@��!IrY}���R:�H�J�EԴ�;�lEz!��-d��Đ��C^��@���p!��:_�n�pT��,�K�4f!�\-W��tZ#��y�k��A�kQ!��=ci�)��o^z��k3�6Q!��]��r���@^�u���ra� ;!�E6l���Q0#K�Sh���Wbҋ+�!�d[$΄�H��>p���P�G��!�$ؗz��,	 �'9�U��)	x!���m����+�(/�$0�*��Tt!�M.Wʕ�������"�ʆ�:q!��Z�b�����!����5(�+S�!�d��g����E[e�d��463!��7<ǚ��N�M� po��!�$ڔ92�)���S8-0z�K�}�!��ХD�<z��V1SL|�cP���!�|���RID�~:��1E�;�!���?���pŀ�R�$u�ǲAՈC�	!4Zp:�.ɯ�6�iHI�{�dC�	%J�8�g�W��4dɥ-��0C��Y$�4�S��c��}�C�	:�02r`�g1
8��ٵ!��C�	bh�҅'�0X��!F!5#zC�I�-H�Ȇ�C*	xZ-0�DH�2C�		R��P�tנr	x�!F��7B C�	�����js48�oE�x��B��?
��T
gl�:r���PՎG6�C�I��5�����5"
q1��5z��C�	)h�����*��Q��^�C�	�@Pl8���U�ܸ�bF��C�I11��q��ϝ�T�r8 �㋐�nC�I�t�	��f?K��I�C�X�DC�ɺ>��i��m����w�C�I�;����7(� !>�����R�A�B�	�d�z):&L�����5��14��L0�OV!d��M�aIH=[����� $�jc)��a���p�.֡
�\qG"Ou�j���*��j$���"O�9����f�)��%vU<��"OV�JqmƑ2���e0K����"OFm����97h���G>�"O�Ѓ��8,"�	�e��z� [4"O6�b��g��`��G��͋g"O(I��f]<�<�*�H�� i�&"O��R6E��#������6@��[�"O�P@O"i.0�0f�2�pL;�"O@p
`K7������%6�D��"O$�۫cU@�:�"�3/�Nq��"O����d�)d�^��q��#0�	��"OP�&`�2�f���]�L�C�"O��!�@ͬ�����"0�	�"O�d��'AbM3�g�����"O`4q�e��Hmf�� և-vаG"O��������R`�;
*)AQ"O~e��DԭByRw7u�^(�"O$�������Ò�?���A�"Od��x�V.Np)h�	[�J�!�D�tZp����%"�J�H��E�!�d�>k��Z)u��q���	�!�ě�I~��b2$խEBJܢG'R�~!�d�U����}��MÕG]�
d!��FI> �q�֏r��,j����{]!�Dω���f�;lK�X�CΜ�4!��:6�	���N!�5�͔>9!�[�#x�A��b�4ޘ��m�-0
!�$# "�!��Q���bI��6;�C�I�)^f=s��H	r�"L���F+gΤC�	6��ɩ�m��b��ͺ��EV��B�	T�N���`��8�E�ǆ��R"�B䉔N���� +%��z2� B=�C�	�:pn]�7)&���Ȳ%ݜF��C�	�i����p�@-�؁�Ac��wbjC�	9{a�1��	j��I���S�(dFC�Iz|�c��R�X"�xH��U9:�C�	7�|�v��sθ+�-%ihC�I-z��b��#M�d�4�KN@C�I$;jS�ѥWe�4��F�W6*C�	�y���r�3P��4��ȝJv C�I;p,`4�&l�� (Rprס�1m�JC�I�i_�r3�D1KkH�2ό�Ab�C�I%o��@�'�#`a���h��C䉞j7$� ��0�P!a
=�B�ɖi'����\9)�6�xV�`F�B䉎_(�Y��H�S�6-�P��8�B�ɪF�1�Ab3s^<	�a�� �B��D�L��@�9.$-"FJ9+JC�	6Q`�Z�	�^2)Rĩ�n�6C䉛"L8�2�C37��SFz~B�I[�~��Bc<1�m�q
nC��)R�a��A�v8\�ũ�G6B�$'�pL�QA#A:��(�"�<B�	�R��E��0�,�8 �U �6C�<���G�'n�����E�	�lL��%��A��m�@�����d�7���ȓ#ZT*�/K2����<�x��Ul��Z�F$0lCT&��n.x��ȓ$j<i�&��!: 1^-|+��Y��AQ�n�(�	���(T�萕����P���A]>���I�	iF��"�
@�E�գH6���΅!Z���jQ%B�]P
��t[��/��|C�E T��(r�M)4�� ������?r�͡��\�h��]��|Ҥ\j��E�m>~��e�c_�?���l_������qA�%��?���J٢�!�$+M(�����X17��w(B�e�,����k܆	K��P){�.Dy�JҫL*���O�U��,u���`B�  �����v�I���3�hsp�O�����O =�l]�Ef�&x�8sAa	�I����Yc�|��G���ԱtoA���'����(�N0x,���R�#y���0ݠ���Of�,|�(p��W�sB�$��9Q@���t$�1N�xi�N�B�6�+ed��KE����ǘŦ���&7%� P�D���u�oNl�2	�O��p��7~�X�愖�)��U�4@�32���,L�<�����V�,�52*>D�|�d�סP�9T�`�sD��7G� yJ"��t�d��;G�|xcԯҦ'� �7`�d�S$*��B����z#��P��f����@�sF�rd��y$�!�@�>�� %�@N8�B��iŜ脧
�\Q��Ȇ[��,���Kr�!����U��5���ȖJèT�`8�P'�G���?�C��+	�Da�����b��?9���)�J�ێh�.̑2�RC�]x�(�aMI*��@�' ��ە�{d�:e�R�J�,-�-O�y�a�U�M09�d`֊3�`�.�:ܠ�U��M�t@�5�p�r�%9�||�4�ƀE����ʕkh<I������`��w�n(q��B(c� �S��K#?̥hw��F_"�"�� ����Xw.֍�1�P���C���a��� ��3MQJ��"��@������Z*��j���:^�EJښ,�ѐ�bI(bӼ�a�]�����a�\'��
�;��R�9+zIK{�ʧ��M�џ��E�[��)s��^`.u�d��R��AV%�&��:��P�V�\%��g]@t��"- �Ma�1����R� Q�q�tAV�B�B�'BL�{T���^�)se�����p���?FX"A��Q�T~������ "��<����2ZG"횁���!���
\�4$�tgI h��Ap�F�1fV�����!L|�(�v�^fg�={�&_�<(�d�O��YHF&��k���!H��k��Yl��آ�l���l�!"@ �"v�\�3�Kb���kG2�" !A)e)�Ex���"[�����(�zƢ<�#�{�EJ�~�)�D�!�&W	�n�?��o�!@&�Y��S:O�a��E�O��q�e�4��T#�H��
(J0HW�Q%XreYS��53����$�&+r(�1��6K@��
�!����� F�Mhr��S�4�f�R�>ĸ@�DZ�&$�Hb��ϐ���e֬yD M�#a_�X��C�7�y�$��FD�ȚTJ�P���C�����/Ox�yQD�6`�R1ȟ��C�	�i�کj�'h4X�d�)�؅����%X�3�Y�������Ɏ�8C����d
W$޸��ɉ(-���ٓD�({B�T���9~����R�O=H�OZ<����7~�0����Z��EJ��ɢ~)\����}��:7�ۯP�8�'�7J﬈�6�̋�0���=%Y'��*j�����2����䊋^e|�5˷OB�Ͳ��]ɪ��/]Z�X����D��HqL�Yjb��ť
5KE�Ղ�D]	Φ��UF��X��BD�U��^�iA!�dV+hB1$ꖸ"@X�r�*͉u����&�U�D�x�kr$�,�ִ��jD= $
V9!HL�*!J�
rΠ͘���'������op  飇[�s(���ɐa´�1`dm7�Y�DB�%����SL�44G�xP�C��h����J�?�\Yc#Dͅ3(��!)G�-r�ಣ�Է2J�D(�"���O�Ԍ�qn�-��H��\4|�I�.^>����8k#�h�F�Uv8�ъRŒ�n����b��m�^�D�ߔ%�`���qatC�~��,��� �v��uKPQ2����%��厝��,�bg�U|�an[�\��5B��΁+��0�@����n�#���'�
P |ʑ��4�TC߾ sspc[�cz^݀ $$�O��@V��'N"�yqo�8V�;��KnlH�����Q�#%q�F��"I�K�D�3B�{�r��2%��@���ΙI,_2lI�AG�22_��EB��1��YЧ\��H��g�-um�5�!Z�i��I�3�&U@�b�#�͋�ɟ&<L����ŭQ��jq�?n��u�?�$��j��}����:.K�Ȫq$�ɴ,8T�����%�ح�M�>s��i�2CDL�������7
Ĕa����'D��_I�d�A�G'�^pa�	�|M�ܢ��'�y��II�-#�.�,��a&�S�5�d$�U�L��b�AEd���OD���*�扚U���邆�l5���LU�KFt?�����"t���ȸ��`T�P��ӑiz�P���^B�[!%��(�4�	ܔ��=]��b�fd�(�N�v>4p�DX�%�d�rc�2��O�5Р���d�t��" �6�����Bt$r�L�3�v�9�_�*�"�1�'���{
�$��y�R��D
j
U�>4�h�%��v�^�O���R"��sCj�c�<�b �j�)��,�s�����,/������� Q��}H���&�0X����k�s�5hq�d�5��*ٛ=�hu`�'4�ǁ ��<ٳJ��\� �U��Yt 0 ȍ9�HU�ea�[̀jE�� �c�t�(�a KD��'/y�$Q��h�KL5C)=��go#,���D�v��ە�@/$������>H/6�G^�_��RRN_�+����9~���%��#��)�b�� ]R���F��2j�]�c*�X�ay�튱g�ܼ��ԯ*�B9qt�7i�>a+Ѩ�9����'�n�x��n7��dóh�i<�FA�o� ]S!H�7>��b�|���ҕL�[�B�׷3X\�2�?��W72\P�B`��>q�T�B}Y&�+!�}qp�B�x�����o�٢�KEK�Ɋ`��lK$Q��A�>�Z,���:\O���M)&T�u�5��!r6x2'�_3i7Ȱ*�$Y�%Z�B�w��-�6�![�Y���Y�w t2ʞ�� N-:�+v�0�/ͰR�dpfO
�@eiF-Tx8���.NF��5"'g�P�r�z�ӻ/��4P���"qt��Ze	�/Ps.��RN��C��	Z��J.V�h�2�cI�0%2Q'P�C2x�q��j8����\D���egP�U�V� �g�>Ss`�{EO�F��灘i���c����S����+6w��V��Uxv�#��Ɍ	��)��	P�X?�y��LK�W��'�xTːXo�0\��պb�"=��K�6
��U����R
^�J���4�C�Wd�D���̿*��-��芿�p>ej��"%P�2�nV�S�p�Q'K�W�(�P��Ĭ$�x�AE-�#t���'%b)1�KO�o8�8�#%~�q�2�B9NM�$7J�IO��	��:�@9$�=�!x���Wr�8p%CHӈq��<ODKP%W�]$���Y$8�  �%�7Zh�P��N؞�$��I��# $��E���DH��<���/>�B�)�sښI���/��4��J0yjFr�C�9Jtzź��B�8�W��P3:���G׭�Q�D�q�/@]��GH��Ą9}�Ą6���1i�0<��r�D*/
Pp3h�j?с@��Ot�����:�ި��T�^@���g�;��~�'��DSG4t���JU8{w\�@,�#22~X{�)�.S)����'���1�;N�|�q/���;5����0h����5�u�#�Eg(<�� ˻z�"	3���f�:�P$x�,��'l�>��*�&ѫ�	�f�����허M�~�bq��=�~�`�3���11$�]*й)`o��p<	f|�l�8F�>P�	'��eǞ���8�j	)u��%AN���H�J�򱋱J�Wn�y�a$��a�Q���u�þ2�A�� �7��M��6}�o��l���V�.z�Y��&��m���&�<oW��ˑ�;4pHw��B6dU$F�p�����u�a�*�o�P��iA�3��K��Ƣ�lM�V�K�J��P��8a�`4� �4j�p���A2� �{� �yG ;[������(�\A�ŭ�9�Px"�`��
AN�3K� T��U����haب��)��
?r@a�`,�i��b��^�L�h�g�f~&��fS���q�N�-��LJ��p<)rj?���B���i?v���KXkU�<J&� �Rw��A����s��Ȧe c�LQ���'.�d)��'��!�D�92��V�S:@0�0O���qmަp9�P౎U�B������9��E"����P=s�틯B�E�F���j4��i) H�B�	�}���Q� 5]vi�J�7-G�8b`'?�(-cVo�$E��DJ"q���1l�@�I ^�<cΩQ����2zz-:P�CyX��$L�/�J�u�7/X|�V�OC�8]��*źPU.t�B��d��y����-�D�S�C�+Qn�$���@�L-I������+B�m ��0LOP�Y�
U�"�8�@HņIc�|;���2({�(�.Q�8�3"�	6`��<A�0���25�3<O2��o��%��x����	Y�.P�!��D�Q$� �X�}�(4�7�F�B�aҎ2�a�7��;{�F��B0�x�8�c���y
�j]�a0CH�C*dy#"�XX���1��Y B�5&:<�a��hY�i$?)��w�­(dj�*c#�xYD�־|�ĝI�'���yd�J<��k�$�%��%�e��EӦ�0��GH�n��F��ѵ+� @��}�@�G$*��w`ɣa˾� p�É�y"�W&}?����FĻWE�>�~R(�,��qPߓ4H����O�>�����۽lU�A�ȓ`xs�敗,�R�+0JH*�(���*[�X�c�ۓ@z(Ӕ�ь^��+��)�eώ�J���\�l�|5��?L�R Я�q2��5CPĆȓ���Af(��	���a���JT<�ȓ%�� �H���@+_;s��$��B. !{��N�pb����4b�U�ȓj�y2bŊ�F|���׶w�������g���̭a�C�VOtI��X��}+�B:�l,�D�Ұ,�l�� L�=y��Y�G 6S5��k���7^4U�@`�+_�&YZ�����Յȓ8U�A1��Y�W�И��^09���ȓ@P���B"3d�JЉ�D&)�ȓ\�`d3eܐB�V�3�b�C�đ��"�&��V�O�A� %י����ȓ|<���Ǝ�/$�,{3ː:^�����l�v�@-W��!;���(Z�d ��6��B�Oٟw ��U,�&�$��ȓ�Z-����?ֈa�'π�NƨU��wةϜcnt�D��='b���x[� �'ޮcB �pt��=iS�%�ȓ	�LuI�iٲ"tP����@� ���ȓ%������Ʊ,/���u��{�f̈́�S�? FD��N�c	��r1M"��9�"O��KU������U�i�\���"O��SD M9]��]�
ێU��s�"O�ZF�3�n��Ag����1"O���g)K�^Y����
^�I�"O����B�T� �e�W�e�By�q"O�l��&4U�p����gЦ8[�"O8Q����u�8Yx�#�:~p5��"O��
�hQ .9�2��8\r�e{E"OZ�� ��oM8���ϞQd��5"O�g�գ`jة���Ů$ihl� "O&���X>�8qڅ(E2"�,���"O�U�һ����U&�::NZ! �"O��*#��O���'�R�HW"O^b���O�������H�"O��zfI"WCԈ�"\�l���I"OR���j�@y�`
F�X3Ԝd��"O��T���/\,�$�а>"��P"On���	8�\	��˄+�X� "O ��Э��1���|�6�ɏ�y�F%
e��P��b�pa6�K��y�*�}���x�ĸW����0���yr@��4�Niү�B:�4��y����J.�(��
䬑 4���y��$Hpxæ��^Zz�QS�P��y�a�*4��i��@�b�I�����yBD?V�\�j
�d�xA�3�yb*�l�x P�G�6���h�	B0�yr�X B.���W5=A24r��T��y��0b���0���"mڌC��J��y�������jL�Vu��C��Py׋/��ĕ� ��l�Bk�f�<����,4��<�?
 �v��a�<ٰJY�>zQ�O�,@���P+�b�<�3HS}>L�`@D�}�Di�$t�<Ʉ��4*x�$�F�I1C:��XF�n�<	f�Y�G��@Dg�- ���@��i�<�G��&>���3L�MCTpR�_`�<)�,�/T�专r�
!z(x<�3��k�<�U
�)Owa÷%�p��(�F/�Z�<�Ť[XTR�J���j�t�x��ȓD��R�� 4svi���`�,�ȓ5����`�v�lL�TG���G�1#4�
� ��V]`��̄�uf�xB��֒'H�TӦ��jt��ȓ�� ��}Otـ�mZ�t��݄ȓ$dҍ�l��c��`JVD�Xz�,�ȓ�ےnS�t���cD�TNV��ȓ9��T;���@�
��)Y �t�ȓJN5��	�r���Ղ9}����ȓx쐜P�&�+q�P�s�"��b.م�4�a9C�k$�P	�i���ȓi$ ��'F�^�~�S��#uȱ��|����*!�0�8q#ߌN�t��ӳ�ޮ�Tؠ�h	3���ȓ+Ų� B#O:Xp�h�S1���((���v5�i�\�n���ȓ,J�����>�Faj'C��/�
����
dD�BA�(�j�,\V���lgNt��U�&	 f@�Z�&��z*ĸ�a��� <�����)x/P��ȓy! 1��g��u��l��U�&�]�ȓTt|�$��B��]��Hm���`22��h=�ʙҐ�C6n}$��S�? �@�$9ADYp4I�0<z4X �"O�\�ƈ<���S.\���Yr��m���ѣON?1�ƭ�`�'�����6s�A;#)Tq�|!
ӓ8ꦍ�Q�:x� ��΀�_Լ�#�'G),9:KԧT)���'��U�f!�	%<��#Dk���QI>��Fh���a��i~��a�#����N�P� U+q����;c�`C��	A�����CN�I@�[�l��(HI1,(�e�ğ% ĺ�F!��q�d_  hb@���D��t �O�t]���6K��QWfA�~d๱��q���҄��ql���&ߙo�N�)g+ɍ�0<����c����7{��ɓ��@R8�$`DV�3���K�/B��e�*cUB�i7
��� �� �� O�] ��%H�Nݩ&.�&:FM(�>����	Gl��n�2)JTش��8��c>mQE% �Fh+W�]~#6�'D�DX) y�B����65��!�ʅ���W�U-j�:}{��&�Fb>aKS�/?��`Կq}� a�'�.���I�g�C��<؂��*�,0P��D��b#"QrSF��1�������
�1/�W�{�@�ҎɇdɚP7�R'CZ��@�"9��&�9+�A�L�]A���b���+��2]�����J�GC��d�ĸa���:�'s�$H�DlВ�j��87�̠.OU�1kO�����1D������b>��J�3�4DQQ���-@�p���,D�(�T�F,!��pcw��%1�ܸcv�K�I�z�JIO�r"Q�L�`ؤ��,I"3�,?1�GǨO�� �kǋ	����Lj�����gv�CE��8-x<݃����:�l!��"΅C��I� <o���㉮+z�= ƅ�3\�}�c��M�ʢ?��@ؖ25�La�N�K(	s3J�i�")'�F�4�eІ*@�SZԩR�R��x"��<��0;Qm� n�Fų4/ߥ��D�j�=s�/?{�Lt�LN77�^H�f�[q�ӷd4b�9S�K��4kvm�(��B��2m����5O�/�����IK�F����ݚY~�H����i��,	T@.��	=j��(�'~&���W�b*�YQPF�,v�I���x},���`�����U
T�*+�8"���t d�1��X�^��b� &�Pj7��-B���g�L0%,���tN��?q2�<1Ұ���ʿg�9���"�� ��̓(b��-D�&�2jP2����N�Ks�T�d	��iKX���W 7���$J�Xk�����h<��G&>F�}�N	�&(Q�������2\ʤ	��ץ�����"Ox�Iu!��Vh�H %�Q�~�CB��R(��%��_�hը<'=���
��+QJ�yO�d�1��e:�K{���F�+/E�}�&��-C��X#	�N*ؐ�j�j�JY�]Ȭy�TK!ȴ@4*=l�Te��CB��4��E�p�,�4Ύ�\[ ����MS}�M�F�!�3y"'_�(�R�+SF�;�0x[3��%vy�=�1�X1I�px���O�m��å�$�����&xl����ɘ|�T��h��Z:�U�U��#m�ٷ��:b�����_��xBf�z�J�cV��
_3�M�5A	!i�ѧJ�^t�d>Eb�R����C�I6<�|��G[(Z�`�a�gѽ&�A�##�Ku����d}�;B &88�p��G��Y�p�9? �}��C�6M� �qV>�u`�ʋ4O*��3P�8�� 8()� ���M��|�)�"&T�Q��.Z`�pS� �"� "�ž~ ����J�`�4b"�@ $+N�k�� &��`@�7J���éӜw���⃂>?!��&:�ꭓ���<3\�ȼ4u&I���8]sN�s� A:(�Ej�OA		����#Q�P�q�3�P3!/����)҇��6��<i����Fd��U"]0%|ಢg  h���$-X*�=3r' �(|j`BFIzؒ��\3"uȚ�ǖ .v�!K߀N�\��U.	�	sb����M���?��V�ةІ��w%jp�E
�1T� �R��i�I7b6�M#�jBeQ.(�S��'�X��kՉe�8)�C�>B�����ll(ڠ*�;5�����}�y�a��)B�Vళ,'W����jO�|tB���Z+b��(�pf��8���gg�M�jv+H�h8����#zy\��To����4� h�4mA?~���bǊ�:|�pL�'��Q���\���y���̾�4q3`�ާ/�ƍΓ��o�CP|��L��T�i�9ِ%�D_b����(^��&Sx��FJԈ/���c-9�Y�o"h�Z��� ��O4d��C�4�y���yb�֙�y��#l�L���mÍ¬!���R?N��I�g�z؟$x�m�(FN,����0?C�ڠ(ݱgj���R�D��(�dʡ��[�6ON4�!���8N� �p�3bg��ۢD����d���*6�T�3�[)dzF G�%ʛT�$�H��>j���A���:S�4��=s�J�Ra�7���v���<!�it��X�����k	��K7IU�2��O�M�&�ܛ\����% ɒi���J[�@�W� B����
�~���kg�i9b50B��+k�L���iZ?7��Ӭ��k�8��o�(jpbm	�/�:�D��
�Y�Z��ϓw�2���3j�dx�0"� 5�iA��î/�$�j�-$(b�Ýp�,̺aL�m�zD��i.r��r�_��9�n�A�]�b)4�J}��O�5�'��p���	�mv 8[��PX��BK�U��1���'��I�Eάw���!���|2IٗWW��:�A�+?�h�N��x��XY7��ư<!�A��()�ҮԤ�&�5� b���ϝN���2��?o��i6l��hN���t��**�Zɋ��a�x%�VdI�����)D��t*ǁG�Řܓ��@j��'Ĝг���i�ތzį$ufs�l�����kL�C�|�`�l@w+ʨ*���)XF�FiƉ �p��(Aͤ]�
דZ8��%Hن�z�"�L36�D���[��IpQL��(�ԀP�#H&]7�����l9���M�65�H�����<	�j���˓l	�j/<aO��ڰ�!l��`1d5Z(�����\	�$���I
G>A��B�8^:����kS#h��8�ҷ_%���5c��>92P���2d�����/����-�R8��i��3�t�x4G�[@%��d�R�U���r����b:;<Rhv�T�,�Q7��:V'̌���E7b�D�Y��Ƀw/
hpH��Ec� �`�����'��<��� �@�� ��j�ID�M����@���*lSp���V�r"���Ϧ(�v��f���p>a��;�,��j5=zn�*֬�������n?��m�s�W�dȶ��'A��	�o>�b3f�m��9Td�)b��hSq���?�LQS)�
�	�/>�RdS�J��ǚ��*3.��C<O@ IX�N�б-�n�Yf�Z�S/�P���J�)q�'	�}��M�^)��Yf%8�"��t�hg�X_;����@� f�<�q�1���@ o\5}ȼX��N�Lq��ٌ��i��a�@��@��	5?�}��mΌN��AX	Չ7M�'��� hS)`�8�V�A9+����Aiй�>���9	ơ�(�/GDT���Y�'�-�ӊS�-�\�Rd�'�ū#	�I���Y�)�A*���s`�?=��e�4V��=`dߚ�~B��'l����MA�����;&�R�
BlA�T9~��3n�.���j�R��d_�c��x4iާX͢	����I��H�&� �K��)0bO2Wr�%�D�-e�
l��'��b����0_�dI� ^�R10 sǓO�`	"���T��Tz���PA �'8b�1�-�~�^Ց�B� P���L�d�����--���	g["aB��\���Mr�$S]���'��tl%3�~�	Q��I�$�sc`2LP"s��ŤX��ΈFH�D��ĉ�4�������9�p��'
ڬZG덧���a�=��� R@)r��L"q+\�pm�����	"�����%���y'F�>���H�w�x�����)p��	Ã��)0��	�'>TT���I�BBH L^���0E�L���8Da�����y����T;���D�H	D\t`Ь������'�<�+s�F�����m���I��&�!#@��5+i  ���B�H��T��ovj"	��솒a"A��N�����W�S3y�x�q�Ҥ��x��N8ke˧�,fZp����I�X&�����V��n�a��3j�����b�H.`�ʀoF�sҢ�h���8�Qa�b�"x��Ly2m*4�l��C�R����+w��/W�8�.�p�͞[%f�*w!J�zY�#�
Q���'�n|�;��R#�� פ]�+��<��O ���-�M���p��N瀝HCfN�yҺ���� ���.�0m��Ӈ�ʉI���8��P�	�p��a�dק$tP���mY
l���������l�\|�g��;{b���"�,-	`bG��lш��֊Y.�ђ т"~��Z��6<O�p1>���Z �ߒt�����$�	8�r��0D8~,�'�V3����s�C������*l�.0re�M�B�f���Y�y��]�j�Ԍ��#C I�RDo�v��u�f��)i;:�!�� G�uH�H�h�҄&?ax�wLH	27�߇�x�8`�ʨOr� R�'C���C�˞O�Z�c��ީB�]d-=����D��?,�:TQ��S�K�N�^b��j�/��9¶��E�*���	Џ D�H�Ԣ��yTtR#
�w�d��¬������hQ����5E���	��	?�툅�ǃ�!�d��vĮ\A�"� o+��j���G�!�$J�`���R�&�|A�mK�o�!�����I8���8
�p��2LR\�!�DW1*�� гb^��b��j�[	!���*9jX "&E9�T�D*�!�	�d_�����\j���Ѐ+�!�D�yr�)Q�jC� >q����"d!�D�GJ�"v)Ɨ���T�O%za!�D�2`���~���jG�(NQ!�]+�:a�4ǎ��p���jܩ{\!��]y�h
�W����9R�5z;!���&��"� �"��ۀ!V]!�DJ�������SK��"���<�!�/5M��a����;�
�!�!�P�B���Ce��S�(@r�D��!�d���4lQ�Us|xB���!�қFT
 qD��
\��{���>*�!�d	�6~�P@�NJ�$6��ʇ#m�!�
_8��f!|lX;���_�!����Q�����`���Rf!�� ��Q�[ƨ,yS���^�eӢ"Oq;򥇷M֠�j�K�u@r�0�"O��@�u>�g��QM ��a"O�B��[P� ���T  ع�"O �ā�0t����"�2��u"OX!�l�	�<�rCPFX��"O*Y3TI�4Ǌ4�B ���.�k�"O,|ѧ� S���t���HIX�%�z��y��K�O��p��x�+�
�L�*fI�.�r �F�>��� �-��I�<	�'֥��Qr�q�1B#OiTQ˓�+���5['"��I�<E�4��KH@��SkY�+ �ta��W>�:\��$�:����2Ox��çI"H�À!�"O�ؐp�@S3�d�4����(�'��9%cV��X�H4�w�r��6̃1#9h���O2(y!L؇cGp�b��9O�!��˞�9���cf�] i��8$�i�~�3"�x͎�4m�<�u�h�b?u��N�g� ���-V�`�ɤK@�@�R(��������O��ؘ��qdl������%� �3ߴ2qO"��S질���
��" �E.R�6a#\�۱O�	�m�v�O���
P,��&P��p36�Q0�'(=�vL8�)�Ӵ"��8�r�	�`���{D����sOB ���s&���eG]/fE�ӀA��7���^�� K<i��~&�����!9@V�;����'n�>t�J;�$ҧn�<ʧ��$��k��A�P�c��:Nx����'�t�ɟCM�u��c����r��&I��0�N�	Z`"Y}�MŹ^q8���=O���~,�V�y�K��5f]��&WS��0�'�v�RsA�5OlpQ9��>�}�'���T燚��y��9�N1�d�Ot|���/�7A�����0|*�y2m���E�(�D4hD�5`��'{�	�Z�d�O{���= Rc��v�xeI�`]+5�0�h��D�5�2�`��O*V=����'�h��J(w
��i�O�5�R)P�1O>-�w�Z1:�:`R%�Q%]��uh�b�O����'��O��j�M2]34��#��� -�-C����s�d��a�|J?��|nZ�>^\1��O &K���0�Uk�6�˫�ē��N�O�"T���]�bͺ,:��	TU�'q���\l� �m�&Э
�'���Am+,h�𬓓��E9	�'`��c�m'��)�Y �ȫ	�'������]�Cb�y�w'�X�p8	�'�<cׂ�) �XX���^�F�(�q�'�\mb%JĞtz�T�BΞ;>Z�Y�'�X�;�a	�D:%$
� �<��'�T� 'G��7������w6�:	�'A��cq���9�����h֩�\�1
�'S�-\e�h9���E���!
�'4�Ek�a��Ш���0H��i��'�4D� �D9ay��� ʘ2p����'��@'��6�bak�ᚹ9�(�)�'�@�Ab-�&w��0@,��M`
�'8�Q��EZ;�D��Ê+͒��'x=i��Gc�=��/T�$J�'}�5�m�B~�Ϗ��y��'E��CԦR[H	#��*Y�0��'p�"R��FaڐH�M NھPz�'��a(��A��+P�K�w�.I�	�'����%�O%$��ˆa�ll
 		�'$��"`�y��0�u v��0�'�8�Ze΄�p�� φ�^GȌ��'���h�A�V����K�]���
�'�,4*�S�3&l��	A�R��L�'���1�
�x��(1G��G�^$�	�'#�S�X�Vܢc�>�
��	�'�$\�ǫ�Y\q��D�=8Ppd��'`�X13��$tľ�)�GsB��'{�aA�R�c�m#w`L�F��|
	�'����k�+�|�GƲEx����'5x<+��/)5�1���9Onj���� ��b�D��:���/bfnc"Oby���:S���a׀�
aeH�""O��
��	���|
!�Ɍ,a�8J�"O�uc�	&gt�B�A2
wX�+"OjQ�ŮT~�%�2��nB�KQ"Of�p���'�5Z�Ju}��*p"O���T��QwB�{���'*�^� #"O��u�3�x`Ti�Z�{"O^���&�\9�p��7*��<9�"O L���>���t�\6F�)c"O��)�@�/t�n���O^�(�~e�D"OX�9�MY og�\�d�U�c��J�"O���EoI1��`�f��*u|�J&"O��D�[5^~����
�'��Hr�"O�WCɧ1��}k ݟv�XH�"ON��ҀI�9>�s���}����"O�q#�c��G��x�Y�H�����"O
e;���4�N$8�M~;����"OD؊���\0��v,��>-�T�5"O���RF4��l�B&]�*!Zqi "O�P��t1���ab���"O9��a3VR�HB����L1�"O<E���F��A9�@�[�Q�4"O��`s�HEH.��a�W�-X=�s"O�d�+K�g���Ј��j���"Oh���O��gdFRE�Mq��"OB���e��;�l`����Q&e�"O�,3�%��9p^�)Ua�'���"O�pU�˸U��u�Rn��
�n�b"O����0La��W���C�t���"O.�`۴'ݮA��
Y�h���B�k+D�x�g��
!�=� �P��	d�&D���4���@y�"C�5 �Y�"o8D�ȹ�F�� ���_d���e�+D�@z��V�jX*�ʀ������$'$D���2����-��0�^]Ȱ7D�d[��َ����R3.3$qX��1D�\c�=$M��8dl�W����w�0D��IŊ�7pb��	wg�ݬ(xC�,D���0Lצd�4Ũa�I�5�0Iի=D�(���*%���*��3_j�%� D���� W8GUVMS�Gڑ_�X�Z#�>D����/n��bX�">�e�gl/D�H�#c�)8���{��� i����-D��`�Da]��"煆,^��� j,D�T�Q*S�ܙ�-�)*���S�)D��;Pn�%jF��j�IA�\k�Y�4D�0�'��)'�ȶ�8X��p'2D���"F��(�b,��KEoH�i�&0D����(I�PY�Y d)E�2���x#.D�d%�C�l�
����ĦA|��飪+D�(����` ����� n%� .5D�\9��S�* ���fl�+�o4D�y�〢J*�U��,����26.2D����.���a�A��^�d��g0D�p���;
vp��T�ǣ+�ZY�j*D�����]+}���qdDFw���@'D�0�"*��pK����c�6b)mH"D� {Q ��fqj	; � ���|��. D��U�2Q1v���Y)��Sdg?D� A1�A�c^��T����>D���B�޵�S��CڎT�v�7D����"�8E� V�^�N��",:D���I�1F,��@��>����L2D�� �	f����tR�-�"Oz�'	�:�I�moᘣ"O��:W3e�躰!��b�~�J�"O��;58a�q7!%=G�A�C"O�8ɶ/ޗE���[0�J�@�ě "O���ж=ȖM;����XMp�"O��à
'�E�5Iѝ4ڱh�"O�+�a�,R�I�����9.�9A�"O���h�#+��t���¸@#p�c�"O��XB�F�.h��]4*1�1�a"O�uK�o̽^Ϊ��U$�)F�uxF"O|�H (�y9��4r���c"O�a�H�!Ds�%yf>%l�ىD"O�q��@t��J&�R�&I<jd"OZ̛SA�%W�]���<8���"O�ܚd�Q,+%ܴ衍ȑ8���"O�Q a ��}��Y����5��6"O���w������0���0V�^w�<�'�)vj@��7�.d�JU�@/�r�<�k��`�ڤH�&�+�<�J��Li�<�S�,8P�aJ��hP��g�<YP@�3m����(H5kX,�c�gBb�<Ie��T�jP	R.�<u�6��თS�<	&Eαa-H�`V�̴E\H�'%OK�<1B�it,ds��/6�Jׇ�k�<)S*� x��8��$äjZ�&e|�<I�B�2���-\D< @�S�<y��0̠|Re`�'x!�X���L�<i��-E;`m���>|Q���1j�J�<���ˍW������=/$��G Xo�<��c÷h%�iAwc½:Ј�cS!�V�<�CR;`� �� _�T��Y�CO~�<AD�N���	�s��<"��l^P�<��B_�H��&��%���	��SK�<	dB@ay�@�ŉ�b�����\�<AE)��b��(��.~�����<)��hH�5:�On|u�2��|�<A��M���E��hɧH	�y�,�nܘDg�<��`GA�y�g�1x� �� �6@Zb���y"ٻpef[�K.�z��B��y"���w"N�&��Ы���y��.�N�8��V4P���H�jټ�y2�P�@Ih�aU�'NUZ��d�=�y!�J���)��:6
�� Ց�y�i����d���4��E⃯�#�yR�Oa� !xF�ǽ)�����T��y�CJ�E���1f�69���
d�1�y"c^(�$�@�F�$y$Q˲��0�y�g��Њ��0_��rb�Q��y���)����d�( 9��Qŝ��y�D\e%Th�$CE�G��#Q�	;�yB�ё$��h����5n���xC���y��V1,
���g�av�x��o)�yBh��P\���F3�L��I=�y�j��_o\�!�(��2P�V���y��P�U�ZݺSb$�ʐ�P���yKݑ�rы�Ӓ{�lȡ�d��y�KõԊ�R򯊱c]�A���y�����+(��}��k���y��MS�bʅGN�u�j����y���z��B!u젼�ů���y"f�BVv%��|J4ȓ�ԍ�y�靿0X
�!��>�LL	5�-�y
� Pl��ELH����X�6"ON�iB���w�!�,�d�[�"O^��w�M���ثtDE�IT�"O��YaML\}Z�G/���"O�����Y)x+jtr���J(���"O�X��-�5�*)Ф�P�xi�"O"���F6Z��dĽnx��"O@d�f$��~��$S��Isa���"O�ijр!��e�Ga_"[�]ID"O,�+�C������@([A9��"O��t�Uc��ur�і-ԚLCr"O��ҥE��P����+�8\��X"O^�8��� @^�����Q#0vh� "O ك�/�)���
@�w��z�"O�`Ç��DԽY���ٶ� W"O@iɦ�kML0��'�#fveQ�"O>�7���Tm�f��=X�1��"O�}Q��� 9�8CB�ҁe*|��"O0�*"M��<�s%  0pq"Oʼ`�*�'(�&x�v#�6���"O2����L�N��L�2-րH��|qA"O�-�ӣ�/Ҙ���8:�\�@�"O��"v�B�[H�+$qH!cV"O$<�a ���[�		1W��a;�"OD�{�߼v��pc��;��d��"O�Q�p�]'t� R&b@m�K�"O��7��=:��|�a�J�B5p�8�"O"릨���C��%$���"O��u�`�[Ђ�b�T��"O�̣F��$�ieGO"A�!qb"OP�@��)ghI�!g����8s"O^��f�!�)��M*	�❊3"O+�H�#I������֩�E"O�X����m��IFC�L���"Od@����s4%�4_�*�"OF�0�d9�dq1UC
J���9�"Op�����<R2���&GH��"O�|;�   ��     �  �     t+  P6  �A  hJ  �V  qa  �g  n  ^t  �z  ��  $�  h�  ��  �  .�  p�  ��  ��  7�  w�  ��  u�  6�  ��  �  T�  ��  ��  �  � �	 �  F  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!����:}�����ZIZuH��Ay�t|�A�/'TB�I&	E���)^�*���č݄�h���.��06p���8W�x]��o�6F��}��If�$��,&$,*D,
���+j�;e��'wўb?��E�����ږO���!{sA;D����7��PiZ�*�ޅAщ:ʓ��<)���\��c��d����M�J~2�'��O��9ri�^px���h�i(L��LIh<��~�ڥ���!Q��3���S�<aG��%:��ʄ�G�.0r-��BM8�XDzb���i"2�Dֶ^�|P�*�8�M��'&ў"|���F�Ĺ�f��(��k�I�f��O��?� ���HSgXm��ÝK��a;B��3|O2�$��#au"�3��&�1*���4LO*M�'�ҭy���qs�.3�©'���y��'��{�339f��"G�Y�����'ͳ	�z2���˒��GlA{�y��N��!��&�}pP+]�/W&������џ�E�����!vX�c�E%u���q�D��y�,
�_���3�c� ��y�mY���IBX�� �H	ys���B!d4P���C�X8͓v�S�O:^���Ac�Հ���kԘ��o[,-*�B�ɠ���Kl]>*Ѐj�k� W\��'��IX��p3#�Ɠl��,�𣝆u�~%r	$�O�OB�P� 3+F�H���k��qP��D;�S�S
���(a�U�I��ȡ+�^�f�<��T>mKS�� � ������n��U")D���A&߁gNLŐa��e�B4�pN1?��v��;`A�f3 �E�^(@��ȓs�($�E�T$Lu2�c�<Kﮐn�-��d.��=9'��H.*�Ђl
�m��+u�^m��L�<��%Q� /T���������Si�<��j��Lc0�;�!�9~����P�<a#��J"�p�" �@\�&#v�<� ��������8Zbp���X�<	"H�!{\�8� X�3(����A�Q�<!"�iF@��@��l����g�<!�Ϛ9UZ�r��C���'b�<I���(Epb$+ ���Ue���w�Dc�<�AAWB� ]���y�A(�'�b��hO1�^P ����C~.X��1A�����>|O$]��Ï�m!���E�IB���8���kX��@�>FﰐR̔7m�=sÈ(D�����X�vZ�i�'f�7�f��#?Y�􄕑l�d��ԃB�=Op�i�k�/L!�ʨ<Q�� '�/(4�l�#�H:B3�	�qQ��|�KY>��0#��I	JW�@��-@E�<��ޮ{�y�#	��%�@٩u _}���=	#E�f{�Y�fH��b�n+T� bq��.FD}�3L��V0����5D����æz��}���[� ~���.D�T ��Q�1D]��`z�/D�LX�[�(R�&�wJ��ok!D�h�i��
I�D$Z�Jf.� DA D�DauϹQ�<9��� $!5g+D���󢇋Y4��ۆ�C3
}�T�6$�4�1�ʦd���'KF�w������y⇕�p�3�*�d�ۚ�y���x0��bpA�֥�#���<qM���'�]0􂋄/�m[!�^�`��
�'"��Ӫ23ʠPr��C�r*	�'����5��$v�jժ!�R�6|�Q(Op��ɷl�x��4I� 50yr��>L0ꓸ��,�~:�On��D�)n86iǏT��d��O�0C աv������@�&f̜ᦊ"打&E
�	{�S��O��ؓ�
x���Ѡ�az��B
\:�d���{�h�x���Z{ ,��DL��7a&��B����Nq%��>i޴��O�H�*�I�06�)�o�`�
�'	 �y���W����� �|
�'��1��ʂ"|�A���՟&o�%�	�'��5�VuAgG�5O�6���J���yB�^7L�堡�^�t�zl����y�/��l%���#�\d~qj����ұ�	��H�)c�s$D{�h�(A��`��������SZLX��@� ���I_�B�)� @�XW���IK� 僽NC|��c��*lO�Pe�]�n��E�sX��p�1"O�����Z��Ĳa#L5� �2U�I@��H��&Vˈ��J[4����Z2Z����4ړ P��@D�?�$C�C-pi�k O� )W�@�jDL����@�{
��дi��<}"2O?7��\�֑
G�L�c� �[����x�Bf�i؟ B�DՅC�(1OR��Qr�j�^�=�}z/O�@�+���ȀO�.tƅ��-J��p>	0P�(����@BR`�eGr;l��WG��y퉐�(Oz�(bL��`�UŎ �N	��#��'���i���Y�LJ�Y��	 ��jGr�'���Gz���צ 6���A��\07�G"UV�I�<	�}��X���<e�Ƹ,��ʗH5�-�HGn�A<�z�$U@8�(*�nǵb$T�s�e�;F�@�C$�O�6�>�el_�[e\��g�Z��i���/[e!񄕼L+.�#3��� L���Q*K��a����w�ĕGKv��s�l�P�&D�����PlN�(����T S�&!D�<�DC�_1L���ޡZ��:B�3D��h�)�,$鵪�*+�t�ɑ�/D�8@�&�3 ���g�Bn,ZݺA�.}�'��a��kȬ)Blp��Hc�ݐܴ}�!�$W�0. ^/��]<qa!�S&Œ��M(n�A3*͏`!���"g�l
�����|Õɦ6J�����)�Q���"?���%I٣(C&PI"�Q�<YD��N ��b��>ݘ�Z	�hO?��	kLT	:���7:�R|˄�D5 �B�ɡR���	�l���{RC'K�LB�	��$��Ȓ}N���$h��	�B���.�Ib(H	bIΝ'��uI��Z�>�B�	�Xy�@�]��`y��Kػi�B�	=p*U�Mϻ^npt��
�~�B��L61:s	�r��U[wL6v�C�I>_p��ŊRd���A!O�\��C�ɧ�~�Z� @�}^���` 6�xC�	�k��� O�p�,ȗ(;m�B�	�f�r8�V��0X"0e:�"�`3�B�I?t�  �D0p\Ԕ�$�Δi�C�I",���Ѐ�B�j��p��O�C��)T��a���j�ֵ�f�D��,B�ə
���k^,}SpHd&A"B�I/1ϊ���ɝV��p�C�[Y��C��-H���P,12��ؑ� Z0��C��i1Jd���3I.��Ն�s"O�@G�ԫe�E�3A�5��!!P"Op%���1u��s�oC�\WHȃq"O�Q��)��(-�(Bsˡq��)"f"O0��E��10x���rĎX�t�@�"O �Ñ`.�xc�b�8{Т$kU"O�����ɮ�.��5@R>c�d��'"O�p��Jƶ�J�6�ӆ(R��k�"O����4�,��F��+8����"OF��A�k����=@�� "O��$��~��׭Hޚ��"O����ޚ,��Y� LF�;.��@"O�����,/b�b�+��J��Y�"O��3���3 ��ӆ
Oܴٲ�"O�QCLO"1��dq0`�2&��u"O�=zŠ�m��(Q�a�.��R"Oh�D!�X�b$@��f���"Ot	�ɞ�T���K�w{4��"O�-��S�-��Qs�[�{a���"O� ވ����;��L�T"O�%<O�8�b�	޾�y�"O`${~����M"�&$�u"O��	��ڗ8��������"O��/;KP�	�@ۃ���c�'UB�'YB�'q�'Ib�'�r�'F�=�č�*^<��˚�(A��'�"�'�r�'B�'S2�'�b�'�^$���u<�T�P�`"9 ��'�R�'=b�'!��'��'���'+FE�V�
:�Z�䎎�I��ĘC�'���'�B�'�'���'�R�'��KV��.|u¸����%��RG�'���'���'�r�'f�'�"�'�V|��">�MY�aY�F0�x@A�'�r�'���'���'�R�'���'e��2MG�4Ff�$K�����'���'���'��'
"�'���'�"�:��S�J�����n�V�'���'�R�'�b�'��'���'ȆD��ŗ�#>���P�e��8���'$�'�2�'b�'c�'�B�'i[dC(|�x�!�e 2~A
4�a�')�'CB�'���'���'K��''.�(@*�W�F�iF��^�"�'���'��'��'�"�'��'���rʌ/7��9�˘�"Ɋ�
`�'�b�'���'!��'���'���'�V� �O5@�r�kHJ��신�'v��'�b�'m2�'�2@h���d�Oh�x���q�q�n\Z��Q��Ky��'t�)�3?q�iFzq��N��`0D�@��D�Ya���r����DO馁��]�i>�-�M{v��6��&G0j�Թ�A
�֛��'����$�i���p}l�҃��N��э�3��{ T9�$�	�~Q����y2�'P�X�O � 굣��N%慰tm�p.��25�m��	��$$�S�M�;s�������'��X�u��P;@�1��i��6mk��ԧ�O�. �d�i"�DU�b����J��!����VT�d�)*��Y�Ԭ��Qb�=ͧ�?�eeZ�g�8�7�B�?�����<q.O��O-o��)P�c����K�,"�(�+�^u To@A��	:�M[R�i��$�>Y�ዿ����F��;�^M��#l~�ʅ_��I����O���յ����I7+���O�����"֗#g�'i�ן"~Γ ��G�KR��E��J��Q��fJ
��D�榍�?ͧ��ɓ������ʟiY�4�9A���r���Ċ�_�77?A��KUQ��hP뒼[�9�#R5�&�ҳ/?�J|���4�*ʓ��@$�����D0��xPLǡ�ʩ�'#�7MF�>�1O��?��D�A���f�� 2�6'����ONIoڰ�M;�'�O%���'��4�Ѩ�(��}�!�[�P��Cc��(a�%ۨO��:�"�&� �8[w��'���b��@�k�"z�dY
�a�!���(�����<!N>��i6�A
�'
��(!��cڴj�f��9x�ß'��6M,�i>��+�M�׳i��-(9\y)r�P:w8�M]�gcb� !�i��G�9#���,�^(~�z�O>�O]dq�֘4P�]���oq�S�'>=`iB�<O,��<�-O?y�r�	����ݰnu�` t!�I��MCAC~��b� �O"� ��R�;7��1�%e"�Բc�`�,�'�*7-�����R�lZ�<�d��� @�Q(ِFh�L�J�7+��9�0O�-���X��$����4����?ivCSS
})��Ɉn��KI��<�I>Q�i�ntK�y�R>��U�<;�1�j]Q��i8 (<?�&Y�h3شQٛ<O �����rD(��͝�@��N�?F�A��Gr?�as�����6�v�k@��sg4�h�/2?Z<�����4�ne�1�J�z�2�r��R�`&��oP�	�D�Q(9tE�A� ���:��A�N��U3 �_�,�t9�j�
h00��`�Z��y�`9��wZ,��$��C|Q��$��mL�ຶ)�/{��q2 m�n��!)�=�*	��*�.�A��|�
	q3+�%W�4�h�Z��H`�/����ӕᚄK�(��P�x�9���D�=%ֹ�D�]�Xe(w �gqv�{�_�g���YF��Hr^��� ��	L%�#Ib�^}�``�9�Tّ�M��iR��;N<����?1O>���?ag�O2��]��hO#Dp�8��@"rr@��?���?���?����?ဧ�!�ֆ�3@�@�d
�!���A�\#:��?q�����D��{I�I���܈��8)	�mWHؑ����?���?�,O�A��%{�S::�����Z��@��I
'�`�z۴�?)H>!-O<9��Ĕ-J�`�ۀ
�2!:�t��yZ��'2T�\!�-�ħ�?Y�'Bǜ9��	)Rtw�S�FAh$⁔x"^�P�w�'�S�t(��@]{�A�9�2��ć���M+(OB�;gA��-Ȫ�������a�'t:��C۴��sj�K[v (ߴ��η}��b?�Q@Wq��p{��04�L4R�${�.�A��ۦu����0���?�kK<y��-��[�Ց:�zC�D�l�����i�������񟄉���O�էĎYߖD	���M����?���>=҃�x��'��Opx�d�'^b��#jٺD�����M��1O��D�O��D��ht�kAbF�*�`�|��xmϟ����6�M����?���?Y&[?A��#�E��A�	X�ڠzg�� Nb�Xm7��X`z����џ��Sş��IIy��Y
�10�Ivf ��I!r�~@�aθ>�+O����<����?)��/�� @�&	�k�����b޳,|�xㄉ��<�.O���O�d�O|��/��lnZ4�<u�K[�`=��R m�M��xٴ�?����?A���?�.O��d�>	�ƤH��)�G��	�TOԼ}�`I�i����^��'r�'mh��~����O~aj�̘�w̌��&�F�2&;jNݦ���՟��	{yb�'�T��SS���%����,mvA#�)�#$(��m������ay�m�#��'�?�����F��ޢ��Y	0Q&$�5h�.0���OH��O��D�\r��ry�ӟҴ�b�ԯq�|�湸P �X��M�*O�yq��Ц��I֟��	�?� �O��8YV�ɑ@��q ��6�'8�*�y��~:fퟥ��O�ޤS�����k��M1L�`��4f*L��ְi���'*�O,���';2�'�ԩ�7�+$&R�R�oD�5YЭz��i`���O��Ģ<ͧ��'�?�t��2߾��A�-�,*s
��2���'>2�'����/f�P��O���O����A�����W�^=�[�W�\Ġ�X���'
b,3�O���O~�D�Of`�mS�r�� �3Ȉ3&���w֦M�I �j�4�?���?��W��SJ?!���1����7LR�+3�y�d�D6-
�NL��p9O�˓����?���?�5��_�Z��s$܅}Z��� �̦k�ʤ8r�ix��'b�'WN�'����O�)�;T(�Y�f�f!jUPR��8��d�O����O���O$��ORU��G�qA��ͺ4Lpy�b�Ǎ#.ƙ p�?�M����?���?������O }Q0�ԥ�'�E�X�R��e��U�ʠ�0"�馱��;bD��	ȟ�:����a��Φ��	��C &�����i�j ���
��M���?)����O���Op�ɇY�|�	@�)R*P l��p��SaG0�?���?�-Ռ8�$�i���'�b�Oh�Bv�	�hD�*�H
\� �7�{ӌ��<9��"��$ϧ�?a,O�i^�KQF�ho�����m��޴�?Y�&�(|���i���'`��O��d�'9R�@%��F � َGq���$K�>���.�������|�K?����͞7K��;D�U?!�̰��Oj� Ջ f�צ�����	�?��J<��l�<��'�P
5Rv�Ob�49�i��Q��������3�L�/� ���	�9h�ë�M���?	�	�jM8C�D�O��I�BҜ�5B��D��R/ךf�jb�T���3���`�I�LsVM�8%.4q〆0%�f�1"��M;��(���P��x2�'���|Zc��0cS�C;��U���PK�O���d�O����O �(u�`���L~1�#��9l݁� ąy�'v�'��'w�ɡ*tԤ���S
ʀ�I �2r�R頌&��������� �'W�p3��c>�æbQ���"�6wô� �j"��OƓO��+e�1�'�-� ��3o���Q�1���
�O��D�O��d�<�@�C;�O	0��e�@"q,���4E�F�[��cӬ��!��<�Q��k�-��%��:2�|p��L?6n�$l�̟��	Py�RI��������2U�ϫ^�~=�BO	��dX5��R��Ry����O��&9��m�6L�Zծ��3$c�x6��<i�L�Z��揧~���ⓟ��"4��%R�����+Խ��x�d˓V�6Dx��TE��\3Ą"0�R $�P�J�MS"K+���'�B�'��� ��Ol��3��ljA[��ŐE"���A���R��!�S�O)��ʕo�
�
1#ĵf�|����M�7��Od�d�O�0P@�Z�I�����}?�Pպ`�3*��em�d0`�R�[�l��<���?���T�2t�p�Ö6��4�O>� ��5�i���:��O��$-���(ҡ��,���F��##�FH�qY��Q�L2�ğ�����'�&��#B�t"�%�t�"[+�$O�$�O��Oʓ6L��[�k C�&�Є�ׁ4��Ř1�Ru��?1���?9,O����c�|��� A��Xj�gϐ ���[$n}��'��|�V�h�bO�>A�ˢp�HI�� $�����s}��'<b�'�	8"uh!�H|�(Ŗ.p��;�
��Frq����b͛��'g�'���7 �.b�4��O� oN������z�z��E/yӌ�$�OTʓV_v����'i��MqV�����&y�,p;׫$::O�˓h�Fx����a���3?"Ĩ��e�S��UAa�im�	�d�(ݴ5���ޟ���3���ώf�0�9VA!X��{��[=��\����[��|&��
rƞ�0J0�E��w��DP��{�z���&�����8�I�?e9�}��^�	�S��+�
H+eFN,>6��oQh��3��̟�cd��5-B�K5��{�n�H����M���?���v�dzՐx�'m��O���WKe))3��*Tn=�ӥ��'� t!�y��'�R�'�j�8eȻH�����Z$J��tӤ���3%n%�@�	ß�&��ؼp���{���=����c�\�g����<����?y���P���HዎNM�ꇨ�4=���r��I��ş��	G�Eyb�,;��Hr�KL�^�������eHb�yr�'s��'��	����J�O��YF��5�¡�ҋʜ5 :�z�Oz��O��Oxʓ$(�i�'��*p睤b-�qnD,+K�T@�^���I�� �Ijybm�{t��(w��0OJ�3�DS��8e�ʦ��IA�I^yg5�ا� 2���͕* ��13E���Q!�i��'g�
otM�N|R�����<v^��G4,<�e�&F�ej�'Y�ɔ[��"<�O$d��%C6��Kq 0I��4��D^�6� �m:��)�O��	X~"-��Lˢ2��'�,�cb[�M�/O�����)���>�eAdcڑ�hi�ڵ�v7�փ��AoZ蟸����h�S���'����E��&5	��յw�i��V��u�5�S�O�rDβ��	�
M?2n�!�B&G��7��O\���O�D�hy��۟x��F?Y�F� +>�@�4I��8�{�I	u�/w6@�<���?���%F���G��|[���_�E:��IB�i6R�۹^�Oj���O��OkLW�`hL��@o� ;�1x�1__�	c��c���Iݟ���[yҎ]�=��lyS�U�)x�d���P�0W|̣SC(�D�O���"�d�<����nD@/��Bh&�HbE&oB��<Q���?�����4T�l0�'0�pXJ���!g�Pi�5��#��Y�'<��'x�'=Q��H�g�S:5hr��$s�I�j�>����?������O�3Bu'>�Y4D�+8nQ)�KB&j�x�z'@!�M�����p<�R��~�xd��Ŕ1Vf`z�RǦ���ş��'�2���a<�	�On���A�1A����UH�b#A�*���%����ɼuސE��>7�|h��J�E��6�<ɕ�8V��K�~����BT��,�\"v��u"[)O�2-���].���'��Ħ+��O>��xbmNL<<L��eQ�[�����M3�HI�#4���'5B�'b���&�$�O`R�+�-FE��*Ύ-;<(���K���}�AE
r��|�<���� ��K?X�`{¤՗Vv$Y�iy��'J�(�&s�O���O��^v�GCݳFn0�ΊNZ��>ђ�O̓�?����?�uL[7��݃�ČT�l�WƎ�~�'T�@�E"���Oj��O����OI��T2ŭ�)?Uʄ�FJS}��̘'	b�'�BV�8P��;ir�JB�M�F�<jS-O~�Q�N<a��?!�����O��D�a��u�uAF����g�^?q��ju��O��$�Of�xq��!�;����E�*�LSSECo����x��'��'%�ɏo���I�6&6���Pu�P6d�P��'��'��R�P�p`�U�2:�b&��v+qf��YZ���4�?�O>�/O,��d�:�I�k8b�y�I�m�$�*�� -�7m�O��Ľ<��h6h2�OS��O(b #%�J�82d�j��JdM���1��O��DP�sĆ��'�T?�w�-��2g�F{��1l�,˓W_���i����?�����	�gߞ�H�Pv��A �6q�6��O���*��.���%;��ST"\8Ct�B�n�R�����{\L6�O����O&��TI�9�!��̆O��ܸ�A�|蔥벿i�V� �'��'���d�i� ��g\�~�YQ��4��o�ߟ��IΟ0p6 @����?i���~��� �i��2F���&kڬ�MK>9��<�O��'�r�;h|�3F�#	➰��0��6��O>�"�AS�Iߟ���B�i��j�֢B *�9�h��+Q��>i�!K����?���?I+O����/�?*�Y!�
&{tk4������'����ٟ�%����ٟ���4�̨�6
��-N�و�+�f]��	Jy�'"2�')�b��@r�OX�����"9�)�G�@�V�D(�O��d�O��O��D�OF �2O`p��j��Hf�\s$Q".-V�d�e}B�'�b�'��a$��QL|j$�=�XI�g��'`�~�F	ѫQ|���'��'���'u4qڝ'��"�*���W�~�<�c!��#I�d�mZʟX��gy�i��o�d�$����
�B�����0�Q�7���$�MO������,/�H�	[�~dQ�\f�Z�l�VO䡉'��ɦ)�'�Lb`mӖ��O���O���"
m���K�H=������m�P�	�7`��Y�)��x:|�FJT-Ba��$��X�6-���n�ӟ��	����<�ē�?��a�=^�PȀ+�X���p�����/��y|����O�x��k�x-�7J�g�ƀG���%�I㟄��I�� L<��?��'��1��I��Ez�T�'p{���4��CX�E����'���'���!;(��x�mɐd<�Z��g� ��=2 �>����?!(Ok��e�V�ċԔ'֊�cg�W1T�	�r�
b�P��؟��I{y∌�X��Ϗ�<�;&V�[�p(��5��䟸�	|yV�\�7�ɽo�>P��K���Ѯ��
b�������	@y�!�$%�5��t�S=@��� G�m����?	��䓲�$�n���9<��q>툽���/p!@�[�|������IJyҢ�.P8:�H53��'K�ލh�Ǻ��¥������	}8��R�DnY�ay�G��B��5!6�~Ӓ�$�O�ʓpi�*4��4�'}��nlb�eM�	�LĪ����O��DW���U�ݩwOT�Y��I�o�V�'�)´1�v7-�O\�$�Oj���0�d$Atĵ��W�)����ňT2q�@�'���!V���'��+��T�~� �J`�N,8�ū����d�zF�i,�,�%M|���D�O���T���O����Ob���a�]��bW��� Zd��0O�ئ��"����Ly�O��OM%z%b��B��&�tc��Y�\|�6��O^�$�O�@�a��Ӧ���֟��IǟP�i�僕n�7�:	 '��8��Ӡ/k�֓O��q1O�ҟ���쟠�D=( 5��G�Je�c�N�9�M���4A�w�i�"�'���'�.��~RoS�[i$��m�KZ�Z�^��M3��R�h,��͓�?!������?Q-�:�c�j.r��'�L�����~l(�	˟��ɫ����<��Vˠl�!�V
�F�tBC�&|� ���<���?i��?���?��)x��@��i0<J����><@�F��p��bӺ���OJ���O��D�<!�oH1ΧQ}�`� ���(��*�z�A�_���I���Iҟ|�	"T4��4�?	����E�f&�s>x�De�9"~���0�i�b�'��[���	�2Z�H�=yf�D�`&�8!��9�Si�)Y����'K��n�5bQIȟDG��'��y"!�PT"bE�IZ�G�����'_�}�G� n#��&CN?���e�&x�(���P�i=�0a�
ƅ[H��AƊa<TE��
,��XDg�,&�zI�v$$�A\'/kd��dü-Eh$����-0eœq���k^�;�D�BL�mb�DW134X'f�6�d���:L5�Xs3DJ�
rĹr�� �d@2'��+
\����43NL( �'[��'^�m݅b�MB2`��O��R�dXb��35���j� C;�?����8l��|&��ҥa�W�4�9)��r����a�Q4n:ƅq�h^�?�둡(�\�>�O(��lU�8s�ز�핒�5���O2�&��i>�F{b�m۬�`'P�b�ɓ�H͵�y�6�H9�U�F>��b�����Dr���ɶ<A����S��M���1ĝiq�@�g�(pK��ҥ�?Y��?���^���O���`>���*\Bw��*G�F�f�X@���J�q)����b���
�O=*�]���QuWQ��Y$�W�a�rPz��*2�t 1�ӨL�͊�'[�C�]'��;3FZ�V�Q��a%��L���̓�c��@�fU''_X����i�޴�?�-O��5��2�� ]# y�Y��Y�i�.���"O����cĄb�JYS�	�<L��Ad�Uæq�	xy�Kk�맗?�dS��Y��7Gg�M�����?Q��G|�l����?��O�D�07�ƾx�yr#��nᛦ��:s8��20"I�qz�AƤ���p<	TM�W�U��Q�}

ٴ-tB��T�	N9c��S^b}��I�Q�,���O*˓ q�xأAN�.��l�r.�1nA�<�
��d��c�
y��X7n��rgv���~/�Ƃ
Y�:hY�d�"n��{�ǁ�yb]�L@v�W�������O���9�'���W�L7�:M�Pg 8	��#�'*�-?���B�������	�|��+I�e&@-Ս~���a�+�]��6-�X��S�w6�p���7�!���5�i_ h�����JH�f�Y�v(٣|��{Ϟ�I9�M{��������2/��8��E�_�6���#��Ә'L"�'�Bx��
$r�pD��5-_h���ś�gg�O�gP�&7�h�
M�w3��ӁM�˦)��џ,�i��JՎB��D�O�$�O�#S���	R'ӎ_��d�A[�O������UU�9i�-�����v�#擢+{x��9O6Y�uˍ#��eR�.Z:T����s��-s��k��;|�h�uL�.q�tq;�J��yr�~�јu"�z��y
��/�7��O^��]�O�&�4��ʓ�?���?����\D�%�'��<KM���T����x�ѨE�~9 ���|�ru.T�y"�'Ą#=)�iW�t�&��?]d��H݊"P`USpM��
f�ͳ	����O2���O���;�?	������T�5nm��鐃N�8��)��%�R[���yW�ǫ�0=�rK��f�mae
6T��հDB�Q�6�i��ݞub�b&��V�����L�����N��u���tx�����۴��'��b?��E�����2h�~�ꙋ�e,D���7Ƞ��Ʌ-���5���)�I��$�<�ɕɛv�'�B@�jPؙ	DB,�&��i�%N�'ވ��'��2�~I �&���f�iPN�%,.�d���|�� � >wR�E�:+
A)��(O�xxv!	�	��&:#+��kwȈ�Dg�H�d-��n�M���o;t:�ɏ���|p�~�v���O����_��-��k����1�b�O��d�O2�D�O���h�O�=sDF�h/�ED��5����On�l��qޚ��ᖊ� =0��I�LG\\��dyr�H���7��O����|J�L���?1����EjL4F�v����㯇��?Y�H1��Xt�R�zaV���\a��2g��L�hi�+��Yȃ�ʽ#��M���&1����А>	���]/��R�"=yP���[({]��� :�e�]�c�����^�`���d[���<[��j�h�%>I'?5�&f(\�*l�N�����N!�I�H�牕1��2R~���Eo�GtDRG *��|"��	�@'�(!�Ɖ3f)й()G��f� ܴ�?!��?�w�B�"ր<���?q��?I�;tҸ���: �l�`�00�1'	\��J#,nӘ���&��#�1��'��[��C.P�L��E�Zx��̴��`cfƀꦽ��̹;Oq�ɧ� t��g��q�}�$�فdl���MϦ�	*O ` ������?�OJA�n;�HS���O4��"O@p�WB� #�(y�#M�E�z�h������?��'���#�Lx����C</��mh�N�3l�t�'g��'��o����ڟlϧ *�*��=ݐM٤��*]#,;b���4�"��Э��{�L���DO/���/�&�|��%ȉ	�z�aE�7��g�Jq��ήg�]ِ%��:S�xІ���(O�� O\<d�8���x�h�#׹:~��s�^�nZǟ��'Fr�7?���D��9��U:d�M�qka|R�|儑KZ4�Q$\��B�zP
ޝ��'F�7��O\ʓLq"��]?�ə{��l��-32e�b����n�^5���@�0 ��H�I�|�k�?;o@ S���]̜m�d9%���r�E+8>$�`�A�f&�-"���.�8H����"/VQ�ԯI$1 �BakǱUH��2�/�,5��f<��V%�	&�MsEY�H�e+P��R��E��Uh������O�����Yk� :#ξST�}��D;�!��OǦ�4� /o"��S�	*^�x�ov��'_��i�a�>�����	5O�����w�t�p�&ר��W��2���D�O�,{RjW�H�"$!�V�E�h6���ɯ|T�ǷL|P@��M5�����B�f��Q.Ss e�C��i��iiuo"ҧ8;8,�d$�2lؔ8��(Z�ﾴ�O�%qF�'kR��ٟ��7�T�W	V�3�؆�bd�Jlh<�CM�5%,���˖�pe���E�Ԛ�􄑮]�����r���牕[��'��}Bdb[���S��H�޸(�*B��y�I�2���{D�Ȝ;���� �9	!�D��
i�}*s�W	�� ��I�&[!�D	./Ԉ��#'M�%6`�$�j<!�DKgLB���H)!���I��&*!�dO���%ʮK�2��pI�q!�$ x����R �Ax���'�9X%!���0�@�qh�=q8�:��$!��E��zp��wq.��C��l!�@0����5iW�;`:�B��i�!�Ą�8;b�Y$@�R�ы'��>q!��.�h�K� ˭5�N�kb�)a!���W{\��� F�h�aa�b��!�DϨx`��Q�#j�}0恆�(I!�d޾Y�TA�� :V��R��00,!�XVT؉�e �Xļ8�eV�!�d�79���b�:FL�Ţ��"�!��x�Լi���;7TaPő	+u!򤞰���1EB�,7n����!�!��	C�L�R���&7�}���!��!} �b� �����%F�K.!��"p�s2����0�%N�,w!���T�Q�Z�喐JC�B�!�P�k�Tљ���L�ja˥��'J�!�q�\I� ��${���*�'N?Vm!��2)u�ܘdɋhN�a:� ��{`!���"/L,i�/�"n�غw�)
�!�#zK���"o��Bր�7��.t�!�$Deu��P���!�>������!�$ő8�HX���4~��Iɑ�`�!�$�<��L���U�T��&!�1&�!�d��^2J�(C7q.1�E��31g�	�L]�T���Oџ(�!�ȨA]�����x�
�"�E��<����MH����Fr��6Y����;	]�)���� 4jČ!R��e��x��-,���@�N�8b(�R���<y�V�?e2a��B�z���n?_[��y�ȍ\�"�`�&�ӿE]x��T�ځrvQ�}34�n(j����V{fi���;�'~KvXc	C�F_���i�%w�A�l�%q0%k�-[ h��)��<1���D�����H����+�LGcl��J"��D�C�O&�c>c�ȩش`�`�#c��55"X�1m��<	BFr֊ZW+��ZS��>�W)�@����Z�Vy�q���s�2�#T�/h��Uf%�[�:9;#!SټB��	?az#B`�#���x���`4ޢ>���b��92�D߯�~��E�v%
 ��]������D�"P"<)�J*e
��B�O:~|����i?Q�`�3�=I�JG�"���@�єB�j@:�R�U�?1y����J�!���iE\Ԃr.S�? NA4J�5\ܦ��֊S�5������0#Ty�Ae�-)-8d[7'�
��
.S|c���-��4��́;0����!U1 p>�۰
^�L��(�*=�R��M+Q�X��!�
)�d	��g_׀DQ���>���68���<i$O�&�"� �<QaH2V���C�2#TX��OE���"gM���>!7J�%y��%��Ɔ��D�B�d�ƍCt�b���"�>�� r��ADAܠ�(�D)��Z�Q���"K�<R�@Չ�o���#<qr��*����b�C��~b�1�Θ��?�ɉ�"�r5�5� �f�<8�t��;��* [�\���zVldr⧘��C��\���9:�lep懍�0��f+=#I�d���E�v��		gƘ .6r�1��Y���*A���T.)��#�<���U�6<X	e������&�]�:��I[Fh�U4HLq�+DJ�^4�%���%��RA��4g9B����MU�0U�	85�����Q�{o@�CZK�p�oN�<�u]?��U�v��$6t8+���O��b��	(Y$e��;�i���Fʘ��1HB�a��#=�;R�%�T	����a�VHgFs�CN�V������k���:f&`��R�i~.�1K�_M���mQf��?Y�Ө!k�J��ү�)#�&(a��ga�OJh��I���(��Z�Z&-ْ���b$�*�ă��,�HW7��@)A$W�O���boǲ1��u�	�2��{s��	���@G7F|�A*G(O�w����c߂T��Ew�U�=t0J%��\�H�aN0G\�G��"���FiE�0QvdA��L�Y��H��I�eF�Y4(�p�nP zƹ
�Kْxs1�Ǉ��
2,�]#܄�dY�y�����i�9�	�<�v8��A�+l���@Ņ�p�����o��}Rt��\[7"�I=�����l���$
7�BՂ��t�věz���(�ByN��+@/�+!7@��C&�rz����^r�]�S8�Ta�L���@G�/$����i_0�i5�ȓ��h��5q�����c�<��{n�P�'l�0!�.G�N�@"�Q3< ��1�	/@�$8`���\��9�
�2"��C�L�"�%KK�~�a. �~��Q��Q��4��#���~�����'�O�@�0Y���$Y*=����'�!Eh�������c��vQ�����b4fu�sh�,I�x8�=$��k�gW%�yr����Â@�".p����,Ub���
ٰnm.ehbo���V-�8()����B�f�`1�2�y���6��#�L����!FT.�.��`Z�X��H+j��˾DE�Ӆ`��*�O��Is�(��ӄȻ}�d`�5 5Fd2���?~͈�ٓFF���1 u��]�x1�Չt�	Q$� ��S^�6-�پ�p��M@Z���
ߟ��'��d�������#�(?��R�)CCW�`���6��'̒�҂NF�~�s�DC�zN>�G(?	 p4!��Q
�8�-��{�l�8C�J< ��j�O��/I࠰Ƿ�
�:�-��;{l�:G�[2x����&vxv@��hL�Hg�E[0�� =@a`�o�m�5�p�J�A�N- T2�fa�v`]�<Y4�� D��邾i�=���w�1���۟G�>�ۆ�۱m��Yzsf�o���{�㓜-��ي��U3...�a��!�\�x�o�0A�^4���D ?A�F�0S>��O�m��.I@^�Z�͟�<�De�f��6:m�@�EH�'^��ɇDD&�y��Lh���D�: ����>�?��O`�SE�yT�>q�w�;��u�0�Y�sELx���E%dyGx���/����6i��g��(�`�	����Q����@C�=�\��fH	1c��Ic��hE�Hj��ܾ�li1���;U���Vl�-I��s˗ 
N^�5�2+E��Ӗ��+z7|���E���!�����Pt�E�,J�rר���B�s!�<)��M�n�bM	Ǖ�K�\zU$[g�'�vD�3�S�E�4%�S�� ��pbW4��'�ў��?Uq�䃤�U:����-7���Q[�^�R��I�/�N�p��j�ա�!O� U�5����.U �!d��O�=E�ġ=O��I����� 2�[�z� iC����K���Z7�!0�K�: ʓ+<��@�%Om��P#} ���'r,x�=�0�?�KSKQ�<�� R����X��?~����@��
� S�M1�N�U�0�C�{���"�V�
,�D������0�������	e�'<O�p��	�6B|�
������G?.x��!�����F�!B��ђ5�Z�&"Jir����c���bT�V(	�p�$��H&^�m���Q-��<��05$�?���ό=~֬��c5%�L���8,O�X$����)0��А�	d�k ;��ʓ[�T����=�)�'7�v	�S8iF�E�C�p�&m%�ԉ��&2aqO����r���VP{��٢%P�e �x�U�ˠ%��	q%%�S'�G�q���Jz���=��i}챟��ObJP�`5���:T��3�(L��@9�Px2�X7CKNt�b�@"s�L8a��ѝa�tt1��Tg���f�PB�'0>D�A��͈)x���I]0����	�Q��3f�|"��������FX^0ّ� I�����vBB��{��i� ��58� Z;
�x!3�?��'�h�@b(�{�S�P*��	MN$�}����I�� &����%�y�AE?Nz�e�fK/q6:�Ss�V�}�qOܨ;c#�^��<���>Yq��
+G�`
�mn�|�#a�!���7�
)�J�r�gr�Y�v�_�)���@���J�v��Q2@�r�DҶJ`��pg&�'8�ay���-�a%�LJ7�U�gRd�q
�yZ�H'��>��*K����"}JS�ʲW�F!��_�C�Ё�\V�	�`��9���� ��QvI$IY�YkPQ
�Pm2��xҨ�T����牸}��R�eZ (��D�"�]r���sf�J�y�ģ<�Oװl[�/֤��PY���DÂ�
�-K�Ę�i�w�'"���,
6�yG��,�B��M�2e�$T%�S7�?Ɏ��>@d�g���G � �PK�"rp8�E�x�';����3/@C ��b���r�OJ����x[����ʓ<^�x���T�l�?�u�X�-DT�h�A���AcV�Ԩ_p�l@�k�4���1a&юp�1O�&D8FqJ���=S��
3�3��'����G���P�P=:ou�v�+}^˓u�{�m�9h.�{!�A�Ge.�Gy"��
��U��%�'o������_2|`����?}ڰ�V%3sV�ʱ@T�a�T+2�҇MnT07o��\�Q�4B@Րbs.杌H&diy Dh�̚ ���*��hO>����<F8�+�+
a��=��A�v��4Ex�&�f��q�S�G:TB^t9@+��e"�+�'A�=��$Z��5�g�ޟw'��-O8��J%n��1w�ߛS	���I,W����C�ZZ�3�Dn���p�	N=N��x���:q^E�R�/���'���¥���T+�b���[U�D�s�m+G&���dE�S=�Dʲ��`���"�� -sQ���2�0�)�TjW=)�
�� �k� A�o8�@.3��O��$j�d{��I�^��0R&-�`�0�9��5Z�5�р%R2	�3�Ӻkw��+4:5ͻol���kK:SF0��A�� Hen���fM	���
�y��H)��=�?����cd.���M�ra9���O�8����#/����`bкw�@-���x�eZ�ՐWj�2�TqAF�G��vT&�\}���<��۔9"��:���*���moj�	5���7�� 1�\ P�TAyԎ����{7GQ��!A��H�K��,�D�*h�).<�	�a�ۢ5ÖM`�Ă� Tp扲��d�$F�,YF	n��(����@�E�nĲ�d�/	��bӊ�9��}p�G._D�&�����-�L)N����<	�o �<�X} Q������ȯ {��7��'R�|���OL�����ϼ�UfM!�l$:�`�m�T���@�Ȧ�����@�L��'�X!�m�c��S�q���A_1L��=Jz�Eѕ����8�td�WL<��1�G(I,T|8�˓MF�<�P	�?&�,�	S�M,N�FUc`
�
���#�~�SJa	N�"�bp(1�
�@�ht� ��- ,��FΓ\9(X"�D��`�f�*�
�8��=ˑ��ǴiJBi�F�0O�I�T?���ŕ�Y��L
�O<mo����u�Vl6%1F/��wIH}X��<n.�'�6��� �g�-`��4@�|وCQ��(Ob�lC�̖�\8�I�^���D�V�l��æ�l-"���c2��$�'liQ��	��[İ���w�Ve���ƺ$<*l1c�R*����˘'"��jT4�(�Vd�D1��|�a�z3L��/K���'��dW�"�r�6,�:otf�J�(�B�:�,)�iʹV�(����*O��#cAQ0릴�C�$ԔM��f��̀�l�0K7�[a B�4�F��f�,(HV�p�ڐU�"�H7�'-�y����43~���!<Fx.EC)O�Q���W�(p�U�&�b)�$副�6� ��G*�V4���9>�Xc#�ԑ���,��I(���w�����W=9Y(��6���Q�(x#`J�:�z�:>���{�HϹ5��yu`��y`���~m��D�P��H�Z�O܋&	H�6�1`WF=�%�@��L�j�W���'��8���=*���sҢиt+D����̾Nw��Q�Y�cҬq�O�{��\��]s���JW�qؤɲ`ͅA!�Q�1/�1{,t9�]�l������n�����HѝC�1���cr���j$`ט.>�Ȼ���m%�<��ڒJ��去+�����LQ!i�,���n}ހ�v�(}*���f�1D�nH���.�У*(�,� A ��Լ�D��J�0aaxx��0�-���>���D/Sv0!���LH��70R��f��v�F��!�^�_"<i��Q�[�`����T m��>��_�bY�$K���6�n
�(?I�C!-�
�$�1z�~���K*�y4iM�)���͑����I���0Ҁ���"~Γm#�tj��+�0����ò%�|�2�]�v���	��,3��3�3�	V�`��IT*j����C`X�&�	�
D��b�Y~��d{$�	%a��X� 
M�$�v*ݗhZ��6!��"�ҠDR(!'Q�|�b�U/*�杭3G�Q��m
'!Hĝ�7�K���8w�	�X_�q�L̉?s���0�Od��A��6w�r����I�Y��@���	�9^d��E��7r��~��kC�G��+#�S߸T�P-s�D4'�p���J<&�t"����]���Jt�V4{�!BEu�<�kB	���cf�Z�?V�e�V���ȓ}*<�S��dj�)'�ۻFͬ%��?���� �¿F(���R�_;R�(���"<l䨃Ñ3:��Ì��^P��y��D�CW������D�GX���ȓVDxa��
�_x
Y(����4��ȓc�v%rA�&{�(&-�S�n-�ȓ�����#B��l����y譄�S�? ���hQ�y7M�+AWL�IA1"O �r0�Àn��tK%
�8��k�"O��C3Y�X�R\�s�!V>\l8"O\rW��4�t�c�ѓ8XL h�"O�Rgȑ�w����ʞ�=�^�*�"OX��.� ����S+ĳ����c"O�J����QYc�Æk��$�v"O�"��	1�(�eߞo��"O���4NX�h�e���O��QQP"O�5R'�T4%"���*t�m��"OD�D��Z�6t��)��i�"OA�@�d�������
^��`"O^d�sLH�&Ą�Y�K�9k��P�"O�x[���_<$��9T[|��1"O�B MZ�.��I��I��ER�U"O~8!c�O
i�B\[3/�#pCd�3�"O��*�)�ٷnK"z$Ω6"O
D�c�C��-�0�s�2��q"O��Q(� y����+7��h:�"OL�����"��$�Ȍ�Ml" r�"O,Q ���!Z��a�"O��7K?o��`R�:>��"O��f;]�x���TO7j9�E"O$X�%I09	#�[�"U�q�@"O��ikʗ2�y�'���]n��#"O��ᣥ�έI ,F�,eL(��"O���R��LI;g�@�`^� �v"O
Y$�Us6��,^�[T�V"O�-�w����=���S�JV�@ "O|qk���`�^eH��\;<�4�q"O�Xv��'KD	ɷB�9�N���"OPA�F�~�2���A�.3Z��bG"O���$B/H)�!��*Ё~G�=87"OQ��hմ2#hػp�ʡb"Qk"O�عe�	�B����e�|C��"O"���R>a��QBD@;�I"O�i(��M�S�5{� C"*/���"O�!C)$��@@�>'*�y�"O$��lQD���&a�&��"Oz@;��>���t�\/h�LkB"OJ,�rK NB�Q)#��15{��"O�X���G���@�K��l �c"Op|��G 5&�ibj��.d�[D"OT�K0��x���R�C�*�e��"O$� R⋩D(6�
C�y_���"O��i�jO��<;ˏ�sOT�P�"O �sAԱ&�P,Չ�%S!Fxi3"OPty��ɪ)�
���܊� Y�"Oꅫ��n7|��A'G
��2R"O�=��0A�Q�B!����"Ov�) �Qr�d�Yp�	��z#"O�)�sG�b>hp@��J	���"O��@�Ӽm��	�oY=�t��"O�1ۀ�	
�2�s�.W�l&y)W"O
4m�^�K΀m	"f���s"O4���Ŏ0;N��x�i_
!���Q"Oz��`a,(��X11��s��<0#"O��/��z���kY�[�+s�<Q�FG�|8 ���1v�}
%��n�<����h�>����B:V�th���g�<	���&!�E2�C�T��;��N�<a�$;#\��	�A��FMn��q	�f�<���>a�bŘp���/N<�R.^�<!�LG�r��4�����t�S��W�<� l��h�' ����ܤ`�H�z�"OԥxA.D35�j�$a%/����5"O��!�fQ��z� �2e�<�"OάAVMU4"%Έ��ZSn�"O\��ڎ?k� �TMF�7�T3B"O�x��ϧAX��s喴~����"Ob�ybǭ��Uy�m��o��۱"Oxh�&���3�hA��9	��"OHd��n�זa�¡�X	��"OtjFV�3�>���!@i�6T��"ORY�7G7Q�nE� c���V��"O�E0&MZd���u��� �\���"O �X�oǅ��D�4��~�^��"O\�
�^j�k`�ŝ`���!"O4���ӂ&gXA��H�G����p"O,�uC��5��|��욲�N4
������B&� A��~%�I#�AJ�IfP�>)��)��]�ty���*aNG�-K�!���"�La����lo�%��"�yC!�$^�O y�� �7
ɾ�Fa�&q[!�DO� |� ��a�J�G�U3t31O�����t8��u��~��I���[�t!�בLP�<���	!1�N���,�C��3(H0B�V�sx� r��=aT�C�	4c����gШm����Ƈl�C��".}�r.���|��)�'�C�I	��`9�Ǘ*l��0�u��4��C�	N!Nxg���-Ґ����
��C�	�+LX��W��*:o� ��,
�V �C��%+�4����H��
�bȶ5t�B�� ^��"5�KByp��lF�U\�C䉅q�j�3�Π>�D�	b�C D��C�I�CN���'�QZ�*��mE&C�	K�,�j�2�хKЪYg�O����Y��գ��a����#�B.d��x��I�2P�Hg� �<�Ay���<<PC�3A�0����I�}�$�M�"�C��vLt@�b 5*�|y"	[;0?.��D���B�Z�&a�x��\�f!̜�70D����W�91�\�$��L;����.D��C�%Gx`���s-F*eG��s2�'D��;&J��H5(&�3'�Dhe;D�t���	/nK��GC�	 ���E9D� ��H�tz��� ,QGAd����9ғ�hO���a!�	��
)3�O1�PB�:L-Ľ��_�,-�[���NB�	(b��3��t����bC6B�B䉍pZ�U�
+�ʜ� k_�m�C䉈A��-���v<}���^�T��C�I>����h��E��������C�8a�%c���>��p�dH�1�B�I���!�B	8y{�����83<C�Ʉ���@���-9s(�B�@��B�I�Bh�p�6�ҽ{��e4�^�d2�B䉈E�D�X�cC�hy����._�s(�C��*L=1� �9t��\��AB
>�jC�?[��࣌�#W�\���-2	BC��h�V�;��Ʉ;͞��լݱ�C�9-��[b [
M��Q�Ϝ�!��B䉕OP�\	�e���=)d��0ԸB䉯t�µ�����R��Ȫ�L�:Gx�C�ɺQ�qB4,�9�4��fL�)A�C�	6:�h����I�^��a�SdC��
vM�2�)A�1RFQ�C�D�E�8C�)� b!x��"p�~ �@�_�K�p�B"Oz�`�/p����K�'�~� "O�hzQ�D�yn�\��'J1�Xv"O.Q��QRJ:օ�s'$� D"O^�`��^���t �D
xk"O��!�h��mCX�1f�V���4�*O��XÆ�.O2}�hΆ`����'c<|�&E�V<� C�c��);	�'VF��&.��)���6!�&]۰�b�'V&�#��b><]����ZBT�p�'��� ��Xm�1f��CA��q�'�@�� $��z\�1 �ޑ3e&y1�'�6�p@ҙK`ũ��Dv x��'a��cME���	z�ˀ�{�(�'+z@�$�/U2�c� �x��i��'�ĵ����+�8\�cE�m��:�'^B�%�4X�d�jr�8X��C�'W�(`̣@�hR�!ާTu �
�'�0�E����fN�G��)�'T�=��K�B�zh�#bY>9gR�I�'�^��W�E74������7?�X�{�'׈��	�|�c��j�岏�� �zĀ�E���Kl���gnC�O��ԇȓ�Y�AA�@Ú|����*;��-��AOvY���$k�u�3$M�|9��K�a#�Ӗk8��1JH�����lJt*"�¡X����*�	��p���i7�<D~r� �d� ���4�����h�4�y�	��<�|	��o*W꽸�(\��y2dZ�2����'NU'�BU�2���yB�C�pӪ�q��/���
��5�yR.^1v��ԋ����L�����y�Y.i0�0`F�]��pS H��y�	�q >�6�D�]`�0c��ŧ�O��=�O��q*s�< �,�b�m�h��'f}�3��D0�,PtO˕l]|H3�'�2�YG�ބ;>�h
$��i�����'|,A�R
J�q.$�"��/�>p��'�@�ԩ޶%����dW 90��'��aS��[��9=:*��
�'�*!"�
	>@N����oޚ/�N�[�'wv���fǮV���qK>$z>��'b�ڐ�
�T�9q����J�'�̒an���ȡ�gɚf� ��'��E3�+�3P���p�@�^m�!��'��%Z��#��t�׌W&�)�'��%��O:
����g�V���
�'Y�Aq��Y6�ca�UݖT	�''�}�y��L�:�Hh�j�"(�C�I�T8�r��^�#U��� խ#��C�	'VX`�%�=$�e@����B��>+�ٗ��;qbza��
WVfB�I�4h��#�Ǡh <���C'GB�(8y��ŬST���� ��o��C�	Bk����h��cc|�{e�,Q��C�	�!�paˆm3
$��Y�e
�G��C�Ɏ��5[�C��V=v� תD_�~C�I�R�b�3�܊�NYj7.D�X�dC�I;X�( �CH�;�MJ�f�
?�C��l�>�c��^��`�*�^�8O�B�ɤ���D�;{&����ܤ%��B��?4�2m��c�+�LA���E�8�RC䉖���{��3E��B&0 �B䉻O"<D������ U�j>�C�)� ���g-+>�T�Za�X�6���"OH�%-V�r��7�R�,���Ya"O�;���/x��H �MQ��e�"OlupW��a6�tg��%a*J���"O�8aV�#s������z��6"O�����I��RnY�Ì�Q�"O±�6�\F=��G�&��"O��qP͞�`�a��e��
����W"O�IWj�O�a��A��d�6U�v"O�q1 _�l%(\�rK����"O��r�
�;-�� ���G��[�"O���` ��F��m*����=0�';�ؒ�(8|�u�,�) �H�'�\�Qp�Z;m������n�MA�'�t%��M�U���d�͚|�RAI�'��R�(ݗ&�=�ԋ��p��I�'N�豤��/�Z��d��$\��P��'A�Ѩ�&"y�y1��՛A��@��'4(���
6��%b���f?d��
�'���cN�/y�<e��
]k���'��a���Rǀx2O��[�d|�'��-	T�5]���1��^-O�nL�'f���G[!wqz�{���8��h��'�X�$.ǝ�#ѯ�
�h���'�KF� i�3�Ɵ�x`���t�<��fįG4�H0�
ݱ "�ً�Mw�<)G�ځ2��34DRr�l�'u�<!�!Ɓk`�`�����U�]n�<1�G���`��@C�Gm�<i��H/i�XJӌ�.!u$)���o�<9&+�&u�����[+�j��j�<I�i��*�IPdLU
?��B�L�n�<�`NبtK�I�MD�����j�<9�a�b�����ٻ_�1[3��ȓ7�����:Xd]�ω'B"X�ȓ=8J�y&I(T���%Ӽi�@ �ȓyl�`[)9X�Ѱ����	�ȓ�hd; �P.xZ�M�u�nɇ�N(Ҩ�t@ZU�z�¨Z_쑇�-���̇+2��1s"�,d��ȓ?P�\rF
�nŮ �� %�t���N�d�7���V݀B
C;!e���y�*�R��Q�4��0#׋�m,:A��S=��"��9�<�d���"-�ȓ	��i���"+�,��@�ؙ�h��ȓvx|���%�� �E���ȓr�d<�����v���J_=f���ȓ"� �b �O�N% �)u�ZZ����v<��O���PzG��?MM�ą�r`�y�-@=:�b�SN�I�|ąȓ�֤!�IT�C�2�r��=:DE�ȓ^Y�hP��޿*�b�:�J :ʘ!��^�́��ʥ{�J���Ԟ4v�	��!iڕ9�Q+�(�����@��4��Rԭ��V�ڸ)30��[E�х�VΔ=��Bߩ?��"v�1�u"O8 �UM#;,5��JQ�<j�y�d"O�uc���e�.�*)�aeX	`"O,��Ƥ�;s4*�J�C�E_*x@�"O<��uFz�~���dW0k�"O )J"C��v�̏~S�YÇ"Oh�@�H��6�^'`��5�T"O!cmoÚ-��c�/f|��b"OtQyUjԔR�
���!��9Ѯȓ�"O� �8��RpN�9"��P�+^ʅ� "OVmkBGM�-�d�(�$Q'-M8*�"O�P0��4������*�0"O���6�\��q��{ `� �"OUCc�R��5�aUGT�|J!"O�.X�Lqm�!�T�Lਤ�n�<��JMD��B����O�ְp@�Si�<9&K�oF�	a��
����"��K�<�`.=��(XJ���cmƹ�C�0��y�������x#d�Ŧ@�C�	�xݦ<!%'$��x����I��B�=%��Ӕ%ԒAؤ`s�eϑk��B�IP��vc�,���A��M(��B��<u����2��r�����(��B�I0�bEP���y�D�Y�&��
�B�	)'HN=��T m�����ZC��;Q�x�Rec	Q��3��>�C�63G��3��O�J�� ���M d�B䉯 �87M�h�ޤ�Dm��>G�B�I�D5��c�H�7A��)F$L�zzpB�I�hbl Ȱ�Z�U 6ݰ2LݡW	jB��=!�^��3��3?t`!SD��9gՐB��5-gZpFbP�E�#���>!�$إj�X���S
$�����SX/!�D�1(�l��i#~&@�#��pv!�$F�>4E[q`	�r$��Ǉ@�zC!��mj�Q��	xf��I�'�6�!�d��l �A���W,���fR,�!�$��B�$��QfC�`H���@�=�!�$��6�JHe�P������ �!�R�I���YcBۀ-��5R`�8j!�dZ�lWT,2��V�[u4����;s_!�$�l�h��ɇ^����̲B!������hZ� ����� �4!�$�4zD�;6]�c��V"�<G!�$��S` �Ċ3x.He&�@!�dռ�%3�͆Yg^�	+Y�L!�$�4+�X�)�l�3t�"a��ρoh!�G�>����S ���Z�HPh!�DDPiP�y��V�L�
Lå瀵}F!�DÒ8j�fW�h.n�rs!�	!�
J龜�L_�c�h���*G/!�D�;8�a�B&',6�p$�wE!��"�tp�H"S{���F5�Py"'��}��bS� m,�X���"�y"�V@`8����.]���S���yR	�&l1AvkQ�%� C��+�y�W@� ��k��D`�핬�yb��:?�ІjJ� �N��y�C��a���(���DP`��U
��yRU.ppx�[$�#6+�!8u
�%�y�.�)� ��1hշ,���"��A��yr�FMtN陧'R'�vEB��'�y�H@]sL	X��{����ʣ�y�BBZ��̂�� Pi�b؝�y�HԾ?qxD�QN���U�P���y��ơ��@�E��}48��&V'�y�@
dQ�8b�ͨuT�1`sW�yr�.�ؘ��(L1"�D��[��y��q�šA9�.!`��S6�y��\>X�؛���=6n�P�[��yb�,S�8	+�ΕX�����y2�ܵe`�%@�E�"bs�)��Ʉ��y�ۢ_� �W���ڵ8���y
� �y"�Y!��1
�.�G�hܺ"OXTA�/�+ݰM���O�@�x��"O�4�R�B9FM���m�$$�"O����ԃ1$�)�r��	@"ONq��h�5�=@ÊQ�*��b�"O��;gO�) �@]�	�D"h퓥"O���4ʎ#	F^�rhZ.'>U8"O$M��dɍ'��D�*яuʪ���"Ol zm���"y����2�h�c�"O$�S�
_�Bz|\�g�؉fx��H"Ov x�bB�@7�THrCY����`4"O� P��.[A&S��6��4Z�"OT�
sɈ7^;�<y�Ɵ�(}~�7"O��K��p��f�=?�~��"Oxm[���*�*����(��9�%"O�$Zco���t�Cǖ)Wh�1�"OnAQ�h-p�^eXakʸ4V`q�"O�p�`�$�<���Q=2;r"OV���dG���m��"Q�	:V�zA"O�Б
AHq�a�ǚ�5$�s�"O�1�f��:��Q�&L uAH�0"O��@F�}y65��&K�[7R���"O�����d�`�e�.0��]��"O���`N$Q�~�r�DmPtS"Oh��-[vl��$��)�A"O$4Ф�N�3JB�0TB�'��9��"O����+vF��Y6c��QG�U�W"O�1�aX�~�D��^�襈AN �y��ݸW��y���$������*�y͖҄L�X#���J8�ei JD��y�o�"�)*腄E~8������y�`��:`�!�@	[�
I&ɂ�y�$Թ ��}i¬P�st�pu�y��P:�
�jF���^�	����yo&R@0��7c�-O a�����yªĘ?c�0c� �1��p;���y�J�;Z p�A��).�ad�އ�y�.��
p���6���3EJ?�y¡ܛj�@y�݌��aa�LѶ�y�b
o(�d�Y��M���y"Cʱ&V,�a�"á�V�k$(U��y���W ��i#�{���"g����y��A�"D��&)I4
�N�8���yR�<�|���ҝ~.�ppC���yR�d�v�xq+�pܤ���,̰�y/�n&j,R@�T���Y0kZ��y"-n��`B���E�7j���yR�ޜ
�8�*��JɁ�� �yR�G�B>��; dK�=�Hͩ�ͻ�yₚ�2�*���~�$E
�@C:�y��!8ZRprWd��D�:h����y���'��J�aBɜdK�MX��ybDX.J�TTKrH�'<���0a�Z��y�o,�dTɡ"H�0>�
�Ý	�y��Y�"UAKю0�X�q���yb̙�ug���O&*09z&�� �y҉�.o�j��U�%;���0�L�y�́8��c��6uf졉� U,�y�%�W8�po\�YkH����!�y�A�f��� !��A�=�Q��;�yRdN��[5'�|�6-9�Ȑ�yB�ޭw�|��AZ9\[<��e(�y�ƀ4�^t������ �A�'�yR�^���Ar �_�>�ԉ�,��y
� �0z&��DY���.g�T �"O@�(Y5�D�h��!]�Ţ�"O2!qEH�=70�\����<M2H� "O��a��M;�xi�)<$Q$"OTX���"�$���
�i$L��"O*�h�JT'(�����O��%�b"O������&YQtL{�&P���0D"Ot�ْ!\Ԡ���=p����"O:x�şxޜ��qd-'�͙u"OP��Ɖ�/�x����g���D"O�����I�8�H1��$��"O�XC�� ���(4�F�ܴ��"O*)�2�� ��4r�Fl�t�"O4c#��[���1�d�����"O�x��FZ=hZ���S�rz��P�"O�h1���2�����5o�+"O��R�jX6(	jiie��~fZ���"O�Q���3=����1����"O��)aES�dp�����6x�G"O>���6W7�@�S�M;@|]�c"O��H#,X,M���P�E7htC�"O)2��M�+�&���P./gX�E"Ozp��č�
����׫�,2Yl�1�"O���w�ŧLM�ܫW�Jv��F"O�<r�-�+Z�Ѻ�1=��"O2��?�5b�ľPt��"O�H�EM�4��铴N��l� kS"O*\�G��<z����n�t�b,"O\��tm֯&�4��&�A1Z�0�33"Ob�c0@8b�(X;���$}��� c"OJCGD-�1Iw,�6�@��"O�YГK7g��``,$�|q"O��ԧ+�P{m��0�pHG"O�(�固b:�х�ҐfV鑒"O����yTMh5���-b�,;�"O�� �Ʈ�`E#��Q^GDxYU"O�S+� ~��"��#+*�)�"O�8���� F.��,����2E"O^8����1_��+�2"��p"OB��a�"8�հ�J�(�T��d"O�	J�8�F�pь�9gO����"O���3��*4f�4�6jg��P�"O�4`0� �E���K Wlp��"O�l�QbʎZx.%�G�.*c8Yg"O�-��jM�cL�,8�n�OR�;�"O�x`s�C�nɢR�B�8=e1�"Oҩ�7N�:�6�^�X��,�E"O�����`Њ��kU�?����f"O�q��[�?�T
�+��{��!"O�d	� �X����ꉙ	?v�ȧ"O�̃��[�@�7IH�1�u��"O�@x2�άUw�1YT��-H�����"O*0��e�w�dI�/�l�a�"O��hġI�]��8[�@��d�hd�'"O~�`Aa�?P*��p� ҏ]��$�"O����@}vr}C /éN���PG"O��rH6,HD��p�1"Oڼ"4�E,E�n\�V́�^�=�"Oν��A�����qa�/hl��Y@"O�M���M5H8�!�h���Js"O`�bE�J=]���`����eb�"O\@iĄǰR��Y�SB����"O�-A��8Ty�@`�nSH�4�K�"O �Rh�p�^̂�l �~�T}��"O� �@�@
�-<8�� � �Zn>y�`"O�ț���N���m
,lOu+Q"ONj���N%rPj��K��@�Q�"O���b�o
d���L�$����E"O�蓀�G+�z�+�1ͪ��0"On]��#�t��k�-�+R���"O<��sJ�N#��A��\ �"O��n*Z]R��!�0I�nH "OBt�2h�2͊�I����B�~�D"O�(�2�C;h0��'��0P~�z2"O��jG�P�MSL������Z�"O�����l�@�BQ��)�z��G"O$���!�$Rz�0%(�X%�D"O�A
g�¿fۜy#M��%��1!�"Oxp�Ү�I=Z��L��z���"O���)9<���EڢP���X"O(�*�F�x�:�j��	8M�����"O��h��U=�=�R#G"'�0�k$"O��`�L"
Kr�b��܌��G"Oĭ0�B�<�h��ć� 6��	�"O�- -�����9�� ��r�<�b�Y��4@�&�Hv���t��k�<A���)cm�Q�L�&�܈����k�<�f�E \��tf\�U�NA��Țh�<I�n��p3�8e��y��Kg�<�a"�6��`C�=��Lav�]_�<��E�\p|�G�9��D��nZ�<ْ�?�ձu��2T�6�)lY�<�cbX� -V[')M9Z9��oq�<�To׺7�pe
����t6�x� m�<I���(J.��wK_�T�j5���}�<a�j���<`V.D�p�\�5�F@�<��),#.�H����.v��� Bz�<)���LC�l(>K$8���v�<9�×�Q��@��$�Gؘ YIu�<�C�4l��b�>0^t�G�s�<I�!	�2x�T9��������s�<��E�1o����.�R����6��q�<!@nX�
r|Iq��qÒ58p�Rp�<Q��1l�dPGڭӤ���Oi�<�pț�h�7hM<Y��%�f�W�yBZ"+�D�	�� �șq�d���y�'I66`T��C��t��⢏K��y�!B�AJ�1;r��mA��y�� �y�Қd�P�R�O+�����yR`�),}L )��	4������yRM�+���xW+���2���y�-�?2A|��I�;�-��n��y�F٨x�¤��	��d"G4�y�Ü- ȩ��	$�p"!�*�yReE9���)5�[�=0 l��yr-5{������h 1gÝ�ybo�j��i��*Q�v���ѢK.�y�@�6B"8���K�l�� ��μ�y¢@�F�x|z��!aZe�U�M��y��{���	�B6V�HBu�_��y��WT�PeYFD��=�j��Ej�5�y���[7 A���B�$L�	H	��y���-��!��$�����yrL@#�F쓰b]̔s�L���yR������*R10���Y ^�y��ˋ;|T1�H�?a�1D��ybߐP�@�#��M�����1�y�����`C�B�m�������y
� � ��B4�޵��,�9n�X�z�"OىB��4lA�I �:d���p�"O�E�֠�%k*hR��Q-G��Ph�"O�H�&�',��v��#���"Ox��錂4F��g��B$�5�&"O�yS�!t�$�t�R�m4Bt"O贂0��=pd�@�L�Y�|�4"OZ�& &0#�$8D��UH��"O.%x�m^1�T�����	A
�
2"O��q��i"�D����l>\�"OT�Z7p��M0N��G�I �"O��X�+d�p�����2a3�"O|���vr�yj2��6-ܴ� �"O�@��*_�n����*1<��"OF���f�{����iX �DB"Oj����PG�t�M����p�"O�y�s.��"�X���扷k�*��"O�����ܞb� z�K��UwQ��"OJ���ǐ�& D��#J�	Gb����"O�9a웿=p�јc)��j�N��R"OP��nڍ*���pC��w��x�"Oʭ����	$$���pG�Mν��"OZM�$Y3;j�Y+օ����3G"O@�{�`J�a�����ɕT
VК"Om +B?Bpع{TCF����"Oh������2�Z�:��J(=�&I#�"O�YP�N��t$J�!Ǉ�-  T�"O�d���=��y��FY�X|j�"O|e��aT�\�ؼ�!OE�2��"O(i�c��N�B���:�Ie"ONl���ÿ!j�0b��R�_��P"�"O�Ū��8~��8��"ǂE� � "O��Qu�_"\�����z�pu��"O``RhC�I
>���n�BE"O*ɺ o��(�D�^�2"O�tä�Is��qun{̲U�%"OM�E�U�u���7�R�c��4`G"O��r�]�n��r��T�h� �"Oԭ0֣̱_��cr��|$:��W"O@u0�k������䔀z��"O���Շ�9.�=AgN�=����P"OTHbF�Q�	Un(��*Q��"OL�Q�	�F� �y��P�9'
��"O�4��E�~ �uW�V��x�t"Ot]���'�@�a���0�"Ou�a�_2]���ː|��"O���׀�5] ���Fɋ���xI'"O���Tl��t��Q���:�L��r"ONQ21D�L���Q�喔���"O�a�sh�*>�و��u�B1�3"ONa�bJ�/� �3��^�Ĝ��"O�X�$�_A�6`��]6>�p�z4"O�(�"�'A��� ձ$jp��"O~`CWC&"d;Q
�"���u"O�p�����p�bܠz2�A�"ON%S1L
$,�t���J�&v��W"O���f�1�� gc�(4ψt2F"O��X4Oπ���`�"�W�l�[�"O��:���(��t9#�~�l���"O�hX���--�Aʇ�1PJ%��"O��ّ�:HMJ��o��9�DcQ"O�p��ĉ���Dwg�>32T�A6"O.娗�W=xD쥡2���%O̱"O�s/=&�<���+gK�Eڒ"O� �Ei��@(5'N�S��=m/&$�b"O�)����
,v�AbV̄�Xx܈@"O|�`�E�)�@�Q���Dhd�ۤ"OnH�5D�m��ip3��nW^�*d"O����	�%�������l`!�	�'��xbwa�Q
�T�bi�5<s��#	�'�D%����d��5AR�P4$�M@�'*���@���pb���'�~ �'M�+�,E2�H	iI
31�0��'�z�)�+�7���bw��-B`@P�'$r��t`���	�FU3�B�'�`�����=<J�*V.,���'����|�Τ�� 34 "�'>�pPTYE�"=C6��\Ӷ���'޴ 'c
Z�(ǃ�+NM���'�4E�l�;?��
�:���@�'o<˶K�mb����F� �����'K��� cB�0��в[&�
�'��]��D�<��%���+C�]��'���R���D����� xPq�'� �a�.��8M�s�f~1��'��-qR�յ5K �i`�Z%7���
�'�쌊m΂!װ�HP��u����' (`���"txwAya�dX�'��Ųa��� ���E�z^��b
�'b���(	����8׏Юz� A�'K�u�g�K��3/�=n���j�'�ld�6���gP��xR��d�؄{
�'�D@���)*>�y��U�c_P���'VMz�bYը��K�Q�rl+�'����U�G�q���M�Dqz	�'锰K��2�1�I]�ڐ3	�'��@�,��B��#��
C8�	�'����3�P�A<�J��Q_f���'�z�bV"M6Y�mIeK�3w
5��'�@H����?�H�Ӥ�c(��r�'���f�ߌra���"h�+S݀ ��'>�Y
�+���Ҽ��`�W�xQ��':����:0Y�F���P� �'�F@��mF|Ic.|)6�@�'N �j��P�L�\��(����e�
�'46(jCK3)ԑ���$d(�)�	�'������w,0���S�U�=x�'��u����^��5�$d�N���0�'�1Zu��9Y��]�t�u*.$�'��pB���	}#h(�E!�w����'j��d+TbŰ�I�4"i�݋�'$�!�U�T
�hV��p0^ ��'�6u���Ѯp�T���؈k�s�'Ғi��"�bW��/!��vC�n�<��DL�O�5�C/�[@q����n�<	d��u{ �f��@T�W�H�!��M0cs���Q�Q"D|Q��Ž�!�D�$l�r�@����|_�ݘa#�X�!�ĉ_^�8R���TJ.�rq�I�K2!�d_�g�&� �G5Ld�s a��!�D��Ld��0��fT��5�G�"@!�$M��V�(=��`��fƲFl���l���瘆��mK�o�<G�	��|�H#c�$�t\�pF_�nø��ȓp>	�e��l�Es�B�h���ȓm(h��R�8��c�S�\m�ȓ9�p��A��%E�X��,�.x��_����q>F��!���Y� ���S�? �M����Xw0��r*��5��s�"O��*�ȅ�!��U�3ߞ$�w"OzR�.�-<�^�#HȈi�!�s"O����
�;#ځ0��7h��!"O.}��C�}8l8�����C�ؘ�"O�y��R�k�4
�@�-�Z1��"O��!e�ā7"`#������%��"O�yC瑷4B4	���z��W"O^�Q3�B�!�R�A�f��Z��)��"O�Ġ�N�:�z��* Np�c"O��zĀ�0�0S��|�F�s�"O@�U�B�j��i��������"O^��t��?^�A�Ac�2\60Z�"O� ��CX� $ ��g��#��$h�"O�} ��=���"��ǧ9��B"O�4P�*ܜ�Dy� �Y���I�"O 5��ڔ0��es�$��x����"O��� ��������71���"O,{6�ґ|ѐM����%�5�*O��d��E�h��U*��
�'���E��x2C`'a�X��'�fPX&��7����
�v�D��'2�%���U_A�UZr��<^����'�h(�B�D�a@���	6S�tH�'ּ��fHޜ$�!oR�R\.�`�'ن$�3�&ax�JQNȅ��c
�'_t��t/� ��)�@��P�4t��'mn�84O�kO��h��@�VT:��
�'<`l�"���W�PH(�̓G(� H�'D>� ��˖i��y˱��B��M��'�Ds뒊r��[�"��>v���'$��p&-҃OS�E���G��I��'�aB��
H�`g�&Jm҈��'�,���%*V���]�$���'^$�â&@�?�D@R�ٶ+��'�P��T#�@ ǎ�,}���'��ܘj6n�X0ʶd�(w~���'ܲ=�Â�2���
Do)f���'��HVeȇ52p3*��1L���'gjI�T`Ó8�6�1�%�G��r	�'.l-i ���_��!�G�Ǡ�&��'w����\�d�ȼb�M��6\2�'0|�'� ���(���,��A��'��=(���	'�v��[��@9
�'����A��5`P�bN��y�ꇣOYXt(b�9-&�Ue�v�<���ۖ!�Vl����c	�͊�&�f�<���X�A���a@�
oT�:2��c�<����2=�AI7.�B��ݓ�_E�<i��61��@�0�t�g�h�<!`�-�N���/�2����g�<9 ��&q���g��)i�p��Qm�<ᒉ�(PT���\��)#��Fi�<��ጦBy�`)��hZ���d�<��%�h��A�W#���"���^�<�)-$9���'�R� 㰅�bEAP�<1 �
X��#Cl�iw� ��f�K�<��J�:嚔J炈 F��q��R\�<Y�%ƺ	-�e[���@�����%�}�<���>��ʳBE�^�hy�T�Gw�<�c'=@�!pi�ADĵ9V�K�<����'J�\,qBΗ?� Y	�fU�<FڤB󶰺uD�(OƶUI�Fw�<ɄkS�-�h�!��; �����~�<� �҈���p�C-�3p�pP"OAa���" �]3gA�o^8��"OF�rk\�-$ްCvB��v�H,�G"O��%a��q@������y@`�# "O�л1NI!@����"`#Z","O�,�!��E�všF�3r�Ч"O��C�i���ġ[�#F's��e"O�XQ�B,vn)e��o���e"O�@2�ՀL�|=���ϡZ�c0"Oq�$��;�J�{	ׇ���"O�h)��Dg�fȖ#Y��X� "O")��T)�uG	뺵ڃ"O^2�\���G�R�v����6"OP��S�܄c��&�&o���AC"O�	�vk^�R����U��g`e0�"Oة��0g��9y���WϦ�#$"O��ʆn��\SD@\166�BSH�<Yr���հ .
�H�A��nRy�<р��E�d}@� ]�b>duIt��q�<Ŏ��a�^�ҋ��OOr�C6�k�<`���
$$W�E��ɐd�B�<YS�D�9V�d���ÝO�2<j��=D���W*�KHA��Lc�@��<D�����v������H~ԅl>D��rN�1�3-��&����K�3�yb�<l@��!��r�	��ߝ�y�W����Zu�P��+�;�yR뉅Dpd���ʿd_~8����9�y�+ �ynm	��?d"=w���y���7|��]1C U�Y�x�`fCB�yR��o�|u�DjU�Iji{��Ψ�yR��F�"�(q�I@j�Q6��+�y"�Ծ�P쁲��/=�t� ���y�Āts���7јFT���>�y2-݌V]�����B�M��3�j
��yR�O0�麐�H��X�X��y���s:�Թ�D\���آ���y"�Y=ib�5��[{���{�A���yb�A&���dE�n1��bGo+�y�CW�Pl*���*b�f��cЩ�y�Q67BH�FbT[gh4Ӡ��y��u��"�.R���0D'�y�gO�PB���d��H`�����Y��y2�U*�ذ�QnV���M��y�e�`U������b#A��y�+F��AJ�d0���)�e��yrO�>T��
�.K�i*H���A��y�c��&8�ۇ)�gTZ�֊���ybn�#7q�=P�0�ʨ�	G!�y�`C44�0�&�O�"i��Y����y��M����W�1��,���J��y"$M�r��/uqX� `�*����0��e��J�%a��w�� ��	^�� ��P�P���"ԒM�z܇�KD|Yj7oR$1������Z¼!��=� ����KcP�#e%܊l�T��ȓ-�0���h=;���c6�
��ȓZ�Z�Y��1O��yT�K��e�ȓvE�U��KE�k>�Yi5�-qp��*a��	p��/v:ِ��(o��	��Vʚ��a�J��x,��	B�1�لȓ1����#��-;�
P�0͛�TD�نȓ� r!�0O�J�Ûr-����.��9� �ވ=���j��*͆�S�? h�9uf�� ������F�Q��"O^Es��i��ѻbU�d.�ˢ"O��5�ޑV�l�h�'T-R�\Q�"O�Qt��!q%,dI��w�4I"OVD	�f"i��6�º(��i�"O���FX6���C�5H���"O�P�f��3M��X��ׅI2�r"O���1nkR�����)u.����"O�;`(4&����qOU�&��\��"O��������y�  �ixVl��"OX��B�fZ�I��-Jv�!I@"O��!'	�,w`,�Ӎ]/'j�lq2"OxX 	�.; ��ծ	�wa���"O(�`��(<U\I�-��S,�"O4�	4OV�<���陆5Į�Y�"O$PSeBÛT����9l���F��P�<9�ď({�hcT����@��v�<ɓ�Ƣ,|a���#|�ĨP���s�<�gF�<��u���$8����r�<I�!�|_�e
6�
� �lrҧ�p�<I!��AL(-ۓ#��G��c�n�<QՅ"*���7�IS�&�f�<!���*��A��K\���PĘb�<���
0n���vH��L�Kv�^�<I��G��d�9�F�F�j�+��[�<iW�5��2��'�x ����X�<1 ��Y����B�S6C�4��7�W�<��űz�D�K��@-j�"��d�RV�<�1�B�9�|�aDC�>G��r���I�<���e池�@\	3,6풵�]H�<��V�R������- �:���e}�<��'�=;��*��L �؉�H_d�<��HH�+�vu�,[~Y�Zc�<�� R�%Qs,�~�:yâ��H�<b���$j(ҳp8�h��_G�<�A�@�V��V�ЧZ��8�e�Y�<�Ù4h�L�����3�v%�3�T�<��
0v� �fýAmF ����y�<q��5
��Y��O�W&�:@Hq�<y5ᜲ{���%Í�4��)3�Ru�<q�g�E�<�!K
�t �@�o�<ٰ�h���5I�>�&'�l�<q���68	t�"�����5�q�<��mU\�r���B&
�8�9���d�<���P�~�J�y�J$y��SL�a�<yM�0�괫�3�Y4C�D�<Q �=Y���j���[^!��{�<�pD�xO�)A�V�#���T��x�<��%H�{qX���@n�F$Ғ��l�<�R�S1K�4񃵀Y�h:����f�n�<qVL���8eP��^B��IW�s�<���*6�@��3CЕ|KX}2��u�<Y��C�h��i+P�K8x^Q�欖I�<��d�7eu��@A��1B�M���\�<Y���;(X-J���H�nLQ�Kn�<y �׸�~}2����&�V�c��h�<����m�(1��)=����d�b�<�F�ޚ���AG��$Ɔ�x#@@G�<�O�2hؔ`Ѣ 8����YK�<�CI�R�� c��2Qy8Ո�^\�<1���'_��)��NÆ	�\ �JU�<1Ǧ�=F��R�T!`@� �x�<�&N��lxq �>N�F(���w�<q���czy���](�أSi�s�<� AT�F
�*��2�� ,���S"O��bcA,�i�5&�A�"�j�"O��`DiW%Y�����'�<�`�"O6�˥P�On8���Ў2� ��""Oҕ����^�`!�2"L4B�p੕"O(%��ӿY���J�%���"O`�S����/����1�
��y��75F��pƄM��jɯ�y��M�+r��/J��L(#��y���)I���A�!
�  xg�F��yRa�.~3޸�I� �6�����y'H�@�X̨P���J�@l��#��y*ܩr�<ؑ #?��L�PNʄ�y��jlT�	+�:�5sS+���yb��>�n�QRm%�X�!�>�yR
W�t,�i�hg^��&[��y��V�*0���oپb��i0 �*�yb��%i�8�%.��xh����y�'�
$�(�
#���",�����T�y����ԑBa%"��A�W�
��ybd�	��e��J5.�Vq�V��y���* �0�*�'���b��=�y�N/8\\�`ȁ�l��&�ʹ�yr�5#�(Pk%�"D�@���y��w�H��G,F�"�2Ż�M:�y�K�݅I'�p�I�Hӡp�y	�'ƪ�8�ɓlk�-�Dȃg]!;�'� ���ڵ&� I!#�L*H�0�	�'1�A��*B���KV&<��	�'����Um�}�&��!/��u
�'�re�E=��tS���t�`
�'�D�3w$��:���R@����'Bb��JJ,c^�mh�N/�h3�'�|� ��֞T��SFΒ'?��!��'��gMѠ\Sz�����5���#�'��;�� u	�HT�&�����'�\��4(kz� ���"^�j�'s�%;��ɪu{�	�@k�&�%��'�-(�E�������!_5^<��'C��jT9DB�c�
�w���	�'�ڕ�ԅ	Fv���+ޟt~*h1	�'Ԇa�"N������&<Y����'���3���0څ0� j�$h�'�@MCVe��p�@�� ^�4iR
�'�|Q ��q���]�e�	�'
���c��%ZYQ�b�U�v$�'�xy[�	90������ޅ_��$;�'p,q)4l�2w�6TpPK�g۾1�'{��sC�z���35#V�]ʼ�	�'��ҮH�8�j����S _��0	�'����,6���w)�\X-��'�J�[ǈC=2t�i;!���H�Qh�'HI�L gz�K1������'��'�IND���3JAR�'����3�آu�>MX�CX�����'Ū(2���tņ r2`�3jƒ0��'K��ڐh�$��K�.�"%x
�'��ݺ�
*D�ax�.�<#, $�	�'2D=�#�S�����2�D��'�Ћ�UKr]X�%8�Y�	�'8~8�u.Z�L�:s+�)�b���'�����U�U玥afȌ"� )�'�v<�ƅ��0�TlT�d,�D�
�'D�ԧ��a��ʤ�	%�f�3
��� �< �b W���s�E$��"OެpAi�c��1��<w7Ę �"O��Di��&D4����.~(lDq�"O�#�ċ� &�qBam!Z���"OЅ�@��"���`��
���C"O��3&E�,3��%�WG22�{"OJ���8A�~���_j)��"O���JݠZY��q���V(HuH�"Op0�I]���t8�i J$�`"O����ju4p���#���"O�U3V�5C��)���,
ș�W"O�!Җ�Ϙ<>>a�� ң(x4`2"O<)ؗ�����Ć]	��*F"O�Ӂ�!{��	@��:��@�	�'*p���ȿ�v)���G~Q�
�'1+�[paZ���z�\x�m#D�`��)K�`�1�G�Q0}G�\a'7D��2D$Hr��9���
���eC��y�07_�,�*�6����%�'�y��՟+��3r��.@$iq��D�y§֖j䄅�  �x����y$ٚ- ��15KL��Y�6̜�y"ő+C�H§F�,�F��=�yR�2��|bR�_0?f��Pm���yb �0|���?���Q`R%�yҁ�$;�
 �Y:�!
�I׃�y����Ƶ�r�_$5Oz��@��y ��(=8ǘR(ڇ����yR$�,��20j���F�M,�yRlߗw��(�I|	�Q�U��'�y�k�)������{�����η�y�c�����eD�y��--	�����U0�1��R;��3��?Npp��ȓ�����k;	lI�C��L9��U�P���nN�|��$�����b^���ȓ-�,���
u�V�>Oļ�ȓU}̭є+�j����+5eV���|����@>�P`���3c,H��U� e�0 Ǎ15��o�Gf���ȓQ�U�"���x��Q�ߊWS�d�ȓ$�,��!)�J�����m^�5���4q�R�.:rm�d�		oD�ȓ��5�����!�����[�#tЅ�,
�L�'mN(e��X4�TPa�݅ȓ_��Ā�ۍ4�D�	s�[� ͅȓq����ئZެm��܀k�0�ȓl����ï��) C��Y.,�ȓ8tl����	P�=�t皌>��Y���$I�F=n�����bM)��;0�(�A̖��>,�A�15n,��Wژ�/�v�x��&�-eέ�ȓr,��"3�y$ A���O&=�X�����́����1)�M���	p�`�ȓ7�(�V8���>�"\�ȓ/^�����/-�6�h��ȼ�,P��]�p���R�-7hh(��<?�n�<Q�FN���m:��I)pІx�S�x�<���4�s"�4�|��&E^�Hh�C�	�%�F����1|r��&�ܜ��C�I�{����.B.Ifo�;9�C�I1VV�����Ҙt����wɬC�	�V��d	<������B�?��C�I�,�nl��.ۛ3��5�4b�;x��B�I����A(�?#�!`�b�r?�B�)� �	��I�.#7�%��^��uXu"O�YPA],;!���؈4�~�s�"OL��AӀ7`��
 '��J�P��G"O�0���Y+d���m�(Hр���"O�)A� [��r�,^Uݾ�!"O�uR�U�a�
������a"O����+�v�d�V�\����%"O� � O1��ʃL�bBU�1"O`����=Z8Z�۴�Q�u񼱙&"OB cK�n�`�(D�2K�25�"O.�Crb�����Ba�-o��tS�"O���K���rP��\�bAf�Z�"O�M83I�&`y��ܞ$,����"O�	X K�<L1jBn�]&��"Ol=�Aᚊ,�F���mB�ZX��"O.e�H3 .�q�"�,u
�"O&��tt�̠uN��\Lr�����y�m	u���`O��j��%�AbE��y�g��OQ�����P�Zf@�Z� ��yR�/� )S׍�!IQ�%yU��?�y�e�/-J.���&�F��X���ޖ�yFY4��1!ϊD�#��y�g�j��	�$ ΁e�j�xF�)�y��W;1ld2d�Z�^h�u&Ŧ�y"�[�LTp�!�*VԪ�R��&�yB�T��
3Q���KUh�03�xJ�'F�Θ�i,���1"�#D�l��'���j�흕e>@�h&��#�N���'Ҏm�l�`�����(�Z�a�'�H 0��?���㒇T��u��'|���%�V4E��8���R�pX�'ؔ�+p-^9g�)��Μ�]��,R�'	J�I �R����S�YY����'��|[��%���˒�R�LF���'�@�(P#!`h��g�K""9*�'�����&	e��#����p���Y�'�4�l�Hn�����YyҸ��i,4iU*�?�� YF�ϰ�ޭ��!�8|�S��| �XJ̳{�j���b����3QjZ
*׆);z�p�ȓ"4��4!��|��}z���$;�n��ȓU8Hx�6
�+H:�9ʲˉ��^d�ȓe��сU���
����*B�`�ȓ@�&Yx��(I_�1�#ϣx.�(���`�R�U;�*|�ת��o�z���~:��dC�aɴ�4��d�2`��q�(r����JP���ԌD��tn�%�!��&!  �Oϯz�~�ȓ\�~q���u@2l���(3Dɇ�v	��V�ӌ2mR2�(ݚ�� ��I�Q��6Z�z�1㓖ss衅ȓS�HaCB.T,�N�١g[j�����'9��s�['%�!!�՝(U���ȓ�8�C2�	�m�(��0����ȓ.4|��ޗk�� Z��0�a��Db��a�M	������C�;���ȓ|R̠S�5 ����_�T���%xL��	�.ά�[��;Y��E��m�|�r]�*�����4]�؄ȓL�S� ǏK4 P��ظv��Ąȓ��<4�W�Y�n��3K�$6�l��5��`�Q'>r�k�ڍ@c���ȓ�@sR��Y��}���
����ȓf���Ȓ`�j���4.��i��y��S�? �8�V�P�(��EX��E"O��w�Q-z�d�4��7��@"O�Ls� ��JW*�מ�@�"O����1Ҭ�Y�	�1�HiYP"O�=(R_�Z)B�9�  8�"O4d�@\HL�#&64��� "O�I�"F )���"&��!T,B��"O���CAʟX쎵��Z��~�[�"Oܝ�3 �kYnP"S��g�����"O�����jDM�,K� �R	x�"O�e�ܰ� ��N�x��"Op8�5L�=\����w ď0�H��"O�(R`��^�M�=d��0K�����I�(h����'C�|�v^6*`�B�I�v���,6:P��ɥL�2
�B�ɻ��\��B71�J%��c[3u��B�32l ���>b���b�M���'�ў�?a��N��x{�0�E�P�!�Έ�;D�0qsN�yd��BC��3�Z�p�bc��=E���&��,@ Z(։�a��!��C�	ɦ�PӨ8h�\LҬ?��Q��;D���
�G�m�g���z�j��8lOh��qd@ǜ6��h� ��LH��5D� �U�[%�^�(0nW�Q.����4?�
�{�N����I&��t	�8`
�t��@}B)[tI H������hڴ%�ȓW�28@�*m�-��B�p�r���Ϯ$b��Sd"<�X��]2d�왆�D)H��_# ��8@l��^�z\FzB�~��B؍o��3�!Ło"�-�j�m�<����h��'k�kdZ�F&Q�<��"�������; ��P�<�`�^��B�b�phS��ZP�<��!�S�����t�@P�GEҟnZn���O�x��'St�WIS�� e3�M�[	Vq�O6����(_Ŵ���VK3� �RK9P���4�O�S7�ܻG�9�b���Q�"Or{�c�#e�&��o��x��}"C��!lO�ʲφ�TJ���д]ɴ�Ya�>�����(v鮕س!I�dBSk�9�	Q��H�,�����S6��ƙ�O�A�"OLM�!	 Z۲���EeG�%��"O�h׏�>yrL�����K2`P���Ij���IO�J�f��I�0
�тHj��xr�	�p�1��eU%���,�&C䉗3���� ˧I8(��c��<�H#<q���?)����!*��т��N�r� �wM4D���̗�v�~��a@{V��Ƈ�O�7-8�S�d�$��T�^i��5`'�1v!򤒅V���G��<6���O���v����՛����h)��C�ˤB(�3"O�DF�٢�`y������4��'�'p�)��xBiW�7���(���T��4���x��'����b͆�����2]�	�(:D��X����5ĺi� �.=��[D�9�	w��r�'>i:��	]=��A�b�03:�m��'
��2�%�!��A�.>\)��ēI<k���WW���L9,��Ey��!��+�<��-^��"���%G�B�
&h��Ε����f��^U����Y=��DeӦ	j#F�~颔Yb���PxI�A"O�X�!�E���{��%
pj��'��'u�̛3	�i���H3�B�����O������Qr\�2���y� a�b�R.!�� 6�qAĕn�p#1
ۂnMnc"O����-?<lP�ToX�4xb%"O.��6d�1M�2�H��0�b"O���4��b�� F���"O�L�@��yP�#C��,_��u3%"OR�!/�%O}T�����p�P"Op�� �ܕpȬ���V����"O`�+V H�f1LҲIXG�n1�B"OX�C�I��9hnП+�>H0P��F{��	ѿH�0-
SE�Nx:�2�K��J�!�$�R�h��� M�e��4X�H*k�!��#
����.�΁��j��!���m�T�2�"�"g{�$�����M�!�Ĉ�(,Ѕ��M�h���ƌQN!�V	<�PЕ�O�I}l�����g��y��I��ѻ�DS m� *�3:C��
[��qA�P�@�.f�fC�I�fs���Ï�c�Dy�N�A4C��!gB� ��6/~��2C�� (�&���	/`��h��ȟ#���$ �e�bC�%-� @��?M����s#��VHB��,|�,�� �܅<XTC�ᇛOp@B�	�)#���ȉ,��uSCe۟dv8B�#5:&�he�
?ҹI��רq0B�ɸ)�aJw�A�'���kpHVu.B��!P���%	�P�	0�l%-B��!jKj�cqǃ99Ŋ�wi�	����e��0��%qb�M��������fF1D��ӣg��d+n-��/	��`R(1D���2a�ߢ�
&��7-��dRgD-�D<�O���-�6}��ż@,���"O�}cs.�9�Ȝ �MF�MTL��"O���dбMM<��D����+��>�I>!�%(��?�)c�A�?���x��L���x5"D�lp&�ǚvE��ze���z���b-=��ȟJ���L�iP��3C��u 8a�""O؛Ąs�Lq9�a� 2�t�w"Oz�����TH�hj K��0.:�z��>�נ;�S�==�6�ʬyв���N>C��a!��.D��s+��M�� �
�0�Q*6��O���S���.Ay�AC�'V�{(>0����Q!���O�� �lй*琁;��Dm�d4b�xU��E{��� p�♯6�(��@�[�D}���'2�'�:�����#��A���>b.����O��Ez��iF-�t�b/��xbD��
�*�'�ўb?i�� sa�)V�ܗ>o�a���<!�B�6���c�63 HD�K�0��B8� �>q�o�`yF�Ȁ�ê%έ	���w��$�LZ�[���m� �+���el%D���0C��Z,	��# ���e�"�		����6��DoD�{NXIQ�-R.����Oz�=E��GE�  �x ��.�v�� C<��=�b�|bCG7-.9��@Be������~��)�'QΊh�
��7CTI���[==�8a%������� ���&,_6������P/d͆�>�,�3F6Nib��5b?:aF|2��-d��L�e���FlBT-W�+C�	5K��H���^�,d����]�6�	����,MAOQpp�P�R +�Nŀ�"OJ��JI<2(�H�3!�yn�Q�v"O̹��F�b�:*B/�q]�B�'���+9��y`�̞	V���"o1�!��:O�fġ���7;�~��	4�!�$Ӱ;�c3.�y�2��UG�z�Q���'4�>�  �QD����a�Ɋ6 t�� �d)lO�+�,͔r!l�q���i�Б� O(�d�g�ʸ�ub�/���b`kԶ\"!�D	�JN��R�)%��ԉG	T4I	1O���$�*^����r�Q�5	J@C�N�6U
!�$߁R-��P"
�*�)C��!���Vc�kB�O�w�l8j��6�!�dӊ|z���k�2�6����!�D]/?o�������<q{@C�q�!��Lje�=z��Fu`�*��ȸF�!�D�*$r"Yg�]�i��$�T��o�!�
�a����X�iB��!�Dɝ?�8�bDm�	�@:c�6W�!��>c+8�s�ʎ�G����� &j�!�β%��� L��i&* �!�$�Є�q(��5̢%Ѐ�Ջ�!�DP/o�I�+��z��FΖ�f�!�dD�F�Sm�,2��� %LQKm!�DF�K^���/�;4����!l�N8!�Q+�  ��'��2z�E�3�6),!�(yVM{��[� �\m��i�H;!�d��'�� :#$�3=hJ@��
	� �!���jL����U�J��l��z�!��?F��3�σu�B�'�8&�!�T(U� ��qB�3�V��4�P�a�!�ۂ���SѷX�h�@��v�!�$��M�)�k�9��x���G�/w!�$	�@L��`,���t�J�H!�DA�ր@Z�X0]ܢ�rt��'hj!���`",p�Qe��BM�&a!��_)Nd��Rr��1a�8��,b!��A�z���J�]`�#��� hR!�$P
�E(b$C�N]z�Y�M�\&!�D�6�v9R�	
�8@�9�T)ϓ"!�D�i."�8�^�#I��'��'?�!�D��3G��� nï$X��u �x�!��6�L]���+�	[�+�!�dK ��hRk�7U��,4��(3!�dC<nc
I�rh�(n!n�$ T,Ʉ�+�Tiʱ��52l�xH�S� ���G���V�
�B;I��
��h,�ȓ-�c��Q��0ˀ'�чȓ7:	`���v$���R�dN�	��#=*0w���K�<��.L:"�jD��~�$.D�a�Ѷm5:���&�8��c�}א�҃�Z(@�p�ȓ;��
t�9ؽ�2$O:3"���'
�����_�{���WB�h�ȓi	�\I�%�.�r<*AM�]��f ST���� ��D��I<`=���^�P���Æi-ZB�8gZ��S)۳$,�X�+ Q�B�ɥ4�`��U%ZA�X0��AiZnC�r���"�Yc�Ȼ�&�r�B�	(!8D!�B�J���*R( N�C���Zڂd�H(d-P�bU�C�	3���H�Ϟ*� /c��C��:���뀊	'�q7��#�jC�1L�N�X��GH
qh��]��C�I �(AQN4/�^0q�� GM2C�I*P(��y�lN:o=&�A����B䉂N�U�'�"0*�'*C�{�B䉸O��([!dY�b�DC��j��C�ɻNS�%Ï�z��Oڇh��B�I�0FH��(�p�(�"��:3�B�)� , jVoX�E������W<$[!"O~Pr kL�"� \;`n�6w@�B�"O���v�8D�T9�eC��n<Y: "O�)At�9=�%������ܪU"O(\�R#�-�4`��ɳG���r"O���D���⭊�%��@�"OR�[<Cht1��Մ*��D"Or��O���$4���
E�����"O@�5�S�c'L�J�(� Ӽ�"O��æ@9G�F�Yri˭���P"Of�2d��7m���C�A�Z�"O���Q�Ҍ1R�Ar�ZmC��0�"O�Q -]��t*��CR��"Ob��E"_���R$κ!!�e��"O.IB5EZ7>������U"�Ԃ��IZ�ZT��*
�o}"]��5E�\�0P�cI�e�.0�4��A�<iT�B� >�mY�N�l��[S�G�.���8�L���O2dF��O�}Y��&"����-ߝdː�r�"O��� Q'Goj,��b6D��1�%�I�Byj�&Ɠ}-nq[ʛZ�axC cs���oR�;�����0=�iz�V�b�#�4
	�T��l
:tB4l��U2�jG�G.Ov����]u\X`5LE�<���D]���&���$]�z���5U�^`�3��, J�O���1�уXو$J�m�Dڂ�h�'t���-Ʃ��=�Dj�uWX鉊y�tU\��=�|�&剷T��8MA
V���@�So�<!
��"�t!�A�6~���
JNU��h��dȵ6M�a�V+�=A��Éw!�T?`��U@��@n l)@�07L�[��֨_�I�a j��ɡ���G5y�x�R��F�:����-(��W�N)ۅ�s�����C���iC��T2\{��!g�.�O�]C�S8 k�L�����h�W�d��nm�p���t� 	<
1٨��йQ��<,2�k��^[Ԛ$q"OB�#��Œ5������ؖv��eX�Լ�^(Qs�O.N��uQ�K�w�D�+X�?���k�t9�L����Eb���T���S���{p�'�� #�)N<�KyӘ��'k�� �)*���_�65 ���~�t; ��OH�х�St��Dˁ��(O�}� �J�2�օ�š�B�R�k����0U�偧�%+7�扆	v []w}�m�P�I�=-J4AʑN�8y�jR 1̊P�s���@��D�'ۨE0v#,B�V<97��/[��1�-څ`0,�
œrW����*�"`���
�1av�|7����T��#������Y�>*$+e J������]>�M�T	
a�8y�0g��d���C�b5N��6-֧-�ܨqQ�~�F��i2��CY�?�(S$M p��̀;\�P�SD��o�]D}bဵ:�� ��EHD~�	o}ur�ɞ$�*,��ԡJ��ѥ0y��Ab�i~���)C��]?M�(Exb��(>:�����.o�1�m���~����c=eq�`~"�_�;��nKd
qoZ�*PH��3���w6��wN*m���".S9bM�!<~⢩��I#tݲBA�,��"
цPa\�\4���T#���8ڴ]����u�jЇSgP�P|4�Bv�Ք4P�s��!*���$�~	N��P
N>L�xaW��G~�tID4f����t�i��Z���)@(��ּi�<�';f�(�Xw�N����T��N@��ߑ|���R�	9����@7�/�����O^���.�+u2�����.o��3��4Z�֜j`C:�Z��H:1�.l�ol��᠎#�O���j��T�����AmR�6����<�q��l~R��(w,��ƵH����S�0��Y��L�c��8�D꘶j��%�^�����p>qV�ѥ��4R��jk�ɑ2]g�M21�i�(A`R�iv�Hs�П@q�R�%�� �;�y���
�^�D#hї�y���%,oHx��́�� �&�D��Y�f�%~��@AX� m��q��%���N �l���?���E:a�S�
4�YX��B���2������>=��:�酑3H��I�-ϩ\�i$�X,C�Z1K��
���Q�3�������[zj��;P4��1� 8zլ��08`t��nO��Ӷ�H:� H���Ta�!��"OHԨbǚ�ڤ��ŹTW�9�鄌/}�%ÀJ�<YU�p�6�}��yC�1PFy*���/�����b�<���B�o��)�����شط��<�foQ���'z���Q-6��l�FF�ti�1sg�],y4�|⬝�v��ɇ8a�L�##�,^�|	dZ:e-H6,�H�@�-b ���N�:n�^���9D�� ½SS,�?7�$x��oŪz�|<p�"O�R��\�9�����/��"O <1�d�9� =Bf���DtSS"O�E��֘b��0�ȁ$F�4q#"O��A�d%I�\4Kg��8�2��B"O���W�ӫM)��'��2F�N��w"OtQEd�:m������Y�P�5"O� ��Rq�dF�&%����C"O\m!G-˫� @�e���);T"O~y����u��B҄�.Ū�$"O�DDB~��r@�ǁ|�|8�"O�|a#��z���� =>���y�<��ǧ6��t@Å����*w��z�<1P�����Q�b�`�`�-y�<�H�n�A���
cjh���Fu�<�%)�<M�YRj�=��yq�dDh�<��^?b��ǚ��f��Nb�<)D�F9䲭�� �<5�(���d�<���8�8�Ă�
�2��"c�M�<Y4A	�3���He��?~X(���@�<�NO�cqN�����[�|M�"IUe�<Q��f+.i녩� \�B��W@J�<��	[�!;�����6z ��w,C�<�Sn#o@�D��kK3j��D�ҁ�C�<��(��b��`
� �N�E�z�<���;-��a���x���{�<�Q���ҧ�DU����&Au�<��Fp��u��*���Q�Nd�<i���2�~|z$�T�X-<|��Oi�<!��=�� ��e���\���gJ~�<eQ
{T.8����{ �q�Jw�<��Ш4�N4bA!F6	��-�Ԣm�<!��A�b@���-u:H����m�<�E�*$aV�K�����4@o�c�<ɡNk>V�Vi��F�[W��G�<����";�&=)�'Е[bT��i�[�<A�<h�����������S�<�Wt�B�p�Ѻ`��Q�QFO�<��$Ȏ�8�&�6B�d��'�g�<�����/c>�yrNQ0"|Ń��c�<)u�Zz��P�����^�<�V��g������O9W��y��.�L�<�T� #��-��@0|�P�Y��@�<�uhU���% �Q�M����J�D�<��땕A��� ��A�uAb���	�D�<�A�1xB����l�#M�¹��E�<�!�TCFҕ���oӪ�2�A�<�D旿h��p�dA� �(6B�<16"أZ¶scP-�,t���{�<���0t���2E�*y� #cmZ�<�u�%p>�뒧[�Y�B��NW�<�W� BB�e���T�(��E#'$�t�<���C2Obn}蓋�< GLmced�t�<aF�D-~]��J��&l��:��Lj�<��,H�B[�������jX��2�
I�<�Qd�26�(��SK��@�<Y'a��7G�5@��Ռq�seJ�|�<)�h6����N�:�RI�,z�<qbɃ3m��hР��5$h^ ;��Ku�<�L�H� c�ǆ3b��ʀn_d�<���H(z�)7��g|0�����d�<�秘1w���'-�'{�-���Ko�<YF�2_F���L�"�%K5.�B�I�0Y����b��-�����,�B�)� ̘	���t�D0X��Y��Ͳ"OҤP�
=jj�db���=^���d"O��g�2�<}ɗK���v�j!"O�41�傫|�a� D8����4"O0]�ׯV;W֦B`n`Zj��"O�	�Wb�p�����E_ⵘ�"O�=3����R}��铗9v`"G"O�B­����P��D�>(�4�g"O(��f�	|Wh`��(2�C�'�L�y���19�
���.x�<��'��M�uB�?^�X�s0��+�X�J�'��"��B�J�F�RǪ�7kS�u��'l����9$d��v%ǜm�h}B�'+��l� �I��A�^�j�X�'��h��t_8�qA�� R͜�k�'��P9gU�Rf��c�J�TBLyq�'�V�!��ԧfǔ��fn,A��1b�'�@��Kѻ^Y*�0g�b�x	�'�����O�'V��fڟ3�DA��'blH�m�5�b��؊Z��mS�'���装˒Up�x�Y!��h�'Y��a�
)<2�y����4|i�'F(�2��{.��Uu��]�	�'��Q�6�P�A�6�Q���h�,���'����ӈh�hpH�c�0E��'���!E�Q��y�!��f�����'
�A뷈�$���A-̖R�� ��'�ԽirM�09D=�֎@!����'�D��1�@L�$4���>BN���'dDA�ǆ�=��0'+:	$��'�8� ��=���t��)��QR�'�4	�� ��U���OR��p�'NZ�	Ğ�B	2�{��M7���8�'���9�&T#8(=���F�M�t�	�'9�I)&��,s;@U	��۵8��pr	�'ö����fWƴ��_�>7�< �'���9*ۨ\r@�(26��'�.Y�N��l"�� �ǃ^Ȉ���'O$@�a�0O�(��Gb�NB��ʓu��a���#x���ݥZ����ȓoI��e`�}��=��edф�_rBL�0D�g�T,qqÐfʶ�ȓQ��P)���mY��|�
i�ȓNy܅`�hg��������$z�t��A���ǃ��v���&���ȓ<fx�J�k��Q3�h�v.݌J-t��}��$R��P1�8ѡ"]�B��4S$�ᢁ���b��S��t�\`��#�2=ȡN�6j �p�NY>����6q��) �weʈ藇��-pЩ��G�ԡpׯN�EȰ�����Ҥ�ȓ*:��y�D��ɥ	�=��ȓ-�Vx▍�� ������H���:�nЅ�ַȸ�EE�;Ӻ��|螰XfkP
+B���
X�~9��s_�t�SE=����(޸n�>�ȓ ~���b#6&G�IZc�Z7#X����=B��CA�	�z$hߟ݆Ԅȓ5V����ˠdgV�2��ŖW�%�ȓg
��:$������aN�B� ��{�
D���CZ$�V� 9��ȓc�\��ĩ2a��0��ɞ�?�����$[���␢N)�e`��"ޭ��&�Bd�⇗�����!A|,d��S�? �4J��\�I�&@�vU��]c�"O��2�(̙[��ۇ�L=�ZD��"O�(t�P4�8ňD=KT�Ĺ�"O��B�Q�D�B`!�ꀱ^f��bT"Ox���Ι�1 �ػ�ʃ53Q�9 �"O�9����	d8�
�7J�A�f"Ox��P�8�yu���$Q�M�"O�h���˘�-{���TJ:�"O!�q��9Kx:�i�7��@��"OB��o�L�6�H��5H�*�a�"Oj!J#�W�Y&0�S�����@9�*O��ys�t|�� U�\�yb�̫X�L�_(�R����9�ʓk�^lFNI
m�FUDjӝ�4��K��t�M��(H�]9���'��]��<F�\;��]�nW�D����H��	.j  �cʵ
�����>�B���� �za�&b:<#AI�?���uxp�ō�]�l��dEX�i^q���$xō��o�Ƭ�� �Q��M��6��q���{��}R���e�n9�ȓG!��jgaU4%�i�Մ�|��)��@i����Y�<#�"D��Y�ȓn�Xѕ�\�P�����vP�ȓ�Fԁv	�v��%�S���{�x��ȓ-�vɻB@]�X��q�$����ȓ^�ڕB��T�[]�<r4�Uת�ȓ4/*�JTlm�V�A0�Z�Cr���fhTiҢM_�)X���%��xd1��C!&�a��>���'��2�=��@b�l ��I��e��@�f�������glȍM�X(�s��<ZT �ȓ�A'.��=�X���Ǒ~����]�`����D ��
Tڱ7&�Ȅȓ	��ɖ��H>��6i�2]�<Ԅ�3#���0���{�����k�>!��k+���lK**-��sC҆A�܄�q�`�h���H(D�ط�������ȓR8T��
�3����FR�fŅȓ@]]�SCBKF0�Q���Z�х�H%�2W��8p�L���%�|ȇȓfs�t�F�[6F�p$,�'_����(T�]ꃧܔ6���/�>���/D��Q�K��x2!c=R�ސ(T#&D�)`����u�u�� G*����$D�����#v$�i��rk��#D�����7T�����ǉ{-�X[Te?D��� �f(\����
W���"(D�y ��/����o�OG�(Y5�=D�Ȋ��ިNu܌ p�l�fـ�N8D��E�b�b%^#/vٹ�m*D��Y�-S���ڱ��YXy�6�<D��@ �ل5{�ض�ے�"r��:D�xP�2@`.��	����2�6D��0]u]0M�g [�>g �"'�Ң�yB
�H�i!"L]�-v%y���y��:�$ a���~a�qA��?�yȇs���"`%�*\Q�&	��y��F#ι0@k��Ⱥ�L��y��V&a˪�9F�K�Z�������y2���l6�d��`�?!�ej�,��y���*xWx�y#��2A�(+���y���B@��)��xZ��@f*��yҌ�4'PY��/=uH�Y�Lء�y
� B!借Ha��7m]�X�"O�di��;j96	�lV�P��D��"O�a�C��Xz|���@ �����"O�P��m!w��MB�)Q;P!�A�s"O�a���?L3$aj��I�z/Z���"O����H�۬Q$�1;-�s"O�(����)]A��	7=�q"O2���d��l�wIEA�s�"O�H0$"H������@-vf�d١"O�82W��9v��A�ʖ!_���W"Oh��A�[(-�P@3�5$FĔ "O���dO�B�����g����"O�!� ҙ%
���Ș�~���#"OL5�6�>g�2a��n�h1�"O��y�ѻpE:�C �N	����"O:�[A*X�a>6���9��y'"O`�KE��<��vF�:	z=��"O�� @<�Q�
&d��V"O���"�G�-�=�4d��z� 1��"Oh4Z6 ��;~eyg�S�{d����"O|�#4��o�
U�R���d�	P"O^qC�۝F�\mh򡓌z@�q��"Ox%2�f�0=Px(��Qb]�"O�����ޗa��q`�L&LLe"O̹C�={�נL b�J��g"O��'M� UPW�o�ȥs�"O�$���X!G�����h�:�0}�*O�Y�Cけh9R���/�1gج
�',LD�dO^)~�r���a��O�,4�'�4�CK	�!�^�sa�=����'P<�����k9��EȖ�t �	�'�@���n�6U�*���cG�f8�	�'��c��.'i�%����|�'��Ր"I����#,V��	K�'�8MSJ��	Y�Q*E"�pV�d��'E�L�"���H��(��n��o�@{�'m^%:3AՏ{0�;s�I�_10���' &���A�N� �����<$�0I�'�0�əH%v���҃1İ0�'�>�jv��:5�fy�R��5�8�!	�'�t0	�&��
�q ��8�EK�'%cP����I���E%Z��'��#�N�4�Ba�$�f�B�'�~�P3��y��a9�*ε.⹢
�'��r`�02�01%����p��
�'���$B�d���
5���	�'�v�����q���7�S103��*	�'Dh�S��H"�!ۡ:QR`*	�'�����3�"�:��ټB2���'fP�ԢW;G�����$׽,��	�'m ���C
j$�d�W�>娑y�'1�aʲ)9rPp��W��n��Eh�'c�9p��n�
���(ZB��'~�CVM��e( A��8=Hhi{�'�0�t��Z�2�U"G�$}��'�D���Y�r�j���-
V�-h�'���a����XP�݀B4Z�
�'��y�7���C$G�:)�.�	�'Er�� �LV�$��'�ּ�'v��a��Um��3e�ΛK����'�d��eҰJ�����K%9hN���'%�� �(�t��xAt�R�:^���'��U ��Iq �:��_0m0�I�'�+5a�2n�B��$�L���� ��s#�
`X��iŃI�>�0�"OȨP@�r��$آ�_8���Q"O��Z@ݝ{ް��K�gv��Õ"O`y���R
�@�*
�g�(�"c"O��{�%
�d���7%|\m��"O �P�&�pL�5�Q!pZ�9��"OL0"�ŋ&k�(1I� C8i��"O�mڕK�iN�r��W�~�I�"ON̪���/�	���ׂ-�L��"OP��ĉ��49��U,�)d"O,�E�N�xVFu���.i�x�R�"O���K1i9(� l�.�<��"O6h���<	�K�3/@U"OfYY���B��MҢG@ b�ȶ"O2=����*v \PHdf�k"R'"OVm0�F�'(Y6�I�.)4�[7"O���r�*!L�ñ{��j"*OF��a�\+�	+��=V��a
�'�*I�j�1�XX��ȎA��E�	�'Xf���ϗ
}���G�t��z�'H�|p$ϟr'�RWC
N���'��\ v���)�bѺxF�	�'���a��	qr��qw���'m���2
�|>25A����^�n	�'�����AXA��qS&��7Sj�$ �'����4�-4અ�$��[dz���'����-ޭ�e�d�PJ��3
�'-�@PSf�&�����Ŵ4�dJ	�'�ʳ�E��ą�=H��'Rƨ��bH�p0T��,��H��'Zhh�i�PNv�2�D�	SF�mJ�'&��#@��P��b�D�TL��0�'B����J�$7�e*7oK4Wɐi	�'�:����;L��f��g��Ek�'��Hcv�E�
dr��G8 <c�'_)@rH��.���$h
44�*��'v�(G(HeK>LbD��#O\�z�'������!�i!C��Q�
�'���!ႌ2����B��?B!X�'%��X�/X�þ�hR+_� �,��
�'r �kea�/D�t�iܚ4*T�
�'d�e�檍;|������!;2r��'u��H"AS*B
䐣�
�?ʒa�'j� KPޅl�@���K:3�q�
�'���Q��+ �5�EOQ� �vŀ	�'A���W�Pq eϹ`�b}a	�'U:t
����JO�3�B�d�\���'+�UVKɦf��D�Y_�,�{�':���tȜ)v[ܠ"TJ�F=�p{�'��Q�`� C�!��p�'���#��u,^y�uңsD]��'N�V�L�
��)됪HR�'z�yzFg���T`���}g����'id�إ�Z#k�8�(5-�2l�p���'���1�3�zh�с/p�jP��'uv,B��Yg"�2���d�T@��'ٰ�x0���O8zSҪ�_p�-�u�ڌ ���tC��"��t���"\֮� �h�H6f=#2:O��C�:��%ʟ��t�7�ԗw��9T��[���y��|NyqaG(����J�#1V�ؐ���T���iZ����)�'"ݬ@�@d�i�01�� �%7���oڕhQ�"2�` ��b����#��ēR�`�'��\}ʊ��4�'R4��
�5L�Oԣ=����(3�G�*�d�XA�Ř>Ô�yp�|R�)�ө�NMr1�S���9n��"��hO�T�?� �y�&�"~�-��bX������'j�#=E�$F�;��� ��O%�Z$�¡��Em��Fy��)��"�6�Jqٶ"A*�x�$���%_��ӧ�7F�xK��x2�ǡ_�`ʐȤ��8�0|�
�E>"�;ԍ���R�B��Z���'(\� �|h6.�r���ز��'��p(t�x�E�OXe�=�~���I�b��a-�3ú�R4�C/�O�|��' �x���"<P�
�Jwb�&(�|h�>�)*�S�,C������	��*��Q�SȄO&-Fz��4���r}tiA��46���S��3��dKZ��(�b�X%��R�P��$ŝ�Tl|����'�ў�~�q�V7J`�a��;x��M�Tn�'�a����!7���圴k�<T´k�3��'�t#=�����I٤��x�mA�2��c$�x" �B���Oy��86������aѮD9��ʬO�@����i&<�`K��>����0N$@�6�A�#�T�«���E
H��T;@����+=|9F�ƭZ��x
/��6��"�jذEk���E����i�	��H[�i�Xx��)F�-(!�D��,3D=�w!�/kA�M D��}�!��X�]Xv����T�c���!�ę����g[+6�9���
�
�!�$�=e�a@��+P��0*�`��!����e�-��� Q��+�!�E����qN�5 �Z�CY�=u!��{�Xk�kQ�w*M�Ee�H!���*`a|A:�F��q�E�\:A�!���%+g% s������}�!�[� ���]/4�ŲT/S1Kn!�䒯M��0`�b���zeq��yW!�$�,*�$(
�ݜ]��Q��j��%9!��N�g;:��w�B;y��%�W�=%!�D�f�r z�hT=G��I�(
�m!!�Ė=�����#
R'���f�W!�C�D�n �!e�7;�� ����<l�!��mX|a v�F��D��*��	�!�X�A�0�I��l����g
�8�!�|���s%Ȥ}�X��gj�=�!��\y����-ħ/�N���鈭SE!��)i���#/Q�L�4����S!��80@h Ƙ4L� �����?/!�$��#�`�S��&q��+FÏ"d�!��|����NX�}e�ɂ'��0�!򤊸q|�P��U52\�)21�ѥ@�!�$W4M��a@��4YxD�I�,��+v!�Dn>���v���ek�	aA��u:!�$_�d�rѩC%_Z�<�A���Py�L	f@e��.���`C˃��y�Ƨr��ےKI�q�t����y"Cؘv� )-�l�
�['���y"
T�bv���#Q��pG"���y�N�$+����G��  [�HѦ�0�y�'S,-��p�n^=�P=�0�;�y�Ê.\��5��睶*�B�WN��y��e��l�� �.Oy8�C��y"���|��Kuc��XP��cIY0�y �f��l��5e�m	v�H�yBÑ�W���x�k��� /�p�A"OV���Ȅ۲���*֪X\��`�"OH$hS��:g��͊�O?�D��C"O���f�,2��*NT���$Q"O�����l;v� Sg�#p�t�7"O2��#�,H��9�p��+_��$8�"O�Maej�&�qѤ���.���"O� ��%���#�h~^��T"O� Ly��H�O*�!�Ť^$��C"O����$yŃ�1$J�4��"O$�P,X=��C�ɮA"b�q"Op8Q��t�t�j�c{k�i�t"O����)W �Nh"�`¿B�Ve	�"O�)�Jʠ�R�Ư�);��hIq"OX�¶���L�sq�I(j{��;�"O�$cvCس;�R�Bn�\h�5rq"O���e��bP�bΟ��fqBr"O�aơNY���8v
�x�銐"O  1��\i0�[�gS�4��C�"Oj��dHҠ"�\�-91y"��"O����^���{���c�`�%"O*���Ϧ-�`{D�T�9���w"O��
�넝e��ta�*'�Э)"O��E�%`8�غQ -z��OL�<	� �F6�5�pIʺcf���*�M�<��'Oކ<뱨�+<x읓�cPI�<7J�"3�}�������㧉�H�<Q0���B���-ю(+q����_�<)S�/bC����GB�b��&�\�<���+.P�y!��U'*�Yw�Xl�<�V��_T����j"u�$�j�<A��Q(O��0	Ε�-#4ȳ��m�<�����"�l�§O�1�J�����t��Pg@@-~ڙ� ��6? r��,�d�
���z�\��`��f��E������#5�b�2p�"C���ȓv�8�"hܧZ�0Ղf�U
�)��:��23�X�U0)@d��w����f�@����3;�\s'��
EHe�ȓ*8J�#nA�0�����L:z9��kk���Ԃ##Qd��/_<G�Y��P��T�7�J��,�� G1S�,�ȓ>1�b�H�mE@�`�L�0uX��J]�e`�`Q"J�@��ë���앇�#�<�j���7Ě��� �L:�@��;}l�p�f��O�^�HR�
�y:dP�ȓ+o�y�v��u��x4%z�n�A�<ـ&(6of������V:�Р��F�<a�c��3�Dڰj@�	Ĕ��'�{�<qTfΎr��0�j$Y�J �'�p�<9�	�=/�,ዓ͞ �*�����V�<�� ��z����Qbt����A�-�y���p����^�c�ҭ���y"�	2�쁣����U:6@��� ��y�� /Vs$P8uL�H�*,"���6�y��Ȓ"L�(���6ᬘ* ���y�ق(��9iV��-̠�p��6�y2��Y�ze�&ݱzRjGGF�y�K���3 c�r(���ϝ�y¢߹r� ���ꊸ}ΤM�A�D��y�戽j:�0��U<?�T	�A��3�y� Z�0�,M9�#N4�Ĵ�����y�C�!L���cA'���rdX5�y���?#�����,Gu�L��$�yR�F�h�-@F�F�D�= ���y�N����6��W���>D�X;���@l|�s%�4Z��=D�:���B��|`Pn�"���D>D�<���غ>�KV�>�n1�ea��R�!�'I5���(U�� 
E�H=5�!�$@43w~D:!��=	��	9V��t�!�D(�R���ꏈE�ȕ¶��%�!�� �XQ��Ja$}�S�]�W�@pұ"O�TQU�ДA����#�t��$�"O>v��ksVX)2(ɰzXr��C"O��	W��$k�:��'M� G9D��""O|H����t,�y� 	�D"�E�"O���bi	2(�P�F�N�Dg��""O����j��A!��!���'Wbp��"O-��i�	�B��T�Z3D��[P"O�ဇ�=P_A�c.G.N"�96"O�0a�f��K��~�6<ɇ"O�+�H�D��2%�`��"O�����C:��s�웱l[���"Ol<� C�4X�� �E�ذ/���f"Of��hHRLЇjڌ:�L�hc"O
 *[08z0�Ԯ\瘥�d"O�`s�㞖D\���I�Vn���"O���2kȉ^p���m��|e:��E"O@�1������eŉ;~��m�T"O�Q��F"�^�"���~�i�"OfԀ#(�Ms4���
��6��t��"O��j���A�l;5�֩\�y"O�Lёb!��	���
b����$"O�(�Վ-����Ј�Zؑ�"O:�uLC9P�H�b3#�4]��7"Or�b�AN� �������-����V"O|�RM�[���,�l�؀"Oj$#Q�m.�4iP�H3)K��"O������=���C����,Dj�"O��ȃ��]v���5P-�|ʵ"OȕX�&=O�L0J�l��*&�$�p"Ob�k
���q����-�E"O.�QB��� 1CٓD�h�"O��6�ܨa���)�Ed~8��"O��ȓ�Bo���@Ls�1
�"O�d+ �3r:�r@N�)g����"O ��c��]`�S����A��"Oy�Ő�_�F�ĩ���d�0"O \���Ƅ]S||�"�6h7����"O���
8h�M�&�\�OW�y�6"OP�@@�ȟ
b�4�F��<j-���t"Od�फ��c��)�#�T$ 5""O[�J�=N0`H�rIF�����"O�c����1��yb�i��>����"O��j���Br�| �j�5��y q"Ox�!�б0!���� 5R-:y2"ON�1�L)uԶ%j��_2Jܸ�"OpW�?8Ҙ�kvhNK�@X�)�E�<i��� ��@����m��`���U�<��2y����m(,d���� P�<�&�=�Y*��)���*u�K�<9W!��u��uK0)�&@�����AO�<���W$b��)x��PN�<����>`��p�づ�rZ2n^K�<a`k֋z���!t�Û ��i�kD�<1i�i{X�1��6v�`�H�{�<���A#6،A�X�Ro���@�u�<��*�	Zt�rF�����Ѡ'�s�<��n�eD8�0��.r�� �Yz�<�$�q�~A��쑨��\���t�<���	��}�f
վf�	Vd�m�<yֈX�$��g��<rnj1a�̈^�<!h@�=޴�!��7-m VF�T�<Y��a̪\���ɲc�.$��ah�<	` ݎR���7�\�D.L)���d�<� �xy���RWB�6�LVIXDqr"O�y[��Ll,�E/��;9��x�"O���#�ʙ$� H�VȔ''d���"O܄�G��0�F0i��K�$�2b"O`H���֠NOH1q4��._%�Lc!"O��iS9��8bG��0bp�d��"O|����.|9�āG�֒i���s"O��dWH��j'E�+N1�i"O,��t�&8�����c�] U[d"O@�k�Fj`���@:;��("O0=�U��:O�0d�p��e�ZY��"O��R�F�<X Q���٣p�8��"O<���FV� k�: ���g����"O�*"c��a,��+�6&��"O���i�8�HD�
˲.V|�0�"O�4+!
�	[�ty'�T�P1�R"O�1;�g�!|�	#(^�J3�� D"OT��"ʝ=QrځP�L'����$"O�q��-���F�G-�_dT��"O�0��艒Hx^H��.޷i&�xaU"O�t�4m��Jխ�= ��0q"O���5+ĩ~ ��7m�=W�Ȁ"OD|-T @  �+4aɔ5�"u�1�p"O�X0�]�ys����ۯ1c
�s�"O�	��͘�ъ�j��	$X���YG"O4���ĵ1L�lkӃ"�@�õ"O\��G��;7�U�!Y�R� "Oȍ�'�����/F�G��ˢ"O������pΈ�*I��"O|���'h���0샙
��ڧ"O�hv�M�4�hk�+�n��0��"Op,�a�TƠ��<:�h��"O�����$8�&���ʛ 0�j�8�"O���@P�{�Yr���7Kv�=yp"O�LhE�ũ%�hD�'��So���"O�Q��So�D$���S�yrR=�"OЄ`F��WAfp�lZ�xm\ܹg"O�hbBRE_b���őV��uy�"OF�䠉#�`����)Ѣo!�$�4b
��O>3jԲ@MI�0�!��O�N�04-B+e.� ks�T8kF!��1dzDCa'fBx0� 8K!�dS�6^x�Y�)��f0Y4[6p�!�Ğ!�����)m�iR`�
��!���^�]���Hm�����PyR+�#9  ����@w���y�d��&�4�ADn��6�K��yBa�?F3P%C�]5��"��y��An�^�
�,Aɬ��%���y£U�
�z|IS`I)#�a�4�A�y��Qj&Q10H�Z.��@�,�y
� �,���܅
}��3J�L�!"O��!�d�+5���(�����ܨr"O``8��_�zX���ky��
�"O��E�0B����u{�.�y�H
L��IS�R	%���õC�9�y��-����!7�jp"���0=��P��b�'�HTE�j�*Y�,X=x��r
�'8ڍ �F��NU�1(q/�9)��d �{2��jy�O�Ow��K3�O4nj�U/Vu��#�y�<��.S�R�
�� 
��\5��)��v�<�'j�8�M� *�,]j^�Y�^r�<�r�(�ʠR`��H��V&n�<��lˢ[�.h��^�L!}�i�<�� ���J�Q�Q���bSB�i�<GX'B�l��löi�\ BHk�<�b�?$7�9a�c6	>�	�Dx�<	G���=�Gǘ;Of2Ѷ\�<�0lQZ���0�f�9;@pP���p�<q��o����T���G
��l�d�<4�	�E2���36�V):�`W\�<�F(�*?gN�R��,��a��Y�<�͆��̨ʠ�U&H<� �C�c�<�&�P�]�:�ӣ�O�7ql�; `�V�<��
�U�iY�	DC�����FX�<�G�ϕG�đp0Ĕ�]n>+�AZ�<Y�e[�y��C�g�Z��<��(�[�<!D�Y�Ҙ�F"�'<|���O�<Y&��-px����E**�u�Uo�<I򭛊a�R��q��F�LJgc�<��D�2@0`�	��H��Y�U�p�<�tMR�j�N=� l'�<�aa��i�<	�P�4��X���"J�|3��H�<����&M�X�Ã�[X��1��Rx�<�4@P�O�x����[*8�갎
t�<�f�@%y��UX��ӛ~b�hNq�<r�%�&�!�O�^M~yѳ�l�<�te�>0L�#ă�.p��b�d�<q��S�A:5	�M�:بdC�a�<y�]`��� �e��,j&jA�<�%�	���h���N�X��4(�e�<!2��~�j�AT$�"!&�DTc�<�HZ8�>�Y7� �`|���P�<	P�N8* � ���F���K!�M�<!�(ԯ$��ժ�,052�Y�2A�f�<�kݫ{���s���fy��E_�y�X�ue�1���D5"�XuP��'�y¤ɾiO4�Yb.�W�|(Q��y����W)�%J��y�Aᘚ�y��t �۠��sNPѭZ��yR��d��l�)Z�&kV�A6����y�3�BXi���'vq���[6�y���E;��20��D����cL�y����j&�	�U�Z�z��&����y"�Z;�`�82l� U���C�'�yĉ6 ��ɚ�"����l�&����yB-�\��58�-����j����y)�I�!��m�$$I7ˀ��y� �^��P�����x7h�0�y"�J�%(r��ؿy~M��C�y�+I_�d�d��R�}T���y�_9�iՍ�U�V<aS	�yrn�&#@�ъP��'Hf(��E�y��ɗ���	S�I~h<y��2�yB�a-DDKs����`�[`���y
� �$Y0k��2�d�C[��|���"O�����:}\0:b!�>33@��"O6h��G�<*V�� ��;5�5�"O�m�W���	`�̻� A@�����"O������ZߢeF���*]l�"O������Aq��E��<_D*�"O �wiq�a�p�<sb` ��"O`a��k֣?Tt�{���zi@�2"O�R�IΤo���K���%���W"Ob������gDz�D3�Z�K$"O�y��F�g&���N6�zUJd"O,p�7��`��AZ'��*;����"O��{p��%Q�V��ё i��p"O��q��?d�^���� b=̼�6"Op�1�_{�@0qG�M�5���y��Xͩ-�� `����yr�
6�� pM�1\�*�kwl���y"�T�J�m�L��T}`bu���y�̍,m���'H�L@bl�4�_�ymEҦ�s�臺,7hQ���ѱ�yr��atn9(�	��^Ix��3Ć��y����c4����W;����O���y���.��`��ti�w/���y� �#6�����]G�F����
�yrJ�(��XGT�%	Xd�aL�y"ᓀ
,�p:4)R�n��4�Q#��y�$�89�H��J'`jR\�f�D�y��^Pu�N���4
�Y��yr�)b�Bh��HΣ�lh��j�?�y����]�%W3��S4P&�yR%V� UB(	E�z"��%��y�/\�"w����z.��P�I��yң�<�|!+R�[~C��i�R�y�#ԿZ�8d��ʁ�v��]%ƣ�y�)�X�(���?wTp����yd�3�e(6n�m���P�A��y����0]�P���_�쬑4K*�y��A�F��MAGBN�_�°h#͞*�y��<Q���
Μ#�B��b�	��y�'G�@�\�E85��I'ʜ�y��ڀV[�qC$ڊ(�8�2�CȨ�y2j4��dR0��sn^���Q�y��ԑ�r蘐OY$k\�"u����y��$�X��c�B>K/��A�(�=�y`����@��]�<��1CŢ�yrK�?�L�t0^��A��yr�Ğ{�@A��k��C8��A��y��+~0����Y�8Wl�I�=�yr�
&��5��)69v��� ��y2E�^��4pJօ,�ܻD��y�Ҝ2���n�� R���b��yB쎋!9��I���1!r�|�C�%�yң�^�J���H"�Й@����y���?�P�j�&f��%��ybn�(�Fh� �O/���i�<�ybn��((�3w�&?\a'��)�yD��(,�i�%B1e:�}HƇ��y��B�~π�H�#?h�f(J!�:�y�Cߏ>q:���?�� $�J��yd�@z�h'H��p�k4�Y��yr���\X��<���I4DY��yR�O�s�b:A+҉2�E�V���yRaÔQlL�We�(*�̡ʅ�݅�y⁗�=+�����E���z����y
� ��2jÿ^Y:�A�A�g�m�""O������uv����p�H���"O Qy�d��b��³�.�4	"O!ږ�D�͒�쏩>��%� "O� I0M�
q|��u�H\�hE"O!�b^"� D�5Ws9��K2"O��ҖX�1N~����]>3b���"O���4Q�V����8p t�r�"O�H7	�q�𼪆�Ԧ���S"O���W&ڠ	��!�0�e�҈�"Ox�"��[�dݒ���k^�K���
�"O����e�9dz�q(�KC "��a�0"O��!&"Ԧ}�tJD���"O�x`��kr �@�G�@��p"O�����w��P �ƷЊ���"O$�'��9QK�9#g��/s-�i�U"O6��%��+B��pc��[�f���(�"O8���8�U���B�j��h�t"OlX�DF��$>A���$\����"O��11��o���j�.�*�"OB�����X�DpgI�# �Ț�"OlG�2H
���Cf�(p�'"Op<q��EeV��Ėw*��"O��z''#Z��cd�]b���"O��C�G� ����B�)Ce.�""O&���LF����[�0X,��"O�7`Q�is��C� �*{�p�@"O�u�4�M� Bx���G�pjޡ�"O�#J�:'~�1H8�P1A"OJ4X7�X%�8L��{06-p"OL� ��@t�� ���d,F9;�"O�� �I��@Y�!�2t�H}�e"O�Pc��]�h�� +��`�,H��"O6}y�͡}���虙J*�(x�"O`}J� 6@�؂S�G9d
�x�"O��r���G�Zk��"6�^upa"OZ��U�9pw�̩�K�'h~֩q&"O*���K�e�F��U���a�JIÆ"O�2�ո4�fyc	Ir�z0c�"O1�?���a�R'_Y��@�.D��XU�S#�I`��S�e�fI	`6D��s��V3���g�O�U�Z9���2D��86��4͜���ȇ� �2�9��=D���k��Y���S@�'�ީ0��;D��yU�vz��b�l�k���f�*D�� �(K�|`�$HB�c�pI�W�-D�ĸ�/^�4�	���?Z0�$`�%?D�<c�*9X�"�NEߨ1��!D��٧K�b`��c]�G���;D�L��G&�YY�F�%��qz�E;D� ��,�~/
��#��L��e��)%D�,���:
�pE��n\	n��LӔd%D�01�c[�8�N��-]����'`,D�x�S`�:�,u�7 ֛a3�1D������K����IՒgT ���#.D��� ��9U$L��O�3�]��/D�`{Ё҈T��01b����MY`�&D�4q�G�� �U��a�c�n�B�&!D��j'��1+��k��O,rJq�r�>D��C!�%t�!�!�	�m��u�b�<D����]�g����� ��=V�(D�t
�jY[gΩ�c,+��՘7�)D��xl2?,��TE��a��*O輨q�������@~�ɣ"O� R�Cb��n��b���<l���۰"O����mV�#'�9�P�:;�~Ef"O����F[�t8
��[�g�zeZ�"O�2����q�f	���MW��"O� jU�Ԥm0�m�2EqaQ"O��ZCb�L��@J�k&PI��"Ot�g�zz�D�|I� "OtY�`Ό�5����m�۰��!"O��)GgE4T�LP*�끍x"$ S�"O����C�0����FM58�ebP"O�8)�Я]?lL#BL�x�՛P"O"��@������!e���I!"O|� �h�:r�2aA�:z��Q�"O��ԊK-kT �A�܁^��X��"O�Yu,I�Z��,�e��9�R�Y�"O��i�ʑ�k0Qk�
ǭ�.���"O6�Q��7Ѡ(PV�C<zA��;U"O�٨�	AQl��M�R7��P"O��&$�!Q�Lc�k�a/�$ذ"O�P#2e�?�� ��AɏC�^�ц"O\� ��U=*K��yQoQ%}�<p�"O���M�-V9�L�]�H�f"Oؐ#�@M.@Z�s���m	���3"O���4�S)
��鐀��Uq�"Ot` ��O)���fg��3�P��"O����6����І�zeԨp�"O��*5`�%8&�i���G�X�h���"OAJ
��w��| � (;B���"O���7�Y�8-�/ҦwM��HR"O|�z�j�,�R0���G�BByHs"O2i�DL���8��KL�QY"P"ON�ŌΏ<.hP���B�z��r�"O��gV�i_B�ᒧT	m��w"O�� v*W/F&0e�b&�FRBP"OPt��¼@��B֬�t�ps�"O�P�eX��Ҁ���3&0�"Ox�J�ҹf|lM���!r��ಢ"O�����C3ဘ2�AW� �:�"OVbN&m��i1 ޜ�T��"O�U��X}g���`ѷ��( 0"Of�d \>[ZTݣ�`]���y��"O*j�L�8
��'@��yO��@ "Oz�Z�$ЎEc�t�#N�7J8�"O��qVښl	n4��Nv�a0o�;�y��D�Q� Z�c�^.89�F ��yR"���p�AփU\~���!�y���e90�Z��J��.�����y"Ā�%����F*֭t讐cT�
��yRX�o� ]�Bo��v��1��H�y���BG�A0���T��ܲ�Á��y�QI�f����F�X��(�Ȁ��y��ԑ<�jD��^`��"���:�y�$O*}�����z.3�yR���'@d3�
2z"�h�3��*�y��?^`�"��E�pY� ҅���y�l�%N"^��j�Xb����i6�Py��`U�-1pI61z���c�K�<�`��,c��� �P�x�����K�D�<��n�w���q����8ˠa�J ���H�\Qp�M�ɩ�a�>���U}���@�G��|A��
14Ǻ��&�O��P��'Q��1�m=�$2��<�VP� ��*}p��+Ɵ5<��D���YSBb(I����8����6�'�����H)�(˿+��I0	kD�ѵ�4���"ڇ�.l��9��<v4k���C�:���G�T?=��S�? ��sb"6ƎI����\���wZ�\8fl�4-�c�"}�+�+G�a�L�	����U(��<�b��6��O�>9S��b�>�5ꄬ|�jE�%#���ڈ)���)�x�=x$��1h.��sM��$�U�}2	F>�E�W$����%"c0xQ���+�I�c1zU����i�+Z��(��x`]��	K(L�I�f� Ĳ4�3�)�Ӗr�@��/�F���H̘?!�H���hTAϹ �ƈ�I�r�D��yJ?)0�ʦ�h;@C������1�J��hBq�*�'��DmR�0�0�!PȆ�R���J�7W�$Q�=i5��k>!�Z�f�`��վ\u���2�>^q��}��$��wD8!� �=h�e��kݑ��I�,z� �?�J��*�������:3QZ�M�E?a�ԕ����D�$41ڕ14�]�N��Y��CqD� ��C��c��|2�"�S��$BH��PG#�	O����p�+�0���S?6�WT��baȵb�����ڍ{�nB��ħ_r\�񢪉�Ze�Ta6J	�H�\�&�P��?EŴ0R�LO�u�m���X!)L��z�l_p��$��"|dC&(
�H­����$�T`��'.��K~�ɢd^(��p�C�|{�PX�!��.D�������`�O<����LE�S&\�ȧ�*MX~�`(4�BB�	�y9��#e~���+9>ꐩ"O\�(��@�t�9b�)e7�(�d"O�`qG&Ԑ�p`�/$��s"O�="���n��iQ�\:
�-B�"O���C���|��`� )ƷP�ҥ�q"O��	uaG*���C�mԔE����"Oh�p�]S"��̑��B�aS"O�L�o�yd��@̗�Q�e9P*O���G��Q4��g�̛xk��[�'����#L�FbA�f�h�'��8��ͭ4���x��X���'NnX��Ƙ-O�`i"E7`��h1�'FɑŐ"_�����^@��'�]��Ò/�� ��+�NfJ���'��f$׭#g�-Y� %B�8��'�jl)q�Y�%�x�Ԅ�4`�XQ�'���%o&9��#�8����'p�u��H��-J���S+]�8W����'`ιR5�,
�r���K�ZT�\;�'q�9!�d�1�f�#D�&R�P���'�
��@L�%Q����K.B���[�'i�(#���:�r���A/;�r}�
�'��"�m�53����N�/eZ<��'Or�ڇ��	~p�Q�@/[[��	�'������1��x;�J�~�IR	�'pv����|�´���֡p�����'Ӑ����Ja>\Z�C�
hi`��	�'KP�Z�'"����QS�g�X�R	�'��u�r�@�5��4�A�žj>z$J�'B���"'��5���9`�n�p�'����.͞V~�SN0�T��'G6�$��EQ�b3�ʹ ���'�J,�t
5>X�
 �O,޵#�'{���c˄Z}��g����t��'ՠ�Sbd�s��(s�EԷ���K%j����F�(�I�k@�q�ȓ(K�ñ�Ӳ\��`�r'�<gI� �ȓu�r+gC
�B�	QeIMe��\�$����7W,�@���"u�͇�o���Ig��DKXܳ���}-�|�ȓ�
ё�Ğ<Y�}{P��-��lDK&��7z��q�WK�)/���ȓ3���+,���|`�G	K�^n��ȓ�2�B�e�_��d0�aB$A���S�? ¨ ��U-8�va	!�E�,�@�"O(�a��I\V�8�q.H���<�g"O����fɫx�@M�q/əV��V"O�4��e�&?]0t8��� ����"Od�v��J�^�0��|�A��"OT��a,óA�,t��$�Zgh��"O����M�>9�\���3[b9�'"O4LZ�#7Nlx��Q(J�͢5"Onx�fJ,�D��SH>D��R�"O�R��^�n��bG�;?'��0�"O֩z�V�k��h��.g��AT"O�����:w�`�W5 h,ق"O����jP?�򅋑��L�:Q"OرQ!���7K�XP�IĪ	KLY2"O�Y��#A��F��V�=
IJ,��"O�K�,�A�`���N,d��"O�Q(@ _�i�����/ fA�x�"O��Su�ݵX�p� �NV>O&N(	�"O:Yx���)O������j "O��S��Żs���C�%D���"O<5j�L{�W�]�3�Qju���T!���*K�l��!&,5x�b�����!�D(/�B)�E1İ`ƥ� 9!�d6?�d5��D̞+v�J�E$]>!򄈑L����0#X�ʛ \!�䓜+�� �DR�_�2P��$dY!��=͖�#���9�؍	���:a�!���� ����*ׇۜ̓�5!�$�1�a�'� E�.Y�&iy1!�$��G���Č��x�ZM�r��1!�Ė=��h��K�t�x��$�2Pw!�$I�
0(�z���.9��Њ6�OZ�!�䋹'4� 8�G`���#q�W�M�!�D*?��<aRa� L��3�N�:X�!�}����֦A��V�x�c .�!��ڕ6|%��ː�c���I$�]�0d!�$[�)�v[�B !��H��!�!�� � �9��]�gs� � W5�!��ў.=@i��Ν<�HH��_�$�!���~pR�k<]�L4�À��5n!�n�	s�+̯B~Xm��\�!��Z�Rp�`��_�D ���$ �3�!��N�H���].��)A�x�!�dx5d�3� �%LP��u�;C{!�ܽC ,$���%�h3Ξ �!�$�{~`�P��?����b`��!��M#>.��#d^H��1W��=S�!�$��W�,�)
���	DJ��B/!��:lH<�W�1R�TBUc�6w!򄞟a}R�'ǁ7����	36�!�8wu��L��I,싷��5Q!�d��8ϞY�&�6.2�xa�fO
B!�DV'd-����퉇$�l��08�!�d	"�͘��A�xEb� �!�܆=��Ai�	N6<	��CL�?�!�$��rp� �Rc���ZE+6�!��ZC��Plϱd�H,���ȿ[�!��G�|��@�ce�*0¨�ʳIP#<�!�d�Q�I��B�'،�i��RF�!�$N4S�:=�C<B��5Ӂ/�!��۵r8�tJߐ�~0���ċ�!�P<i䞔zq/I�Bw���a�V-hl!�D��?���ƨP�v[�9�4�͒V!�ć�I4DІJB?~��DJ=<!�� ��B�]1)�R!� (0 �pc"Od�#��&/��bfD�O���:�"O΁�#!�>\\�[���4{\�<@"O����#iB�u$)s�xi�"OaKe	�a5��X�c�4���(�"O�DX!��1�fؘP�֡)H�%��"O���W�҄�H����?#/��2"O�(� H	Xް����,��q�"O��r��ɿk��@aV�'΍��"O����Q2Z-$5Z�O���U��"O� Η;HC��r��h�3"OtiR�� QS��sw 	z�ڍ�"OtI����4L����A��n�B��a"O��r��R����N�<I����"O^`Љ\�>��]�G�O37[�"O΅�VD�"������0.���"Od�3&�0GI�B$�v"ju��"Of�B��E�(�R�>s��d"O����K�8��$ڦ���B�j}�3"OIs��Ɔ*Z�j���$�H�"O�x�gCY5jvu�b�ӝ`��DBQ"OTp ��#T�*��f��~�)#�"Oh�2�
E�u�v42�T>Pl��"O��ci�3V�B�W
r^�[%"O|��
�i$>�
��\#E�� "O
QQɃ�y�z(�-ǕnK�Q[5"O���ʎt3ڠ��n�����Ȣ"O�����Ϝ8�T(����1���"OZ����͖R�8�j0�R�l���0"ON$�!��C\�=��N:�05�0"O&��`̅�;P]�r-/�
�H"Ol
��I q�n���mܢ>��A�"O:��T
���b�{��U�<��a��"O�D�(Ç<^>@Q���)RgbxK�"ONQ5M_3���K�#9~K����"O 4�G�WC������-����"O`��N%|��MQ禄� ��@�e"O�ݣ7�ۧ}Y�����Y���@�"O���!.�2%7�5ꡩ��1�f"O��82�;E�]IC�&MJR��4"O&�5IS�"����!R>��"O`���A��C���0���i��V"OęYb`�8l���)��C"O�PT�H)8�>}�F*цs��4�#"O��9`�H�z���r�I�I��L�"O���C� %�����O?�nIJ�"O�iJ���wv���W�P���僅"Oʰ��W�5&D,���3~Ě�"O@��C��}02���֙*Qh�!G"O�I� U�S�R�k�%cH��CD"O�@�"gZ.Qga(�(�G^J�&"O�q�H�"M� ��J+,�X�U"O~l@f��eu*P�c��<�A#@"O�%oR�1,&�[�QM�4,�r"O4 (Q.	;��y�,וzu��P�"On��ËW�Y��3���-x�h�v"O����	Ԟ_�&��(�;.��РE"O�T��Lӟn0ZY9���80"Ov�Ȱd�0�Ҽ�`�Y|��"O�� �%U�FR(��R������"O�uIB�ϟ688�6/A��E��"O^�a�hN����4Nèv�����"O�Aێ_��T��n'�0e1�"O�ڱe�/�R��nZ�6�"�a"O� @��uf��u�`��Mכ|��ы�"O��P�ζ\;�7ď�,�|)b:D�����3�L��sℝNl!��_3��yB�!E ox0Ȓ�jǭ�!�D�SU�����Q�]��Ҫ�/\�!�D�.X�[х�$G@a�����!�ʯl/��0E�?�a�'��N!���b�����B�_#8��׾A=!�Đ%Z��L�s�����]0;!��\43���D'逐�$h� f!!�dV6
�s�
�$T(����Bt!��ޮT��l��e����Nڃ"Y!�ď�:���T`@ܪ�n
�J;!�$��l�h���݀>L��U�Bw$!�Ę7n���1FW.Y���p��ҁIC!��˵)m\�h5��@#FI�H�!� �mHP�I0n׭�8�p�� �c�!�䄙�.�Qt"WEz"E���=~�!���:-xjy*��N!@	p ㄋ��!����?+�E���c�T�ȗ�R
"�!��BPn���[3���e�Jys!�$�; U��#��y�*i�@�oc!��&VC��+��;s�\�7 � y�!��\.i����g��CV�])��$�!�DЅI� @  ��        �  e   �+  r6  {A  �K  U  m`  �h  �n  Ju  �{  ف  �  ^�  ��  �  #�  g�  ��  �  1�  t�  ��   �  ��  ��  ��  �  ��  
�  M�  	  H �   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b��<�ߓ#d��t	H*"F��9S�U�ȓO�����0U���6�*hU��zЀ�L^4�z�׈�/Ae��?�-O,�=�Q�A�
�b��҆��Й�I���yR��)'��S��ı>v&�c �&�y��ܞߌ )0Ֆh�]�G	$�hOb��I!k��̹�0Q�A��
��u"Ovm�� ��q��&@?1�,B!�'�ў��s�\�=����M�2��l�$g1D�L��םC���@#
\��0�$G;��hO�Ӕ���N�\�jpT���{-�C�	�3Ľac�tX<1צ;f�c����I	)��p�C�w�l�:�ʄWg�B� /-��b]�c$���bD=_��ʓ�0?	�#])m̕H��S��20Q�X�<1a�D9�%���ѽipfH�Ѩ�<���9{���2���2r&�#��G2��''`"=��g�����P2�Q�eB�yrGäw7��b��"A��$��Φ�yB��$����F��h�t,�=g��!C�NP37$6Ʌ�M����;�|�3E�s�4$��W�<9@됻0� �S�%@�=>��g�Wx��FxR�
r���K�w�X}���m�J��\؟�k�U�W�� �$!��J$D�X5�f��x%�)�T�Jtf�4Lڴ����
�\>@�ȓ<,�dKNO*�$Kr�ֳUY(�'�<!���#X�j�K2��4W:�"P�Y�\7�C�7*M���]7���$��,m�B�I6�$QC��N�s�ڄ
�+G�r	tB�)� Nu���\.N��cHF�y��![�"OV��E�R6L��-�!�� �"O�HX����mZ%/�R4��P`"Oֽ
w��4B������~�x��D�>I���P&P��4SC�@�l��ɪf��*�~���OD�ԨKX	�U P��fV� g]j�<��&L�8Y�� G����f�f�<)@��C��г�+�����rN�j�' �y/�9&ߠ��e��2EE��pv�����e��(����Ej�;Z̹�g�N��-d"O� 9P�+V�d�B��P�6v�K%�'X�R��?�"(��gć[G�m�@C��S�!�O��кצ�c+�|XG�� ��
����Bu�ӺK�yBʗ)`ZD|�b��	�Ą����&��ޟ �?�B�Hի-�9�%K�:��/�)���O<,��I�:�n�[f��8J2��L'd�(M$� nZN*��O����V=Z�� 3ac��,�Ex�MN*	9����'��5@��j�D�FA���y�g˼<q��d�(61O"�P��7?c�3U%�,�:'"Oj�XW�0Z��*掃%ub�Xƞ|¼ii��>���lF�<Y��"]�9����:D���W��21��Z��s\�A{���O<�Iʦu�'�axfP�P����)D+3�>�16H�y2�	X�1r$ֳ&VJH:�/��y����h��,M���)�y�0������?�2��f���y�ߝRtn�I���8;�i�(��y��T=���C�*a�TrT��y�`������֏��5���rb�N1�O*U��IEh:��g��6:���J�,h�*C�	� g�()Ar�����EndjB�I�Bf|��� �&	�����ך@�
C�ɲq���M׮T~�l�!��L��B�	a�Ŋg�ɻ~��4�lQ�)��O��=�}
qD
�#LRHC��JL����HJ�<��-�C��@���jG�]ҁ�QH�<ٓ� ��P�{c��D��R�-�G�<�J!>�4�槛-l��	�!�K�<�tj����΃,y��Q1l�M����?wN��d~��4G_(����B�r�'�ўʧyN���@f��S��Qzw^Ѡ<��%�b�:3�K�m[�E��O�V	�ȓX�֨k3KFQ	z������K����?!�Z+ta�aJ��1hN؋m/�h��!x<5�D�Y�O���z�fճJ���ow؞�&�x����5^�J��&�_�0g|q�s�%D� �S	 �+D�	�E�H'�R9�R�!�~����a]�	ʢ	�%ސ�����5Y߉'(ўb?��6j_�>(N8�����lU@�H:D��(��� �|� �ʧ�pX�� 5D�����ҿ]�j�(�ɌQ����`4D����d��Z��Y��	A�>����0D�г���o�ȁBB��6� V�,�����'�B���U�X�X8�s'ʡ�m�ȓzp�L饆%WLJ� t�Z�a���Dy��#�S��G����E��E��I($�W��y�B���6�J`퐁"
���� �y���(I5�x�c֊/B��跥�"��It���O�ȫ�-O%O�nD�q���4t�O,���8d:,
�8Hwj�q��Ì4�!򤐘�6�BƁ=`��d�X��a|=O>�+n���ЁR�MI|�YR��A�*ғStax�jПm�UXM("��p�+ğ�'*�I�<��I\�1|dݑwo	�%,����+�!�� n@����� x����
&'N� �]��'�`��Id�N��U �u��i���O�~C��(��a#4 ��]��"J��	ey"�Il�ɋo7pI
Fc��mz�$A!#��B䉡[�h�rw��&�h�BŅ:��B䉋r4�3U��.���ǹłC�	!%5X�5�9�@���#w42C�	>?H�a��f�4�X��#p��=q�A[r�kS"�}��
�%�N�)�ȓ:�օ1T-X�ǀ �1���P&��'��}䘶ZN@������vqp�L2�O�#*QG
-� �Ɓƺ`/B�7�:T�<
 �� �H�X5O� ~\�Dh�0D��j��'^�f��(9=&�x�)b��G{��)�)��D�46Ba��E�qO6���y��i�,ɚv�pmq��{��Jx�$�vlZ� ȍ`��0Wl\A��/���E{���^�G�ڬK�dZ;��H�4&k ���S�t���aD�9F�t��׊ۀ0v�$�dE{����D�'d$\ui_�'"��-F�'�ўb>�C��<X��[��ٽ�`H��*�	az��E�f�牜�Qg�I���$�O�\�剾)��t0D�����H.O8���Φ1�6�� �x�#!��RA�E��-�HOh�G{�w>4�����9J
���!�X��
���yb;an���t�K�I�(� m��y�d�>X`�8C��^BB������y�J�E���5�ڟ��� �.^r�r��%�)��t1T�X�s�ڱ��� �;z�
�(;D�L�ЈJ;8d2�p�Y(�f��w&y���<�O�$�$�V;:�H�u�L�(�!���'��+�l�`hS+ �t��#*Иu	����	H≚(��av��<U����D�?VC�ɋ��q�	j"���<E�B��$%��P�1aJ5#�>ɀbퟴZE�B�� �p�C��
}�([?��B�ɴuKڠ��-�	g��P���%7@C䉔�V�?�a M�_W,DX�'�6ٙ��6�����Ȏe�0`3	�'/��0n�=?�Z�C��N(�vt��'��	�k�0s�X���W�QJX��'@d��i��[����a�ӰB�V��'���uG�9\t�L+B.�)Z�ŀ�'m�a�4� �<Yq�B�<&��M!
�'2L��Y$w Q ��I��&��'�v�$l��*�����':�i���x�� ����\�@8�
�'r���Ђ\>$����f��Q���
�''�H��	H�Q���a�� ;
�'ږ��m̀Uk��2�ǒYl(I	�'�8��*��0<����B:he����'т`�V��d>�e���([֘�'Kl��c���ZL�`c`@�9vG����'2
���K��L��!��8K�'X.�c,�pF�%�e� ���q�'&�#O&��lJ`�D�~0�AJ
�'��X���<8�FH��Y���
�':"$J1�O�}{$9�R
�+m,��'7D��bM�'�*b��[Y���'�D�J�a@�8x�؂�کNe�=@�'�n1�Ԇ� qx���F� Hr��A�'��q�/�*x�T�Z�Uz���'�����kf)q푴<�f,��'�4X���;�����\#7J��
��� ���n�?>�H	�J�as@Y(�"O�arA�\�,&yc��Xб�"O�I�h��+�pi�"�l~Z�H�"OԜCgi�9��pE��0~Ab�"O�3��^t�1葊�.p����'�b�'���'E��'VB�'/�'�:��Ga�0i3r0y��]<Y��C�'3��'���'A�'��'t��'f6YRV��+�)a�)N���k��'��'�r�'p"�'w2�'Z2�'�����G0F�8tLݨn� ��'$��'�2�'S�'r��'�B�'ZPK[i��dp#�P	REFTȟ���ߟ�����ޟ��	П8�I˟$H��Η�q�E�V� ��P��h�ȟ�����H�I���ß�����	ğ<�e�V�����`� �h��#��͟d��֟�������	�X�I�d�	ڟ���Y�d#v�Ic�ZY��Xş��I�t�IğL�	��Ɵ���ȟt��Xg"���� O�PL3#�ɟ��	����Iɟ�����������I��p�E�H�1�0�~EPq(���H��ٟ��	şp��������l�I��p3Dឿ/�<�k#�W�ke�u+fW�����h�	����	�0����\����<�'��J�:�RSX�Z��aC������I�(�I����џ����H�I�4I��8J�
�8*I���Y3f�Οp�	֟��	ݟ��I�l���M���?����g��=�g+�-8k6��$p��ퟨ�����Ĉ����@&��9�2�Z?1�B����f�eɛ��4���c��m�ቚ�)��ݸ�G­+p�5�$�֦��7Ĵt�uE%?��n�-I3ⰰ0�,�$a��H��� h[�5qp1R �6��'p2R�$E���ˠ!`�at��3.*V���׍a�.6ʾj�1O��?y�����șr�R]�T	H�\V�� � دy�½i��<%?y�������6+*�a���WI��싶+|uD��0�v��lǿj�2tD{�O���ѿ#d�1R����C ʖ��y�Q��&�L�ߴ:�:��<��	$�6\�/jFvER�lD���'�l��?�ߴ�yB[��X��*�2}��i�<z���2?!��	x=<�P�/CşR;0�q�OE3�?y�Ú�wg�Z7
�.XlD�b�2��D�<��S��y���9Ң�Q����K` ��́�y�	c�v�:S���Pݴ����4��T�P=9�iJJJĠ"!
��~��'R���'s�͢������<#��2/���BG+"Ќ���Ա�޼OS� By�*E��M�plμ>�e�A����:�J �޻��K�MT�8�DRtM��Eu�}�@��o��<��E;{�l���Ҍ;8�Q[V��%�xl�� !g1pu�Ba�?q���y��O�|�*V��A�M�F��TRq-L�z�x�1+� Y��y�D�J"����Z�0tM�R����.K�f�$���͏'A\`a�5DK3�d�I �41����=nW�$���E�
d��SȄ1m�C�FN'�4t	��
:-� ��O͒n�����Z.5dr�1�����&�0ծ`�ӂ�֩�M���?!��zC������W}�T� �Ԣ��}�Sd�2ʓ@(�(Ex�O��S$L����rX���I�$Ll(
f)Cڴ�?i���?a�'K�'�`J�j �x �O�>p$�W�̃g�7�ՙ���3�	̟�hïJ�'�x���1C�r��򏈒�M����?!��B[-����?�.������I�A��qE��#�� H0��&��'�h���9��O�D�O2��n¤�� a�a80��@��A�I�� yK<����?K>�1y4^�_8��㛁8��@mj}�����'���'��_����F�%0h��!n!^͸ToM��y�}R�'~�'2�ɭD���E�ٿlF����,G�kg!�I��X�Iޟ���џ�����������?Or��%		�J3p�*�Y��M����?)����?!��$9s� ���7�T�,@� U�	e���ν>���?������J�ҭ&>�*� ��9;Hp�.E0PWtQ0cě6�M�����$U2;%�O�*�R?2�4Ez4��5�Z��1�i!r�'���'$Z<Jt�'e��'i��O�u�@),�~��U<(�^�+��#��O.���"w��r�T?���iUfM��	X�W<e���}Ӟ˓��	�Թi(��'�?���)��� )��1ciߵ!RZ����'�6ͳ<�6�TL���O���v�' n���/�E��}{�4,�j����?+O��	�<1+O*`��GR�t�ȹ"5�$[��-��Ʀ�ʵֆ([�b�"|���TU�)�T�\1㘸�e�U��$�i�B�'��H�#�X6��O����O��D�O��G�<`HV@�7~��uN��4�v�'�2�]�_TDઘ�������$�O����+$X���ϛXx�-P7��O��!d�ۦ�������	�\b��:��%#bElTP�Ȑ�ba�
l�7��3\���?O>�D�O4���O4���O��ݪ bn�ӗ$�Bnb 9�G�+Or�1��Y�������	֟|k��pʓ�?�"mE"0e`l����#��=�d�g]�E��?A��?����?�/O���ÄW��H�NxY2���;Ϙ�� �k�
��?�.O��O6�$(Zj�$��#�R�H�'	�K��l��`|��3oi�V�d�O����O�˓���U?���
�*��Ai]!W	8��!��~��4!ߴ�?�,O���O���VtM���O��$D1,�*\:���v6�T	���-n�L;���O����<ɕ��~��џ�I�?�T��o7����ō�)rY#C�ʍ����O6���O4�*5;OX��6���π �IcNpD��#��m���7�i-�0Q��@�4�?)���?q�'}��i��Ab���MPv�8u*;Um:��$hsӎ�$�O�H��;O�OH�>=�"˔����k���Wfx�D�rӎ�H�	ݦ5��۟���?���O��E��0ck��c��yc.��H�x8Ac�iP�I��'lY�<����Rm��fN���Ж�d��ڥ�iJB�'�B�O�^C�7m�O��d�O
�d�O���0D`��%K�0�� K�#r���'�B����I����I���$�Oh��K�1��A!@F�0�0�6�Z֦��	D(�ٴ�?���?��m:��w?q���\ x������TSM7��T}�(�/�y�X���������x�I	ִ�h!*T�_� P��͌*v�8�(��4�M��?��?�R?u�'E�B��\��7��)ݓd��3�q�'e2�'�R�'�BV>ipR$ͻ�M��$AV��*�+t����G��;{�F�'���'��'+�	��{V�z>�𐩁/8J�1��<E>Lm*Q( �M����?���?	DY?Hba��M����?�g�/d��ٷ����q��K�R���'�B�'��	��i�bi>��Ii?9@��2y�^u�#퇜F���:�����}�������ן�f�5�Ms��?���r����7}>i:�Ǎ9y_�%�t�X̛��'8��矌w%u>���|y��M����H�еoD�E���9�����IɟX��n�M��?i��"���?�_
�"�.�y��L��O	⠴p�O��DU�AH�$%�4�H�O����ͅ7A�D����+��Aڴjhl���iw�'L��O��d�'�R�'�u ��$
�!Ќ@0;��2��d�`�`�O��$�<ͧ��'�?��W.b�"��J��#��8��.�#\��f�'B2�'�"y�?���O�����(��M�Qh!�/I38(xz�0�	�x�b�X�Iş���6JV�� ��zD���Ȝx��yq�4�?��hDU3�'��'�ɧ5V Fy�8�0�`��e���aϠ�����3�1O���O(��<I���HL!C^� ���n���][��x��'���|�Q�h����`N�� ��������:�c�L���(�	myr�>mj�����Z�-��%;uę%	���?a������3��'"�*��c!a�A% W�3լ��?��?�.O�e;�ly��J�5#��Y5]Q�F�W���ٴ�?�O>�+OHiҐ�Q��Y�*P�{^�� c� ����'�b_�`2��1��'�?!�'���c��
�v,C��R�ɶ��6�x�P�����(�S��%V�2q��z�HU�#��r���M�.O��`��N릩x��x�D�~��'�TU�2(S�2������X��Q�4��H��b?1�1DD;9f�4S@Ĳ z之��q�0iQ��ئ���ޟ �	�?�	K<i�2"��,�y����á�-6KHiQ��in>u����ß!أ�m�R�N�8{x,�����M���?��I�>���x2�'��O�Q!%��?!�:yc\H[�a����P�gN1O��D�O����A&ސ���i����ݯC�oZ۟�Bk����?����Ǝ�"F�)�Ч['b�,:R��o}G���'�R�'�"P� �W�:'��̋���'B�ި[�W�$�hJ<A��?H>I/O*�� ��?*V$֊ٝ(�L̓O�$!�1O���O��D�<Ѳ�?e��X�U`6@aD`�Yt��	��޺G��I���I@�	bycՓ��dE4o�<��'�I�Cĉcƻ6��'���'�U�(Ё���ħo��<k��قt��xR�ȆN�:����i��|B[��:��3�ɭ)/��%�V2<��0k���6��Ot�$�<af�c�O��O0�$ŗ�_Ix���ʋ�aY��� �)�d�<��Fi������E���5���Wj��:TlݳS>��X�� ��Mk�S?����?y*�O:��R�D�F����$<R���
v�iZ�	�R&#<�~�q��}�^܂�S��]�4�W��5��	�?�M��?�����q�x��'1ؘ� b�`�$�*Q��G���HA.x�H̚E�)�'�?�1�"qFhH��P/1l��v�2A��'H��'���+fO(���OH�ĺ��s˙:�ZrKB�Ԥ:�($�	l=��П����\�����r�L�I���`f��2�lL��8�MK��"�"�t�x��'�"�|ZcN��b�cT U?�]�RbC�O�-��O،���"���OZ���O��&J)�盼a3Q�B�[ (�u��F�v}�'�'��'�	+lߞ��%�-/�|�!lB�@�
�w,,�I����Iܟܖ'��S�~>��r�C�3IaB��P��X%�2��O�O.ʓuD��'�AK��H2`��U�s�I3`��O��d�O.��<)shؾ~v�Oђh���bj\j ��A�v��'�l�B�'�d�<Ѧ��S�D�Jѓp�F�F�V�hUG2W��o����jy�/��eM��r����
���!��7n�������3%�TD�	Ay"hS7�O�i�+
0\u��!ω6
���&�-#���o�֟��	,�����4�?�*�8���m~")6Z`0�w�V9p���T�V �M�.O�����)���H�d�Le�|���(S�'�>6M�_�:�mZ��4���X�S5���?���r��Y�5��&u��y��A�w�ƥV��O��$�O@� �BFa��Z���%d6�u�"�i���'�B.N+)�O���Ot��f���p�N?h�V���	�^|�>Y�Nh̓�?����?�#@���$����/�"�Z�#�V�'���Yr�3���O����O���k�/@�:�T��f쏧P�:�Bg%�y}BdI4��'B�'=�Q��Ҁ�'`ĠyĦYX1T�A���Q�H<1��?�K>9+O"0�S`\�j�b8���%�����rT1O����O���<�S*�{�Ɏ2H����+�+W�1�L�[�	�����I�I@y��؇��d@E`�]���5TY� B!LH�9Z�Iß�����ȕ'� �D+�)rb�
�(��5N�����'YB�mZ̟$&� �'���}��[XX�A�V)]5�d��:�M��?!-O��a3��A����S 8QYtG�Fnj��g�ŚX�$O�ʓ_���Fx��Н���=1�r�d�4Op��ҿi��	�hB��Aش6��S؟p�����B<�� �B�^��M!�aՂ(훖W��q!�S�'Ny�H@toGo���:( 6+�7�ޏ:���l�� ��ğd������?ɂg�q����
9T���iԮp��&�+�O>�	7� ���L�\e�bN�p��ܡݴ�?����?�a
P�_��'���'��d�4��j�5U%�u0��5v��O�c��d�OH���OB�[DF��N�D��"��!e,�bd!Tܦ���!9�Wp��?�H>�� �fxx��-����KŨj����'��$Z�y"�'���'+�ɯ>�����hFp���p��!H&���U/Z���'�R�|bX����N��\\�p�(%z8��֒*�@b�8��ޟ���ey2�+]���=/[�����߯}D����� �JO���-�D�<��@L}�ǽl��A-[2q�BE� �K4���O��$�O�˓r�nY��d/[�1���yFǘ����#���.�7��O��O�����>��Ƈ#��qz%.H� :Z�qa#��)�	�� �'Ryy׍#���O6���f�91���~e|�i��_�:�5%���'3 ����T?]BV-�4a|X`8��F6�~��R�iӨ˓T|�»i,��'�?���L���Fɞ��f��R���Y2�6�<A���u���O$Ræ
2��\�@�^{j��ߴ	hu�iV��'���Ok�O��d�I�\@hI�i��ً捑-t9��oZ$@#<E���'.W�F��L��������A�bp�����OT���;��&����ǟ�[�J�[�+C�R����@�-N���>9�o�Y̓�?	���?!��FG���e�	n䀔� �ԱX���'�p�JA�<���O`��&���"���F�)A��-b`��t����T�|"�<�	����Iğ��'w�X�A�S,�]�`ā���)�""�ROp���O�Or˓j3�`R�dL�'
L�(��oX��+s�{��?I���?�(O��0���|���N���%a��U&�����L}�'��|^��*�!�>A@��Y����N�gr,M�q��K}��'FR�'�ɀd�`|�I|� ��`�̕ ��F 5����	Q�l���'$�'��	�L�c�8Y��ǈ0� Q��"�^MZ�/u�d���O4ʓ+�R�ד�D�'[���Ƕx�r�M��Z�� K�G�O��@�V\Fx��p�@��	�j����9H��X�Q�i	�	�ֱH޴%����`�9��d��O�� ���G'�P���	H
��Y�Ը`�#�S�Ys:��ՅJrx��%�$n:R l��%9����4�?���?��'C�'(��#D�����]!���):!| 6M�Zk���3��ϟDK���W\Ո!D;�-!�(@��M���?���k�9(��xR�'fR�'V\�*�|��� ѱK"Dxa�>�	63�Lb��I��I�<R��d�<]D(O�%/�l-�ݴ�?�f�F�}��'�R�'�bY���#���R����qZ2�	eȅN�D�Xt�<���?!������t¹����7W��!p�F�-`�!�'Ck�I��D�I�'��'q`$[�#��T�|��4S�4�:|kA����'���'&B]�0�sKDQb�c��ZNQ�կDYq�D�"F�V}R�'E�|BZ�@�5��[?�䬎"P��  G	�HL���BO}�'��'�	)l�,%?�񠧚~a"��%�)N/D��$A��M�������d-WT�@����<1B�IU�%Z��"im�|���O��P�l���'�?���45�#��>r�\������ꕸt�x2�' "c¥mb�|��\�v"5��]ٱe��-��k��i�剂_��0�ߴ��ßx�����4A}�{ �۳;v�3��K��6�'�W�x�R�|B�� # Dٰ�S.~� ���%C�����%��7M�O��D�OJ�	�r�	ğ�H�~�x�����6"̝Z���M�s�]S�����DQ?qڠA�l �yQF*Ů͂Oirmm�џ�	ȟ�x��L���?����~�G�Yx�y��G�?���;0�F.�M�H>�T,]�<�O ��'��A�B�����R�ȸ���[X �7-�OX�1���Y��П4�IY�i�1�ǀ�OI�� �sؐM*f�>��؛�?�.O��O6��<AF� �]�׆�i  6I�-�����In�'Y�'�'X�'��<b�$�i��ظ3R�$*�:�M�.|I"^�T�I���xyr�M4T32�ӫ~��Y�hޭ6Q02p�������?������?���SW^���C�����]�-pL�Sȏ�yrH�uT�t�	ȟl�	my�	�q���x�Ȉ a`�e��q���ぉ��	h�Iퟘ��@�b�8�U���N�*L:r(J�x��Q�AwӮ���O�@P�j����'��T�S%-7�e�NI�Pll��CU6O��$�O���	U*E��Z^�tu��Q��}]n�Pyr�1aN�6��e�D�'C�d�/? F_�q�	��i\>]�@�Aȕ��������F)�ܟ�&�b?p6*�K�. !/u mq�yӀ�+�i
Ŧa�	ݟL�	�?��H<���R�� ;��S48�x�AZr���$�i|8a��'�ɧ�2�DN0M�Ra T��.[j2�1@Q�@mZ��4��ǟ"S������?)��~�!�����^K���g����'��x�Ғ|��'�B�'� ,Ir�;M
P�:�]�2���y4�x����Q/lH��'������ %���V]D*!|)�5�BoǦDj��E��yR����D�OP���O�˓\�H!N 1�R,xƠA��A!'ԃ8�'���'a�'���'�M��ҍ&a*���\� �f0c��RY2����U�2�^�{r��Zf�-�L~��
2��,
NO��"ք�P�<� ��@j�O�u�� �!�eܓdK����-R9$�8,��œ�u|�3���
u���"�8��A\�8�zE؀��9!U�!)caC�u,
�
ܡ5a���xdPs�	�<��$�U,�P>��aD?s�l��e�`��@:K7�TJZ�Kܜ�V�>z��� 4�Ù-0T'*�1W�2J��&}L����C�O�*��؈U����L <3@��G�ON�$��Z����0��i8N�K.Ѧ�qZw��]�R>]AF�.���:�N�4̠���i-}rK��D�s����E1��i�ם� �|�mi��"��,��U��mݨT�x��O��b�'�������FK�!-�ؽ���:�L��dA)D�$+v,Lذpa�j�?6 ���%O�Ez�͓b2쉄L�DU�d���=�>7�O����O2����%�*���Oj�$�O�nG�_���h��Փ{X��p��ɕ?|����l@�_�����45���1��N�g�I9rF��fތdvXQF�_*0y�)d����uI*=;n�#�h�
�q�2]`d\�\;C�f����,체�a�]�M��\�|y���O�I���[&�����b��6_q��AO;D����ҍJ� z�b_1�0:m7?��	"�M������'`���"�f3�du0�b�q��=����pb��d�O`��O���;�?�����&37��bq�C��}�BNU=I9�Xz�eU�!�� �M����y��X�@W���"O2c�4t��nŸ*���C���4	N�u��-��y��4d��Т�l[��!�g�7���C��?i���!�Ɍ% ��K�bֿO}��Q�[f�C��7a8��#k�&?fd�EM��b���O�ʓ0ر��S����L�Yu'�0�40���W)C�̀��՟����Bǟ��	�|ڇ��#n̙�$5t��Ċ*S&*��.E�y�h��֪�+(�xbmG' �:�f�8^bl��A�Ԑx:�D�C�G}5�܋r�X�"Z"��僼]�\Ey�%ʕ�?�����D�K� ��N�Z��ܪ�M�{�1O���$H���t�W�(f��,P��8E!�ė즥�W �J���)w�_Wti�C�b���'A��f �>9���Ɉ� H�[2N40(�u�6;l᳴��p
���OL-��$%}����DW�|Y�T>��O���Rd�(-��C�Ӛ.��QYH�(��둼}4Ѣ�d��&6��ҏI�(�#0�?�YQ$�2��Q5ˋ�Ybm�҈"}�
���?�d�i'^"}��'Y�*Q@"�����N�('� h8�'@ِ���5��9�'�/\b�i)Ó+j��@a!'ѯT�tK�b4c�p�@�M���?�L��#��!�?)��?A�(�n��1$��HJ��б��ſʔ틐QQyb[,���R��L>)M��f\���T�iQ&!hȱ4p�b\�t�W�:�q��'��M��U{�;u�N,w�B5���~�N�'vf�C�S�矐�I�8s���w du�D��eǴ�i"�N{h<��D�7]���E�a�����O~�:�S�dX��8�dPo�N�Ȁ�Ùp�ؠ��Ŋ����Oʟ��Iߟ��I��uG�',�1��x�Tf�15@t�pB�\� 5"��  ��X��H>'v@R�+:$�ax�@˟y��QjB+Ψ'�xT��]�͛��?�:{r��!ư���<ˈO�qⷠ�C$ �B�PC�$����ourir�vM&�����L�?���8`͘��1�M�7g����w�<ag"�[�(�i%��$[�\��H̓=���'���*W�U�ش�?���9�L5���7���P���i~�����?�Q���?������D�&k~\�����(�8���i$�[���0��)dP�z���Z�W��d�{9 �2�L��{쾍i�g�@s�TeA�S'"���k��o��D|B(�?I���� �!�� ��@��d V�D�!3O����O0�"|"Ån��if@V�"�D���NK<�4�i���䟖W#�3c��<gn�4[�'~�I�>t��)ڴ�?�����IHT���d�<���#҅��0V`�lC�h&����O���p��'���t�$׺d
�|�(��	�'[SB�P[t���а�>��!��9ȜA�pEK�1�F�"1̅I��%���Sf��LD��È&&��<�O��:R�'�\7M�O��$'���O�#�,R�9z�e�p��� J�e�O*���Ol�/<O���0��=jћ�-�5A��s�'2�#=� ��q1J5��lM8u�V<X�BS�Z���'�r�'��9i0�����'��'�֝�f�t�c�ɛf��b�㉶��ʥ&
�D����4sJ�33m�y�'EJF�z��`���@�	�rE$2��8z�2U��,��0q� �BM�t�x	�v�R�n��>�:T/�M��$Ԕ2�T��u��{�ƹ�ōL*ي)m����E.n������?!��7AE�׈T�k+�|��Gĳ�̼�	�'\�#%��<0R��d�"0��OڅGz��O�rZ�tJcb�6}/&5�dЪZ<T§-&!�pq*��П(�	�� �	��u��'��8�"�S�
ѐg�Nͳ�P�]\M��'��	4)ش8���{C�Y�� xB�܋�(On1��+X�4b��P�gB��A$'���:�� ��m�� ĦyʗBZ�TIQ��R���k�c��ZjB�d9��S�S$���]��ݑڴ��'a�b?I eR>M����h�15S ��@!D��"Q-��ݖ�⥇0D���/9��4�M����]�(o�y�'�"�4z���pfLc4�;�㝜m��'�hUY��'0B7�xe��ډ7N�pB#d�>Q4��e��]9���*dK �b�Kr8��2Db��W��a��,/�Ʊ�!C�U���{Ԍ��l�rH�Q5|��xB�Q��?��i`�7��O 1*�d:���eM��r���BC�<9�����.Z��/t��GַB��	J#O��m�cx	�5���`ƭ�W&$3�<�	NybM����6��O��$�|20`Є�?Q�� .���Zv�C�5���AA���?���mt��ڐlх.1��C��Q)�*�Rʧ8�sS��E�M�,�j5�O��5gV�
-6Uz�AO �8I�,�Qp�O܌!*�蕰]j^��(:�x��J��01��On�n!�Ms���OF`R��O�TR.<�BB/���+�y"�'��yoV�Y�d��V��&-J�`s'�U��0<1�鉶%F��8BK�hAX��x(�uS��Y̟(�I֟�R�ާ���������[Zwd|cԹ(���B\'ee�49��Ϳ�����D�kA��å D�Ce1�bO����u��H�˜%
�L�s�4P�hSD����S+��wq��O$D��GN?q&�D�� :q	BɻDT�	�/OޅK ���t�OO�OvX���� -���$U���t"O����Ȅp�|�i5�+t�N��t������?�'% ���@M�O��D8<�� �@�
<�`���?���?a�'�?I���?���G�:����K߉$Cf	�D1W��
�'w\u�AN�1a@���N53$�JŌ�8-Ī�Ba�M�hK���P���9b���3��G�NnX��'�<6-Ȧ9��^y��'��O:t�k��u(��m߼`�Ze
��!4��U ��2ҫ"��9�������OPtm
�Mc.O���Ū W}��'���ps-\�yB�Bg��I��%�C�'��E�r���'��I�H쐄+Fh o���r-F���P��恒P���%� ?"�`#b�"�.+�� �#X�o�f���L�?��T��	I	�a��b�:n�ڌ�GA.��O&!ж�'@��'��)�~.���C��
��d�'eʌ/��Iß��?E�d�UR�t�%��9B��!@��x�Cr����1��K�zl��eP	Z��1Ovʓ-��9V�i�"�'h�S
zF,��I?U0�agLB��;!�
���Iǟ��Ʉ�%�!H��'ڹaG� ��I�|����pmC@F� ��G*{����^��Y#f�^{�(+]o��}���^ 5G4}���|p4(�,�w�dO8Rzr�y�T@nڟ���tD]��v5��,�9l���"�r̓�?aI>Q��?�)O>Ɂq@�	QLqgl
��U�S�'��7M_ަA�ɩ�M���;$�u�V�~�@�aF�cTH���?��"A"�s�A�����Q�.b�%��H�`��fě��kq*"M����+��1Rd�]�Z�q�ꁛ@�هȓ$��@ ��G�$�:�Ӳ���R���{>d!F΅C���J�� f�X�ȓ�}�s�I�UBj�����o�Թ�ȓ��u�V�̒-�2U�s!#8$��E��l�d�DYs����*-A�Q�ȓ��31
�D����e��&$J���S�? ��:G&O�FHk(ʿI��TZ�"O��%"[�:6��6)[9��H��"Oj|���A#=Ѵ�H@'é/y�%��"O������t�`�&q��)4"OfXP��\@<$q�&��|Qh�8"O�l+�
�D�ª�  9�`w"O*�6i��&	��c�L�S�"O� 4�	�>���ؔ��=HZA7"O���Ҁ�Eガx�fE�iVD:�"O8|S�Lu��`����S�HI��"OD
 !^�W'h`q&I_�+휹#�"O��X��;_��(#����"O�U�g 8B�B�@��)bT����"Ot$��A����p�Ä�}���y!"O�GѲI�M�҉ޱ`�X��"O(z���RS�ܠ�O�=�B�u"O�L�2�(K_����-�6
��D"Oȅ�F�t�ddJ֋�LϚT9V"OR�1'T8���tm�.�>�X"O yL�5N�vMp�KVt��"O޸��d@�$!��*��u�	�w"O�DX�c��3�Pz��==�(���"Oh�zb� H���V�O,_c�5�ԏƉ��$�>iT�/r/���sӆ*R�Xf�Z)���R�Z�UiX�b%��bb���/��֝�r�L� P�bޝ�E�T�a�=�E8����)�L�����-_�&
U`"M���a�_�0��Or���&��#4|̙d D�4P֖xb�ȥ]�Pa�O�tyVD�.=�~�S'<
�O���|���
�#c�.옂BŠ|"���ҽ4-�:dǃi�T��/<OM �I׊ю��O�O��qʦ�� a2|��`�ܖu�H�d�ң��,� �OYT4�(<��6@�|x�%�4�j&�ܺl��m������(O�S$*�<AeoX�3�H���'qzD�v��3v��9�a�����8g�z睶[rF9������It �t�6�d$�S�O7�0��1qv`�s�h-p�k� �X�1�g�;z�����qPZ�O2��E�[2&���@1k@��J�\�Dx�%	3Bs|��1(�)�J�C�A�
��lKcC�9����@���Vl��'�t8���N�n}�5bՆj\�mIO>��O�E�Q�'"Hp
���\�x����'��z&��P�\q���=l��D
���O�O�U�Wl��{�h�D��%��'_���T�iChTyA�?yEp0�� ?
LT�2�V��HO�.��?r��b�;�F���îr��"��N;ĸ�@6
O@E�"e�yJ8<�e���
��hKR���'Z�U��ꏴ}��(��,��B&*��O<I` ��RxpB��7z����Ga�v8��I��=b_興F��-[B�.��n�����3mT@�A6��4��	�-]<�8�B�9$�X���I�Ԉe�7�X�'n�p+�	���'�ܩ�R�$M��4)��
�lz�����ģL����UƁ�)!�=1`�U�`hHC�Ipw�I�-H�x!�ǚ�h�sO�1\��U��p��"�ϊ�C�h�]&.({�lB�`�pH
3h�ZC�	3W�Z0[uV�m�Ĩ֩�;A0�`@��V3L�~�b��� ��)�U�C;7�Q��bǨJ'0�K$MSJ $�`�=�j׈
�0�I ]?�!���%/z=��ލ$V̵y�F�Y���<y�N�w�X��ǣ1?��Jf�L����'9498�.�'��,���f� 1@�K��sm�}`E޲-�\\��+N+��b�ݡ��"�\̹�JAk6����N�i����,��|RD�jU
�>F&��^5-��I�-J���IT~��O숑:�Z1hH>pAN��?��4�N��R�<9��>�lI`A'ՠp?�4ZB.WEF�q��ĉ������䨧��?��j��*�&y�Յ�Z�R���� m��I�� I���jy�a�']X`��'h�2MJ5�~�`�¥+H���P3�+�W L,�$�h���M��~rᚦC҄����L�(�Sh�-817*�>i�Lʓ}� ���h�H?ц��!E�
�<�萵?m�fNߟo�ވ"$D��MX��}��?]C�\� kv1S�iN�z�&��$��o���nE�#>�QϤ\λ��a�2l%�p���牙#m���	F��H�^8� �#��8r�+��9�d��&����O���G�ns�jG��bՕ�H�mE=���cN��N5~P�m�>	C�'���gFШ�~Q�e��QV��@kL7_��ayG��o�|E��a�O4�u�!D�7$���r�G�Y��)����{�	�<p�p#�*�Cި�SOP�$E�P`��8`�6���>.��O� MI���1\�d	�^�<ӗc����'zr-Fy���1��X�v�:�b�(B���D�	13K��k#��
r#=�;j����'�fމc!�սh2L���D�|-#���OZ�=E��JV�k� �Eh@ %����AK�]"�LEy"*ɴ+2 �A`P e�����I[�����
��պ����v�ޤ��#��:b0˓�Oj�J��S�&�R��ET=qV!��F&u�l;r"��3����6�G	�dіc�r(9W�+/n�r�H5^�'��Ɏgڦ��d^�A��|�2��U�>�d?6����޷is�Y�Ӯ'ZQ��լB�X8�x`pO`�
�1���M�TF{�O��q�H��� D"Ƅ�$��0+TB�9'�x�UP�HO��OȀ�cR0�,9���6jx�'�ԇ%�4��G�'�ў"}rpR?0����Ԯ_��Q��Ecc��jg�8}�Q�F��;~x��6���T��`��d�{�X���PM���e��`��&;X���@<�PxI��E)�V�J��M>l��MB���mQ\���aՈ$;������DI
��?%?�d �D����3,�	#Z~tC�5}�oH�Sƴ����S��@���'�Af��m�>����i�1� �	-�a���ԫfʂ�Q��1�؀
��:-�L�h�$=EIX���؁���y��� H&$w%�7[ۨ��m8.Y���l2�)��,Ox�*Pś�e|��g�׹�J��?9�IM�Zٞ��Q��K�U�UǚOy£���d%Jɪ=�f%������I�d̘��'�O��S�4#Q�x���Z��*,2<dH�hT�+w�[� ϛ��rZ�\�'�ΪD�qO�>���	hR�4�@HY$���K�h Hܓ X�$I0��x�V��ق�Á�o��u���_"*�� OԵ��^)(T��� �e�tP��S�9���`���_%0�B|�M�&[�P��ǀ�PV���d�1l|@I>�-��J���b�.� Tj�I��ǆT�'�U��C�'4��e���V�$���ٍvC
�$�Hڷ��[mqO�����E�>��HP(�-7���bQ��k�hU�aqO�>`A��-r@�k�K��b�Z�a��a�+-��ZA��x�I�������L��0r�	��\��'��<E9��k�'&���B�Y�a�	�'�5}��h`֣�md��8��@��u�G+z��Ӝw �a��AQ��	D��%���
6;��⟢Z'�x�j))��� x�6u�ag@�`�[h��b�������R��@%�`�K�S3$zB��?{&6�v�����%��s�S�A�S�f	9DK�����(ПGk���Ǡ.L�SDm�<`�{��1\�z����ا��O�������1�W;��3W�>1�kH�6�&b���39 aVhI_������1�/-oV\ t`�s�`�*E�	�%Q��R���R&oރR���Q#Ě�\#@4*b�%r�<�5}�ԣ<��0+"r��0�N����edItk�d��Ĺ��'*ў"}HEX2�(�MN�@H��H�H��"�
�H�PH�B��e2U���n��ɕ.!}��V�-"L@#�����e����,�Q���tn!v��0Q�$=42lkc��j���C�O�9��W/��<�bZT�����ѫ=ur<hg�j��K~���y�|PNJ�d�憝�?�s�اau`���CF��n٫��I�'��
 *Bx襣&��P�ڌ�A�'��O����b��?SD���u#u��<*-ȇͅ�q��(�5�K��@EzZw�xUX��+�y��N��[�E<[����,Ӓ�?�y�(ۂ{=���&DFm�'X�:LJ�!W�(B*���MH{��	� �1�Ƀ2B4�r0!��=�	��.�a��O\	$�̼�|:�k]0~l�m Ĝe�^�F�ص���?��Ӈ;���N�&R�\ �ӗ�A��ɏ%P4��L�yZ>|kE �A��ZMC LT �O�Os��3}7t	�#Oɥz��p�G]?~M��D�������	)
�t��ç�'zn�QK����'b�LRc��r]����Udx�#�:���'gp `Cmz�d��4Mf��t��/Н&�������c��^7~�kf(QJ������/Ma��	k-J�+��̻I��� ��",���$}D�aL�X`�L�Wm<b?YiUB[�L��Q��	ye0賤BG$"��OT�@슖TQ٧�3\r�a�c�>)��E�jQ���_�kQ�C%�&�V�'n!x�
��擂.5�PHǧ�B(У� [�nO��x&!�8#��\:o�T�I�'گ'�ҍ�4�O�x)�"]�|Q� c"���j~� V��jd�d	�<0v2��\�ڣ�O4/^��@�K�@?y��>���<i� *?HTUyr&Ц:�d`���ޟv^
��'�u���'�������
��n��P��Z�@i{�*P:C&UBԇP,�牖w,�7�I��Pe�O�]iq
˔/k����"�t�C�''��`	R���e�A��a���P�'2t��:ф2��(8�IP�[o�(`0�Ï�(O<�*ь�>� �ōw�1��'H8�˓k�R������	�e_�\��V���a���8J-�AZ��p���]�a�HH���K{}&ϝ<����r��;%@_c>~�������'�~���ɛ3y!:I"sG���$3����?
�z�1� �����V�n>����N*I~�CD,�p=�1a�'
��J!N�H=���3\�����>)����\�r�oz�� �0��1�h��Pg�g����rC�l�Z w�:O�����OHX�v�%Z���$j=�G��<u�.<�FL4�,��f��	%��3._���ъ��E��,��}�l�a�8��3�t�x��S�Z�$�h!���*��h�d��*)��I�!1O4	������:�/]��� �ШW�G>����T �Ɔ��5zx�C�!Z`�ӥC�/�����7r����IǒH�~�ś.3+�eZ�2' ��V�8�N�4V2��?��ƟHlbY	�P) $�Հ1�D�q�!�Dބ[[|4"��	�C���r�$G���L���Wr��A:p�8��?�p�,W�Z�ψqz���f�L�v{t1�e�}��d�}�~��K.��!��]�\����C�#�\�x�'Y�r�JA�'����	 XY��Ō!��Ȱ�����������'�9�L��eIU- �� #[�B�����uX�əuI�\���_n`�[�͈�ā�ō�+EAB�'���'l(J�f@� \3�*�=/�DX���C�3-����jZ�e�l)D}B�ڵw�䌨 /48�P�-�t�\Ex����DӢ�'H��k�dSJ���Q&E 
�X�p发V�6T�`�X{��u�D� b���*�w��)W)�0,�C�J�G@�p�����'}(�BF�{e�y���E.@0���
�]ɓ�D�!1��B�MW��Ä<��'j�� �A�W�,�� D�k��&�=�
4{��4��ɒ�O��I��� y���eT<h���cP!��/�x�i�N�8B�Fā�F�B��րW�fl�㟒�.%�cGH$4�P,S��
Xj�ᖗ>Y��T���"�%߅D��	���j��%�6#a�6,�X8"o��`��\[&�D���0|
����`}0��\g^%ca�P� `*H���'a�ɉ��O�^$ae�@��r�K�i�����W'�!I娃�!��������7/�F�bu@a
P�`��L㟠�'(��/��*��6B�
Š�<14�Q`��5A��֔�
�3�ؓvy��I3t[lL�'E�|:R��!_Ş��� �QNh'N�^�2(!�]�+0�'�LH� Q�1�s@�w+���'���m�<D�=I��:80ec�'2�Ix��fŶ���OV�*I2��'[�Ĺ�j�vtL�b�_�md0�`�'p��&�>�$M��Eþ_�H��'��xp�(��}�J�ʴΕ2]
�[�'jͫ0���c��k�ȉNT��	�'�*`��Y�O'�!IW�V�B����'�D"�"P(M���Ɩ'd����'��d���üx�{E���H~^�{�'D�RS<DҞ�W6�L �'~�x�G�U(&p���|$x
�'��M���H�U���Ѥe���8!�	�'/x���`�<a���N˔�@	�'o��Xw�ٴ2h���cn���h�'����Fa�2&��zծ�+�'ܲ`���m�&Y���D�v��t�
�'Ռ�w(ݷ+\M�` R
l|z}A
�'`�Kf��c+��@��ٽW�r���'��T@�@2Y溉X'�Z Y�89�'��yjeM>D �	���9XQ���'���ťQ$UF�1V%E�����'$} ��C r�I�#�v">��"�H����;5�[>���ȓ�L��a��O�}�&g��pw���ȓg�(��6���"���#JB5�ȓ�J=I��+\���	�KY>H�ȓ(ft�i^�?�� �$�,=�`�ȓwfvA9���3��|���VKX(��%m�E��&�]�bi����z��8��mF �I�͟9������%
Ʌȓm��1 [4}l���16.�\�ȓ���Y�B.���q֭�+,.����y�(ֵ&� ��C�ys�E��a���pV���yڣ�+�,�ȓ_�0l���Q�Ei<�)G���)ÒЇ�Yʢ��@(5��3GC<���ȓU֎��]t��������S�? (ͣF��<���8d�K�|��0��"O���%E����ܖj�Lr�"Ot]���3Ulҭ��BV4dI�"O�a)��5S���P��
�q��"O`�Kd���gmn(s2X9���ɗ"O���w�A%c����$T���8E"O�����.�y�#�>0���*�"O��[�.-������@�Xt��"O�Y��;y�!H`��,�0"O�pk��߉t�Qh b��	^q9U"O�i����@�"��P�Q��"O$�z%펞Z��x��\W10�C"O��0�O�>뼵�''@%Ӥ"O�Q����!	��P��Wb��A"O)�	;lX0}j�D/��=B!�J1d<�	z�Θ5?�YS�%Q�!�dńxg�1� �8Z7��R.µK3!��Z�wqрDZ9[%-�� W'!�$ũ	���K�nG�."��bR�2!�F�7`����W6r�8��ހ$!�J�P���uTz�0��	,ZT!��_r����B1<�Z��R#N�N�!�W<��b��߃-��D� `��z�!�$T�f����غa���R4o�T�!�$\	'?�[��)Ӑ�#FC�h3!�E4^� �	�Q.i�p�sFdJ+!�Q�,?�h'ˑ�	6hQP�&M'!�$!bF�� ��(y<Շ�{�!��
�$�l��G�P 6\r���\�!���+$�XZPo�JCj�С!S��!��τ'1����	S:H �mA��!���^��q��ǳ4v��ՎТL�!���*J��]`v�/h�H�kd��O�!��@ ��B#
-��Q!��ֶ�!�dǘ.YLș%iG�,�t<��� �!�d��\b���5�H��� �!�~�P���↱
�(��"e̓ RC�	��l��X�Q3�s`eK�u�*C�I��
UG�8ׂ�b����48C�'9�p�!A
Iv�wI�?��C�	�G��qk��u���׮�WZ�C��fb��W ��k�b(�
D�8L�C䉇s��1�v�E8<�,(�R*5��C��&<�"����?sh�M�.�FC䉰Ę�5� -QN�u"�/\�5��C�I�Vbm�e/G�c�ȅ�5/Y�Y���D,�8���Qp,Tl�Xl����C���ȓ/a�YA$�?6L ٣�̎	lx���>��k&�	%G8�lK��ɻ$��`�ȓB��u	�C��YI^����PA���`bB;Q����ǓK�ҁ��yP��j�L�.Zi�ݻ�N�7w*1��k��<Qr��d�:��4e�.���\�:͉Ŀ+��Ё�G�J�:���C�p��F�:k��ե��kO����|@���NP�w;t��!�$=��	_}�Gͻ0}Rx�!�.pQ���Q	�y�L�(�V�9�j�+l,0��
_��y��n1�:�`�;4�
��℘��ybAա1�>���&4b��$ ���y��ȡ6����G���S)Cq@���yR��	T}T-Q�З}�=���L���$&�S�Oߦ��b�$,�y���#rInU
�'��������f���$[#ԾA��� r	�t��B�ȄB � H^qA�"O��� ͨqX�Ջ�Ȕ�?��Y��"O���������$Ȟ�&���:"O� T�)0ȕ��a�<=-d�a�"O|�Rb(�;�����F�6`�u F"O�̐�J��H�@u0#[�
U6�K�O���fbL�ZY(���5P�L	H#�/���y"�5D҄�ac̴z��mQ���!�^� �𑡇�Y�*X��Z�h�^�!��R�v�����I�\qzU*#�
��!�[+!�@�s L&Y_ �¢��[��O���䚯D��HS�K�7�ȼږ&p}T�ȓ2G�-j��xR��ke�!|��u��':8�����n�4��W��G�����'���Z�"�,�nx����>�%K�'R-�X�=Ȕ�!kX�6!��I�'y(@�f��?��]pk�(��1:�'�r�`� q�P��^�.���'������̄mO�)2��J�'�)��'K`=k3�#;� ����U�^��
�'����ta��$�Р�!'ھ=sҬ"���'�,����|+�T�_�!��'Tֽ�D�� 2bGIrd�	�'%rM��ܲ���r���=���*	�'8x����20����̭=����'��4�Ľ �P�����1�Z��'q����'C�~�����&1z���'�X���o��4M��h��0H*-K�'VlYb -4C<ţ�-[m;�'h���AY*i7譓��$<(��'N������zk�yJ���2�xXj
�'M�dK�j�8�@��ӑ/:��K�'���Q��҄h�|����.^�ܲ�'r�%*�D˱+M���§A�8B���'U&i����#T{������jN�u�
�' ���E��D$�dz�F_
��'(,]`lG_���FN$]�&E�'�0�+Eo�7� %9N������y��^7�D����2߶= pb���y�G�r� �q�� �7��8C�'�(O��򤜣j�J�Y0lؕ?�H��fB� C!��B��I'J��nҰ0���%�!�D�ES�y����c��a��)V�!�_����C��/�^�ࠌ��t!�$�*i{�9�����궨�$�!��X��; ���� ��i�^�k�"O0���ՂG�(�Qʃ�*��R"O��8��ڛ0���K43v�*�"O:#%eK[*fQC��Ǆf�$I7�x��'՜���ם)��+ BK<���'�ҫ��U}|����c}�0Q��M��y�C�7)�h���
X�h��rH�y�
0�p��� ��Q@6�k����yR���p3T�[�C�X\��K �y��Q�eUܢT-�=���5E� �~2�'��]���3wqT}�ɼUv�B	�'�L�%!�	 ��ɠ'IIje����2BÆhI��2�	�"�i�1�?D����\�?Ɓ�Ȟ34I�e#��!��hO� ��D�TKҤz����vCZ�1B䉌L�pꗬ�� ����W��65��C�IM��TcX4X�M�&"V��C�I�p�$P@%QDu�����F�K�|C�I�kT�]��A.|BV��C��	(B�)� 
p+�K�u�� ��mV9�"O��)өX	�)�-Z�#��4��"O �)ӘZ�>yC������P"O� :�GN�l�KE%5u���
M��~��)�'�6���L��Zƀ��èz�d�ȓi(و���p� �Æ�A�"v���ȓP~����7�PE#��I�<���A�� B�*�2h�N��0��Ah���^A��W�܇	�d\KP
s�@Q��l�L�qE�&^��0�Ӿz^����[��1!��4'��Jd��0�Fa�ȓ$1`H�T�!3�(	�V�O�b^�ȓa�t�%+Ӟ�^�R�H��4�ȓ� ��TI^�_�)ꤋ�U8 %��!�\���ތab@ۏK5\�ȓCO���UbY�n~UI�ױ��$��G{���l��o�64h ���d*���yRE��4�}�E�H,� 7aԎ�yV�3J��`
�	lI3ƆX7�yRCYL{~%���*l��Rj	��y��#,OX��Q"Х,���A���y�ޝGF��1g|�R�l�0��m��u���b���`V �Aա;�D�ȓ�Z��P��0x���V'�؇�xQ��x4��Z�`��b�ΖA)欇�3� D���_�Q��y��芪 J͆ȓ!@ځ���R	M'T�6�@�+!\O�b�@�Q�]c���%gL hLy9��=D��۴
W i*Y!e�ߔv(#	;D�p;��DX��b�f܋{.u2#�<D�����
*4B֨W�}��)E�9D�8���N�dH�%h�0����$8D�� �ڊ	��Qa�/�&ٛ��#D��C�mU8_���8!P1d�s�'D��C��:/��B��P�<�;cF&D��@�����V\�;� s�g"D�$+�o�5in���Ԭkr�81��#D��Q,�/�
���'��I&򙱄"D�ܢ�H�5Dq��:]��EKUi D����?�����~��!B�F D�\qf�Z'TtDaZ�˔���1)r�?D�d�(��1Ŏ���bR1A�!�o?D���v  1r�����D��K�?D���wa���(أF�+3��N0D��ئ���V�BW	��E^�Ԋ�,D�$¢ըg��bQ̝W�$ZSH)D�4CPJ�[ ��b�W$�>��E�!D��B��ؾ�T9@�a��~ba�7?D��!�OD���X�O��T�!a<D�H��C��j�v���(?s��@� <D���%T���e��v�����n&D�Iq�ڹ%���B�a)��[UO%D�����9%�Pi��T�=˨3�%"D�T@pökA���KQ��d<D�P �O0f��|+C���WH:D��ʥ'�?���0�zO���+=D���I-x�JE*0
��q�S(9D�С`g�)�����х<E~!3��"D��@�AQ9�����`�w�,�3q�"D�(�D�09�� go��t
��:B�&�f�'�ҡ%R��R�R�|?.B�(>ҕ��S:RnaHC��,B�ɚz�jX�倕7s����.��4.B䉉Y������G	lC��B�"]�"B�)� �i��l���U�3�3"�ViH�"O%�&$�"?�&��㉟�d�`�z�"O�!�i2=1YZ�Oup����"O*M��c��&b�ã�-=\�!zD"O��Ɵ�)�2�s�͏6h��y�"O�<&�4},R�C��ZLY��r"O��P�@%X����U�X#Z7�t#"O<���ˑ�S��*bߴ^.B]�r"O�ɳ�J(}��g�^�t�b�d"OR0���Tw�,�C�	.Պ��"O9���WY$���9)�"���"O�\K�I������MVz����"O��@�66+:,2���� ց�"O�]+W��#C�ԫ�=d�� v"O(AY�
�j\P��
X�p;�!a"O$�q��OH�i���4���""O4��2�ڔ~��+Јߓ� -g"O���×)%J@�F�p��"O��1�"D[|����Ȫ�J}��"Oڔ�Y*)?���ƜtsrQ9&"O�@��o��bn��qe[A���j6"O*@�4N֒�,����hHrp��"Of���c�:b�>��ݫ,$���"O�d9�/ ~�P���B�$��x�"Oژ9�h��(:������4.���"O�	�㮌,f�+C���h�c"O&���F�e�Ĭ��j[�}��K�"O��j��@���b�gL�[fQ�D"O�=�lǓ	'��y���BD�}��"O8�;���\�M�=*<P`�"O�!ǎ�XL:�h��ßƠ`e"O��� �(1�,|���/�	r"O����\�dXՊ�-=����ȓ�V�i�
4C�+�-�%򐙅�z���ǂ�.�P݂�dƢftq���Dc��4Mv!�,�83�4���jU䌝>�	�Q��Kߠ`0�"OT�E�-D 	2lV��p,(c"O�1р@&��2��9¦� #"O��������i i�
u���'"O`���@�9���ݢB�tX�"O�	,]�&A����dZ�#�-W��yBK�96����b�t��t�Ȃ�y��:'DkBǒ�a���$f��y��R�	V�3���*G`@�c��ybd 97*D�JUb�""���f@���y��R)J/��3F/�#f-�e&ä�y�\9h�2��f.�? ��0BU��*�yr�:;��E0�Q�y�\�c	�*�yb��m>n��cޮ��b�ͫ�y�j�7��kgeX��ə��1�yr�PM�u��N�Ǡik��*�yF�pD�����}�X`��ۖ�yB�Ҙ�bL����|M��e+H��yr��"���c�s���%$[��y�'K�S�,���9o����Ɯ�y��a���Pi��d�j��®Q �yR�5N��G��Ҽ	ӌ��y�C<b�l�r�,���IWL�C��B�I+lq�W�E
 U��+�
�LB�ɪ~���ðh�S�Xa�a�0B�I;4��'W3ڈ��R؄{tB�	-j	"0CƎ�8� ���D��C�I;"x"���.z��Xp�o�/m��C�)� �ucg��4sذ����}Zv���"O�<sp�A�E�q`�.^�O.G"O�I�w�+P4=�nA6@M��"O8Q4*�/
d�{6o� �h{p"O�p�rg�) Y�H+Uc���"Oa� �J"Z�5�m���s�"O��
�m��,�Q�/\O���Y""Op���6It���q"�,g"OΌ)F	O����1L]�M��y�E"O��s��1\� z�떡(T� "O� �@ϵ8Fl��@ZMx0ES5"O
07��??��� i?`[�D�"ObX��P��l��d⍉Z� ��"O�8!gj(zG�e��ɤ1���j0"O�]�G]N���{�*T�VVe �"O�UH�'/b�&�Z�<o0K�"O�dk^r�@p�aA.\X��y�
Ѭ�yB�ǿ
���H�U��Y%�3�yB�[�[/d9��	�P�<9aT��y��(U��9qn �Wt����%�y�"�V4�]�vaC9損"-ʟ�y�'G6F����N& f�R�yB++wF���gG�@�p%��C��y2EՊ:Sґ@�=7豲��'�y�aC�|��
e��	F��q����y����e� ��b��8m��PN�y�H
#��W$�85r�dB� �yR�نh���uBU�-�����?�y��['��
�I��p�1�
��y��&D6� �б�p)�����y§Q
!R�`��Ǖ6h{p���y���P�(m`�ǔ=h�ؐ�\��y�
�>-̎����-P��)�	2�y�Z�$	��G�#��Z��4�y2Ó<�|]1tMh(��$ր�y�K=g}�D�w��"mX���.�y��
�C
�Af�;]�`r�h�6�y"���= .,��
"2�&��F��y��ؐMy��@7`�;w��2/W�y�i ��q'NL&�r�i�`�1�y�N��"�S	:
t0'�?�y���eU"d��	*�Z�'��$�y�_D�Pd��l9U��Th提��y2��q��)�� PP/J,y��ؙ�yBi�qj�혦3���%�<��d�ѡ,���i[0"帐�ȓz�@uH%I��� ��fV{�ʈ�ȓ?d�*�i��]| ����u[���ȓ:�NɁ� ��8{'�������=�"ܺ��Z��<#q
�&F��ņ�pG$A �M��LbN�j�h"�D���}�����B׹(Kp�@��E�X4���Jp2sM�8�1Hw�ǜ��Q�ȓ4��ɚ�l���ct��i�nE���p��G�3G%%��˪#p��ȓ�|īT��g��mh��0@f̆ȓ#����F;LD�Bo�(%�*؆�P\@�U�Cg��x�J� ډ��\�,�)��H�QXP�3����$����  �p� �QV�ȓ^�ex���2ZGx���Y�2��]�ȓg�65
̖�a��ZE�âv���-%)Yuj�ha�9���	0�R��ȓˆ�3i`�1E���Ї�S�? �p�/��EZ<I8&Y�t-�Ęd"O�-���6}J��V�D��R"ON���E	�܅���L�R<��"O@Z`I�u�N�S  μ7X��"O��i��9Worx�&.?�narw"O�<�'
/V���-��3�IQ%"O�y�ܼZN,��lJVa� �"O(L	4eM�EI�a�ҋ�>2��""O��r2/�."h��l�Z2X��"O��12Ę�F�\�Ӥ�;*JUJ�"O�E���؋@~*t1�,�R��&"Ot9�&��g		��듿s�� �"O8�Ŏ@����`�������"O.R1Ny��@(�HH&,:h�"OJ�����A��غG"�u�G"O�{�E�Y�$=9�i� �F ��"O��tcN'\�}X���4Kz8�"O�T�sF7e�$tx�C�O/2W�y"K�3o���&"ӅW��9��ǈ��y�ЄV�1����H�v�p ��y"� 	$(���#P���j`!�,�y��B�p�6��o�v+��1�����y�ꌂmd�)H�h�	�ŧ��y�	Xj����q�O�d����@Qx!�dZ:`�(H�,��	v�Jd�0%�!򄘲w8:lr�	>)�yٽe(!�6Y��b��{r��
o!�Đ�K_RA���S\�� �*�P!��%1���G�ƈL�DE3ժ���!�D�U�=��\�=at੃I��d�!�i1Z�sU�3ALƽy��-4�!�$̴%�ȐQ����"g�U�$і�!�����EC�T�|����Ӽy�!�D��@y����@�tcP�!�׏Z`�� c�!V�ȱ�!�_9�!���1��!�
�x�<�4ߒO !�×;�XP�F(�x���{GD�o!�D�'R:��P�����ĉ���%!�Y��@i(��r{����/�?^�!�Dһsuy���G$hl�)�Wo���!�A�1�V�ae��(uZ��(�Yw�!��W�Ri�0��4Ii�d��F h�!�ՆO��亱#�=NB��3�KS=�!�$܌.�Ԩy���:���Dm	$�!���O�V��E"�)
�|�c�L��?�!�D�:�p�ʡPy6]aWM �!���h�����ˏ�$I#b���!�$�]���B��-}�b��yw!�DʭG��$���</c��P4j!���L��(W

5��-�@��.g[!�D]�0��.%;X&�����>!�	B���I 7)��7`҉(\!���;K��@����!@��w�W�1�!�دQI��C��F�plˑ�ؙK�!�d 	�h)a��X,3�4x�b��3_�!��A�1��A��,�y����(y�!�ėo��A��!X���� ��p�!�D�>�p]�Sl	#0p��C'��X�!�9�t��U$F>A��,ɐ[�@G!�ą�7�X��p�Lks�,JN7A!�$�Pi�to�un
YW�Z&x�!�䖌"{�!k�M� MY81��̯o�!򤜜ֲy� ��/�H����x�!�$ݠn�8���X�^=K�j/3�!�� �E�ʖ��9R���d/���"O^�@n�
.<d��s�(F�)B"O���� �)lzػ���M荳�"O�D���G�(j��+���3"OP�g��L��	��`*B�R"O�E��Gn+@
~ڲ��7�;�y2��*IsjD�g���%[�k�zC�ɽIˊTx��Ϭv)H���"�?RC�	4U��H"�'�J�j�b�;HC�	gwd{C;��p3�"�qC�	�d�'�A>l��ʁ�.��B�ɺNX
�QO�O�X(��P��B�I�4ʰ���LX^� ��!{�B�	�TH�2�Ո;�T�HG�
:C䉻P����W�O����J�)K(C�Ɍ8jq��%M�����A	>T�B�ɱ	c<,�7�U�WAV!����}*B��?:q`�C�A< Hm���Mm�C�I3jY�ɡ�I[u
MYg�]B;ZB�I������4������+K�PB�	��T� ã�Qz�UA�lX�h
.B��!ZF4�����-(AB�Z�"B�	�!y,q�/�
������6F��C��,7!8����E��O��jC�	)Nx+���gBT��Pi[)
C�	�	�>(�G-U�tX��|��B�ɛ"��$"�(�����U��k�'X����L�i�bCPKE.a"�٢
�'j�;��
\�3�G�vX-��'j��q�@E@Z�E���	#��q�'�1p��(E�<P
c�v����'�(:rf�A�P�Q'Σh���'0��RoW1� ��f�G-b�!	�'�Ri(g��&5��*�Yt�	�'���*����/	�H�����'�vYj��C�!���+�X����
�'V�� �!ڍs�4�L��S�-�'@t%:�R�D,��EFԺy��y
�'~*�9�C� �rm*&��'�����'7l�����%D*�	#��N�b��'�bDٰ��4fD����|�2�R�'J���$30�p�$�IqԄ��'�
d�f�D�(~�T�s!�	i��@��'���� �/��p�c�"hNP��'��œ��R/֌ٸ�`�sm� ��']����W<:ŎM1eAi����	�'t�X�L ��cH�]S QY	�'��C�n[�J�9"����*
�'אl����}Bd�!��'2,�A�'h�r�ʧV��Ҧ��l��Z�'�҅�5��&!+X�6ƾ">��
�'�f���B�J5��s�	����@N�<�`K�6^.&\��ޮ-��B-TA�<��ʀ2)�Bq@'J��?�|p��}�<QX8mJUOнQ�6qJc��=Bч�-��L�B����5 (��d��B�I��&�FR���� k�����谢p��	zv��6�<J 0�ȓ�
E"%l�� ���5J|L����\�DR�+q���ʒ%v��ȓ$�|�t+@tԄ�c�[$w֐���5.�	r�؄TIhMZ�ˋ"o� �z�7��>4���N̤e��ȓsT����KKIBl�r!�.�0��S�? �sA1h�l͛�ϐ�sy�Txv"O.h����>�JMp��
�-x^��"O��CG.�8N7~4� Ōl���u"OZ QHݖj�]RV&P�R�PT"O|Mr��'<�P�A�3X>EIv"O�8"c�ߍ6J&m���_&*�)�P"ORŻ�&�6d:E��M6}4a�d"O�Pb�îzĊ,�֮"VD�`R"O��0ҎЂ[b&<����;=Ѵ��P"O.�q7`�S�J8(ፐT�*`��"OL5�π�`�m��	�;����A"O\�q�ؼ/6^m�	��!���S"O�1���T-ko�� çK_+:�w"O cώ".� m��9�!�"O���rm�e���0�W�k�2���"O���'�N�ATy���<q�4Q`t"O�1¢�6�7�Ϯg��q3�:D��� �4/���C�ϋQ���,D�0�t.	%o�1	�W�f	p"G&D�L��MR�6�mS��8)�I>D���W([oI��ʤA=+�x�C!D�L
��U6/,�4C�뛍`ܴÔ/-D��QDk[�;w�|����z���AK)D��s� _�f$���@��Rhu�#D�8"B������I �^�衮"D�����hT�e��	/�@���!D��jǁ��MȒ��f���X)�ͫ& 3D�T8
��T@��H&ۀ��(>D��ړ,�S�XQ�+�T�V�H� 7D����$^�|��$e�j�BТF*D�p9��<��]
�a�d� <�Fg:D�R�B�3��1�N�"�HA�@9D�Ă�l�8b��m�t�O��ph#3�)D���F�
�ϴ�H3%L�D�N,��A'D���m�7ɾ9Q��/���R @*D�H
��S�,��p3���R��Y�(D�L)LѦs�*P�tC�U���&D�(k��Q�z�#V;7�]�7!D����A�K��=2�]3tqxѨ�#D�,`G`W�m��������Viq4J"D�t2�cߵR�V9C���~|��1L$D�ԉg\�M���C'�B�v�q�).D��w������+v�:-9�(D�,
�烤&���5B��\�N-h7�&D��´hDS�`��`��F�&�@,%D���A�X9�,5RV(^�e^m���5D��;H�3~��
� �j���7`0D��A��S� 갍��蝖;��u�)D� B�MS0X����YaB��J'D� ��-�=);(h4�iԶh�d!D��J!!U;���A��"U�؉D%D���R+V�<$��c��gX�1-#D���$HD�y��])�'�$Z�v�	��#D���S�
	�r�`�� �����#D�xQ�fa@�`Td��@�h��B�	�B��a��"�`]L�yе.��B�I]0c��/�)Z��I�?"�B�	pTj���8&8�Cf!��&`BB��%?� M�����𠹣��B�	/�'�s`А�S�љsɢC�� u�Jੀ�1-��T@��?Z��C��<B_�U��k�>#���u/�tALC�I�mC�@��"V뮈�V���t�"C�	�wh{ѠD8(��8%d� �C�)� B���h��!2DE�`>\��"O`�D,Z�P�F}�&�
�H9F<i5"O@�����:��\+�	Z�A(�b"O�7��5<��+�Ȋ�U�\�S"O��;�J��j��Ģ҅��,^��Q"OR\��A�+�h�4�Q��,��%"O��	�JS�F$*�r$@�O��I"O�$�R��=��(�a�6.��Q"O"u���Q�N��Iȴ���.�Z�b�"O8�ː�W";�j=�G��^��2�"O*�r�	�=j�� �2}�i�4"O�H�D/�d�HO��w�c�"O��qG��6ҀY��� |%g"OP���M�w~D�M�3�d��"O���D׳?��"�këA�&�s�"O �� ��Tv�i�vJ��5�j�[�"O�䙒$Y?k�d#�� (�����"ODmБ� �'�z�a�Dߝp¦���"O�p��I�L�qQ��!�X�I�"O��yS#٬�0$���0 ��"Od՛'-��ځ�F+���h���"O�P
$��"[-z�{#+Q�a�${�"OP$���Ȗ~&�J�i��y�ZL��"ONX�_wq�I"T)�;1�8��"O��1�� �z��h�.,�B���'�h�" �'��0�$ȏK�"���'�9���!C�|]�"�\�X0R�@�'��R�&�ô|9BR#�z̠�'}�h���X�cq�=Ca%�&m�
�'�)#��I�:��3�Ekq�t�	�'*(YW��^�ZhJ��]>f���Q�'j���Cl�(}�h��p���B�'Fjt)W�ɜ�욂c��cF<��'�ҹBR�����R(O�E�,�@�'|Y�T��	Vt�-D s�:%��'���8f�>Y�l<�����:����'sTqcn�%HN[��N�>njQ�	�'���J�!
?͞�U,ҧ1��k	�'Ĥ�A���8�ni1$�9��	�'H䄊� �z��S�/-���'�nxn0Y���KC�sw�u�'T���DF^��c&���q}L�
�'�����CD<pnXkEG6l�@�r�'B�t�Ӫk�����5�)�'QMiC�C�#���Nd��Ub�'�.<xv�B4B�����U�`8 �;�'��`�
]
`�ƫ� V�Z ��'��ٱ�̊�Hi��CC�Q��y��'2�����*7�M`�.P'Ķ��ʓh>�A�'������\���D�ȓ(y~!9aO�#"=*q@!����g�J��q�S�Prs�k�L\��W:�m�K@7F/�ţ��Y�+�هȓ@ �i�H��9)`$�U���P��h�ȓ\�0�Ah��!4H]����ȓqNh3")�3ry,���T;(���U�1��]"ȉ�Sn�&F�L��]#D���E��=Xz�.ɹN�$��/wJ��S
F�&P��We�9_w�Շ�>�BXI5���Y��	�!N�4]�ćȓy�X�"d䟑2�0)4L����"O2HP�D��]���CHR.Q�2��"O�}�&��,�-I@��rQ�"O,e�&�ƾ���ӡ\A��3�"O� �IAO�]�a�f�D'3I*�"OFqcp$L"L	���ډ^1�8��"O��:4�H�5izux�d��O�A��"OPX��e�ah)�6"$QH�U�v"O���0%�W��`��#�<=�p�"O�X�"B��pt�H> <�z�"O���f��L���Q��0�"OBq�p+������1�J���"O��8�
�.(��d�T+F2�h�Jb"O�\��`�0��*�_��Z(��"O��Zm��+i&,{娀�(��<�"O )s��5y�@|��h;f@��r"Oz�9Di	<���p!iR�V�" �"O�K�A��-@���c����"O�I�C睛Hm�U�JNj�J��"OlD��ED�,N�	 
Ԓy~��""O��K��T	ؕ���_-uv�y#"Ol,
�AP�V�iID,�(y04"O�i�vg����B3��u#J���"O8�2D��F��)�W�o�����"O2[�P�d�s+�.N��A+B"O�ɨ`AZM��c�i@ r���"O9sQ�< ��dI�	�7�l��3"OJdad#�o{\h�I��ve`�"O��[W��V�,2�	Ÿ`φ5��"O��'P�^��P�苓Vͪ$"r"O4sp��� ��5aHʧC�~|s"O&����v]0-�%'�)6*��%"O�Ј��t�4a��=�R�3"O&�����+��x `���š�"O옻�O#Cwt��tIH�H�
l��"O���U�w�X�W��d���xf"OLx ��:J��0֠���Đ�"O������/: ��eBT�9�p!V"O��C�jN��t�����;�*���"O���#ȃ�a
j�xN�=iފ�"u"O��uΈ�rJ�@���mh*���"O�@˓È�M��$!F�ߚCW�|�"O�X���Z��Pl�`��	Vf���"OHmx�m-:�&� E'
S���e"OH�AG�LY%"W��E�9�3"O^]{�J�+M�X�ϛ AF� IB"Ol�%d�78�E;�HxC`�a�"OB���ı�pk�-O1:|�Z3"O"x�!l��/��Mj��T�#B"O(��W�ľy%�5��&W��
x:"O@I8��$z1��@�rB(�y�"O40:#�[�+�2�- �f�+"OT�p���D��(A݆$
�͡$"O(�Sk��g�.[�kT[�D�z!"Oĉ ��Y i�1D����"O��,ZPv��%N� ��"O��s���	��ǘr����"O��Z�$�F�Ω)V��U��P�"O:d�ebU�1[��߯svF<)P"O�0ا�A�?���x4��wrJ�)f"OF�c��K&}�4��̅�,b��"O�җ!�$)��IA�k�a�p
�"O�PŅoc�#
�X4Ԣ�"OT}�� O��hi�*�?M=T�ɦ"O�Hi�I�"�,����/V�z2"Of��C$$EL��  �a�H,��"O��1C
K���󉊃Z�,4k�"Of8��#�{^�4��;��H"O� �2�BՎ (�ؕ���n \pqU"O
� �,Q.|`р`["\p�"O^|�DݢT���.G(Y8\`"O&(j��ZF09�M֮V*�ty"O��*5
�16�(�WlL<��EZf"ON`� !B�,�fƚ5���Iw"O�"(�#=�:������wTL5�!"O0�@b�<�ؐ��H<oNv�"O�Q �o�k��M���FԘiC�"O���æ�98�^)��oD)�>5I "O�5���<g'peH1`ω]���!"O^]h7犼	D�9@.�va��jg"O�����-%� �R�BU6���"O�P"�K*U���җ�ߍk/AȆ"O��!�jD�s�h��, ?;2N�!!"Obh+4!�z�Tl����3��C "O�t١�Ccv��F�_F�2"O@��p#���$���'F�E	�"O��q�K��*�숣WgR�Viĭ��"O���aaQ�p�0,��P/`�\c�"O��B2:h��N4C��3"O�ِv 
k�h�
Q!����S"O�����t���2���3��I�"O�!���*~s�����2~Ƶ��"O��!�92Y�ț�m\1�P%��"O�M@�`��BBex�l�Zb,��3"O����V����3�\�r2
	��"O�*6��.Sz��W�U�A�"O~`��O�H�d=s�JI�4��"O��P� :9qL
BɁ�V�|�"O*S��$*I������>A��"OnH��FD�?4�ȧ �.,����a"Oܽ�dҥ'6���v�B�x�r���"O�`��.X�/TJlX�nD�]s``�"OPPJ��A�kg28�$�t�S�"Ozie
�%jb��1��mkh%H"O(���׃;��;�k]&Ne�}bE"O�+�J"0J�\ri̳.Zv��"O�M�P��88��"r���ñ"OV�y���gN�\X� K�o�,��"O�up�G�P/6�;��QO��b "O�\@���+Y;:�24�_ d��q�R"O�@���)ߚ��t�@L�JQIc"O���m���� (4$K��2�"O
EuN	�;�ޔ�㕧k��:�"O�P�f ��ږ6D�7W�A�&D����nW-J��㲤ܩG^:лƫ D��:A٫N��[�F�f t%82+=D�<�am*�ʅ����2F�%��=D��q�*�{�	VȂ�$u��'�0D���!n]�\;��"䇁�7��|��B0D�i���)�`�m�.&舒s�0D�<ӄ)�W��lh@!	9X��)�+D�x���N�`� ��B�R��Ҵ/D�`r�
��T|�,{G(�l�Ȩ㇬+D�4��H�,��m��2�8���>D��Z��@��XSꘪh3, �=D�|#� �{����V�8�"��Q�:D��3�e�*�*�C���e|�0�$D����)U/�~c�5CN�z6	!D��v��-��(�iI�y�X�s#)D�d�l��B�4�G�G�`�9��&D����Ӿw4��:m�!���Q�	 D���,���J�'���|@0m?D�� �,���n�4��5����,��"O"ip� 	;ˆ @���}�R�S"O����D9���� Ȉ4"���"O�Ԓ�GL&r��f�Y�)�P���"O �(�DP8X^����Ԋc�.0�"O0�	��VL��-�6�˝/k�x��"O�D���$ic��"tm]�-�*��"O*�AAKʝ��-L�v����3"O�I�⢟"s�ڙPuؐlI
�"O$L�Bo�.^Xأ�K�3Cm���"ODL2@�>��	����d���U"O �A�K��uU���'L�$oOp�j�"OX��ƅ);��!��u�L�1p"O����94�aY k��xs0-�"OR��WḺTY��!I�Or�r�"O��T˚7u�(qjDF�	wT�ȑ�"O֜1�D\����@営VB&D�R"Oi��_x�����X6/>.="O$��cK�`�6e2���I�X��"O���ׯS�w�����y��	�"OZd��!�6�=��+�1�~�5"O+�?�r}�񊁷�$d��"O���f嘆�th����E��Dag"O0L{&^�X;�H�Ed��C�e��"Ol����=�x1�5H� \Y"OZH�K_�{rP��c�0m����%"O�-۱!�0���0�L�6�Dy�"O� 1�fӳ@�`d2�I�)$s�%X�"OZ��.g�pyY@�!xp� ��"O�� iH�
���n"pg&]��"O��ʀZ��p��P���3�"O:Ƞ'`�rMZ��H�V��y�"O�Q�&�ʬ>�Je� NK~~����"OZ�����1B%�q�2j�"Pv4}�t"ON񨦄��V�>���k�Tx�aY�"O�=v���#��A0l�A�"O������[�&����?�@
"OX��I�G��q�2�&c5"O��(Q�E�UҨ�&�C/����"Op�l鍗 T!����vZ| 9�"O0l��ł�{ڌH4��e4��K�"O�j% �3sK����Ӻu$l�à"O��R��Y�s`$���3!��0�"O�Q0���%�0�kT�Իu�'"OP8��-�Q(��K�_�r�"O��I"Hs7���"�׸q��Y�"O��XU�h�x w�ltR�"O��ðɔ#P��%�k��h� "O� 0��̗{V��k�,���0��"O�M�TF̬ҊS��8�̡"O�#V7ܪ|��)��m�����"O4�hfOĐ))��p�� ]0�9�"O�K��<\5�UC�Mq�D{�"O��Ue^@�9��*X:L�^�#�"O ��"���k�z0�G"O�)aC ���k��
HX�"O\pѡ	�h�\-����2G�� A�"O�In҉vS��8�ʲ3�����"O�W���e6n�{#dBx��Z4"OPsAL�(t����]ɜ��G"O��`I���܁��NE�4|�"O$A��(�TX���uM�%{�'"O�0��ą>*+�XJ����f��"O:x���/l�p0NH;0�����"O� \�k3�wr$Xْ�*p+�D"O�m{��L,oz�m���"G`"O����֕F�2��C�^�( ��ɓ"O���׌E�A<���b�ް
����G"O@\�e�Agr�1�$	����c"O�(�� ]�X&t�d�*�,l1t"O�%#F�0�J�i�ME/��:5"O�����-����F�O.dM�T"O�У�oI+}$$���FX'L�z4"O��P1��j9�gŞ�:��"O�u24�V�)���̟i꘍��"O�����ަa��P3�ԡ�����"O�q�r�,}���Y���?9���� "Ot��ӢU6�}@�Hwڲ��"O�m�ׯN�Dr�i�6��	#H��u"O6���B�p���V�ĵ7>2\��"O��yU˧S�(��K�$�E7"Ox�[�S�(�%Y�9�\��"O���	�$]�(�!�($�4�a@"O�� ��/�~����)�¡��"O��U�ͰF'���!��R6"h�R"O�Ƀ䂟�z�X�@R�~;Ь0"O��*��S3)z�a�`[�)�	�!"O�	k/K�Bנ���R
B$2<a�"O y�%�'+X8�ZI0����Vh�<I�DV7z��#ʡdn<�!��Z�<��+O�er�*!IݜX�����o�Y�<��,ʊD�Ɔ�/v-���@@�<������ya&0�r�`��<Y�ƹ4'�ȶB®OS8M���Bt�<�iE�&���.6�A@��Yl�<y���EbP�;v��q'��;EO�m�<�Q٤H�aJ���,s}��+�P�<1�OF31Yꋁ; ���eYJ�<D�j��B���1�D%0cJ�I�<I�d͸ղ]�!�T�}C@@�v�{�<�p&Q�7���q�J�&((a��s�<���L�$MjP�.ެC72��UY�<ل I�u�8����Q�<�ܬ��'_W�<��
�ht��¢��@���SW��R�<!�9|�X䙤��(�f���%EP�<9�,oM� b�eƪR�.���B�<a#$P�c��,$�� a���V�O@�<Q�l��`KU!A�kVɸjN~�<��ٞk�2hQQ"�$���Bj�E�<��i�"5�^墵��U�>PH1��G�<��ՏU}��s�>>����0�E�<QT �� �xA��&��V4"�2gPD�<��	I�}���F*H1[�Y+�	�z�<�M���Lc�F�2%��|9��y�<��n
pnܱI ���*�)yT�@�<9��N�O�l��-@}��M��Ff�<i��P�� d�9]�8���`�a�<��,�2j�L���lx��FGE�<QV�&S��-�+�5p\4��'B[�<Ѧ��Sj��q�@�o���2�.]�<���D����Y,y'��%��r�<!��:<�l�`�U�S�x���K@C�<ɴ�̊v��B���r.����[X�<)�gF�:%v���Hݛ|�B�($Ǝz�<!*K.f�����j$40�I K�<!��J�[=x	%j��qF�&��E�<i��ԩ���`퉭y�&���	A�<�Q#�w���b�42�|�Qm�z�<� L�b ��>h]8uv��g�p�"O��7'm�Ry3���6I�dm��"O���uK�+�=��n$+�&��"OR5hQ~��ِ�n[g�R #�"Oސ��H��h��BM@� �~�c"OƤ�!j�+���4�;;�"O�$j%˗�W�� ��g�ƴd"O�q���I96��I3�K&����t"O��
2/�!��Q����2o)�]��"O�%B�Đ/����rDLuP1��"OR �D�У�������b�3A"O��[s�I�H{��P� ��"O�)���L�[�hҶ!��D&6�[�"O���3f%q�� �B�lj&0:"O�UY֊�].
�� �+��\T"O����P/U�J���� ����C"O`�ї�Η4d���L[�Cw9�F"O`�Q���:fb��J뗆=_Ʃ��"OB˱�[�aꨡ r�l(���"O:���i9d��ȃ�!XI�g"O�l1��K�}'f��W�"9X0k�"Or0Q刯Cd�)��5v���U"O�5��*S��h�'��t�Vx!�"O*��M�m��v%y�|!!�"O DN�9+�XI��L�'�̥�$"O��jE#�	���@qa�4p�C�'�ܡ��k�4$�����A"/�d���'Np󐬋��<��W���0��)h	�'O�MU̃"�ncv��:(����'2,�zֈ��<-X ���'OK�O�<ɰOL9f�	���'�h�0qk�M�<I'�� D�*��be��,���0�ZM�<�A�Ū`��uze`�>f�@x&��~�<�f�����ǆѶnR�t��n�e�<	g� ��]se�ܗhCf�b�<9uGU�)}��(�,[Nl䜸�l_�<I�F�M�bL�t�A��%����a�<a���%t���NJM+Va�#RW�<iӦ�7M�@Ȕ��Ι���y�<��)�s�*h�Ώ��Z��i�<��M�=\Ӧ�����r�J��d�<Q�K�-A4�,3!��1W�4U���h�<�&�/;=�ST�̫�<�R�eZ[�<�N�:F�	B�3$����#�X�<��.�*RY�C�5Oj8)8u-p�<���@�N�"��R��3ze9����Q�<)�n?��K�T.t�T�@+J�<Y�cܠ" R��"̈́�U,8R���`�<�u(��,dUa1�:<Rԁ���t�<1�ԘW&��N2�,�'L�m�<!4e2�*�Z���2x���ae�<�F�	�K���8nd�r�Ca�<A�s0:�K1#=Ҹ1#[�<��Ʌ+�{�dM$T�����[X�<9Ӧ��C��S2g�m�T�e��W�<���6&}x=I��M�Xph��J�<q��0h`����"9�.�s2�B�<9����^���.T%z��{6��<�'i��=�F�2@�p)���f�Z|�<��e�26���T�K#x$ib�s�<iB_�PY I*h�z(�W*Nl�<��.� bK��B����l��D�P�<��ѰA��¡�<7���P�I�<�ì�P)<ݱs�8X����ƫz�<� ���
a��)�D��#}�tA�"OFLz��T�@��q;0!ߨik���"O�I���G(h,Z=Y6�Dq���"O�M�3i3u�J��!�ӄ����"O�%�T��7j��l]8�^@� "O|����j�-����<6��D �"O�Py��RH�Sd)^����4"O�U��i�L�aB�ٴN��u�"O�`&B�ut�r&G>q�X�"O�X�i`~��%�}�>�sE"O��{�.�p�����d,�Py�1"O�hX� [&�Y�g��J�6�cd"O��9t��4� IR�?k�lr�"O��Aμ"ؠrCgE�hy�H"O��y��U�r�T`�b&ڂv��Ũ�"O������Q���Bv�2��B"O�Eq����n�D�*`�G�*�!�"O����R,L���cՆ�)\��!p�"O���%E���0e@��z1R�"O<��@-ĹxH��Ӷ�"b�����"O@II�ж\ٶ� �%�j`�"1"Ox�p��,dB��pO�}���s'"O��K��a�* ���C5�T�(�"O��5�J��ԁ��(� dە"O�$�d���RD�	�v�]�z���aT"O��D��x���0�+%��(q"O �R���10P[U)��8v�D,�y"i
��õ
^C�4t�C-���y����x2r�3l�n��@���y��8�2j�g�*�b�!�0�ybg�]U���G��*j�lA�i�	�ybM�8H�XI0��.��D��K�y��*E/�P���!��Õ)Ĺ�y��P�|�N0J����j�Y�6.��y�O	zS������D����y�БL09���Ӎo���3j�y���R�6%J�aU~X�E�+�y�aǏ����灙yc�=�!�"�yb�ٸS�h��A�;&�Tp3���yB#0"�Y�CL J��K���y2��=	V�*	!m����&X)�yBf1������r,�٩�.�=�yҨJKP�ya�Y�B�6�Z&�޵�y�O�g�d��D4|�`Kb��y��A�10��1���(�&yCƥΔ�y�j#2�R���
R�S�h��i�8�y��̞s��aS@mZ�F;���fR8�y2�_�kgri�bB�0�����i���yr�	*�΄z
�72Dư�5O5�yr��x�l�hSI�9�!qu$G�yb��-'���C�/I�;�B�t����yrI�ޘI�K&0�������y"o\9v-I���˥T�\9���
��y�휧�x(#d�N�Nu(53Q�yrf�[Ѻ�0�gL�LmJ���dՖ�y��^
��Y�Q@���� o�yb��|QLE
�'��`�b��y2EE4L(�y��s�H+a��
�y��Е��P�Hv9bl������y�f��
���C��,B���C�����y2�U�H�B��l�&�֐�7�F��y�$��"����<r���y�ʼq����h��b���g� �yB�Hm�<ra�+{mT��!¶�y
� ���6��X��	7/�T�0�"OT`�%Ɗ G�ܵ� Nܹr�dM��"O.	�a�gN���	����"O�%�I̛.���cP��nژ��f"Olxc�T39���z�F�+5�Ơ�F"O��B�`� ,Y�}�&�~�4 D"Oxy���ġR��x�Sz�8T�&"Oh�!#��D�QP�� a� �K"O�M��
���	����+F��0R"O�yp ���X�W/H�b��"O�Ș`�]�J+>�0��'<�k�"O�#���ݦi0��=A:�ݨ�"O����� 	e�����sV�]�"O��;1o^�EL�#j��IY�Ly`"O�(Z��A~s�Q�2���F�� "O�p�Q�5в-������֦!�$G�@phZB`B'�a�.Y�H!��M�$�hQ��ޢw�$z�B��!���!.$Qa.�R5�� ��L�8�!�$\9n�da���~����b��<�!�d�o����E/ ~�� 
��!�d��VN�1�(�{��c����!�_X�*	Ku�]9Z�jB�bt!�DD-%.ǅ��2���T��-v!��Z$���d[�u���&�L<[!�$T�	$��rl � ���%�*U!��Ќ:�)�5��70�l<��M@E!��t���#��~�ĐY�&۰T�!�D�qV�Ѓg��#S�̠c'#2!�_)o$��*��C�8J���`͑�E!�D�2��Aa��:1&�1W�=-�!�䚒3`�D���ʥp"��y'
 5�!�<C�-� �1;�՚��'IX!��%p��,
 �X%���Y�hE�d!�{���[�o]�f�Ą�(�4V!�D�gƤ��#9Y�p���=D!��%I8~1�Q���`�[Vn +.&!�ͅB��HK�Z�L�U!�ě�V���#�D\�Ku�N)�!�\��dc�&�:8��r���!��
����ӛsj8�!�$,!�D�Fd.i�H�U�^�1��10�!�d��
�ࢧ�ثx�R�OB!'�!��+� l����{���CĖX[!�32���Zd�� �L-!��30!�+m�:�`ä�!dҝ�G  7Q+!�Q�S���6�E��[��a{���6\h~A�E��R�H���J!�$�.�$�z�LU!U��Pj�(!�DC�.z,i�l�;:��ai��v��~�^���@9ѨP����9C���P��;ʓ��<	�k�-,�n�1�-��*R�a�u�<��D�r��8
���4e��aH�<�F)K�*;���゛LSn��e�C�	ןd��	 �1�䄟x�� �Ö;IC�I�(�!��������D��
b$#<)���?���,d��IC�j�����0D�4�$ćho6��&٠B��d$/D�$�rDʛG<}��g�:EcP��	+D�ċP/�?8W"�B�o�KRB9�4�<D���`<=P�qѰ��M$�C�{��C�	|?��{�m�j����b�1r#�͐��y�!_�Z�����h�j(�H{t�W���"�S��|��K$���Q1Ǟ4�<��E��y
� b4�1�9y�tj�
�!�Ԝ�""Oΰ���Q�fܔ�W���i9��	T�OO9�te޿�2ԩVhJ	~��)�:O�7�?�O� ����W�R�ĉڣ"O�ܩ#*͏Yu؁ !Žm񑅹i\�'�`�����E�P4Y!�9#�TH�'��B��r[F�2�f5r��H�'�\�P��7E\�"�)��- ����'��b�oS�%�ܑ׫ޟy���'@8�K�NL	X@�� p爵r4~�;�'���a� F��Q''ɨ�,}՚�8�'����Y��� �2;��
f�W��
G)2D��)CG�8}��ِ�}��/D�<a�W� ������؎����*.\O�b�� u�ύ@�RH:�Mđ,��qi�g'D�0��Q��M!�$��OQt���8��hO��¸�cL̂^�} �nU�,�hC�ɜ6<�;Agʹ2��� c�Fp��dE{J?i9E�׵|�t�u�	�!"�raG*D�{1nޝH�
���Ƅt1U���Gm�'@T�D�,O��YgŊe � �AF2jv�� ��"��?���:杒�@VM��3�Ǝ�D�~\��j�2}z��L6a}ܱC��M9\6�ԇ�8n��1��Qx\���(SX=���ȓ5���"�܀��ɒ� �#[�B0Gxb�>�M~Z�'���a��$5FNةT ��O��"-O^���*�h-�g�<'v�q1Fڀ:�	C�'��6�	MsPS�/G�+���@C�%:�6B�	�\�P�����5�����wr�	���?я��\� �"R��Ӗ x�K�p�!�@$@l�̛�"�h�\��eL�k�!���O�Ya%�T���ӡɛuO�'��@�<�a�=_@Є�N�PGAK�< �͂}*T '֧'/I8w$�I�< ���9���N����*D�'�ў�r�'���R7
E&d�JL�"cB	Q1�0K>����F�!��9�*L��`q��+N!�Z�3��O�i��O:8�!���[��B�䝧{��58a��k���=�O(�HT ?(�""��5��<�"OƘ�"-T5NA����=e�Hyq�"O�b@Œ�7��(C��2GD��ѳ"O\)�b�A�,�������)1�406�$,�S��*
fܫp��:U(8(��:��B�	�o����)BY&(���^�*�PC�	/x6N�fh܈.Rx�_�q�
C䉓aĊ�mۘs�>� ቉�o�B�	Kj�\�@M�u{b����"c�B�ɚ93�����X���i#�p�j��D&�_��1daK�F�y�Q�G�WF:$���|,�P "?����M+q�R�ȓJHa�f�V�y(���e��;�t��e]��k�!�(d��ي��$1>�Γ��?	��Z}���c-(!WD��1,�i}�'��2��O4[�h`�w.%�����'X�Azd���_�y{W���� `��'ӄ4q��n��[bK?s\JqO�̱`CZ#�XY��BX��<e��O�ذ"H]D�\YZv�I���q�!�Q|�<�d�\�F�tH�ȗ4ռ�V*ZO�'��x���}wd�B¢ب!�RU8�'�M�	�'�r��B�p��%�d�> �FUY��<,O&X �J�
$�e���+(�x�"O(pidu����'�~L!Ӓ"O� d�itM�:9��9k��Vf�Rl�4�	h̓��O�j9c�Z�u��} &��8t���Q�'�eCrH�;� k�4q|���ӓ��'��X���Y����n)`0y�'�P���Ǌ5${A�ؐa��`�'�l�(�
%Z�^i@���e��`S
�'���C'��^��3�	�Y�,�H>������!�V�K +!��;��i�!��77�������`�A��_�4�!�$�$Z�n��W��"C���9�ŉ+ps!��#`�0AG�(<�V�+Ez!�䈘N~Vi"�Z?�,X �4y!��v��' �9X���6��$w!�.�v hg�ĲqG$Dc�BH K�����,<O����-oX���C&)$Q��I�#�'1��/\�u�@С� �s�e�ȓ3=�(����&Hڠ�s�HKP$�Ez��ieў���X��L��0�r���ӹ|h!��C���a�-I�qs� P�nXP��=訉�Q='�I抑�#D؅뉓��M��_�&�%�")B�=0P�s4�HV��8�O���f�%,.�@��a��ޢ����d.�S��,��j��}��d��,r�m�I�#|BB�	�(�"ĒƊF!~`HkaLI�f�~B�ɼؔm��(��T��� ^�C�	���c��un:�
�a�
���D𑞢|��͐a����vh�JP2HաQ�!��C�(pnp�@՝j͠�
C�Y�x��'���6�S�ĨQ�3�L}"����	�@�y5�Š�y���kؔ@S�׆	W�X�7��1�Py2%.`�I(�G�Xyz ���܈5�6�FyZw���у�-���]Δ�p��ޚ�Py�i�)Kv��#�@�MO����D��y"��#,O*��d�E�$sDq���R(��8��'�@O���d����1À��V��X4��,LO�8S@m�+*)��爪1��3��_����۽i� �Qc�3+d(��uh�&a!�D�%D��MH���>7Hʁ ""�+lԠ���)�矀a�%�f!��7h�0�(��E���wh 9�#�%z�xL`d�7mn���	b�I�km4�i�n��aS�fږp�B��>���d%���V�%O�K�L�<�'�ayR����S� �R-��aP:Z�XP*�'bJ���2-��	�УQ���'���0`a����]�F��F��	���*�z�Ҕ��Ň"4iV�V�T�<��Vl~�2	�)�4�@ �S�r�ȓ^2��I`@��H��!8;6��ȓ9�����⎤1 z#�2F�X��x	�Tʲ��4a >d�π�2눨�ȓK,�� �O�'����rȄ�{5\`��F����K[�����.>d������~���#����i�ȓd�2}S��-2��!Ñg	�Z�ȇ�<t��)CD[;NCڀ����>y���<f�lx���:�칒g�8D��=�ȓ	��XQ���Nf}plW�E�����p���XfR0f�6�be;܄���]klɊ�"����l:��Q3
6��ȓe�=�E�"�2�o��d��!�ȓ�t��ZIx,��-u-�-��pٸ��"1@�"��~���ȓz��S�L�/4� ��,یY��ȓ`sd�	ĦG$�0B7c"~_�p��S�? Z$9���cY�e�P&�/iz℁�"O��8�ڕO�X�X��(c��-a�"O��1�ݱ>+%�׫ٱl��A8�"OT����9��I+u���C�@mU"OR	pG�MA ��"*Ȣ �*��"O>���dƗ �����c�5C�6��A"OJ�h�/F�V��H�� ��@kD�"O>0��-�+Et=a�J.A��L�t"OB�c3�E
�& �p�H�v4��"O<K Y/,�^��C��_I\���"O\(�����;�JT��&�:Q%�H�"O����U�#ĕ!��U6�s"O\��I�j��Z��B�?8�"O4�ab�_�g�tp
�>Z�l�"O�i �H�D!
!K�� (R8��G"O����+C .�N��1,��zʀ�"O�@+��lmq� H�o-�d"O����Dm!3�0����D8,!�E�r8z0�ul��,Kw�J�|NxQwCƠZ�x��1sXaz�^ܚ,��D�KΓ`
���y?Pa��h�u��Y�,{�ȓ)g��IUa�*yϢ8#��5a�r���ɾ堄�2v�jeg�6B�����c\��	��È�H���HY.%����K�"����ʘ����D��G ���i�fQ��\�#~-�S$��<�ȓVy��Jv#��x���㋌�P^T���. vh�g��>emHT����k��$�ȓD�b�-U�ȱ0r@�ņȓ!�����%��=�ԂȂ'����1��K�"1>�8��T�+{RT�ȓ%���B�X
�6aH?L쾙�ȓy���B�[4K��6nM���!��'�l��ҬG�+ʸq���b��Q�ȓ&'�� �zy" 	K��K����ȓUqPЭrglځ	�&���}cBX�WNS�(�
"�M 6�ȓK��	�a�	w���ꐣ�L`��ȓݠ������`�iƈ| z9�ȓzd�-����O����҂U¹��b��1�B!Bg�hY�N�#K&�B䉈hXƀ����.��i�F�.s�C�ɓ(��ep"ʇ<N���bF$"� B�	$-���DݯBU޴�'ř��C��1��I��"^�.��G,��"�C��--��=�W�����c�GDPB�	'���2tJ��$H �GbN!hC�I3ª�xbn��$	��N�'0C�	?z�((৒�bh~("���IC��*N����PnœO�H��U8
&�B�	,`��	&%�#�N�@��+ �C��#J���t �`�a�΂�cy&C�%d����"n�퐨�E�C�	)Qs*ƋOFj�;���U��B�	�5?΍"�J(� ��ma��B�3R���)p����b��"O��I,
�hݔ��!�3Y����"OF���ϊ�1^*��3F���%"O*a1q�aֆ���fQ!��TI�"O ����:.��b��8�V4�"Ox�
b�>Y�4����V H�"O~h��F�:Ɲ#���?Q���"O���FK��S��*r�ƎJ"����"O���ȏe
j�Wo�:ż��T;O��p��&�)�g�? `��6�G+ �Dxz���,c'���"O�CV�\(eѰ�F�� �`S^��	4�[�ka{�b�\�t�(VF��a$9`g-B��>A�C:.P7��1�ʰpCA#�L���CF�)]!�D$�l@����^�>��sA��C�ў�Cѩ��T�>���OM,P�# \�|����wE:D��i�iT>��Sf�?EQ��Z�)�ON�qPCO�丧��Fqp�#Yr�h����ź'�f=��f,D�x�w�D�y����C͂1 �Py�i�<�7.ϴÄ��� e��Xa��4|������#/9a~⊑�l���鸗dΙ}�$,-X�A��3��	R�"P�s�� �H�D�d���0T�ɱs�P 9όep�!��2�����e;C�ۈex�1�æ[�r��܆��J�k�˅#)ʨ�V5	���ȓ!N`�Šܠ~�ʈ� ��-W�2��ȓ2oJ��7��o����qIʗ,������X@DK����.�q�h�ȓ�|y���$������� J��̄���тKUW�2`�cϙp&�؄�y�0�����"a���"��=����	��[F*	Q� 3&v����W,��"�Y
p�l"0�,<�q����g@��@.p-��F�N;Du��l5� !?}����v��v-����M	���LCN,��)���J�H`q�DQP�)���,|\�u��z&P%!D��ZL��D��	ڊ�ȓF��ˆP���mӱą'���ȓ�"�����r� kq�5p���ȓ\�rLI�M�z��0���c�H͆ȓ,\t�B�ȑD�X2�БZ@2(��E9`h�R�?hĪTH�"�Y��l����ȹd�����Ə�y��M���ř+��\��P�(�d`<)�ȓ�8�I���*`F��� Ԇ0k*|��?0��2�`ܦdX�HRnۦ�z)�ȓk����g�:�\���/��#�����N-�����0!�0J�Gp�0�ȓ:eE!�$���`��,N>��ȓ/��=m��M#B\[dB��J�z-`�'i^�X��X�Z����Sf^�>R��'k�<�Q T!y�0��O�(F$��'����&(o�$�-ȹ'��-P�'�Ѕ�Тv��l93����4#�'R$D���0�� z� Bjd)�'�X�yq]�b!
X{�h�F����'��Y����R.@����J��١
�'.raB���w� aQ���q���9
�'�u��Nւ;�N1��űt�h��'=*�kP���s���;���u�<C	�'����7���b�Йx�F�`)����'xVa�D��9h�p�#ê��/���	�'5&hI��"hdy�Q�*r�<Bq#�u��(�Q��q�H%�g~RD�x��e�D�W���5b����x��<�����(�Bia�\ |�t ����<��A�ri��z2�Ǉ���:�I�'Hʽ
�MV��p<��ԧ,�|0	��6[������k�xlQ'M�9��V��� B䉶&�ȱ�P/Z%2U��k�*g���^�Nl��g�#W�F���A�8��	�]w�(����``�-<� �`�B�1}X`��'���h`P"N%΄!���/��+�u�=�4"�`Xd��R�H8#UH�p��t�x�	�z&�r"@8��P1�ƛd����$���&��2&�^���x����O�@X�_6Yb>�+��;ft�Ô����u��C~8�x㓏�s�a��#L�(	�BǢ2?��������>[�ƕ�I�3Ƭ80��݊I���� l"7E8�; ��?oxLsu�@&c!!�d�7)�*Qr�HTz�\!r,���;E�j�[�
Ȑg���85�Z^�$�kdJ�=��W?�k�Ì�D�4��n��#��O$D�d�P��y�>y �F�?W�d�yQ�4�~Y�G�l�C���-�d�@ޟ>�P�Hߪt��ʓP�
�3fW�x��$L��7k���퉸�y�&M��X��_�RU ��)Ñ)��H(��\��qx�E��.�&8�«@]�9�@�>�]^��2?^�8A2��4rb��?��'�� �w	Ŭgv�!2ׅl���!+���m��P�7db�Ka^�^�x�@�NQ����z���)���r�YfJ�]S�ڐ|�(���V�`���e	�!ѷ����v�QN?)�sJR��MAr��uB9!�+D���%o	�"]��+�$���<#���\���Kb��>WH4-�.!4(��y��pj���CjR��c�������9R�؂G+O[l���K�/33EM[O�X���~����V^1NDkB�P��h@���-<b��U�Ĵ'�Q����C�m�Je"�-�8L�#�r�v��-\+(iT��B%�O��Ix�����Eu�5y�$�(޸Eن��L�R��`g=�On� jJ����$'��G@(y�A>O��9��J�Hz �!�$�t���JK����g����� �FE0f�J�l�|���UޞC�ɹ0T��e�[smⰫ�!R&J�:��ㄹY�i�F;+4I��)"zR.uS�$O���ǶK}����2k:%HcgE�ta~�BW;9�A�#��\���=�xP��o1>I�� �NT>Ӓ���8����D�O�'�>��-��i�<���>j����$\�T>���E�Յ2P��s�8�]hŃ�J�b���Pt6�PP!.�� �Ƭ�p?��哟wU$ ��$�O"���#��<qw%]O�0��B�	;�Q��s](4��DO�O!��O�����Ç;f��9�i��3^Ĥ9�'�j}E�Ƭ [����� �b%����Ux�B �\�]�)�O���I˸#�
�s�_��~����^y�m2
_Q�. �1NA�p?Yp�F�?v��G��حPkU;Z�Zd�v�:#z��;��1�F���,E7m�J�#��ɓ.���3/(Ab\ݱs&Ef7�>��ɋ91�(�"T&�8`\�X�N,���@d��VJ�x u�,���JEB�9{��'7������3�B�㮙�6
=Q�'�X893N�8�1[S@�&1���	�F��g��'Zf��Q�F�?�.�����=Z����I�<���+�>���U&m̄�)���0Q�D����	y�R}��؞@O��#�I5{��$?�3�'��I�)�E��4;����g�1}m>���j<3TlD��B�:a�\(�A��8r$��d�-I(��pi����둡G�K�Ђ�2OT"?��S�m��h��&Ő!�@?] ��|f�}b�ƫY6X�p���2 ��Љ.X��(��ʪ-�� �p�S�k��C�	���*F印k�>���l*���Z�k*g_����	� �����*��z����O����᜛��$:�lLE�n�A�2��Kc�������`��6�R:D~%p�Q<H����@K�:or(˓G�"�F��O� �4֭h"fMX��4=�8����Z�n�|��e �f��0��j��DQ�X1`�n� ӵ��V�Z���&옋��<���W�a(@�'��R xe{A�V�*Vb� &�|rC�j�3�F��ƂF,T\��)YS�B�D�]'0ה�t���񤒑NkRe�
�6<�#��v*���դU����0��Y*@�Mn^IR-O�O���ä/�t�`=ȰaI�Ok���ۓ<0Q�ɍW}ҋSJ
�yr3d��)�z8jT�[��y2h�%����`ה9@���T��O����'0����y�ԉM�m� ۞H�Q��`���L:����7!VT�rń�+��В�ˉ$_V	B��4c+p ��^, ��C�ݐ4Bf�ղ]����K��];S�\.|����.���ȓw��8p�
B9��g�"X�\�ȓ x����=ƍ�-�4(N݄�p����NȰ_#�qI+�?7ތ�ȓ[N��ۤ)�4��@��J�nHhȇ�L��0�A�bT@&D0Cy�$��:wp�I���.K󾩳Se�
]Q���'�ք2W`T�aY�����0{���(t$lB�D���Y��G�\˞�ȓr�I�Ƈ�V�d������9��_�L��#� �n����eG� �ȓ*J,�&͈$��'�-b��ȓd���Ӕ��(@� P{�͟�w��0��S�? �ͳFbE�[��}v��dY���"O��[�LP1c؍�V�'��:a"On5�JV�"���7���N*,l0%"O|� �I��	L3�/��*z�%Xb"O>��#��!=�ƨ��R�va��"O��`4f��|B­�Vl�of���q"O6E#�ʐ�
= !���SM�	�"O��j��C�Z�����ׄn�l��"OX�Z�M�
!���3��9�lX�"O��6ʒx� @DK�1��iu"O�A���[F�09t+�-�I��"On��m�]["��D�L�\�pI��"O���
/Tv=IvfVúI�D"OX�B�ա4
�y���$dߔQ��"O�:pB&[x(0��|��Dғ"OV�{cJ�{�qY�kο<�"���"OU�f��P�TE[�-�
n�>�i�"O��+� ǀ[��8��-%��:�"O0�+�
�?Lze:AM�M���u"O\�6��^���-ېz��e��"Oh-���E:fy(%t��r���"OJ5+"m�Cnr���V�-�x�<	��6��\�2*��B���Zfj�]�<!TGȕH!x�$������Ӣ��_�<!��'H����w�
+z�it&s�<�d*G�$��\�S`��=�&}�!��b�<A�������ƽ0љ���a�<��������	4��QƧ�z�<�T��I�)p�(�^ABqYg�r�<a�*F&U!@�@� So���2�l�<q��˳b�L@(+(F����h�<���-x��5)�,E8����Ŝg�<A�� ��t)��D��s�NIc�<�J� 56�Wf�s���c�B�^�<��䔮g.�4�P�qOj�K�b�Z�<���9e�x�df�Y�ZQ���Q�<ɠ�d���8\�8<��iߩCa�B�I3X��DBќh%���UC�ۜB�ɫ#ƒ�:���g��u1���NB�Ira� HW�&:H��1�G�+� B�ɷ\��b��Q����6LQ�w!�B�[)Fq�b��m�1X�A�9S��B�I��I���:$��d
�,	�C䉱?j	�VI@�+�&=+�
¢C�Ɂu��DQ�E��J& -z�
\uNbB�	�LRl��J��L��I,fB�	/;B��G�O�'x��s�O���C�I�l��X#��U���;��ݳz�C�I�F�dh��LN��1^�ix�C�	�L�!ӲFJ�m�릂
0w�@B�I�n��UR���N3�-��B]�r�fB�I
�(j��چ(�z`!7똕b�~B�X�}끏�rĘ(�u�'N8�C�I�i[�pxrLVxKZ0�
N 8C��#At�i�@�̧=StY�b	�(�C䉛���h�F�C`�[p��:T�B�1xt�(0%���Y;�Lx�ż��C�	�	�j��G"0���q���9�hC�I�RS�ͻ���h�
�a�>t-&C�W�RթԎ+
o��hw��,t�lC�I�Wi"�ZD3o&�X�����&C�ɦ?Ұa�c`F�zz�X eZ�W�.C�$T�9QĖE-���g�n0C�ɦ�@T�'f�d���2A.@�6=NB�)� n����$�`��㐒7��`�"O|�9 ,�!k$��3��Q�:�&t�"O$	+2�Y�8B���n��e�'"O<I���uB$��색2����v"O�e#���P	f,�	N��9�"O����E�:"Ն���I_���zS"O� J�)�.�0�c����}���A�"Of�1I�Z��T�9J֎1h�"O�
g�I�p;���3M����t	�"OX8bv�U�=ȒL9���1/�Y�"O�L+���'.N�)�N�ZŊR"ORd�.B�/R(1���� ��,j�"O���O�r:�d�Dǰ���"O�d0�F�<G�b�f�j�4"O�Ixp �[�����Q��$"O ��(-$��·G$���C"O�h���0�Zpj��^��x�t"O8��A�hY�Y@�]6.�H�"O��c�CO���r�U�]ԙ�s"O�]ҒA��t0 `$�'4	�U��"O��1��]�#9�\r�dR�d�Bxa"O�tb1#
(֝H���<<�"O��`f�,3�m��%�.Ŝ��"O�5����.K��A`<��R�"O^k�$P����S��T���Z�"O�%���;�YA��[?LV���"O$	Z#3���ABL�i*:]��"O�ͺ�o��4^�b��&Ft4���"O�����y�JS@A  =�x�B"O
yd��!N�"�A��m.��c�"OԄ K�b�<]��@�C	H��E"O�!��)ea^RW�	�%��"O��w�=@����
�{�*Yb�"OJ�"V "y��kTK��C�l�0"O�huaU�9�A�VI/Ǫt@�"OV�Dϛ�.���A`��s��p�"O
I��K^
�&�R!E9e�!s�"O<�Cd�`,���R �ҡx�"Ob�+�Fƛ0BL�"΋ %pő�"O�!��J%F��pԇ$>�"w"O�	��Ȧ5ch�+�!�/2h� ��"O"��� E�ҊT�r=���d"O�U�8���y�nN� 0���"O�X�⎎)�H�b�L�J"�$+�"Ot�4+�H�p��˯t(��$"O��t��a-)10hraK�<�y��/(M���U5P��ٓ샟�y�B�<i=�͓GE�G��ɱ�#�-�yR�!@�2�a�0T٨f�^,�yR-����Mȡ 
#q`l]:#�ڦ�y� �T��P���*iI@�
�&��y�a1:;� �Qo-��k���yB"�r���0�!N@��H�>�y�ʎ�UC8��p�A���/�y�DSh�0	�$NY��YBƪ�-�yb����aA�/��)�uҮ���y�g�!2�9K�"�X�Ӓ�y��
�0�x ���)��������y'�*�n��;���3O�/tf!��Z�w,`�% �W�~h�`-�'G!��0��Q�ŗ*-�&�f��;J!�DA�
��L�$h�0p�e�w���O,!���09q�	�kضOc�pҀ��i!�����sNZ�I���:��^�&I!�� |����ȯgӢ���G�`���"O0I�#A�PB|aç�<r��Aj�"O�4+��ܲ, I곃�
w� ��"O2%C�m�J�^�����36� �a "Ofp3���^j��&�<%�y�3"O�Y2����b����>5QY�"Or�񐎘3]�<�5j��0� i`"Otщ�Âc��X�	z�208�"O���#ԓ?x�䯌!6�-1�"O"�Q��@O"��6�$����#"O}y���	������������"O(����X�kn�� �@����a"O8��5��f3�����O�o�,1��"O�萊�_�$s�jM*j���5"O�=S֮_(��}�q��(���5"O���`�rP�W�U�<�a"OD0���ڭ�l(�E���7�=f"O� '�F�Bv���4��O����"O6,{�kٞB\�M`c���_�A�"O�,�a�C>���k� U�7����"O�@1�I��U:�@Z0���"O�Ѫ1OR�a4��E�z��cF"O������.i��gCK37��J1"O��Sᖇ	�9
���|	���"O�Y�
�Jhp����%Yn�D
"O� h(�8't�-q��&HBe2P"O�%YF<\�8y���/@u�"O���Q��k����Fխt� �"O�Q�'�>F���hĦN\((w"O@ p���>vz��d�_�G t�f"Ob�e�Y�{m�[W��.��Q�"O�Pѭ�6<��ѵ�ďN���"O�qsw���� �"͕}�0��"OԜ��ʚ
<u w�]ߚX0$2O���c� �OJx�b��o`(5��K�#A���b�'x=KT���DM�
=��!�O�Q��Q3�`P<<�!��T4D��.��τ�����o�qO�ݹ��5P��#jr�ߐHc�x1�FB/)g�<"�.�e�<q�J�vH0�+v�J�#����J_�2�*�Qǔ|Ҫ�]���#e�鐀B['���W.dU!��xvD�B3n�{��L�AX��ק��1�X]��	
U"@#F�=
t�KÍI6j����@��l[��>�#6lFE��@�K&(!�a�y�<�Ä
�> �չ�@]��xy&�q�I|� �V���ȟ��Ҭ�*}��U{r)U	3�!�"O�x�aLS�}.@�r�)�(��IM��:E'�����<1��-j�z֎+|�$(
��g�<��E�5������ϓ[�t�9P�̞Z�Zc�/H�a}�(��F�p4�gE�'����s����=9��?px$��'�bl���+�`�	Am��4�jh�
�'�pfn��Ѻ ��(,�r���A�BM�d�(r���KROD	#�T]PqDW�<I%�)#�*�!\
\�~9��k�o�<1�ɳ*�R�Iu��?뾴�v�i�<0�Ųo���P�hA/up��P^�<�r�F�bb��a�	ux��ZV�c�<IpI�/�z�s�(�2L�8���N\�<i�"�9؊��d Y�<!,�ӳ�p�<�Ƭ�����"/t�N4�$�^T�<� �"~�LTwǇA;@9���W�<���]A8E�fLr^8���K�<)�(�<�>� ���`�
��)�s�<i��)�̙��hK�B� ��T��f�<��/�0R� �Ñ+s|F��"�f�<�  a��g[s��3C$@h(��"O��*��O�h��۳ɞ79�䅣�"O��ۆO5`L�u����x�|��e"O���DG�n��<cFI$D��eP�"Od]B�E�{"�= wj	�ƌ�"O�����J�R����L�Fr�cd"O�5(2�ϰ2����LQT�Q�"O:!$e�;:y�,*�B
-�
��f"O���H�s3܈�@��!o�x�Ѓ"Oz��B�q��$a��~�AK "O|5m��E@�G�F�z�C�"OvɗhZ�3��Q�aE؇F����"O�xAѡBkH03���/M(��"Ol��͐$���m�!]`k "O�`�d&�)aj����+Bz4�"O����C��h��!�7�ӕ<g`���"Or �T�J�oJe[�M5F���"O������ �C��7�`�"O�j��0b �%q�NX4$>D��"O��$��� ���k֍X�ʀ�"O�QLX�'�1zKءH�<� V"OX8AF��?����%
�/(��ؚP"OnB���}Ll�`h�3���Z#"O���o�	z`�����S �=P"Oz�k���P��R 5AV��bA"O���,˔	�V,�ĈG�4���"O��� ��pfPb�ܭt(�m���ݽ{w��&ae��2w�'`����� PT �����h�ߓ��'����V+E����ゎ	/A���+O�=E��CC�pw�M2c*�3>y�Ш�?�����+�|��-�E7��0�!M
<J �=�çA�X�wAR�|��DV��G�5�?���i�9��H��V9�}1��Z� )���'xPb�9�=O��	4Nɧ�������J"IK��ВD�*;<��e^�LR�D$ʓ�O��/�*TCn@H�� �ԑp�'�ў�~6,�!
T��*�^���m�'�a�d
������%L�,������'ў�O�����'��#��e��⅋��QɌy��'��T"��Tk�Hz�H q���9K$���@�b�{G"��?���Bz�SI?��J�6N�1�`],!L6��F�׹��O��>1���Q�BQ��"�tu�"��H�'"a�� ��X����$MMi�c����'�ў�Oe,Ͳ&��6J��4�C��@٠��M>�����B�+R�U���ҤW]���M�*��F�'(�|�Aiʤd�t	3eT8vmpyrA��O�H�����O����K�L1¥Y�d���`退Dz$$��T"2�2�+��Y>�p��+�S��I�+�}������a�SG�'�ў�>�����=�l8�'Ձsw��23ê<����Ӈ^~8!�%��%�,�[����v��3���f����!��<!�<�7�*�a��Ea�hL-�j�R聣x��D�1�����+p�Z�0 n!_Z!�d��L�Y��疴Zl-#/	1S!�dB�9�����]�P�D���W�P<!�4RqV��s` �kF 4�h�1[-!�䂗fh\��u�΁ -0���M�"+!�D@�#���򇚕&��cBl ��!�<n�Vi���̧j�X%� �(Jj!�$�Y"
X04ٌ}��W�,�!�N'֬Hrΐtw��K0,�\�!��x{,�yCjG� n�HH�¬�!�dѢ4�捫QA\�nW0���C˫!�d�) �=	b��^p2�Y�b�=rJ!�Dȏ���%OO+m�؆�5R!�� �󇇐�o�޽c��kª��"O�}b1���6�	R�U0�"Ozy���d�����K�5�ĳ�"O(��q	@<���{�Nǚf�@C"OjH�-C~]�1`��݅,�\ �"Ox���	"$�n��U��Q�\���"O���̜�;Bh�vؼy��"O��D�YW�d0Ŗ�"$�Ӵ"O��l�i�P2��`	��C�"Oz�'EI4������2�<x�R"O2��:�d)�r�����z�"O|̓"*R�'\4�z����d�"O��:�D�+T�(�c�5݈�@"OLP�a��9K	"�HPDHs����"O����mV�7=�dR7��bM��Xc"O�[�L�� ���o���!�"O��x�,�H���C�
�H��b"O���0g
�n-� ���%��U�v"ORTr҆��P a`Ӆ��E����"O��dK�'}��{��٦o����"OB����X+KU"�H�dMj]��"O��x�Y<I�~����3pAz �"O����k�E� �ɻ!���0"Of(x���9��X��^�A[�m� "Oެ�s����T C��o���a"O�
��*v��q&�N����S�"O$A���>\��W���r�@;6"OD(�Q͖�څ@�c�%U��\��"O�	@���J�N-��)��"dqS"O~��m|P�p/Uy�̡	1"OB��C06��4rOH�*��<`"O���hU�A���Kܤe��"Ob�p�ΔF2�`�o>��a�"O�]I&�S�XD	U�G�K�> У"O��b�Z���s&�Ñ��	ؠ"O�X� �@�Kv���4��Tz�P�"O^�s䫖�s�8Q��!+��9�"O�죗�Ä3@�i�S�].H�2"O ز�^�^򰈐�G�A���{�"O�ےg��`�����Vv�|�"O"��f�+�&�Q&\�!����g"O��i�n��S� )#�>�^���"Oj��&gW�i	5�m�޵�#"Ol���A�2`�������j���'��@9��+*x	� �I,�4���'��,�!�ўjKxd[u*�.&X(`�'ZR'��&��M�B�V�y�'����jW�A��B1V����'�M���Y#!,P���!R ��'O>��p@X�|�4S櫍�3�y��'{��{N�
T̀�u�V����'w2��2HG:f�H�s�FXl��'��q	�
CF�ч�ۈ?K��q	�'��ys�AR5C��$+G��3�L�b	�'u���V �4bX2-�SO�* 6m��'�����],X���/��pfI��'�:�:��'Z�<��b��2k���:�'4n �Eo�p����Z(����'�� yǩ07���A@�ƁC����'�v$���ͬ4� ��j^ �ЙR	�' ��%ܾ3��q'��I܀ Z�'��"v.U�OJ�����'Eg�y�'�b<�'źH���μ5�\�	�'��-�rk�A�Lc�'��
�	��� ��S5X:���	ցZ�~ L,B�"O�q��L�}���d���\�[v"O�PDK��O�v����o��(�"O���Q��wj�$)`L/$�p`:�"ON�[���g6��H�O���Nԫ�"ON�a֡H�7��=�A?����S"O���G��#bi�A�;^/����"Ox��6mS�d�|�atO�*d�<�"O>TK��ח��l���&א��T"Onl[�A�c0dk5��:l����"O�;�( ̸��5
����T"O���&L@ =(u��i/�4\��"Ox!��N��Q���k��ݾJ�X��"O��ƥ
=n�8���3椨�"O���C��$����1�֜5j�"O�ə�#D�N�R�)�hA""W�-x3"O騵H��2���t�]�Lu��"O}��h�1zU&���e+PԢ��"Oj�9�%��H�,\s���?d�x%"On Qu+���L8i��LC�"O�)񌙒]ZB�e
Ɨ_�!0�"ObP�����H�X�h�>M��$"O��"�bC������6�Ie"OnA���8��;�Y
�:�x5"O��`DiT.?�Kڼf�8���߰�yB��{����ÎJ&aiRQp&�ְ�y��W^�4��W��(��y�ɻ�ybh��'���P��H��x59��A��y2LL=:�Жm��ܒc��y� ��;��ܐ �8�nI�w�#�yҋÕp6es�d�������y�HU6J���z�����=E�:�y"��j3A@�)=� fK\�PʮB�I�:���N�$��S�r�XC�I�r(�P�P�-3����!�+o8C�T��H"B��\D��i%�1�'���B�@�C4T84%Ѭe����'���i�*�V���e^<cUL@��'�x��'799B���ӂ^�L`�
�'�.hp"/B�l`8���*z*��
�'!����IM�D8�8�n�.��M�
�'��\�^�RT�Fn�>`G���%��yƤX琈ؤ�v��U��y��=מC��B�k���rb^��y5?2���dD�p��`RW$��y2�]�cf�.I��4%���لȓc��H�H &wS.��흮������{���y��z�AW�R�������O!�$�C�f=���D!vD1b�F"!򤉾8�Us��Y�]{�I��+��f�!�mc���g(�h���X �C�	�0���k�<+� ���ٺbpC�ɖ{��+k�7���u��H�HC䉙'�$ ��� $����%*�$C�I*a����a.�"�lY�E`X�U�C�ɝC��� ��`G� ��`nB�	^v�7N	<w��*�e�qB�I[rU(tƋ����,�	s�HB䉰J>�x�D�U4+��Y#��Q�|sB�		�V,��+SX����ڹEcC䉉~�5@ �$e!~1z%,�2:��B�9%��arJ͚v�x�SQMػXC��W�� D�99ar��,�',��B䉫MV�p�F�W�E;P��#,��?X�B�)� ��Ѥ�J]�� !�!j<��"O���rə�m��x��Rl*�2"O�u �� ^�|!�����v�C�"O�p��t2)A��U�-r��2"O�b��E7"4(Q*_�iz^���*OԽ�b��X�E	��0���'������)Rܚ��7C	�;? �0�'K	H�7z�(�"�f�G>�l��'�����-�J��KȚ4�:5��'_��2�lϤQ�v�X�m��,�=y�'=�����(_<l('K
eUE��'^����>S�\ 2��!d�<��'aZ	Æd��.LTQ� *D�T�d���'a�P�\(j�YI` ն"�t`�'�������0!�̙#!�x`��'�n��T�<	-�ݑf�[�EҠA�''4�xW�Z�q'�	@%�<���'�������^w��!�L��/��! �'ޠi�B��p� :!ʍ� }�T�'�d�J�]�0>�c��΋SӴx��y�he��2H�)kt�=Y�Nx�ȓGvmV��;�0�8�+ŷWi*)��.Z�TR �D�}H"�P��
3H��h�ȓ?ذ�p��H�-���0��.4�$T������&^�uQZ-a�.X-Vd����+�v$�3�C���A�T�Y{g���ȓ�j|���ݎ�D�ŧM�H�v��TE�	BS�G1.%8�(�-|y��'��0���5���#f�V�T�� /@���+=�F�����aw�y�ȓ�x �����a��`�q/�pd�ȓ���S��!S���Ѱ"�'�	���ȱP��=Z�Rw�ͻ��8��Bg��:h�#��@�&�ҵ8����ȓ�B�`���)#"u��B(� ч����)��B�G�,bA��"c*���g?�9BdJT�SY�$��GU]"����a�Er�oZ�@��M�d�O>����L��d��K�|���>ṅֶȓr(���̸HA��ҥ7x���>�~ܹ'�ؔglx�8S�2;�Ḧ́ȓQ�|��	�*����(�̘u�� P.:�c�C�X!,}Ⅽ�G�<��i[=l�z�{1�Ǘ\�Z4��ml�<	���3nu*|؃��)Tn�a�#�M�<1���):���K�F����O�<�r�S' �&�����v����e�EJ�<d��;R}�]�Cb�E�X�R �CO�<9�!\d���ʏB�b�
�-�J�<鰪��K�p1��D���B�<����[u�1��B�g˺��2��g�<�M�1h�T)���#�lp�A�m�<IW�(^n�9k��z�#�c�N�<iD�R4PԪB��9Gz�cd�M�<�p^�D4�I9�a��Z5<��NVB�<0i��PtUz�����|�<���   ��   �    �  '   q+  7  �B  �M  GX  �`  �m  �v  M}  ��  ��  9�  z�  ��  �  E�  ��  ̵  �  Q�  ��  ��  �  d�  t�  *�  �  %�  R  �! 
/ 7 _= �C @I  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	�Ɠ����Ԭ��ll��vI	d�*���'�5��/?px�L���]̚i��'�RM��cR�l��$C�̐�r��r�O�4r��6e�mJ��˭.��(�"O�\:&�֫[��
f� �i"Ob����	�lK��uc�Z T`��	LX��YS]#��ť�򙡔-7<O���?a���P�	�p���0�x�3p�<!a��,M�5���?�*u��YA��O6b?�BvMR�X� 9@ݻeL2D�d�FlW0VJy2f��>{j��AG/D�� P��P�j���N�?.��G)� n&A��)A����0��xXׁ�3\�R�<G{J?=9�Ǎ�|ɋ&l�*	``�'L#D�� �Q�O�cz�|B%b?7�b��R�4��h��dA�dj���P����)����{b�䏩.Q�����C����:�"g.���`OB�I(\|�b �:0 -�t�' �'��yh�$e�(%����:>� �'�B%O�5��U��Ҫ]��!�'��!�O3SN��fcH�]\|�K	�'�����05�ІT6bP�	�'6��9�-J�~~D!)�A�Tl�{�'��F-X���Y���;K�vP0�8$�� @"$kmr�NX�o�"m��l2D��Q���#�T�6L��@E�B<D�p°�^��|�7ZU�|�3f8D����G?z�R���ظ���@�l5|O�b�|�ըH_A�A��>/�b���E2D��3�1X��t��=#�z�	�.���GxJ~R�_���2�˅�L��������K�ƅ�s�Ш$G�<�$�%s�DGyr�':*}�EĚ<gB�G�<JK��
�'E�`�̶='�<Y�[9T��:�'Ѷ�C�E
4���A�Ņ�7���ډ��#�������!�����GٛcL��p"O|�@'c��HQ�@�'	�RDԨ� "O���u�D͑���|&�e��"O 1�  �|�x:�D�%�%Sr"OJ#b�^�L�J}�
�0.="O̙C����0�`\��X��Z�"O����o1y
���1�)xـ�C��'��Jph���B0c��
�T� :!�ךP���B3'�,�1���vz��=Q�n��6��k�'�yש[;�TsREG�y3�5(����y�_Ozd����1�5 �H�?��*�n��~��IO������Y��6E��b>����/�d�"��� �J*�6q�Dl���+�|LGy����xL��Av,�%g�|��`*ԗ�(O� ��<7�B�@�m���w҆���6ᑞ�㉦e��� ��X��03���N���H��}>�#0��e&ܑ��ċ;~����#�9D� �V�жk1�a���ʳj���T�3���'ͪe�O(5P���C�8�J��b��E
O�7-
�p.U[`
]�/D%`��r��,�D;<O4("�a�N�|�k��N�L�d����U��z,�F�X2���g�b��[TjL�*�iOB"=E��4�,�Z�#� p^�Qg`U:�HmEzb�iC�I��O�<��'��j��r`���STy��[�L��I�B��4�AG�&!L ���<u�=�;O���s�Y�F�_z���ˍ=�i�3�Ot�	(
��v�ZA���d�5$c�h��	>
?r�;ՆܔS(�h ��a�!�$T�8�b���U�.H8��wB$=�!�U>
yF�[0n��5ͦ=9�#�3z����k�ӧ��xw��C셀/��ƓF�AH΁s&*��6@�8P��a{��(� v���o��<v��?D�t#!W4(��d�� m<4��"�^�����d4[A{�*�2> v٠��$Z�a~2T�(2u�����8��n��Bb��2�Lc�@6�Ea��|FzB��=D����Zݦ��"���hOZ"<�+��8�g,�%6B��4�'EN���R"O&�a��ɋZ��4K���= Uf����i��-'��է����g��aX���G L(�b�ޖ�yW<�1Ĕ�G|ظ�(!��+�	s�'�� h��/@ǚ��������	���+����ӧ�^ɐ�) �
)��Iv��h�� V���ŁA;��
�Í/O �l�P�I�ژ'�1��$p��E����qA�R=#�Yh"O!���N/�5b�&�56���'���.�	P�'4�]jdB�n��M+Co��vaI����d�±y�N�.G��+U�ƛ$�	}x�d����8�RX�BE?M(���+��=r}Q�P *��U9b,��6�~�b!B�U�Jt�#�'e��=E�bR�Q�$K@�T�дt�`����'[N7�$�Ĵ|�Q2�{!
��.��ܫb�#/�$D�ȓ>�>�A@�+����Pn�9؎�5�g?���"K�bM3DK�%��R�j�i�<��͉�8�����*#��Z���p�����#�S�dmJw�@� glէH���Xa� �y2�ȶN`���rlA-���@�|�<��+��n��`H4%r�l3�l�y�<IG��jN4�f���0�����t�<�f�A����l؍N����Sq8��Gz�]=$�PԀU5���K��y�Ȗ,3%B�Jd��cJ�Q��&�yb�ˤ[��KQ�}��!1���y�
�0%B��E��D�� q��@
�yB�;@�N%��D�O��M�f�A��yR$�i&N�J@ �K��q�K��y��H	I��	)�,�E,x�0[��y"b\�o8��˃i	�8��eh��yōn���[�E/>N�y��͏�M�,O6�O?7�]�Ad`��Alz��GM"5!�DI�C<�ˁ_^�tu���
u�!�$�:7l<�M��o���'B/v�!�M�
jA�0'K9o9(���Z�F!�	
n"�B�v1�]�� ]-nC!�۠H���jW=+�ȼ�Aoπ�!�Q":n�-ð�_�kl�A�ȁ>7�!�D�L ����d�L�1�F�,!򄐰P��؋�
4	�l-�u �5�!�d�?4v�b��?�(�2���;7�!�Y�R-��	��ʱuJ`��Ù�^�!��1;�l�r�!&Eʷ��!�D�(����ܤi�y�C��u !�B�8d��{b�޾}Qڸ�+дj�!�Ɗ{"�	���1P|<�hE�QI!�S�32Y*�5e5��)3(�
>!�D�T�l+&D�/5� �iˏ33!��^�d�@�J�h[<{x�!AȂ D�!���d�z�[�LW�r͜����+"�!�D�"Q���ɥ�7N�n0q��\�9!�N�Z�$�1D�h�cD�'�!��Ϯp"݊f,P�-�,���O�&3�!�Ԋ;� HHsF";��4i�[�!�z���vi��˖3sM�e�!�D_�~�*��Fe�f�"�​ٍG4!��Ӈ:�VӢ�L�xy�= s(�0 !�$�7!^�;��4�N�eH�#!��Km���%ͼ�5{Ԩ��?!򤓭,���W"ʶG��p���<'!�\�ȰK5�ه_���7��c+!���5�@��W�ц �|��#$C�!�� >?��K�h��HȂPy��˩3�!�D����ͲH�t�6�
$
!�$"B8=7���,�`P��&[!��A~�b��ކg���BQϚ�!��\2t�0Hj`�W�3���EoE�#�!����x	���	�7Ȩ5���9�!�ћe"���i��Q�t�ە�E&�!�� �Y��Zj%��!�0r`"O�uC�a�oYm� ($!��Mr#"Ol��aӊ>ɠT�0��-�Dt��"O�I0��Zr^Y`dF�k���F"O��(CO;{�.���"~4)q��'���'���'���'��'���'z�X����y2Tk�f�	�b��6�'b��'��'���'>��'��'OX��D =Ur�(�P�Խ��'��'���'��'S�'Ob�'�8��s!2h��q���ҩ��Pb�'�2�'tR�'P��'IR�'i�'��q1T�^6 �{Q��
`��S��'�b�'��'�'��'kB�'�xYBg�N�zC�a���
V�8B�'I��'���'���'|r�'P��'V���R6�H � �ƐXb4(��'��'�"�'���'�B�'�'	��bę<g������_�y'�'"��'�R�'aR�'���'�"�'�<ᮩ;>YȇMNMf� �+A�,��|��֟T������	͟|��ڟ�SP蜙�x����n����Iܟ��I���	ɟ���ߟ�	��(�	�D�v�>b�(&��A�EI��z����� ��ʟ��I�������	����I�[�xĻ�f�$1� i$M��v�Y�������ԟ��Iԟ���˟x�	��p�	�^.����Ȫr���U�Q�wP�����X��ğ��I���IşX�ݴ�?��"�"@S�(�g�ȑ�͇;r(�1�RY����vy���Oqmڈs��l�4%��UBF}�C�Z�|L8Ǭ(?�ǲi|�O�9O���	�lmnm�@H�	3=5��ʞC+6to���z�H����'�6�Z$��"�����&��+��^}ȠS���q��A��O���h�>E���I
&(�d�3	�PB��禽c�!�g��v˛�wD���֤��r��� �C��kD 4[G�x��l��<��O1��y�u	cӒ�I T�u��L �!�SdZ����֧mo�(� ˑ
ӈ�=�'�?Iqą�xz�CÇ�Ym�r���<�/Od�O��lD c�h �ㅞ<��0�$HO;NA"��F��?[��.�Mc��i�$�<A!EF�Y<���N�A�h}bD3?���'�B�#`�N�'�V Xw8v�$���Ddq�l�8-��9{Ѧȭ(Ґ����O?�I&��ͳנ�6V@���'װ���	��MS�H~b�h����S�A�R��!>���Ԫ�?q��ɐ�M;ҷi�"�9'�����8�@�!{+$>c{��&!�-d��]C�+RX���G{�O<�u�����2)��pŦ!1�j��^	�����ǔ���';񟖤a�B:ބ��dM:*	F��M}"(t�d�l�<�I|�'�?9�B�$�h�3vG��;W�̒G���4���S}�g6* �E��ź{r�>����10�Y�:(и���x���RR`_ڟ0�'��	Z�I.�M��O�<i́�~$9;�fQ�_������<���i��O�9O��o���M����0�- �2���4'�Q��$c1+��Ms�'���2�_8c^���T"��t��43Ѽ�L}�v��$�͋eo=k>��Lw���	zy�S�"~���)����df�>C�l0 DQi̓N�f���dNΦq&����Ňy*|���'��`{!FR�<��O=mZ�M��&��|�ٴ�y��EI��,��RqV����6}�"#�DB6xY�v��<Z�'��i>��'7rɛC>���p���zT��kB��y�|�a�NyC�|�e��l�̔:��9O���/L~���>��i\�6�y��%>���Cf���G%��P{�Tgn�p�� 1dlr`�8�";?Q��&.� #Yw�(�O���-B0���y��U1Z.� �VO0�m�� h7�Ÿ�xX��+	��;�+����8�MK��`�>���i��W�4| �Dz��\�{j�S h`�V�m��,0umZ�<i��tt��ee�5�El�My�B#]xT3���<o�Z��s$�FG����E0i���(W,6k�} 5Y5qG(�s'��6{�*u�'�Zo�%�g�SSf�d;��T�*k술��A�a
��P&�O�y veI�G��D�z��XN��{F�Q�>S�h`P�F�}"�Eg��l�D�8�A1����M�sD~Tp��F�]�&��SM�n����gAy�dx��D-�lH@&N�gl.�0g����ڧd��&��l��$F�+:�@�쒯sVNI����c:d�
��V	�&f��:�֌aq'A�?����_*q)�5(�E)K��½zB]H1��3�Mk���?����:Q�x�O����@�u�LQ:�d�4u �C��q�
�ie	�<	���?a�g��?QQ���R�Heo�0XM`��O9u�v�'�"�'��g�.�4�����Os�aJ�`��ԑ��=Y�Jy���VA}��'6�4Ԙ'�'�"��#o-nq�aҦ3аM�1#��s+6-�O�a	u�v�i>��ΟȔ',n�#�J��k4.Z1�t)�5�~�`�d�~�1O4���O��$�<)�Ak�^�G.��h�}s�CP �d��1�x��'A��'���� �ə�D����B6r�� �"�E���
tN<�I���	�Д'r��z�Dp>m�3���]�6���H��y��ͳ>���?������O���
�3,��5�Fx�㗊C}�pPt�Ի;��꓈?�TQ��'��+:.UJ|*5BA�kk�˗ρ�nZ�͠2
5:�f�'��]��������+��&vb����Q���+u ��7��O����<��"?E�Or��5FET�g��`l�� ��tHsI	��M#/OT���ObhYC���Ol��� l��
�R���"�N^<PHҵi��ɸ,N�(�ڴ?]��������d��U��q+7H�[x̹��ƈ9���'�"(�&#T�)��g�	��J��cEP�z�����i���7��;!k�nZ�x��� � ���|JV��-k�<�bݐh��Uh�B�b޴m�~� ,O��d�O����O��K�l)�����X��2��צ���ß4���>��A�J<ͧ�?���0��V��
�ݑ�ɐ:��Q@U�T��ԟD�s%#�Iޟ��	��+Vc��2�I�KRw��  �R��Mc��T"	�՞x�O���'!�I�K��k%)�#M�4��̰u7��0ٴ�?�4�r��?���?.O���4?�A���@-F�s��ilL'���Iן��	vy�'\RaK�HEl=�@B�)�>�K�˚"V��ÍyB�'���'%�Ɋ�x�A�O0q�&���6"hD�',�*9�����O���OP��<Y���?9�gn��B,U
���懵t&�p�c�����O����O�ʓ�����$KU�T1�-���S�<�XC�"�4�?q�����O���V2�����1)�yĲ���!\=x���ix��'W�	Xb�y�L|����1T��ʂOZ�]C���@J�f�m�Py2�'SB�٭��b��i��@9�@\��D�q&ʏSC�Y�۴���Xt@2�n�3��)�O&�)�i~��$?����#�`u ���R/�M���?i�(�8��?��3��	�8�Q������y��d�j^<�6��O��D�O��	\T�i>��q#�900��KM�`�(���M{q����Oz����1O �d���6}i��KM�����H8<K��m��\��ԟ ��d�~y�OT�'���رU;�t#'��Ioj�P��� }�p��<	"� �G�O���'� �CXT����w]:uybHD*P�V�'�A�_��������{�uq�p��΋��  ���
!<���'�1����+����O����<�c����jڡIXlF"	2red(�����D�O����O������$@"��3��x'. VB�2(@x(�k^4G�4��?�����$�O�@8s�?���᙮)��c�P����
fy�"���On��5��͟��W�^�� 6킭��M���PkiQ�a�i��	��Sy"�'>�,�Z>i���~Ӽ{#܄T��i�䌟t��bڴ�?�b�'�v�8RI-��kҜ�(�F$tᐥ�/P\��l�۟H�'���N<aO��쟐�	�?y�q`Ʈk�T<��I	q,�������'�ҠQ�DPب�y�����Q�L�j!�ן[���S]���	7@�� �I՟���韀�SfyZw��8��%��RS��`OH4��E�L}2�'�옰M�Ҙ��Oi���ϠLQ���٢s��ٴ�t�1���?��?�����4�V��ڞ�H-�2=��K�nrH�d`� đ�A��1O>��I)��� �5芅�"g՘7+r}yߴ�?����?��`B*��4�����O��ɲe\��cT��S�J�a��א#,6Р�yr���>�������O���:0a��@��tk�jci��U[�7�OX a�O�<���?i���'�:�ч�+"�I:i�-a��}��Ou"q��7���ş��IWy��'���cƄ>�F��ާ?*��tn��/�	Ɵ������?9�H?��qA'��Cz`�� ^����e�@�h��4�'���'��I� C��n���1z���A��Y�(�� ����������	P���d0��&��C]��fH�^y�@P��
��D�O���<Y����L,�D�D�!JG�C��H�R�rp/�:6�m��?�,O�U���x�4gb���f�G�61��j�'�Mc����O:�YEl�|
���?��'�g��)G���P�CjL�Ie���'i�IV�X#<�;���KS�MP7(%���E~?ʔ�'n��b2�'���'��4W��]x�:t����}n���玃���?a2�L��r �<�~bRh�}��L&m׺Jw ���MǦA4�VƟ4�IƟ4�	�?!�����'���b'��f�$���Z�SR��' |�H�@)�/L1O>��	�H&�P��7q���c��ҶBj�]#�4�?���?�P�I7��4�����O����L\����=V��u�aȈ��42�y��י x"�`���O��ɪWNq�p�M�x�z�����6~7��O&4�.�<���?���и'���[V�N�JĬ�ۥ/	�p<|�c�O��� ���I����	Ny"�'[��r��}1��a.��}��q
�j��"����D����?Q��g�b�Ђ*Q!Xl� ����m��N�RW���'=��'�����0K�l	fJN�w`t�D�;(�4�rM�M��̟��b��?�H�Jc,|lZ)�����l&�	���U=����?�����D�O�"��|���^&�!�M�8r�pKwM.q�Z�ĳi���OE����6G�'Ӓ���nR	�-��A�&�Śٴ�?+O��D��uY��'�?q��jC�ބv��yh��2%��;D�-B<�O��20K$D��T?I�o��rip����f8v�`ᥣ>A��aF�t���?���?y�'������a����WJ�*���ZP����>r���`)�)�SM��q k�**�q�	�>7��7�K�(&���O$��O��I�<ͧ�?A.W�iZ�����K? ���C����_Λ���7�B��y��	�O�i� �m�p�(.N�QQ�>�|���iAR�'.�c��H��i>��Iן|�3��tX��G�x9t}#d&&=BΑ���DƳS0l'>]�	ş,�y�����-03�ħG4\�l����*��wyr�'���'�qO蜚p"
�~��thcc�X��d��Q���S���d��?	�����O~��rʅ�vZ�i����w#�5�P�?�~��?����?y�B�'�$�d@�EѶ�W��!/�^U�S��/V�ꥪ�O����OB��?��N^���B�5;	2�ۃL���8����M����?y����'n�M��:Q+�4BD"����Ɉk�j�h%��K����'ar�'��	ğ�m���'@�;C&��$�W�á�]K��wӠ�$5�Iԟ̒�&��qx�O��ʥ�@�	�$)y��ί;t�Q�i��T����&�z�O&2�'���JM�W`��bBϐ�Iʬ�g	X�A��b�\�	��}�d6�~��#4Ut���<>�� �a�S}��'�DXQ'�'�'�"�O#�i�-k`˘�2�怰���V���	p&�>q�dX�="#��S�'G�x� ��h�3��F�2m��?8`�h�4�?���?q�'h�'���v|0б�DT�@��T�#EB)R�P6�ͼ����O��$�O����O�d�OH����C�L5�qBB�ͭD,o���������T�M>���?����~��.T���G�9�&�J3�'�M{���?	��m���!Đ���'���'�P��qbC�4hT��,� X��d�W�s�L���+f��'��Iϟ��'�ZcF"�qs�Û��]y�!������+�$�O��$�O���O��>�*xr$��?p*�B�O�Ny<�Q�d�#;A�	Xy��'e�I؟t�����S�Z=v�֔�B���y��p���G�"��I˟��I�x�	󟰔'��aq��h>��Фن)9v��wB�ugJ��B�sӊ��?�+O���O��D<H9�DH3V��Q&�R]
P�1L��v�o�П��I͟`����)X)IM�]o������1#>
�Z�>O��F�0{��(�4�?I��?�)O��$J@�)'}r�oa��&1��� ��8N�8�޴�?���?���q~�����i�B�'1r�O��c� �|�
��oEh��!��x��ġ<I�7�6�ͧ�?�/O�i.�	��!~��PL�,"���4�?9��u��IQs�i��'���O��$�'��u36�X�?���w�.lZ���E�>!�X�h���?�����-��΃�.w��[��[f�J�ѳƕ�M{�/�蛆�'s"�'��t�OYR�'[���?�z����L�%�,��l�w�"6D������<�Q?�'?��ɪ^�
��@>;�@�"物h (Y�ߴ�?���?��!7��&�'��'����u7mB^��)�O�Y��������M���?��a@��S�d�'0��'x� ����j�A�Hf@��g����%f"mZП@�Iڟ��	���饟���,�D��d��=F2�h�>�W��T~2�'
��'Qr�'��diqh]���W':B<�a�a�}��vӴ���O&���O2��OH������*�&��)B�O�?�9�&�ɷ)���	CyB�'���'��'�ne�rj�6�`gQ�3YN(y/���x��ۦ��I˟��	�d�I`y��'I��1�O�z�Ȃŝp+����J�!$^��\h7M�O$�$�O��D�O���8	@��oZɟ��w�t�����MÐ�H�l�x�th@�4�?����?�(O���}�x��~B����E���C�s�$��3�P,�M����?A���?�B�O��' ��'��t�#l%�y��\�{���ǆ �A�(7��O˓�?����|���4��IL�Y�pAV���TOd����MC���?�� �H���' R�'����Obo��F��A(G��%��h�j=���?Q1���?����4�T�O��W,�e�,u�S�܊o�: �ڴc_�ţ��it2�'�2�O�T�'���'��A���-T���tgh3t�Prk���� �M՟��	Ny�OU�O
�]�g��UZ�d�~��5���?�d6�O��D�O�t��E̦E���l��ɟ��iݑ��B�3^�.1���K[�,��5�o�R���<ar���<�OW��'�B�2 (�)e
<.u8`J���|�6�O$�0Ƥ�Ǧ����������t������~0���)$�0D�,��������?����?����?.�HyZ�쑷*�|b���J�
I��i�>��to�ٟ��	�H�ə����<���\h��JUΝ(�����`�
М��cM��<))O\��Oh���O���z<>Uo�rz��i���'^;@aI��	s�1*�4�?����?����?�+Op��/M���N�{�;թU�Sî1wѐ)����'��'��'��@�i?6-�O����?p������O�8 �k`�wЄ�mZ퟼�I���'�B����4�'C��ӥ��E��6��đc�5�V�'���'s�"ͩC�7��O���O`�iB�g��-e�
�%�[�|��Q�Skd��Ġ<���OU4aΧ���|n���pD�v�P�Ji��3Iۄ46�<�u�N0ٛfD�~���¤���:._�SҠH;!+�C�̬蔥`���d�O T	�	�O��O���}�'�,2=�q�#UF�Ez�3
&�F�i��'���O:.O\�d��BhL( 'G�f�(�$��]oZ2a��IEy��'5�3?Q� �"bቼ<��9� �-.�x]�a�il��'���c�JO8�$�O��	���@�g���X-X��=��6-7��D�%>���ϟ,�' �ʭIU�E25=�P��i�&POf�n���Lʅ�E����?�������T���h&��H�c�_}��0�"W���I�� ��\y�%� "�4�/�@̸pf^)Y�$���g��<��'���'i�'���'AU�S�S�''>����M���ʑOΉ�yBR���I��p�IIy2#����Ө6ʝi���N��@��P�:��ꓗ?������?��+�r�8�O�@�'압�0e���R�3�0�O����OL�$�<Q,�2�O��5"wj�5ځ����'Z��gcӌ�D"�D�O��d��d#}�mƑ2���"�]aF��D�7�M����?),O���7�Y�����ӕ2.*@j2e�?H)�@	,s�R��M<Y���?y�!H��?�J>�O�Y��b�L�x��A�H�ش���;6L�l����O��IO~ҤV\
�ad�]a��󠣘��M#��?)�/I�<�I>�~ʀj��t+��Ӵ�&}欅`���Ŧ�{�m�>�M����?q��P�x��'-�,8 HTP�8){V��1p*�
c�u��)y�	�O�O>E�	1Q�rQ�� 	�U��\�g��8u���ݴ�?I���?!�G��'R�'���Z4{~�H9��U�C�d�pdK�+T��6�|"+�`�.�d���O��䞟����LZ8��Ek��a�|�mß �J	����|
���E1&	�Â��"�ؐa�1]���'��m#6�'a���p�	����'8E{�NP�DE��K�o˷TG�)!��K�/O��d?��?9��Ҝ@}�\A&�J�+&4y��P=t��x(���?����?���?�,O�U��|���S�wQ� �5fȊ�ʱ� B�_}B�'ў̓u�֤�I���`��c�9�p�@�'�gF�۴�?���?9��>u�S*�P�Ox�!�6}=����Ŋl:*�Ӡ�X�I�7��O>�O���O�M�����'�(Z���=h����d]V��i�4�?a�����q�ڠ%>�	�?UZ�
��R�4!�-�5�$�1��C��M[���Q�ꈟ�fOݝ+S*a�e7_����ܐ�M����?I�7�?�������d��Ok�׶#}PU�`�Y�_�:�l}�f�'�$�/`(|pz�y��D`�0s��*ZV�t��d3'"�m&T�A0ڴ�?����?��'tE�'�)�#?]�1����9�L�C�
�)6�6MI�?H�"|��>���ItN��o��D.�&h�h�M���?�7!th(O�˧�?��'�.h�2�R�j�� 	Ѿ��YV=]4�O��'�����1���!hP�y�oFGa�6M�O�8C%�J�i>��	����ODd��i=M�X��B� 08b�V���0O<�	ԟ��ɟ �IӟCvMڨP��2�"bb�a��Y�Ŗ'�R�'�|B�'b�
E�JA���8us�U���%Ti+%A����OF�$�O��j9bhI�:�Bmza��Y:�9�_�C
^��1_����ɟ\&�����<D.�>�5K�=m�
�� I�-��,��Bv}R�'~b�'�I�B= ɺK|�sOAas����R].�����^ɛ6�')�'�"�'؝��}�����B�)񫌇ȅ�>$v�Y�4�?�����$�!>���$>��I�?�H�@2N4�<"��ڭF̖eH�L����?��rr$�Dx����$�1C�-�0�ʪ5�Z�Ѽi��	!_sv��ߴ
��Sş������b:�� �Vv�bH	Ba�V�'�$!�O���x�bW�N������=h�ER�i�p�v%pӞ�d�O����^	&����)4�Kv��5�.���Y.�lDi�4C�VaGx��)�O�%�T�Dm��l�C`QPXۥ�ܦ}��ן �	�}����K<Q���?��'�2]ѐ �+o
jq����{0v�}R ����'��'�bE��v�z��O��k��o�"�JMm��0�/Fޟ@�I�����OҒO���B�=�6`e�S3ÐP! �z}ҤζK`�e��O
��O��$�<���JC���e��)*Q� d�0:E}`�xr�'��'��OV�F���I��Jq�%٧i܆VV1O���Or��O��$`�����/���#���4qnl��M�Lx��n�џ���՟H$����՟�q��	$��6���WL��`��Y�82|�I	 �	ӟ$��ן��'�b��)&�)�.��PJ��JBt��Vk��5D��ozm6M5�$�O����'<]�O�0���Ln>�[B�	�8}�<PE�i"��'J剏|P��KN|���2�l߸?�d�0wAѐ
���օR-�'b�'�-c��T?�*d+�4��H��H1Π�@�+b�n˓?h��0�i�"꧛?Y�'tP����&����k�r<��eT�4�6��O��䎼?��b?aJ���=���%��/g0]"Dr����������ٟ���?�8H<�W�J�pB<�hx��b�Izb<��i��)h�����a���6E�l k�Û�Zq��A�Α*�M���?	�oE�y�R�x2�'�"�O�	c��&h�)��)Mu���c����O�1O~��O,��ُ-�n��diR3e��L��V�T<��oퟜ �.�$���?1����Qպ,�u��$�P%M����w��(�<	��?����?��>��IQ-G.e���"��QFR�(p���?Y��?��?AM>	���?1��P�Z�V�����������o ��@
_~��'���'��I*A;\��O�@0r6����D�G��;C1:���4�?���?a����'�
�H��O(��H��p���+PE�>��W�������ϟt�I�]��������	�ǀ �8�$	�$�����)�v~��iѷi���|��'��b��R�X�I<��)¢3��5
��@���TI��M���?�,O}@�(b�ߟt�s���぀9'=��S�a�,%��p#bw�>��?�����>�o?̀�-��txri����.�tn�Yyb R�Hp7mJg���'��j7?!�Kʰn�
��0I��p��a�צM�	����Inyʟ�OfIQ��[��y�dۉ���"��i�\���x�L���O���'���2Nz��pN-�F\YYtf	A���ɦ�'��F��'�"pA'�'1�����N�jfܬ"7�d�d�D�O�D�F���|R���?��'H�{�aS*!�xuR#g�c��Iطn;v�O��'����,l�,��Ԃ#vl�l� �C�
��'�����_�p�I����I{�hA�%��H /h�'Ň-�}$�,��5?���?y,O���J�}y�A���4�Y������<q���?Y���'j��
)v���e��Q��XbOD�_�6������O���<����4���O�����U�$��]qM�xAA�ݴ�?i��?�rS��HbqӚdѲ�ƀ ���ꇫJ �E�FZ���I��'[�J5S����HYǇ��U��e㐁D�N���(�:�M�����'V�/1�FO����чi"V���GC:E�2�X��iRY�,�	<Td�l�O���'���$�^��4�S�is�e��s5�c���'�0�M��u�)�d9�q��g�3ڈ0X��.����O���G%�O��d�O*�D��Ӻ�P��{Š�[$H֝B"X��'%�I}U�L���5�SⓝiD��3�JY�:Z����$�
�>6�C�f����O��D�O�i�<ͧ�?Q�Ǚb�z�V��G�4�J�䐦@
��5@ #<�|z��D�4�3�F���p��=�՘��i��'5r닻�i>�����H��z'�4��*`T�ň�~B��Z"Fv�'�:�����O��Ʌ6�&8rw�		aiv��h�~D6��O&�� �<����?����'Yb���h�/���)a���]�Hm�I<I�-�z~��'�\�h��Ǝ�u��3�L�"�@� >����Ny"�'�B�'(�O*�I�Euԕ�N�w������Ϳ\0D6MQ&��韄�	sy�'�Kӟ��1!/�'4�E�#�)r_�p°i/��'B��<�5��ݺ��%�E��74��d�#�>�"�E h�T�)TB��Dg������3^a�Ǝ����8�HB5VC�ɨ'1ޑigb��2��J���!Mh�ɤ1R�A7�V�"��<������Q�Gz�RU���6 ���,�
#Nƀ��b�#�t	;儩@������#*@~}��Ι�M-�H�7,�66`Be� �z�㉿l�
�Q @]�[bvb7.��N�	v� ��f��%�%�3���k��M1�  �V�!��n�$Hܤ����?i��k����@�?V�(U:@�b���9��&,yV�V71 �@Y���cL\zA��֘Ͽ녪��5��i@�b�$r�Řb듗^� 3�ɖ�L6l����>�赯�1�|c?�N%A��p85�B��41�,X]�@��O���.?��]��?�F�6.�բ5�'g͊��<���>1�jїoo���I�(�(!7#�h�'�#=����?q�B-��,I�g�m����"�?��.���Y�X�?���?a��k�ߟ�aV*ڐz	�ܪ�c_3�^��Wm���Bs�Z(��9דlX2͹�(� IN]��M^�q�p��eC��k�l0���+� ]P��qR��MV���l��v� 2a�I@,(�z�~�\Y���?��S�'��V�d@�J%l���#d ��`i"D��9�;	������8�$ �HO��'����8Q�oZ�"�o�[Y�� "�ݾa����!.�O���O����]�p���O���*V��a���
���e
�mʛg���C��Ҿun�-�5��f�z xf�#4^�I"剰utp��6
��v�P�����L��T�T�H���
�nD�}bb��4)�
N��1�gNϷw��($�,�gN�O���΋Fz�� ��$>�|�o�&���=1���Z�(��iˡd��xp	�*uax��ɘA�ޕ3G�T~ָZ��gq扆�M����$��>d�O��\>Mf»>�f8�2�����@Cl�y它��x���t�6��`�z@����҈QS�@Ίq�0h�"~CH)�'�3%�4hD!	9zH�<!u�иI-��$A�+���QG��%I- ���B'qAhw'ҝ�h���G4i�p��*���j���	ӟ��S��A,�c�,�kddi���<Y�V�|�r����U�\X��(�'ў��� Fҽ�o����(����1�^��$���_�(�	X�4��#5r�' �F�y}`�륨�u���A�;~�������h�r�Q���y�W>-&?�ɻ������/Ӭ5"r��
V.��bMǑS�d ��V�&��c�
 �h�Un漐��B�c�%�ǌ]�v�Ra�V�'�LxӚ�7��H��%J��Y�˕�A��)z��{����Px�,��N
�`�\��D��$��=��x��%���ݴ+<���|��O��ԡ�%Ze�ū���&5�`�wD�'.>b�'�d1"a�7z@r�'�'=��ӟ��I+Z�J�G�~E�:1f�T� ��a#дo�p����H�%��iF�?�r��ڦ2)1O� (=qD�D(T�P�`��i@��7��q$��K׍q�͠�FJ2mD�I�lμ0��yB%�%k&d=�� \(8U�)�C'��\b�r� ~���D�O\�D�Op���O�QZP%3fH,d1��!�+W(D�!�$�O,����J�~,R��@/^���3l]�' 7��OR�E��*��i���A�@�u�D	�E�׉֮����'m"�'�"⌿Z��'���1@�4�F��>�>¢��4�jI���W�K���r�
M <(���0
�K���ɏ��F�� s���<c��CA\�gH��aB�o�i���Z�P~�R��L�-R�����b�O����'�(�{K�p`E�R&x�h����'����,�?�OS���u�K&a?J�����E=��Ó�hO�9�!o��m���	���t�r�"e1OXlٟ�'l�\�d��~B����/<��p��D`�t��,і*5����OP�D�O2e��&\H��1Y��W��1l�;;��#�7
~]��KX�2s���T�̣<Y�*�-e��ѕmT�#�H��4T�\B��L4��r� �+W�����/U.�Fy2��/�?1��i��b?e��m]-R6�h��+ �V�2!´�v���	vx��;x�rt�iH�=��P�0f6�O&��{��Lr��ՙ"M� =��<y��r��K���MK��?9-��%�r�OP�$�O6����3 3$����DPxP�h���h�d2�|FxB�CP�u{�']�A�R��f
�3�BPG�)��PA ��_wLIA�
�+#WV�)��
�68�����S��?��Iο(�<�6`�*%�N��g�v�<���P&Ҍ��VJ�3�`�q�'��#=�O�f���".�`:$	!'bqZd�'�����[�h��-6M�O���S身�Ӽc���	�����5l`�$1@��<�@I�3�,��e`"\O��
%�O1�:��d�gL8�xs�3a�����ñ*/�`壞���ɒ�e{�O������8Wҍ+�ڼ�6��O�X3���O��D����<�����~� ��cHΦWѲY#���!8F1O���$E
_�<49��т�b0Y���cB��l���MSL>ͧ��(OX�س ʦ	��L)#
�؂k���,2��⟘�IğX��,v��ʟ�ͧ>�,�� 9�x|��Q�J&� !|�0�#�a���$� *H��L�Tk���Q$�1s�mA��?��ʤ@��p=a`�OɟL�I.o"蔲��1 f���R��!C4�&���	���?�O��/�@���7wݬyy&U��G{���H�|ܩw�rt��+�%�*���oybgȏ\R�7��OR���|�E���Q���Y A�)y��%')&y��?��P1�QKQ@T�g�(]��y*���k�,��;��au�/��i5�	
f�2�k��S�+��`�&m�/&�6j�&�T��D�
Z����#����t@�Y'��'� ����?�N~R�Z"������z&f�X�!��u �?����9O �ڃ+�SҴ���ԅ�2ț�'Y�Ot01t�L�g���J���<AD��0O�Т��]즩��ȟ�O����$�'6��'� ��!+C�P��mʒ)*>\1R7hH�.�ꤑ͕��"��X;O��(����'��;�/�4.�:�@g�(9�E��Ӑ���ʡ*O�C���EV	F����	kYB�J ����E��P�j?�d�wG1b��0��!A4ms���П�*.O����O��a��V*N���o�II�YB5O|�d;�O���@�o�8�)T�X/b*�Њ��	��M����J����{2�z��鐑Έ&�*����?��*�`���8��?y��?�����$�OѴD�Z�A�#�#fFp���`�MN�����[�<lV�c砛�	f��� Y�y�J2�0�%�jݚ��5h��
 �b酀^H�L�$��9N�s�OJ�p��=Y��3�^�Т�eV�����@�[�����䢟؈�o�O<��&���O*��<Ӧ�a����&���0�DC<1��؝��!˞�.����Li��i>���^y�.
�44
7MC�Z$,��R[L􅙁��k�"��O��D�O�����Oj���O��0�B��xp:�˱���d���3�}s�BT9G�nԺ�IWx�0ҡ�٢t���B��	�,pAD�oy~i8���/3e5p�
p!<���Aٞ*|�U; ���<W�p�	ϟ��E��2������+C�(��mR����?�������z>�a�&]�)<�HY��݌r5��o��"~���X���x��M}���2D��?���i2�'��6�<i����0�x�*�`N�MB��v�U�^�X̅ȓp��M�3E˔1�=@�)P�(T̅�P�Y�� V�x%`�?#e̅ȓ=�l����[�-�0��Ǝ�&�l��ȓ&���+z�̍�0)ȢDXȆ�$����g�N4wd��q��#2̄ȓW����k*l�� �PZ����de�8��O�F�HEl�)}�⥄�S�? 4z�ɐQHl�C���.Z�>�H�"O*�y3�ʎGC����(�)���6"O>|���8�d-��� ���Ye"O�]��@T�¹pT���8'"O�q�� ]����Ǡ�`��%"O�Q�4`�\(���"��� ݙ�"O�2Ө�2����A��	�Kc"O�l��O�v�k�!��]	�"O�ho��nBL��`��[w����"O��:�eW2���H2��z��"O�}�g�>yPT�k��̴y�"O���d�����k�1:��kv"O�,�Y�/dX��J�{ƨu2�"O�x�wm
�Hq��3�#q�
��S"O�5h��1+{�u �a
�
���$"O,U����r
D��/�$\�^�9"O��h gN�l)T����s �{"O"���G�5��B O�wn�� �"OtHY�.��4�Lq��OIn_���""O�`Z�#ϗ���xG�%n[x}��"O�H�!��%��sd�%P���"OČku��;�j��#��vW�Mc�"OpI�fd)R�=+A�%�\D
�"OT��$�
��u(�(��Z\�b"O����AW @��s��"s�y��"O��+ub�'Kj ��ϳ?pʬ�P"O�����V�����${B��"O:�@�N9qZ�p
# �/�܄��"O�h�%I�S�1��ly,�(t"O @��G�zSƀ�T��"1L�I_!�$�-g��I`�@<y��D���T!�D	�z 1QdHN%4�i ��$84r 3�U�EK�&�az)F" ���5O���Ǝ���=��!G#��ٓ5)B�R6��A���HT�0A�T=�@,�/���N�Qaڨz�(���P�`{�O� ��ʎ�{F�k��ł���>��&�*2ڔ���/	E��F�}�<��Q>k�$��B>>Tx9�� Z]O䱒FZ2�����~�?�.����I�A���n��y���
Q"Obq(Ў�Ab`�����qs8��aZ�,R�Ï%������O
���m�:\�,��J>y �6S��A��B�5�����*Xe؞XJ�.B23�N$���y�L� `��!|�5����~�,$+A�O��3��%]m���ϓU�(	IK�%�	���
`�Z����`��/��� ��J����p?��<Q�OJb��Q�h�XlC2��6�Z}I�O�t���Q�Z�P)s��4�&�ç�^*���u�O`��1!m�ʧb�n��<�k��~���t(׈z� ݠ�Y۬���ɨ:@ ܢ�([���S��{�e�6$6�@��WN��FTK�?O�%��Q�ᴟD�exe���*D\�I0$#�`�壘�I-|ȳt���OZ��c�F��8	�l�;,?|�51O>�!�ʏ�<˜����.̪60��It�)�~r/܈4�V��Ug_Bx���G(I��-��̔ne��B0��>���g�b�'P���ŕxG"���ՎÖP��Baˁ���}bÑ�Xp�"�(�-ָ�eD�)Tȇ
��̸'fH[p�|"���~��<��3ˇ�� `ej>Q��D{U�3�a�f�R���C,L,�#�(/Jt̓l/桡��\�/]ى��k�����|�	��~2�Eg}�F�^t�I:sZ�s�oX/'��:f�űc���	~���t
ُ#�^9R@O3��O��z򤡟��4�V�,A�1V�U P��1��~?!a
�y0�� ��'<O�Z3K�D�۠)�i"q��ȁu3t9µ�xb ޓ��	�Mb�%>��0HQ&[�}��hΟrk̽!V@�jx��#RH�
M��&�� oh�[�e_?"��Q�aӔ����>!�V�ʧ�����o�~H�˷2(������/S{��H�F��`�R{~��ab߳W� �ʆI�OP�Y"Θ-'�bu��P�4	c�{����U�jK2=�g
���Ĉg,rTY��)�5#�^��q��.1��T2Q�յ{�:��]7���'eX\�à�c^^��O�U0Նė?�Dخ7�\)�()o�"���W-A���I�iHx���d�����ƞN�ŨcM��y�����h��� �J즉�7�Ѳ��'��b���R	U-m �(�M���h��}�<� P�Ɂ�I�S�A�KP�[]`%:V�{�I���'a�@�C��)_c�����"��%b�X���8|O�-�M^�Q�� �PT��)P��*�`E{�'
�j��A�Q�T����~Zw{��b�u�R��8��X��1sD�6VxE|BG<GvB|G�ģ�I�u!TBΊ*�D��eԙ�y2hN7�䭪��'��� %U' ��E��,�Ek�e�+N��	/N�X9��ORt ��M$?��S;n���g�p8@�%Çb�\��1-��<q�[�OEl�"k�~�A��N?��ykf���#��� T�<-��Q�'���l���k�'*g�'���U ��%�;�A���2a|O4��%����"�!Ӵ�p�K�?�t:x���� k��Xǯ w��E@��G�.���=E���*˼E	틗~%�)��LZ7*����6�J� Q�y�S��2mN�u�F��jK��S��y�_'.iL��d'+L!4�2� >����{�X����k�|���ӾqM�%`'f;v�����F�oP �[W$] rj��}���5��"�ޟ��x�¹K�o�m���@��w������'[4<
q�-kfp@q�\3)�(5�
�@,x!��6B�eJ�ɺ>Qj�+yŴH� Cb?����r�I+�D�Q�5V���fߣSN��'�P�ē'�1UG��Xrځ�$Λ=��y�'U}�%�*M�Vu��ɋ/A8@�����@�Mi�lEw~��!�o>���iǎ���M�8�@e�$�L�%�"���*O��5�W E�̥[�$�UG����]�x@��Ԩ̻C����i�(�@ԬD7Bl�'#�Ac��&��`��I�8�
Ѱ�jV�
��	�!�7v�J �`��H>��'.f�J$�	�d�"y�'��DI�KȟKĺ��GK�YbpH�4<O.��cE$f�����>4�R���`�#vΆdZw�	V��$C@��<`�dH�5�0���m������O��d��OR���M/e���aOYTM"�%�0ʗˎ�D(�ER7�X>I���d�?�I&�y�͚�fu�7!Cpq2m��ܓ;мc��#��/�jY���ϤL���˰>?�BL�,�`l����zL:��S �oD�肦�4jfN@�ìC�}��D�l�)�T�C[`�Cj5	��ta�f�wE>��F4!&P�Ģ_7f�LrS�i�iQ�K��@d`p"�^�a�|D2S�6�y�D'�<�`DI�6ˉ'�����i�
ᢃeR�֚iR�H+YPQ�h�� z�&�*䥈d����w4R A
��$����b�4/�`�$0�y�j	�(~i����-�����V�V0u+�iq@���(:�'��r�A4�ER�*mP�15%>?ɦ4O��rV3Y�B�R!@&c��:$�i�Z�"��U��{&H�`c�@٘NJ�`"�D���"N` �'D�C��R2T��TX�0Q��%caH�t&>!`^�Q��9���C�戯8p�q���NKa�Eo�8p��ȇ�8Ca�0l�t6�E}R�	���"7� u�ĳq��8#�0��d�#
�����MuNTA������<��IY<;D|;D��N��̉����O���Kԗ����P!ؼ�k쉿Z�Iq-EdH�ģ�O��,�'����ǡ�4Q����C9*�����8��hq���3?5,9�&
պr�^T���A�7�c�0�d���n�c�gTD�XS&ū
��O��[vIM����Rˢp���a�߿a�4��D��(+]�J��=B���YrA.|���Vۂ4^�˓KIfԒ��p`�Ѱ�]�*�P��lVy��a.-;az���+&��h�!�>{s	��*wB��"��ۯ�����"%�̀0#��I�'^�Q��Ì�'򶹡�i��h�P&�RyrD�43<"-�cC��t��pKF�-�C&�P�����`��tRT����r���գ��a5�C��^���ǁ~�z5�2�ƃ9�L �C+3:�(�ѣ�F!k�z��ϥ�?=��	ȮRk�D�rH�)� 1�ύa{2�ƀC���%�ɩ��R�j�	1dNZ�Ya������~�8$袉�2�ە�I)?8�ɫ�V>���dF:g%��35	.i"�3-	x�&D�&!b�c�S�A���$��e�N�%�O�<Q��_���g�ҵXHa�g���n�~p��A�;�>|��;N�8���g�'����W#�%T�hͣ�(O4Y�1@�<Aq���<A�h�5�u��O�$@<᱇O�8e�X�E�5��(83$��_�(�c�
\����c���wÂ)��%;��+$,�w��
�v����C�j莰@�*�0�ڨҥa�I$,���) $�H���(Yv����S�*h��U/;�%9��M:!�x��7iC�4�f�z5g�>b ��i�d�6�ק��'&�$�:~O.�!Q/ŦyBzPX�ЉJ��s��BLڧ�����O�H�I5a�ry� 	�s�6��GN0"Wf�Y�D�&l��:�f�?d4!ve��?����ȵ9��$S�'d�ެ�d�b���32%٣#��%��j��c���gۂx�i"h�G{2�B�e9f�vA�+��JEL�cE�P���/��EتO�)�ʽ\���$Ӕ�z�⇦߳&v�����ɵ3���y���Y���v�N3Q���{ga˾�hOޡC�kN&l�0\��DD�ju�X�1?�K���7#u* F�F�J�.��7�ѐT|1V�Cf<|����;�,��g��D�V�
.�S��ܰ�Ga��~/��q'�O���7=�%�s�^�M^�lIr�92p(�s��U��)ǔ �s�`�9���E�vk쩈�$Wc��ӧi	�o�L�+7Ɵ�,�b�r�h�|rէ�:?����@�Ы�c�>`�U�l�5ΰ\��ϓ8��٫��/.ם!(�z��s$�',v*��I���8J�W��,�^���g٦P"��J�3��Z�uoȄH�2���	8m�Ιx�� ����L+X�)�d��c!�YF��-�t�"��2�� ��xd��d�I�7�@8uBY�R�`THqNT��*�C�Š�ў�P��|�½ӣV�Nn �]��ȋR���}J��%�ʪ���d�'�Z��s�՝YZ��:��O
����֫����!�ڊW��� ��[��K��J<hv�Y�(��Q3��{��Z�z�� ���F�:�$TkK@�GM�1��,ҰÁ1~���&��G�j1[v��4� <X7�֯	���8T��a?xm!��a�$�A�D���'��9ˀ/��l�|����z@����ć�Hp�H����'/
�̪�(�+�u�$�<��@��ɛ�c3�?F"Ml��cJ�@I��4�3�A��"{"�`����+�t��ٌ�d��hĬ�eH��*�H��@�]�^�htKԊ:F����O����'���s��� -Xh1!��	�~���K�p�� +���ԯ��E2P��@�N�'����޺,��h�h�,$<�X�0FT`;�cD85O.��� 8��ug�'�F�Qw�ó���a	H�4NDAykU����]��_�g�(	ȃ���Dm�G%�Jf��+IZ=	ԃR8}TL�i�d A����P>Q0�'��qH�e�jk2Ѐ&��N֐����6i�2.l�.���H/y�p�O�����Wy"��543r�#�Ǟ�E�@z�o,K2�]@5+����UD�78���ZwW�˓�4A�	<krh}��:_bh��U�0u;�h��w-�RT�hB�'����"퉄FdxL��a� �tM:�C�+1�d��@Ʉ+��	�R�L�Lr�pYC,�)Y����tJ�&]I4���1���h҈��<�$Q3 �
&�2�C 	�fў�#G�fH�`�5��d��'WD��3Ɍ�~� ز�E��};��+�O��)ɇj��̙�eO�o*j����K�6�l��N~�`�H�F� 	�2O=8.@�6Ut~�m�:�p]��e
�(�G���=\�ԡ�
ٸ5i� 
�
�7&�����X?#��F�t��\!N|�.�2iNʓ,L��Q�)��c�E�5V����ƈѤq�	�nr���D7�>�'B��I�A"P�� ���pɆ��p�P�@�t@�G�#4r��Hdٮl�=1&�&���B�/���eʼK\�3�3�~ ��pـN>ͧ\6�òmϫa��8J���)-�� :�Mm��:g�%x$\�V+�#^Ԣ=QK�0N�c)WĲ�I(V[�M�pB�e@�S�GZSd�S�)A�莠y��ئ#�iv6dz%o�@����jaK�
�8�(u�Z�!z��P�>� ����6�N�ȟ�%K�DN�\V�e��惪a���1LI�t��5�a�O�<ܴ�������bH����h���"���0O���u`�I6a2�0[Q�|��e���͒W�E�	U�ْD
�;���u��9^u�Tm�	d`|Gb(N=�jeA���HT.��NS���O8����z "P����W�Ә5^$0�D�	:+����ѧǞ]�[�M2��qsm��l)�XKƃ�Prj�k�!D�@�j�0wހ���3SkP,�Ń D��§�� `��ؤ._"_�<��k D�|�b��>cεs��Z�R��	tg1D�H�7�����##F�����g.D� G�E�qt��©D7mM9�J'D�����A�p�q!Ag��C4�)D�䩐d�d��]IV��
��a�)D�@��/Ŵe�=�U�[?������:D� i�Bd�q�f����-4D������J;8)f*^,7z�i�?D�(����7�H@p�Ɂ�u��E�E�!D� �6�O�(���G��<#�Ʃ�q D�8��@P�,Y��r�A�'	��"u�=D�`�� T�@T�G�Z X/�`1��=D��{��ԨX�u���G�s�A�<h�W�5�0*l�i�bK~�<QR��n_b�"Q�0���Q��D�<١�^���F� 6| ���B�<!���/Iv&���dj�tP�g�C�<Y�'�:0aT�����~N6�(�g�W�<!�H�r�.�YHA������P�<�A"&-���0���� �:�(@�MI�<Yd�.Q/H}�E	s��k�@FJ�<��`F�/��cL��E���c��O�<����IO��;��D(P�~Ļ�I�<��*)qR���uV?>�E��Qo�<��J�m�pH���ͽ)H��idf�n�<��C�OAJ�sD�6n&�ۆkQ�<��J�#h�� �6=4]S�#�I�<)�L/�D�S�3�:-[VaHB�<�� N�v��'�\2cJ<�����<Y��?@.�9���6)B$A�f[Q�<!4����X30�G���,�®�J�<1q,�+V<��]RO�Ekq��A�<��
�)���#��	F$u	Va�B�<���J�հ����[9�1"��U�<� X[���!9�u��$U����"O�E��^��D`U��hW�E�f"O�`��Al�d-v��eZ��K "Ov%�Qi�F� q���C�bT$!��*Or� "OF�O�L�V�� ���	�'���0�kͣm��d�aƇ���a��'�H�yrl��;%H�V�H��r�'t��bW��n�2�K��<��@h�'v|P��dTmv/�7;�V���'@ �%2>D��fY*b�"�x�'���
�c�_ ���c^�R�2D��'@�HD�֤J4��ծ�T���J�'�F�;w�Avp���u�F�D���'��сL���:U-�

I l��':�ySr%`��J�Nٚ��9�'�J��ˠ"L4bSDǹ�jQ)
�'�.���Q+v�^����	{(��	�'x���A5c*v�2�N�B�Y��'�����c�X�T�m�%9�]* "O���d�S$��2F��f���"O�eY�$�94+�嫓g��K�(A�"On���O
bN	SD��(xi�"OԨB�H�C%J���f�tŰB�"O�x�B�Z3L�eycHz�l�ڠ"O��
R
F|tK�ߪ3 �"Of�*UhȖ*�Lɣ7��q ���"O Q��;ij(���K�@6Y�B"O`��Ҏ�ki6�t�#R0��z�"O���"iK�;��TBA��q"�̠"O�%��V�/'PU BY b0a�"O�}��&e Е��i�8ͮ�a�"On�3&�	�O��H
B�>�2D�Q"Op��v�رl�5aL�4�2l�g"Oa�1���?
Xa�ܬ��"O@���/�*Đ���ܐ(�|�[�"O���RN�|Q�A��^\���0P"OdMp`���%�NIRҧ��:�����'��	�
�(��O�Roڼ0�hQ9�.B�R�Լ����'f���h�0��C�/`�DX��oE6�f�Au�/D�B�I�q�՘f��=AxbLk�'T#��C�I!W�x�*�$���`���aC.C��"C�2����:c�`d)e	�"^(C�I�H|��ŇJ�������B䉟1��ZQ�E� �ح��!�rC�I�=wZ���U�.��S�`]�B�I��^��A��=�UH�,�$��B�I�:B�1Ȁ��PgE��]�:B�.[.R�!�D!����ʝ�A�B�ɺ]B~]�W�M�9� �Z ܶr��C��t���C.Y�zZ@ᣫ�(e�C�16�2���mV�NTPӡ�!��"O(���Ì�(�}q<O	~���4O:"<�����i���q!G�6#�J(b#��&^.!�_�9vDq"	���Xi2jD��%�)��<�W���,�xT�%��f���Rm�<Ɂ-&l!����E/0���ѴJ�e�<���&H����r(�(`Q�`�<a�Q
KS>9ꇣ(sr�X��WE̓��=)�F"rE��x׎Q�t�$����<1m�9��J���-;m���dK|�<%�H�Fl���)Nޘ �N�|�<��(��}�P�,%�:�cQ��{�<��hסJc���C%\Cm�h�p�<� h4��ǥl�dM�"�2X��@�"O�m�A#�����H]w�h��b"O����d؉�����S�J�Ҍ[r"O�@�@�
�q)2{b�#+yv��"O �a�̓�&rr�֔
�'M&(1!�D�:$��A����A�P���%�"T!�Vrl�V/�[@l���T�!򤛯J4��a�L�($qb�
`!��V�_�"����d�P�Y��^�!���L�n�%�ȩ�
m-�"j!����v�t�5�'��J%ߺ2_!��)=�����ܹ8����R!�ě(<�F�S��U�\^><&��2?D!�$ՖK��[��C�MK���'M��W�!��M" �:y� ��!<���e�<k!���p�6zYJh���b�+��H��'f��q(�]+ l� �<��1C�'m|$�茁G�,�xul����X�'\(���ĮHi"�^;S��j�'��4��ߠ0����Ѭj�����'Z��[���Xs�+i�1\��:	�'(�$� ǆ�j��3T>2 ��'�H,�S�\�w��]`��ͽ+*M��'& q���+H���f��,��M>������I# tH$$J.+x�U��Q������P!p��!��'Jc���=�
ۓ^��Ph^i�cDPM����`��?1�&G/|��嘂1��e�@�UJ�<�Ǖ�Q���y��;$�Hu�g��q�<���ۘZ�n\�wh�-.Jj�(f!�k�<	�%g��ȧ �� Ǧr�&:@���c��t(&kJ M���JïǙf����ȓ�b9!��+tY$|J�� 	�nP�ȓ[-�����R�$M���^�cT���ȓl����W�'l�|A"Tf_�M7��ȓX�����	�K',|#UI�&M�E��B�n(�F��?�'5�-�ȓT�~�{�͌�]��rf�	1^��ȓO���C�J�U,Ly� H	>p���,�$��P��ܻ0�M!5�̄ȓ�ɒ�K����3q�W�Іȓ>�\�Lê6�*b�ʔD;�u��IR��A�]k�4�0Џ]s�|��?�X�H�ȀQ>x`�b��
�'����@�f$X�4��'�l0�	�'��P���!v�����G�
E,mX�'+й;� �_ݾ�y���~�(�P�'�"���X!�e��!ξDLC�'��䃤eC�<π��U�o����'@�9J�c���{��̄��Ա	�'?��E�������)mZ@�
�'��bD�9J�Yy�H�/��H>ي��i:H=Z�1d�wq��k#�Z�!�$L#�BMx��;h��#EȸS!��9 ��p� ݝL.$i���0F!���\9���#1��ГU	C�4����	�M�Ꝋ�@� <�Tۓ�Ͷ_��C�	=#r���V|*��*�Лo|�C䉶��]��E��Y��2H� 9a�C�	�[s�Y�Q��P��bL��C�IJ������13�,���֓cZ�C�I=yB��@ Q<p@���U7\�<C�	�lt>�kq�QTd���	#�:C�0![zU�I�|��C*R�~�O�=�}� `��kT�S�z)�e/\���v"O$���"['�N�@�꛰ �Je�d"O�g�ݪMf�X�΁�!~��"OR�Z㎎�f�L��_�
w�s�"O�D�` +X��M��bY�M÷"O�uⱨ�Yv]�-�|B~M��"O$��v*@G�5�,�;,�PHT"O�xj %�0'����Qʣ���f"Ov2�/m���"%oQ>�@��""O����M?�X���N��1�|��"Ot����!C��,)�݈z"����"O6H�PD�%LB��O�W;~��"O�	`l�(Q-�]
sB�"��`��"OTp��ְQ��(�W�������"ObQ���!����NL �b�9Q;Ov����+�ƴzCLȍTϾؒ	Lz�!���/^d����N|s%��$�!�� 9��5�.W��� (�lC6�!��fI��0���o��ay��v�!�d�o���e ދ#L�1s� 5W�f�)��5$��W�LY[`n�!f��س�+D�(�%ӢQ	)�`I�%�;o(D�p���!|��%X��A Ixx<� <D�LXa���iRT��$� 1$����-D�@�6��p*2D�b��
w��@�U(*D��A��I��*ΑqA�x���4D�p���˶H���0��Do���C5D��Ӈ�%z�V�� L��w�D,JQ,4D�4����XJ�@#��Y?a��TG=D�\�A�?U�D�P����|Z"�-D���w��^������B�KQ�\�P�/D�xRF�Ƚ;6���$[�>�b�R��.D�����0d��]S"˗,cHh���0D���S�3��LȔo��|
0\�g�.D�|
C� ��~� Q�+:�Sk,D�D����12����n�?;mT�[&�(D��J̘W���A�k�.=��'D�d�$�	����ބX���c��$D���C2Q��ȃ�\_䎔C�c.D���?=h��ʅ�ShN�I��,D��q�K��%��	5KښJ),}�5''D�p��K�}�t�@Sx�����$D�|��fA$t~q��ӱ[���X#�"D���qK5~:(��dЫWQ�\c2�?D��x 풘x�<�0�͞k��4h3l)D��A��ҌQ�B��&�A�k$D�{��ɘWg��(A��+�8��G�/D�h�À�'�\`uꇍ$�b���� D�D�%��g�|IhQ�t4����?D�;�C�UX6b2��L72�1��>D� �Aa�.>�(1a�@�&eXhy��1D�tK��G�@z���舃7��Ag�.D������t�F��y����e�*D���e�:v� dɣ.P�|:�qK7�:D��0�;]�L\C FP�H
T�SR�3D��!�ʜ,��	*�1!j�07&-D�P��Kӿ%���� DƷEz��c�*D� �o�*-��ˠ��(F �
bD<D�P��)
�4\�Wh� t����g8D���3��rDN�c�V�#���� �6D�(�u�F�"Z��r���P�\�)A�4D�|�C**Q^��4gS�TdcS�2D�ȹ��^;B�ڰ�S��eR ����.D�0��c1k�F���*��!��X �9D�� �E��
! t�TB��0͜=�r"O�5D�:�T�6����&U�"O^�
�Nu
b8�$����c�0D�@1LF�EL@�j� ��2�JݰM)D���ָ�pM	�2�6�؀g<D�Щ��S�(�t��ť�y���"e&D����d;j�؃�C+ ��Cq�#D������_� � �B�8a&�� H/D��֠܌=��Ѡ"�^/�xA��*D�Ĳ��'@���>'����*D���p�׋K� Lh�1�����(D��؄  �B�B�# �F�``l���;D����ş�/��Q��[^�C�;D�0�ܠWbvQ�c�-`�DR�>D�|zV�	�w�0�����$Vy�e9D�|J�!Pqdq�Rg�Q��ik��!D��"��t����;5�����?D��k3��zͲ���6Hh�,?D��� [��t1��_?M&윩�/D����%=9
e+

��\�v.D�@�Ù�U�n�GBG�=,�@�-D�X�G�L�b����AW�Ĩ�+D�`��B2l6�d��5f��%�'D��K!jY��TH�`إ7�
�'D��������ǯTX �ܲ�?D�"PAU8rڹ���)'(����?D�L���� b(d�T��֕a@�8D������ D�ڥ��(��4��=�*D���IצjLB ��
Z~n	1SC6D���A��8ff!�A��}�P)�Q�?D��E�DIS%A�@mZ�d>D��0�S:�4;���k�*��e�&D�����\6��1t._h6|	19D�t����)J܌@��}���*D��:���8m��� ��G�P=��X��'D�K��;U�S�`�?hrf�լ!D���茟v��%�`ʗ%�pp�4D���D@Ո\jN��w�/n�b<K�#>D�����F��|�����Z�R�Z�c>D��z�ɕ#x�~uS�	�+H-8�*@=D�lR���s�b�)P�J	|ᶍ<D�Py�ÜR�
D�"CL�p����L&D��Pѩ�:`�-����*O�9k��6D�P��d�=����cʚ���(�e4D��	���2g��Tұm�vJll�F+1D���G��U�2T��!�ch +��-D��(�Ն��!M�Z�\�A',*D�8c��Č}̰���
��J�X���
(D��L RN,Q�.0Q0�1H&D���띢sX�15j�3�����`"D��������*��w_�4���r�!D�\���#D�)pC�ȓ3����R$!D��n]�#���1�x���#"D�<����@�������:dHDG D���6��%@� Z��*,]��K0D������&nt!+�']��P��.D��Xg'�p�5�������8 3�)D��RDi��{�P��1��Y��,D���Ԭ�-]�~����o=Ȩ2��,D�,�+�7e�ű����)�䩒�0D�pБ��w�r�
�*����v�3D� Sb�^r��&bðwp�TQE�>D�0�ת�r��p7�_�p�h��0D�x���]^�У4��~h#�	1D�� ���B�TUǸؘu-� |��a"Oh��Aޛ��{f��v�8 s"ON��"��S m�`A����0�"O�����ǸS�R8)3�9��H��yrc�	"���"bʐ �.����\7�y�F�>S}$�p	�*.����V��y"�D,,��� �z��|���&�y¯�� ?N8��	%�0�	�����yX5���� �A�'�P"�y2���SbȐPԆ�(#�lm�v�_�yb��m����d�3rL��ۃa
��y�/iΦ���Ίe�F�A�M
��y"��F|����b��m9�Ҵ�yM�)M����Q�U�E#�D"$Iھ�yR@�o^�k6`Ű�k�=�yRO��D��}���&���W��"�y"���<F��R�%Ա/�4�9r��y����T@��ׇY�?o�8�NF��y"-CT��@��;?y��Q\(�y'߬X�jD0ɉ1��j��
�yb��@PQk0��*�Dn�y�Ǘ�!S�|(H��7����݂�y�"Z>;.	��fH�K�����y����K��b���8�
��Ñ�yBh��"�˶���.�}#S�Y>�y�m�p����q�ϼZ(v��e$V�y��N�(��(���~�|k���0�y�bKp�P�7%�B 0��y�G�,yR���=@`W*V,�ybl� �R࠱��7o~H���5�Pyr�ߨ*���`S,��>B)�0fDv�<�PE�;�����G�br���aJu�<)�OJ�-�á ,'���;�&�k�<��ѫ
�Ԙ�6�+4 ���קLr�<�A��2zbe���8K��1��l�<���^�y"�/q��"��3mj���&n�B�T8n�v,�U�	�ȓ.��8#�*�\���H�h/D�x*2�Ȩ��c/:?>0��:D��8a�ß;��5�S��"v�v�S�8D�L8'MS�W��` �"�5�dIзk5D��P��/,!�ٴa�.UV��!*6D��U�H�<`�*Îϔ�"ջ��3D�8�.�6	b�	�W팕�`��1D���v��q�0�K2ɉ��*�h� 0D�8x���Z�(ɱp�>N�L qd.D�H@�Ά��bl�ɜ�w¤��+(D���#�W�\� Y(dٗt��a���9D�$v'ڢD����C��Rz�uXp�"D�LCONJ~X���<,��Q@� D�4�q�=�N4ӗ$�����d,D���1���� CT�V*rF�4x7a)D��W�L7qrś�"_<P��scd&D�ș��7V. �xGG\�h{� ��$D��9��]*���`%��rK�G%D�p�#��w�>lk�d�7?�!c�e/D�L�E��:���c�8�D�a.D��3�	\�����E/ZF�
%���,D�0Z¦K��M���� D���� ,D���FjU1|��%J�>R��*�$D���lJ#x�<r6眎.��;�n$D���G�b�(lb�n�	.z�3��!D��� -m��:S@� h�!s�!D�Q� �Z�%� B֯T�2��!D�� q���g��cv���x�T�"OD� GU�p&� �4�W6`�&�e"O���=�LxSc싟Un��&"Ob�b��A=M�$)rD+ՊY�A� "Or)0�_5WtD��۪N�`"OF��%�!�l�9F�ŶZ��z�"O"(,��-˨�Hc�*_�2;R"O��A�
n�d$� `��
�`�D"Ov��@h_�����=KNI��"Ox ǎQ�29C���E�	�7"O�Q�P̳r ��G�� |��]QC"O�1��J�	?�̃r�͍@e��1d"OJ  b.|Rls�*K�y�(���"O�)����L`H���cP��t"O*Q����+��9"o	�^A"�	E"O:����>'"��'��;F��qH$"O0Yb��W1@�Xx�/��}�v�KT"O����#�D��M^$f�0�Y�"Oh�b�כr�T{c��th�U"O^䣷DX&�@馥

��4�f"O-`�jG�bf���V���"O��f�S4.i@=P��?���`"O(�� a�2F���o�l�<�"�"O�$���޳���ڶA��֤��"O� �e�� a"�&�40v��R "O���_�hu059�K�+h,���"O�%��m^&D�r���,���"O$9���7�hU��E��j�k�"OH$Z���f( ��� �����"O8�(O��|D�F�ĺ&��9g"OT�%�!E�di��a�;9x���1"ONt�bk $yN������h��1�Q"O�l١��Vr�1���S�}�&$Q�"O&�뀭�0H�R�� �\k��,��"O������9�*|*rȒ�S���@�"O���A�"M��D��<f��y7"O�uB�H��?*�)� �M���Z"Opx+c�Qq@\q�/�8(��"OL�*�(�� �pM2w�B8� �G"O�`B�Ôf�k5$�>�Z��5"O�d����j2��K��" �&p"�"O�z�A+aA@�RsH�=����"O�-(���. �0)��~��U��"O��3EȺV�z�p��ɕs���a"Od�&���\�-u{��#�D��yr"9v�X@*ܺx��+Ӭ߄�y⭊��v��q�H��A����8�y/Z�Q�8�pp�Z3DU<�!�����yb�&H�0��8?4�q!n��yRM7fFYI�K(����@�ܷ�yRB��"��ri�71�q�
L��yB�F7z��� 6�t��R�ybc�SWdp�c�_Bz`QqU�4�y"g�&.Pӵ/�M���t�O��y��N��K��^�,�fK��y҆�Lx�/;;
���EJQ�yR��g*DEiUɕ�i̴�ե��y��ψUO�T��.�:3V><��D�"�yB���n��G�u���QC��yr$��}�R̓f�N*t�L��c���y���62����6D	/C_<��2�D �yB���1���K�o�
�@�W��6�yb��y�K��-�L��U	C�y�a��1�6H�'z@��PV�ؕ�y
� ��5옹�y�h��%����"O`��H��N�ؼy&h�	?|�`5"O�z�«��M��'Y,��)t"O���'\E[ \��eA����%"O��s&�PP�p P.Y�@yf��0"O:F�tj����� ?b���"O�M� �B8�PI"E(\�sJ�zD"OX��L�l����:BV0m:0"OT!���S�4ix$@��j��k2"OD��E�M*�8����Y�h�
�"O<q(х�] ��y�g�{�R�`"OXa�h�5/:dU���S�r2ݹ�"Ob�;aD|�}��oG>��aq�"OXE�bh
#~�T�V��;(���"O`�@1*\m�m@t�AZnԀZ�"OX��$R�����@���"O"$#A��8J���˗Ĕ�2�	"O�e��+t��-�Td�9&(,A$"O�a%H֎���C�̉48ɩ�"OH�j��$��]�qbEM3XMi�"O��׉Š]�*tʱ!�
!>���"OVQRc��&C��#'��
@!�3"O���7*��C���aኀ0���"Ob���"OM����'G�
S�x���"OD`�@�+����w��:tr7"O��8`��8\ˌ�`�j�(
�c�"O�%c�M�?K��󑯉{�Ќ�"O�a�B�J��a�N�1F�&�#"Oڥ�����"姊�}~X��"O4@h�ü�*@��GL�AV�@q"ORpل�I6I���z��%("��"Oƥ��f� F��W腧|< �"O�����&���U���h`-��"O��d�S��t��$ t� �"O�,��EX Wմ��O�6x<�E"O�ɰ�	�������8s�"O����I1@��Y�GV��`"O�H���#X&�1FkU�LND�XA"O�\@UȆQd왨���)sJ(աd"O�y(unG�RR.9겋Y2=�P؄"O���b�6ն��'��	�Nl01"OJ��&FB�y���\wT�{U"O�Py���7��C��6CBX""O�I�1
��zŐ]B��í=6@�`�"O��ڕ��T��yɀ��7��a�Q"O����I��=�c)8O�<M !"O���ł�*w�
�iT�� �"ONI�D*�!!j��!�gL^	b"O�qӦ��%eaYy'� +E�eH�"O� �kG�i��tgZ�xPdy`"O��$A�N�e��$���*TB;D�d
b�;��Ë�_D���:D�t#m�2h�(k�Ӡz!dW�c�!�$$c������ͫSk�d �	�s�!�Q+U&P��C탂m|���r��"j!!�d/)W�\�$蟍%^�1Y��O��!��X�|ab "��b\d=Q�$ߓT�!���g�l�8�߂	;��Jri�/z�!��e<]���D,��GS�!�$�<�j��_f��|��Z��!�$�#ݚH��"2	b�r@��+Y�!�V�4��E��^�|;�
�)�!�͑e��Qҕ���%u�u�l]�o!�K�.������T:�:Eˌ�z!�� ̅A��#^�h�[��K�p||�"O�`�2�O3ad*"�Y�H��Q"Ot�;A� �N�N�A�*�)!����"O�<��AώZ�h����q�4�U"O�XB/&F��$#sݰ!�"ONa�`#+u�|��e!!i�)c"O%ЗG,V�QC�]�8X�ۂ"O��)�a�c��$"�`�4Lx�"O�%Q�KM�P�,�91&��(2��a"O���Q�},����4r��d"O8���� �sJ��'��oO�H��"O�=S��K�G�8 t��/10�]�3"O~�ICɑ=\��:" �W*D�%"O8m9w�D>U1��XR�]�n�<�2"OPl�Qƨ��@h�*C��<�"O��;5��v��ܣHɃ����"Oab���L�*)�2%��~�@`�"On���ZI3@�q�Ѻ��X�w"O4��eLF�E�hU8�����	�"Ol9��)�԰sQ�h�M��"OBI:@�z�h�8pb %c��C"O*(��g�F�J����^Vp�"O,T��a*YRlۙ8+؜�"Ofѱ��\�bTX�g�U� ���"OM@��:���eR �:��5"Oฒsd_���3��,��"O�8�E�N��l���	 䪍�p"ON�IQJO"naL@���\�7�����"O�K2R�x���Ee�Op��Z!"Ov�X��z�p�9�E�Zj60z!"Oܐ�7-��v�e4�%Bu� ��"O:L�-�s��L��bѻd	�8�T"O�Rv �5Gh`����v�6�"O�L�%w��XQ.σ'Р���"O ����	 �u�ӍD�'���"O �˕GG`�D���&��Ly�"Op���Q�+��҅M'@���)�"O��`反�<a��gg����`�"OV-$�~�,���f�3�zE�A"O�X���Z�P��7���d"O��Y��ʳ��Ifc�'�<ĸ�"O�%�4�[�=#4��F�VZ���q�"OM��L/Ab		��E��X`��"Oj)��ߚ:̤�¡�;{n�D�"O�5 d�[^o&1�WA��P�"O�� �Q���G!	�)��)s "O���&��8����(�8�`"Ov�8�l�-��xq�Q�.t�$G"O���!F6�@pUn�#iN�*�"O��!���; �h���I>���W"Od�1!h��\�ӁG��t�0!SP"O�Hy%�Z"r��1a��jv�Y�"OL�с�T5'��X�e]�h�ڵ(�"O�1y�$
���k�M�$h�)5"O��7�ƫC�n���Ꚋ-��j"O��KR�U�)�qH��T' E!�"O�L�E�G��#��@��q�"O�x�`��"���@f�L	�|��"O��S%�J��$�!��n��P�"O<\paB�W|��T�s��)X"OJI�A�P�@��t0�(ΊJNq9�"O&0�L�D�,�P���?^|�"O���"��Z��P T&�!AҀЦ"O��􂌜�f�j`%Y2_՜X13"O� ��7	�!|rj,�#$J�^F���"O�LCv �P�X��SM�=�|�$"O�H� �S&D��� '�ʄ��"O��A�b�zY�]Ca��2Y�2��Q"O\�!K�vꨱ���B� !��"O�-�E��Wߤ���Hǆ��"O �P��_=f[�в �O�*��"O���*?G1ȡoQ6F�RS"O�[�e�H�.i)7��[l11A"O6tk���\�SG�t�^`"$"O�a��=CJ�kl�e�̽Q�"O"��搾6�E{ud� /u�(c�"O PX�H=Xs���A��/U��%"OJqQt)ƖW�H��b��9�i��"O�ٺf�q����ŋ11�^-2"O 4� ��,h��Y�ЦޯPk8M	t"OZ��2@�.?)�<�'�D
R\d��"O�!�I�V��}b�	<8-�ݳ�"OP�a ��
HZ���Fd�\��"O�����)�t�%+У	�1�"Or�q�ɔ8Mܸ)6k�Kb�Sc"O�B���:֬XU�S�5�2"O��GN��U���b�F8�<mK'"O���o�[��D�Ǝ"[*X�d"Od������ -�$�.Xj%�4"O)c�)�o��]Zr	5Q��KF"OZ�;�ؓBᲰbt�÷L<
�"OH� rk�����g�2N�[�"O�l�!F3N�((�@mG
S%�U��"O䅛wa̒:��qzg��3?���D"O�5a�o�I�6���uz�q"O�<�6��8�`*�'
=o�A:V"OZ�	lZ^w�x��Fwi��z�"O������Fx.�XD�`}w"O ���[�HA^]K7F�7�P"O�dcԩ�=�x�x�$C0g�eI3"O&�YVjW���y&��>���� "O:�#C��
,�-�s�,?
TYV"O���2��C����݅{ ��J�"O`|6��Y�~��!Y�Y��h�"O�xh��]��x��E�;�|�ӗ"Oh��d�=F
=��+BM, "#"Oj�˱���K�f��NPnݙB"O ��rF�?�����"ٮE\�S""O��i�M�����˿.��}Ӧ"O8�YE&�qx���[�<%NT�"O\]����5�D�@�_@8�p�"O�l�רC�]�>$�`B%$Q�b�"O��G��/��u�VAW)G����"OT� w��&	>������I�"O�1z�%��9ə2���E#R"O ��� a3��Y�J�5���+0"O����I*kQ�1���:"͂��"O�]s�A:~�tգ$.K eÐ�Ht"O�YK0H�_���*eɁv`��s�"O���'��?�"|3���2S�Tq�"O}9�oI 	�cˑ�LI�y�"O �kӱO�|�R��*-:�ԉ�"O( ��ԆQܱ�$\�D!L���"O���h�=P��;��;1T�"OX`yA%ӗG4�t�J.n�2�"OL�k�gK)&1|�sֳO+��"OsT��u���(�)�8Q�x;�"OfT��S%$nLأ�[a��Z�"O� ��d�wPBh�)�	�R�u"O�-�;�p@�Qc�����u"OT8Y7h>(���k��{7ĝ�"OA�q&��th�4�P�`Q�"Op�� x�2�J��t��"Ot@�tσ6%8iG�	�4e��hE"O�SV ���sŨ�0CN���"O��1��g2�K$.ֻT3�h�"O��ѳ&�� ���&�W1a�023"Ox�)E��0q�9�`!�4V�^�g"O�LAT�Op���5fK	8�0�""O�kR� !{d�e�#f /�͢�"O�3���#d"E2�J2e��"O�mÆ � U�B\�4�(���g"O���R��Ds�g͋V��Ew"Ox��P�͙^�����q�4&"O���mЭr��D��_�!���z�"O�|�H�+-
ڐp�V55EfD"OzК�@���ʄ`�;O.:t�"O��R��I��.��1.xz�!�$�Ff���_�qK��`�KL��!򄎧-{��mD'B,�2�6"�!���wp�ò���Qn�4Ȋ��!�$��L\�Lp�H�6��pআ�S!�$�8`\�4�c�LC*<3��śC!��s�.��f���� BDBja!���Z�Ha
��� S�ES�AC 8�!�dT�2=���WOO0]�ry	���-�!���-GBZ��]t�Q@Ǒ.�!�?�<olc�)xF��M�!���<F�P+@��88���U&�}!��d���� %U&������F!��S߆H`�`:e��Q1B� #�!�Ă�\�~�0�$�[!iЇB	#�!�ڳ/�<�g&ώz����N�:w!��êq��-Q�(��v�L9
�g�;r�!��
�9�(�`�)܀?j�dz�兌U!�DI�n�2u�܏b��{r�ܻoY!��O�B�+&B]P����R?!��\)Q�``D��WAl� ��$]�!��W	I��3���HWF40��ڿZ�!�$�`Vx� @:J��]��@[08y!�d�.�(!G��-���1��2Iv!�$3�xEA�z��<�6mXgX!�D�w`�9���05���ԌL%8�!�ā�&�``��D �4���k�ai!�d�Na�t(7"�g���ɧ���v�!�$P�E�j`*�ǝR��Eq7����!��=��j��B)G���"Cz��"On�SU(�?W��8�-ũ^�T-�G"O��i��V�~[���t�c���r"O��YP�2/ڽ���Q�6`���"O`]���U?i7��X��ƩYZ�ț�"O�q�k�)!
��D��=��d �"O�]3�fI�.���6h݅x���"O$	ѕ(�'zܔ����K�`��2�"OLp� �K�H��i5�ޱw�PD""O�B�#Џ)7����%���}��"O������ZxYq�Ս0s$�"O�Zƃ�
2a�Q����Q�px��"O
�S@Ք!�	�2c~'扺W"O���lH:8��٨�K�{\�`�"O�4���8��m�檚?\l� "O�ㅧڸh���]��H��y
� L�0�F��p��R��(q|�ɢ"O\���O�2l\��o��Uj���"O�����ԡ/#:V�E$"O$��o�x`:h�	i X5�"O�� D�3d�8k��W�:>�t"O��k�'��g'~�&��.<� e�q"Ov���Y�EP�!Ƈ�EAhI��"Od���-�::d<!6G��%�{�"O�$x���'�<X(�0	*�"Of�"Gj�"��}X�V$v��E"O6�4C2}��53F�?1y�%"OV��؈l�v�h���;
���"O�=�� �L74p��װ=�~e8�"O�i�e�N���qX��l��j&�yB-�``:��U�h����A��#�y�`�J#N��i
h]Z��i��y2 � @��-�ԎZ�_*�� ���y��SL�"�(�$�VWZ)�A@��ybG�nr�8y`)�:L0������y��2:~���4!��V�p������yRn��Q`��#��$UA���Õ�y�ܶ=���E�u��k޵�yBĉe+��s���/P�2�-���y�&ѹTwҍ*��?~E�ui��yb-V�>����H�מ�P%O	�y߮t��E�D��S��hq�5�yBgP���Ƞ+�U��T� �(�y�OۦԶ�����]����y�� �s6�i�ƥU7|���2`n��y�O0T�B���
^,-@�Kƿ�y�e�'f�n$���
 Y�e���[0�y.�R*)SJʈ=k�(iƊ�y�BQ�]v�#� �6��,�t(���yB	�D��]�����:���sm�y��]'�2ј�@�5v"��1.��yrcҳ�t(Q�'~��T���+�y�g��8O��I�n�rol�H���-�y�(-+{�e�@Mԓg��r6��%�y"N��~��$��mh�9 ����yB���}�ݨ�0���!�g!�Z|�L��!�#�@�8��5�!���eV�xx���m�Z#�*
gz!�$b�����#L�6�`%��Py�A� c6��v!��P�lݪ�c�y"��<p��
Q��,ʨ��"N��y$�#����Q��{ ��/�yR�GP�"��� e���W�G��yҁ�)��y#ҤZ=^Pmi���y�;I.�!�/���IQ�0�y��Ȇ*R0
%�H:Tfsp�.�y"�ǩ*��m�c�ڭ|�D��A"�y"�#b���7��;Ⅸ�&H��y���9��mRA�w\rȀ���2�yRh�2	Ø��h�mg(�jUE��y�oY�&A�ԪS��cf|����y��,ZBv��$"Օ`�^��t�$�y2��e������R(�@��o��y΄�P�nА�+�B�P x5�W��y�����$)^\��&��yr`&v*�[b���P���U�y\��Z�Q��?"z\Aؐ��y�ƈW�a�V��c�Z����yB��*����g��1`�Pw���yr��#\HP���<Z�JKfI��y
� "��f�/h�x�K��jǼՉ�"O���k�k�֬�3)�&���"O�#B�5k���Q�������Q"O����b�2u*�b�i�+8p
u"O�U���!�������OJXcA"OZ���-�1Ɣd��"�Y��0"O$t	�V'o�t�0�փw+�0��"O���k��>�2�Éf!v�B�"O����E��.(<@q��$z%� "O�Y�l�B42	Z�Z�7���W"O�I���i��"/�$Y'�d�c"O��i�+$�v��QM��cm���B"O�-�Ӏ	6F��#���Gq�h�p"O )ԃC�P"�O�4q�01"O� ���J>�D�2�� �>�D�["O�t	D���-�1�շ�D���"O�MB��/t~�e�W�3=�$hS3"O��qnV:D��@oKN8�sw"O�H�j�q5X��%jf�BГ�"Od�oĸR�8��Ȑ1���i�"O*1s�_1�2����� 	"�"O�l�)�-��DFg��4�A"O��U��H{j���$\��X"O>���+��QX>�^��B"O>h1��
4�8���ʼ:q���"Ox �$�9%x����ភ)n�E�c"O����i��횴�'g�-ou�]�"O�a{�&��I��eϺ��ؖ"O�p�5��$�Fh���<{�5A"OFm3P@0=eʐ�$�!0�z�P�"O@0�tEX����!1�� �W"OF�"6� �L�������\BU"O�4� K�(�[��ߔ��`�"Oj�I�O茌�͈�@���ڔ"Oh�b$�� �Bl��e��f84ը%"O��e��m:�!�[�ą�S"OD�kQ�^z�`�	w���Z	��a�"O,p%�>	�
| �&ӢX	�M�"O-3p.>
0��%�{ ��"O����?5iA�0�ބ�6 ��"OpĻ�B��W'h��#�U��ܕ;4"OL����?q��!��� $"s��s�"Op��$Iߒ�pA�ڂhB��P"OJTK���)!S���W(��Xu����"O�%��� h��}��%��vVz��G"OJ���YPM4�/TqA�}��"OHm9�k]s$D� /�1=NH@"O�!�e֟r� ��pnO0b���"O�#��B0Bij���+0=�t��"OfU9� ֎0F��T�Cz(�"O< �Bܫ}t�C3l՘���T"OVI��gP�p��5�!�&�kV"Ox� �E���H ��4T�Lp"O,3���)&!�bIX�#Ȱ C�"O���@�4Z����@	�p����"O>�2s�V9��M
���f��lb�"Oܭ�V�`����MQ� �"Ovђ�VL	"V҄~J �{�"O�(�gN׊U�R��"��{�\�+�"O�I�Ҧ��+�P����~��x�"Ozsw��z���;R��0��-�S"O����G�v��H����w�.l"O�%�jU�
��"���C�j�Q"On�QH_�	���!ْ]����%"O� �y;�oA�=� -뢯O�DE�D"OԜ�U�
�5�X�ۡ�0*�"O:mQ7J_'|�p�<!�LT"OXE"�*1�|�K�|�!��"O���r�F"��y��J�/zj��T"O�M���)�jv��Hu���"O��C�eI�m^�p��c%YdA�"ObM�5O�1� ���:�NX�P"O���v�2>;���b?slx��"O��+�
Q��%�[�� ��#�!�y�]�y争�	��/4�ɲ��$�y�n��/���Q��ݫ��[c��?�y���"�tI:�a� ˠ	RBk_>�y����0�2ᔂ��H����y�D�0>�hl��͏ ����	��yr��)��y3 &@�M/:H1b�֨�y≒B��<�dk�{��ђQA�<�y�%̿}x=z�ꍫ_��Q!�-�y2%��Of��!l�&X[�� j֫�y�c
?�*q��Ih
8�iV��yr�߼[��(���U�*��W���y��? bd��׊ІTE� �F��y"��&M�CGBN @@j��>�yҨ��a8F��/L��� �E��yBX�,�,�C-Tm@�g��yr�?_݊��&�<L��۲b���yR���hS�"O�:�2����T��y�ڕC� �C-	&ԣ���y�!F@�FDId�)k��b�+�y���B����ɠ>���d���y��L�#�0q���+z?bı���yb���Ir*6t)�6��!�dȝ��9��)\�uӶ��^|�!�V<g�̕a��4!����Å��3c!��H>�Xz3�A�=6N�Xd� eZ!��&Th�b*I`��7�]�Es!���KK,�p+��8􍣡�\n!򤃭&���5�b��`�I�,5!򄊊@W.�Jw�P���t��C*tT!���l����1��)��̳�׌[L!���Ux�K��ո���ţP0x�!��'�L
���4�MHP�R	E|!�d�,$*j��"�ř����EMԏ0Q!�$�E������ؖ��L �D�!�G� K�%�d�T!$L��!�ρB�8 �C�S^b�X �
�}!��DI�h#�J8GZ,��gغuo!�ĂA<���CiJ�lN�-��Hp!�
%ul0�3�IM�q��Fn!�$9Y�bT��-��d�a B�dk!�$�w�`&�%I���kGAX�!!�$�G��$��>Ĺ� _#�!�dV�V�"�"�䕞4L��R@	�\�!��*ϲ|��n��JH8(I$��!򤔆S��%�P�3z7Zm!"�
:!�C=ܴ��I��-:q#n[�vO!�d�>-GZ%ps� �dـ���$2I!�J2N�92�b_���{��6'8!�d���e�Ū'e�@8CA]�@)!��UR4�C��?��Cwj�-$�!�D�7\��y�� �o��8:�NO�i�!��<5�zcC�sz�|2U���!���	Np<qEB>t��r"��>�!�d�
j�[��*F]@���<�!�� ������V����?���p"Or�6�J���� ��P~���"Oz	h&�$U}H%�R�):Pz`"O��r���)�2`���!yU"Oz@�d
˟^� �FN%>�H��0"O����b�UXTt�@d�%f�U�"O����J|������p�"O�%"�A�.�NQ��a��@x8tr�"O>Ӏ�]�[� q6?s8A"O��9Ꮗ�ESd@����?P����"O@�Ǖ�j����ad�T�""Oj��֤�7l��CoǈFy��"O�`���I�$,�"o>a�I��"O0x��A_�zc���6N׊ZDɰ"Op"����s��#F��pH��Z&"O���o�lռ�)���=�L+1"Op`�7l,m�Ј��M��,�p�7"O$ A"џ�ti8mѓ�*�p�"OP��Fi6Ej(eKX3c���"O԰����/-�4UbD(�@�hLR&"OTYs���;E�sT�<�*���"O L���	�P��uO��=`rA��"O�|�DKĠi'��2 �9c쌢�"O� ;֢��g[@�cd�M�'�
�q�"O:< uG��:4m1��	8&O�H�E"OF��%ɘ%a�Ę�P�&L��9�"O�p��J,^��`ɢ��(AA�ec"O|���:y�$t*�g�%Ӻi�"OlȈ�W2����RѠ �"O��:��D�J��r"VVJ�"O*�F雯W�9pλ�،�b"O8A��fجs��hcPF��"Of!	�����qD_�q�>�:�"O�kT��nL�F��B����R"O�%�4K:=8� wA��&�V��"O�8A��� �X]��
 Vlz�� "O��x &��xL�cJ��T�pe��"O��y�蒥��Q����Q���"O���&��+��y�+�R_�@4"OxE	ǘ@날(�	  �b��6"Od)` ,�P����i�	-B\4!�DbMNj�@��?���s��F�{ !��I�D{�KWb\�Q|RتaDQ�!��X ����,B�8���J�k�!����3��IL�ڄ0)��3!�X�7�2���0{�V��g'eK!���.y�Ը"DEG�����'!���v.)�چW��(��!s!�Dңj�Eb���~�ЋpB�i!򤈆ckdyB�!D�BxZ���:I[!��K�q��bD>I�c�� 1X!�'v
�¥�V�Gxq�U�$�!�$�,֜�!q ҏ;�ڀ	�l
.�!��yb~11�
$dԽJ�+ڐA�!��;B��%!��t��	��s�!�dU6;�<�c.ڂ���]j!�T��� �e۔&0��DZ�@`!�$@/=@��:X����󃌠kD!�$�/�ĕ��o��X���ۡd[�}.!�d
���� 'wN�bٜ+s!�d	���]�C��.b�1b��6�Py2Ν�Xۈ9+ 䔿w#���5����y���@F��mp���j-�y��	P�se�c@��ڒΔ>�y
� �0��S�,9 �S��Z��p"O`�S�,Dze����I�0��'"O�Tta]�������+,q8"O2h°�r{~qr��8����"O@LS�*T(���X6Y{h严"O�D�1"�e�Q�߰��I�"O��a�^0G�	�b�$^i4A�W"OZ��lTx�*S��*@i�"O*A�Ch�?vtZ�0!�vA�x�f"O$��$嘘+8�T��-�/<��L��"O�y��"�8=����ʓ&��T"O�k� �~1B��ͥGc���@"O�K�� CܨU��k��GJ<`�"Or'�H>2��C�l��Y�r5��"Oڐ���R.l}�P��;����"O�(B���>1՚�	��K���1""O�uq2$�R,$D�G�%զa��"O4@�?���ЧQ��L%;"O0�D�O�a����@��W�|I×"Oμ�p�J ;��{�l��~���S�"OB��R�U�1k
�Nu��"O�H�$i
�(&r���(� rJ�(��"Op礎�����L�2<���"O����vN��812�ݺf"O@M���Ÿe���7
�Kf��"OX-� �3n�n;���&�z���"O.�:4,�7i��,r�J40���A"O���$�� ��:)I3B�V}z"Ox������ɘ�5���"O��QB [5@x:�Z�a�'6j�q�0"O��!/P1%�F�
a�˘]���"OPك d�<�0��/U����"O� ��+̭Qn���r/�_�D�z5"O��ȷ�Ӊ�V!cNR�z����"O�]AE��63`~�E�&?߆��F"O� �ե�%%�"X�6'X�a�BII�"O�(3�:$|Z���@I�cݚ��"O�l����W�&UX���*�l��"O´3A'^<�>]�V ЃE��`W"O��a`�*@�Й��lP�}�"Op]�%�ϐ��Q˶$¸q�J�#"O~�('��U�؊d�׻&���zr"O��(�m��
%��8���,��D"O�|�����y�M��`ۚ�Y�"O*��h5�<����-�n� "O|03M/�VMi#��?��Cr"O��a�F2k���u��8{�*A��"O�l�e�ZD}�!������"OҤ+�ӎ��h��`���R"O�h�f�1M��pS�m�=@ZxX*�"O������l���Q/9jB��!"O�R��7t�ޭb��	��\��"O�a� 	@S��!a��R�� p"O���ذ��,����"O$���� K*XhcA^
�1"O�]X��E[��&��D#��f"O��K�D�jT���5Mg:��"O��R�K�.�e��ΐh.��9�"O���Ģ�	��µl�$z)�؁"ORE�V���J2 ꡬ3+�>'"O���3#��%,p@����;c�����"O��S'�،�H�;�L@�K8j�"OɁJя�Lx�Ce]"[�řF"OB|h��K0F�4%aуW�h\�@�"O� ��2W
(:�����K[���"O�ahP�=-p��2����wI m��"O����\�Bs��#� M�[<�m`�"O�8iRNS+ t�ɐ��2_%�}p6"O�� �Y#Bء0��)���"O�,���H/4;��%M�Ptj@�Q"O���pi��N��K�n�y���Z�"O�I����>8�dN�P�Rk�"O�$%�S�U���#��]�\�l)5"O��Ri�-r���`�2(���
T"O�p	C@`В$1A!O ?�d�b�"O$tჯ]l�!�So(�>ȒA"O��ڳ��(,����!C�d$�"O����@&z&& �$�!����T"OV��D�I��|Z���Yv.��T"O��� k�p�Rѣ@!M�Cq0�@"Oj�ҕ=j�~�RVO�,z1�r"O��3N��Bң�'U��ۣ"O@ٹ�LL��Ȅ�L>ELH��"OtT@%�E��<S��̀ng��s"O� ~��0"�3E��`u&�3!�d�=B���]�W<���`�B<�!�i
�|��N�
4�2Z$ĕ�^�!��  ��M�vM����A�}�!�$O�|�A�'ۥ 4r�W�V�"!��
U0��9n��a�X	!��ݻs]!��?�,�r!�܄�8K,��q�!򄈼Z2�\p�T���8Q�T��!�d��54x9SC��A�|�Z�)K�y!� _��$Q�b�7[$u���f�!�D�	j)2pcsˍ��:Ԩ���f!�d�6۰|q���V86��Ǔ��!�D�5&lJ���!6��@1���$a�!�̼\���� W82�
�����z�!�dC�n xQ�삣o]"]q�%�!��ЕKS����ʹ3����ǆZ\!���H�;iZ%F �e��[[!�D�"9^i{q����HR$!��-RF��7�]�n �	�=>!�D['V���� �"*�<U2Wi�2
!�tP���J�|��1�G��BK!�ę+!�x``��dڪp�7���D?!�$��n�.�1lԀ~��Hg��M�!�d!&-�����T��mx���''!���@M�q#��9	s$\��� C�!�$(8af�SEW5{l;`��	n!�.]��CLҊ$`r�s�ƍ.c[!�DN�s��IR˃�6I�-��'�!��g��ِ�ѲY�`բ�f6!�dF22������e��sD�@7�!���v���8 En� ���!�$���|�WҩK'\�3t�)k!�$B=:O�G�R �uy�Dشw!�B��n�3��_�Z����㔂0?!��X�x� b4ʏ>`�Q7`F8'�!�d�=lE����bK�Hߠ�Q�
�;�!�D�1($� �8Ҹ�y#���J�!�d
�B?���QoY�@�^�
�f�J�!�$d��	�`�l`SB��8;�!�ă &���0d�&Z�����2P[!�䞚�
D�d��0����w�U�@k!�DK�u:ԍ#�h	;3�tdX`d/�!�d��w�]�㊡`�Ұ�m��e�!�@�%Ĩ 6cҁ`���G��-,�a~�S\?� �Xqq��+�t�`��X�jY� cq"O\d�A��!��}�w.g~�p��'��	XyR�ہv?Э����Lt�0sc��q($C�	*�r��D�m��� �ݙQ�V��$p�6"<qS���R�����8l��1��Il�<at/�#�L�bk�-� 3��`�$S��HO��00��<]� �H�"@�J�P��IR>�c�bU�(n��o��-0P�9D�x�d�*��d��SІuB���O6��=Q��>���^-4Pθ��#� �����f�<)��>�N�R�*xWH���̓^yro xX���2�2T/���$	(_���Hg�/��~�>�+�r�T��O5��B��?�1"O��('� �@{��K�t�u:�"Of�*պJBx)���4t1�a�"O�P����	� �QÛ�/�щ��i���=�	u�	Z��B�m����K/L+�A��U>G!���"�}�!A��Z>����k^�B!��,X�t��v�N�
��Ԣa���/A��G��,��I�&U,Xm-9E�� ���"�S�O�r5CU͕/��lx�j��KUf�	�'��f	V Lb4�@��*IJ�9��@��y��S�. �B�G�N�U���?���$���(OLjC%�o�@���;	�G?D��S�GT��HR�ץEW�l�sL}��	V�S��M��EE4�n9��@�<4��6 _`�<��!L����±�ϛ/zB����<Ɋ���}:й �@!�1�F��'!�B��/|Z��7�?qo�u0�`�-�XC�I�x�s�ͻV�2��@�T�K� ��G�'yў,H3I?���A�dP�RJ]�!�$D�jn ��"��G,��_a!�$r]�(���B�f���"��-`!򴧖��v����M0,�J'�[�<���S�&�����g�&\��քr�C�	�Uـ�`N��@ a��M��B�	xh1����A�j�����;���<�����O>t��Kíwy���T�+)�5c�'�T��c��P`���mτ� ^ 6�K'D��dl�:y3���/ҁ.��CW�0D��u���]�4倳��i��X8T�����D+�O��Q��D�]�-��E�:9_<��\�����)�'�(����{�	����^���ȓ��� #v�2I+b���YC�'DDyʟ��w�و[�t;�
�_T�+��'���� Y��|���)	��#��(J+�c���6�'f��ۂ��G��TL560y��(O� I!�	(�D�i�P4�`)0��I� ���)�9O>$"��J�LF���5C��@@ �'Oў��6�F$.80հ���-��]0#9D�{��߽f��+C��1C�x��`�6�5�ڸ'��1�1M�-��a�"+6��ۓ�y�1O���J�q��P-�&d*Uώ�o�����I%w(�D��愀>��\�BGɝBu�OV󓓈�����J�E�h(K���d-�yĀ>+!�$I�
�Y��tJ�!�J�)�?�F�Ӥ"׬j� Q��	�I��'5��녆ݤh�i`G�m��b�4�~b��s�.��ҧ���@M�6�C�L���b"On��`�ׅ*�I��̆� t"O
�;�&��{��tRH�J]i��Ig���Ɍn8B���IđC���D8w ��h���:3K0j��l"gl�)�(����>���S�tU��Q�����a�ML�!{@B�)� 0}��D�^hԀ�,Gxo��{䑟p��X�S�O��S�K��K�� �fk�t��'~�Y{�g��G�N$�e]�a����'����E�D�u�#��P�k����
�'t�tB�xU�\���Lw�f<ҳ7O<b�"~Γj��a P���F_p#��	�`}r���"Ɉ�25��N�e #	�2>Z��� )��"��44R9�2� .[\<��I�<�O�Fτ�+.p�����B�"Oj]��A�X�)�.
/���Q$"O̕�$ �5 ��zӢ�$&������"��F�'p�6���*ӢGQ�����a�qZ�'��$4}J|�>�W�Kbm;��o�j�@Hc�<�d`�|�����-P�� �B���y�<�C��B��\�G�	�kD�٢��@�IN���O����T  0�j������ۓʸ'��9Q£M�CaNlJl��O��DJE6�
%`��t�����"O��k�&R�fx��Ӣ+���yv�'�ў"~�5�d!V%3�b��E3��	L���?�V7�S�O�2��R���0�<8���w���@e"O4����	B������'AL|��p=q���)h�� �4"�pe2(*���x�<�5�ͪlB<XS@En��L��*P�<���4D���e��1��`�<P��*�ޙ#�DX�K��� �̓٦�F{���iP~���/X�m�$e�V����޵��'ժ�@�o�>�bMд��8.,���'�X�+b�:D��8u��5R�A��O,=��pe��S�Z�8�Ӣ⚑����!�rC�'�����;�ɐW�2-�ȓ4���*Wj	\$��C!׵#�~��ȓ%��r�n�!�b����N0j���}����L��q�h/� ���4���05G"��7Wi��'^$��
O\�x0D2y�z�B�CĈ|TB�I�c�
�z0`�>w�^%BG���w�#?���)N7"����F�P��,��*�+�ax�W�@�<q��&5�ޡ��� 9h�#`�S�<1`8@ȩ
���oBEj��Z�<�a���O+H�)"�O�"����Ũ�U�<v .E9s-ߟM�1FR<1D�iY����h�	hܨɢs`I�3���	�'>��Q�YlY1�/S-���0��$-������^�T��� 䜙P�Ҷ�Hqu!�O̰��COT�X�r���P,s!򤊃uo�p;���E�@�����VX!�d�>��q��M�1�V���dR0;�'0�|"cH*��*����S�`!rGB��y2���Qze�F,�C���r��Q&�qO���Ĕ0b��0���lg���r�)(!�:!�"9s��áw�"𫶉H�4�!����0} &�W%g��k��Z�S�!��3ێŃ��+TH6�a��_��!򤜑@��P�$>^>|��B�F�%=!򄐚6��A�w�-�t�7)7l�!�DK�-F �R���Cƙ���S R�!�����zc�1�TgC�F�!�$�8rB�\�F#V�HW�x�LX=�!�$U�R��q
��4ni�a��'�!�$EH��s�%V0y��5�P�VP�!��Utd4�r!� ���;)	*	:!�$@�;q�q9��C��m�Јʵ=!���/��G�_)@t�bgE�R�BC�I$#;��A�D�*X�2x8w�D/|�B�)� P�����+�<�SP�ҥ�z��p"O�y��b��D�^H ��A������"O��5pQK��O�pmٰ"O�P��":=r
M���:Wt�G"O�9Ȁ��g����#HX�BD��'"O��A�I��
�'�0�_�f�!���N:��Z@�M��|�#BŽi�!�/0&$�c�����e�Z	�!��f �t8P��#Hvd@�GJ�a�!�d܆A���"���:�Ή궠��!�&J����)F!2�bX��%\�{I!�J�w3���S���B��*��ЩeB!��5%��l���6�`]�wcOy!�1G����Hs��$ң �[�!�d�lm��Ba%	~|"%�R$�/Q!�ݯ�����:�\,�s�6y3!��>Uzt�ϑ�	�]�|�!�D�i��HRES�xUc�''v�!���.A(�ѥFB���c �>{�!���L����.��
C�!R��Y���xb��8��뢁��CŠ�j��t��Ҵl4��!�'�ö�:7H2D�lr�Ȼlu*�g��7mz�ӯ=D� �a���~^�9U�ËT���8D��*E% i[��n��U�ԉr�7D�T��nE#TvnH�q�A�8�"(��6D�4H��=A���S�!�\m
ԋ7D�;��_2X|�U��01Ӈ'>D���DS�W(��1v��^E���j0D�X���N$c�}���F�T 0�B2�1D��qmW1�0�{��F�Q�F�*�b-D�� ���6g@:����s�NQ�&
*D����R%0^<u����PmHy�%D�ʧ+8�̉�7m�.ysdd!D�0+���U�
��U��n5@ђR =D��z�m<.H@�`��*m
�)D��BN�)2w�Ex��Q�R�:!J@�:D�$B��	S-~a��d�&kF,��/D�<Hw.�>Y�"�`���?\ĲgA>D�p���˺e�:��UO�(`A�4��9D�d���<02���(%��G��!�U�w�b!
�eÝ?��vnF�d�!�$� Jl3Ф�4�f�p�׀&�!�d�5y��x�LԤ[����ѫ\�!�Đ<��c�E�:d�.����6�!�$N44ކP��3h��$b� �C!�$1U���'C�)9��	x�o�m�!�]$�9ۃFݦm�e9w�$(�!�DS��MR��i��y��{o!�D�$B�d����eΕ����!�	)N����IK�S>����2�!�dɣe|���5�	'JE��U�/W�!��Nm�f ��ƚiI�A׌�R�!����5��(I�%��S=� �*X~�!�]p��YR�G-c&��rĪ��!�g�� (A�\#dţ��U��!�䖆`?��J�D\tv��k!ˬ�axr�֚%������3	Xd��(��Īݒ�Ҳla<��B�1D�$����c0~kթհ|��Õf�>���+O���[���.5P�z���(|~�3qhX�d��`��� nϲB�I�#�L�WeȆL.¸��F�C�. r���xT�`��B��xi�y�n�?ջ$#�I$AR��#�,F�����s�����^��N�[t�#�n%��/���!aeǮx$��6�#H,,��Ѭ�Ur��I  i�Q����Q�H� �e�P��i���C܌/�L����m��9��A�.�.�j`�R$Q;cF&	K���m�!�� @T��cE�Qz~lB4�\8[2�ZԌĄ6B�H�$A)ޡ�1B�@�Rt����	јO�󮒣Y�t4(@&G&�(w��::�Q�����#Y�?��T�>%��ڲC�31�>�0C&ԋI�:�#��[-*6|C�n�6mP��B�&���r�Dˏ{/(,ۃB��Kx���[�-������2<*@l�O2��(���ĴT*A��Ot��)��	�����E#^u� �D�t��1 �k�z""BTj�t���f�Y��O��M�*M��(S�!X5������E��DQ��10��(c���LdNH���jvZ��S�I�:�`Gg�8QB�zB'��L8�͡B��qH������G��A�P郃?¢(�:��ᔆB��i��I� 9ɶ	��ҨN]PT�>�뼳�֏"j��g�1[�B �&h�a�M"l+�͑*�p�0a7§_mdyx2i۫+�;�Ǔ�R��e��#����"�;Gs*�sU���?}hb�*(�ȑ&lYBK��"A	�2~b���Mm˂�q$���t)���Ld�b>)����;Na��ن,�/�X�Rr�ץV=@���䖜B� ����/ mly*��T9N�zrnI;n��hh���zb�Q���8)搠���3����f^4\!��Bn	;n��`p��L�}b�e��bA9+��ݺ5�xEd�h��p�Ŧ^�#���$�4E~��:�\+ع �.���6'U@x��@�;/�H�z��Ҡ=mS�D6=
8�����)"�>⣡�v�''�7�ǲ,�T�3#B�*L\԰�D�Ș'NZ����EN�f�r��11��idG�"��u�e�X7)Z�)5��Af �@�\��a���U��yD'G���}�U� *d��}�x5-�-{���/~)Kc�њ�|�d2U.��!7�\�Bbb�!f�V��>'P�*�2b"EH�M�!�^�K���)D��s��a����dJ�?����Ц�5!~�-���()'�|�shX�
a�hsR�#i萪��>���P�J7#~���O*-,�T��C+4٬q�.�e���)��y�nC�g���֤Ϫ�*�j��¨}\�s����^U#T��L8�jX��E뙈v��1j�*#R5�sJ��T���P׊�#�HdXB�����Dh�1(:,@�b�u�D�C`� ��N�$�@� '@Cp�ezv�G���D� ��T(��gM�<	<�j�^*/ܪ�	�@$)�J�KQ��S���B��eiڢKT> (c�Ȼ�l�7 y��?.ށ��Ĉ���HہA�5Yt�x�'� ,3��F�A�f�ac��s�:Q��159�%�杆��1r�E] k����#��	h�A�1(ߢ5]���ɰ&8�"u�I�)�റ+O �P���OEq�G�?]t E*�~�����Qt����Q�`���y��V+G�NP1Eǆ�8��e�Z�\s	Ó:4�T�GID.^.�P�rƛ	r"����J� h��B�(p��T�?�0���@�i-��z7h��A�$D�p� H�H�b��s��+$��2�X�`�<G�ȓ���M�X�r�N�B~2%�.���%B��l��g�{W��OX��8I-d *
+�Ż����Z��4b����P�ݾN�lYP�:L&~5`�LШ&��Ob����ď��I��#�/�ea���?V^�ȇ��%Z=H(�H>���\2R�0�&z��S��!<��y�A�: ��gȦ#j��3*['W��#���}�`*��1AxH!�5��G�𰢞2XD.蛷4�D���M�/��$�lH��h�T�{F�z�����$��e'��`jN�+��Ũ~�ir��q�'��0��+x�@�H�"��OK9i�/K;^&�fBX�pO�l�4+HT�����ák#�b�L�J���Q%o��_&��B��tF�x��țW�����C
��E� k
NTZ�A_����B�����B�1�bty�`�d�>(�m ?��"A#�@0�ș���!�5�L�UN�7M��5F��#�@�a��ɵ93N0�,�1g5{"�T����|龽�u&ެ+�<ĊR�L���A��Z9Zm���¬B//��Ж'�v�������`CCk�/p]��ۆ��+3$9�S��?	sV=�����MKSF�%zx����)bSl�
 m�5TQ���z�� nX't�\�z��޼�(��O ��" 	��y�`@ň��M`��9}'\���i � �!W:Ţ����"!�������Z.��'�
�<�)��_�DG��SEO8=�B *����4h!�˕!֠>��t[6��\�Y��B|n	�ë��dⅧO ���W�m��Kw�J�Uׂ�+�6#�򂦑�U:0�'/ڄ�s�D_0@�`�Զ&^܂D��>���Y��KXA3@��8+�+�8��6�ȩ"uVԠ*΅X�P���N�*n,��ZR�D�?��@ȵHD�	� ��F"Ȩ!rFh��VK�f�69�L��K	T�ʄj��z��� �(!u��`T�I������	�y"��OHٺd��~���H6�Ĉ?-@���IYjUr��tJ��3U<E����4�'CYt!G���:'T��O��Zr.�p���4��@Zt@��E BX|��!�Ir Hx%��h�]�p\[���뮆'W�J0J��W�{���`q�$CvI���h̙!�Α$��PX�G�0a�D�#��&?��,��c�2��'�Q81�������\!F��
%" P�5�
�(pK�f	�7����\�5��M6n��y��Њ% &|��HQ�
�$la扜2��`�KU�I�a ����z0�9P��?�􀝇s
��W�ÙFг՜H�q(��x	6�) �:�L��t���u=�3l�i�x-����%h�޸Cg���:�*��V0|	~I҆.8q��L-j�p9�W���n�ĈG�E$ �"��cA�!1��Q����7�\@
�k��;�����q��LHOE&�6���!<������D���2
�Yk1�+h��,#�o��O���z#��4�`��V���$���Ô
Llyr*�)΀���o�C� �H�'�!E�0bG�7d��cHR�VtV5
�K@�u@`Y�ሺD�$�H��T#@�*�ė5f��C�蓄PUk$o�>q��a��U�e($a�p`�7B�j�G[�����T���Uo�q�"�P�Y�K(�C�?<�r@z���8R�eiw&¥==���#����T��[�wj<h����>=�|L�Ͷ8Q�]GƂ$?;mC�.��qA �F!��6lU�M{�7*�4��\Ō�J��EZvyò H����e���0v<��D�/n�:�쁉E
�p ����HG"y�Ҧ!v��(� �5r
 �4D�+i�"����F�P@�i�"�򷣓������J05 �y��Ҫ|3*!b�L��W�0K�#C��6��g�"�M�1j�c#nHxӠդW��	�X��ƀ�~n�p�N���� �~`dȧ!�D)� 9`Q@~�/�@�Y��������/\�q��� ʕ�4��yPi	)h��m#W��	�D��N�?e��Z;ST\ ���:���9,y#gK�r�1s��[>�Z����s���'6�8��N;v�|��3��<e�&Q��@҉uU��@��C0=��+5�L;�ŒE�#  ���]3V�ֈ��
���P���0<��-c�,͸���ծL��M� 0@��"���%�"�+u����'.��i�NP�](���GK�|J&t�B��)��)s��ٷ��9'H�X��*��Y��Z>�4yy�F�	@��:QKI���l�glP�DZ�x��Of�}�'�e���lpr��`L�.t�qc�P4Sѡ��Ŝو���4�ASP�jn산X#j�Qcж �$HmC�x�B���L�t�Lp�v���w��=�\��'��M�RekĢ-@�L����?�M#���l�V�����2t΍��/�����f�D�Y����;w��%RJ�8�F$��߄)�7� �@����b~P�pm�T�fCҊ!&���Q�\�Dh��
(̂Pf!*r�O8���J��H*E��@�%W�'��Nǩr��!�j1���/�t4z�㜘~^��1g�T�2�	rf�e�ƝV"�T�ׇʬ�������Q9̆{~�Ȋժ�;~ �ECL�L\a���^����Z<�D	����G�ayRh�zҲ�Ɂ(Q�]%΁��� �f���-����%�9Xl(Qr(8xբՙ!hP�X&��O�@-�� ҨP8�3V�*61~TJ��T2��>A�(�3}:� �-�T�E�g�:`�YhS�B	�6�U�i��T:�,A�e��'k<��􎘃}�ӓu�4`��LS�+��0��\-ǖ"?���$`�<h����L�h|�DɻP�	���¸$����@՚\�$`v_�/�>�o�4��j��^�D��Oc.a��7}""؍0)�-3���j��=���B��$Y)�d}EзS��8!�����&>q��2`��R�Cuohp#�"a�&Zq��*0� 7&Ǵd]*�R`8��B��֞2>zI���؃B0pc�-!f��#xX�)0���1{��V�3=|E�����js�=�U��$Vl���%����������o:ę�ԡ�"JU��oG;7�nԑ�+Ldp�At���Xg�|�pË��.ť�|�)��G�S˺�0u ƹb� �5�	9T8�F-�9�=�v@��E8[�!��\�.H˱ǔ�E�p�⎙Dȕ���r\%S$N�<Q��Y�(�4�4ON��jt%^-d$�C�a�>ybe"(�x	s1�� 	�LzV�ڦ&V\�?���OP�2t����Am映;�%�O �	��G+L#t�ɺ�<��A��h��ԎF1;}�I��-ʤL|[W�N�b��G�yк`&>�8�;/��i�T郭f>��QR.�9/�$�N����<�ON|�nV�[��T��b��F��aT�L�Eҁ���\#~hz�dB��d�P]�\��t�u�&���Ñua��/U��[@�7cj!9���&�����g�� /���q�KH�"�"�g�V�|�RU��b֏b8��AƂ&��H��5Z(`�0��ӌ��I��Y���'���R��O<�ҙ�@-Bw�0��O6�����o8����>K�x��`'\��u������ �@��mD�y���qb-��y�LĮ9�Lб���&��y2�C!MOH�GNݸr��M��'Ȧ/�*8�$$U�z���s�M\�s�\�J|w���o8�4�4���@����5*�^�Pmz�N�M4���YI���çD�U�:�C���H��������\q!"�=1�<�q$;F��pHT#�>�S�-� D���B���u���o�����*w^��W��V&)E�g�"`��Y��$ߋg�@	�t��(q�I��ц���%0TEa��ռ @�,1cn�8EZy�Q�Ք�?"���0�a�K~�'`B�K�DN5)��9��L�V���A*O� �2GD1nTM��fU�D���K)@�1��~:s�7I@�@/A-�u:�����y��	*Y^X����MBXՅ㉖�"\XUI�pN�����~uiAhC�P��iD/&��L7�	�SL����٭(/
Yp����R�<)f�!rD㑮��>�'q�`�1�z�'�:�2��A=`��T�Xjl��S�*3�!��:H}�M�q&�,g=<���#�D0`���Y�fv�Z�����C���%���1qo½L,@�D+<V^|D"�D���%)���?��tA�:T��-��G.� ��S��<�d�Ch\�,,h�BQ���=�K��ָQ��5�BBG��"�
M�R$�Նv��X��!T��}��d����'^�59�љTʕJåӄ`3Ze��~"�`I28�l��`��������0P�,�s`˥ �Q:1I�>��;%���")ǁg�BX����z}B���pO�Mr��ލE�T�h�Z��DǤ\�$���īE�r���M|��(V�{�YK���-�����	?$�A�7-{p\�u)H�\l���c%{t��r1�^��,G~BNA�L�`�;�� 3'�I���J��$V�BO("�%9)T���(J�v�{T�ã5&�E���O� ��D�ܗr�jl����,�b���)��a��v��(�s�
�t]�%��N+.i��I�H�h���BK"Z���Bf��1��TЖm�r.��CSW���Ҥ�iEF?����ˡ	^]C�.O48�t�5��L�',�r���5��@�|2"EM L�JH���KBlA0eo'U�����ARK�+|�t���XP$§y����jt?��ƻZ;�T �>�ySIJIyhЁA2�<�=�Ӡx�1C�1���>z J��Z+l��Qr̔(f�4��B��)T��" &˟#�X�Z*}�'�.!�gA �X�SA���t@�<��}�E]5G���D�p
E�%_��戶Y�
�[�%<hqp�d|��mV�H-L���q��#_� ��+\rj*`c3'�q;&���	�^���h7��40x֭P��B!Y�$���wc:xK��$�̻D�uP`㑈6i4���I��]�b���fP���X+_�R�r)M��V8[�Ś����Em�1.��h��o��?��AH�*[�B4��	̗z�D�I}��	ͨk� �&���l���рSi��s0-֟u�	�	N	ff��S�#ݠp>��AR@Pt��@V&?7=�-Jg#��')Q�����K��Q!� $8�^ع����xS@� +����b�ހKv���SN���^ *����CX 9������ǚ*P,��Vj=����&R���Bɜ�"��� Ӈ)'g�i2E�=-��2B���2x�jR&[&P���i�  ���˟W	W�([�U��X�
�@bÙ��y
� jx�D.		V��(���<S"ȡ�7��ǟ�p5��-�*�;��
x�S�>H����TH~r�نYF�]q&.D�V���Y�O�,�Px�LC,=��II��:$Q�D�D�� ,�!�CI�Ty)�)s ~���b�^ݺ���# Q&��W�A�-��C�)*4�`;�й.�%1�H8ngB��0G�}iwĝt��8�O�+K�C�ɓYJ�9�UFɨa���c���*y C��%g�΍ �YVo�,�5��[C�+&�p�B(Y�l�bҒ!��B�	��|8��CI>CH�R�M	��B�ɱGed��a�
ҭ��%�B�ɾwQ ��S��6:$�y@(�i��B�	��X��J�;��� ��ٚ�|B��38h.2�F s[�=�m��%@:B�I?Ӕ-
��ە'�졃�
a�B��49�$�;e@��-u����N�1,�:B䉡f��<�Ξ2C�Xjw�.c�B�	�v��h�ȏ�����W#�v �C䉅���d�#?�����k��Q�B�� ߘ���*-��� ���2�B�!�%����z޾��! �I<�C�	�/�h]ҕk�0w�ҁCrAC>m/rB�I�����Q��	[A&A���*D�8r��_�|���J�D[)�&<�/D��`��$��[�d�6�6�{D�&D���t真+�V%�'�W8 ����8D�����(D����>Ŵ����+D�(m��RhJá]�ؙQ.)D���\�A�Ġrd����)D�L�����ġ�D�$?�x�1�(3D� �t�UW�Fb�-Io��^C�I�+q�e+��B�0i�5H��ۅm��C�I�k0��3��׬K�z($�2m�!�$YF;��V��;y���;Č��)�!�d�P�tm�1�Q7}q��x�m(T�!�%�E��-ߐk��DJ�*8^�!��޺R֒H�!�D�V���U�!�$�a��!�բG�z�� g0�!��'?�F�"��ű��|2��D==�!�~�=0�aE�zWVq�bJ�i�!�$�f��A ��Nڨ�ŉ}�!�$� B�)���)F7�|"�ȤX!�DJ*"�nd!��2}�v����K!�$��j��G�ۙj �x@� x�!��*[� ���0T���-ҵ2�!�$��Nu��'�5G�q�a��+f�!�B�T.H��PX�g���Vc�@�!���w��2�iA`P"�]�!�ܨcc������|�f�j��@��!�$Z�j-�V·xPpqy���"s;��ȓ*�����W�a3q�Q]�R��ȓB�q�
��JG/�� �����d
E� '�έ
c���a�ȓ��Q��;D\��ُb�h���DR�\C3�A�ZP�e�ad�4�� ��7��	Pqm]�,���8�IV�@���G�Rx�f�;^abx�!��Ivl�ȓ.�qxgCV�D�lp� � m���ȓa��Yi�D��>i����D�E���ȓ䈬I�f��+}���si���Ԅ�	4YHT�.�J��� �O��Q-���>y�;Lnp"O�����څh�:Pir(R�?'�eA^�@k��B���)�MS�s�t|��i�%s�N]B��W;7)�CAԺx�!��~�<ʣ��Aڷ�Эn��7��Ex�Sc�J�� ��-�?9ڃ�8�)� �H��=j���#2��m�̬1��'��xc6��8$D(��a&���b+��pL��3$ϑ�u��-�/)�,�d*lO������݂ ̓*v\!���� ������Lx�u��]��"���u���<shl��ą�-�Vu�b ��yAB���.G�'ƞ!�Ӱ[(��QGϏE�`*���*%��A�9{���|��w�Z�Js�ޖQx���1aA��Eɍ�$�]�^�B��)������ (2�,e`�(�f�K�� a�4���O U
@��R�O���@rf���'�`�ڧ���J��!������I)|�d�ԩ=}b�����A,1��U��(۠��&/n����:b�A*K�p�h	"��#(�ġCד��s�*�<qkhi��ʈ#J��n6tMR�w�M,O��U	!�I=U(P#w�T�|���T�K���`�6tE\�`�I�>t;���b�	��L�",�HA��=�i%�� �8Y铪P�0)�@`��P�,@9���;��QC�8ehE/×%�6M��b�}c��ٝ�<�4��/$[S *�I����i���`�����?D�����N$z��sh#d��$)��.�L���β4�>�������`��y�qO��&��'@$S��_4�x���#J�d�X�32�3����W�O;1��M��;M<��R�,��.�3��["#�\�-;{'6l���Z:V�
��O��p=1���8wh�qԀU'2d���Eɽs� �3�ALQb#f��Q��+����pi�Q� �$2j���q��<r���[�[���J񋜘r��#�&�d�azZq�|����9��]�!�X�:��C�������
��1��Pg�N0@���H���%���Z ��p��;N�O̧u�7�:O�`�⣁\-!����S�*�'�������c�ꙣT�F�?���h�#>�䆡/s��i"ɏ����h�!1KBf�bg]�"���^�"8��{���|�xh
5Ƃ/���$�Bc.���-F�Un8���'Nt̟$�@�C�Rg��b��~�b@I@�V�,�a���#
C<��6G-�� ��2=r1�דK��=HB��/D8`��� �lcTĪ�J��!<��:�m���F���I��=0���-A0`�V聍kiD؂�*g��V�-���ea���u ^nx�(ӳGV�E<p���c�,c��� �Z�n�Ή�CK��h���!s�%g�Q�ƈ]*=�"=���]6��qj&�&m�̅�s+�i���93*Z$�5��Y�>�)w^ �� ���G�<i�'�!"-э}u�D����<�H��'�t��Ӧ��Y�>M���S�5��1#�n�8wh隒"R(�8�Hs��1&�2�;7a�- 6Y�B�Ҏ0��k�{bf�; ��\�D�hϔ���n2�k�H/Hj���\�����  :U��E[1`�V=�%$�L��Rw��yxy�nY�~$,݈��B/v@Hxq0ǖ��W�'����be�a��R��I�L|?!�Bw$��$@a�����n�0�2h'�R)J��@�	^�
��c�끒+W~�c�h^�m'D��D:O�T��C9@��Es`�"�������D�J�C@��� ��I�c�B�D͕�:�@�(�20A�nUD�B=��@���4+���g�Z�a�mM&�&y�U֘Zj��JwC�
��I,0�ؐ�5���ʍ���R%���2K>�t ҋ�ά�t�	�5ܜC�7K7���AM)N/��"�L�3DNP�$��
�ڀ¤Ȩ0ƨ+S�>�$�ʕ?�8fMK�#t�l�&
\4Io�t�sHS cҾlg*�$ӡcФPy��l��]��拗]���А�W�!)���E'^\�5�Ɍ��]� ��A��pD��U�'�`-�Q��jX�qT=b꼑q��Π��a�7M��@��(��M�)0���'�60�����͂����(4�䬉=�t����
:�t�r����ᷢ�8��yy7�ҏR&&�qG��6�*�3�n['eu2#(�v6|l� �a�M
0��'0���aw�G6� �sn�`yC��r>lx���8()Q��{6)�7!?YbL��.@2�/O�HZL"��� )�t��O�����\�C�p��t�A�Z�04���M#@���f1��b����QsnO� �z�@��ׁh&��1�
]}BnP�`�AO�!U���s��3>��J^���O�Y����]�l0G��x�FL��j�66���3īخ���b��Ȇ9�V�;v��&�6��S�����ع�� \7��GyZc����uFY� s�T[��%_�Ԛ�}?�b�4���f�6F��2��=L�	VoSȦ����H�]e��h�G� x$�ApA(.2p��	}�g�8C�J �B �S%HT��/�P�C��K��i�Ŕe(гa��#<Urp��&�THYf��='�E�O�����y2B����F"����ş-����3��%��x�'~���n�1$��KB���?d��1Q
(%��,[�$�>t������T��#����Vψ	p��1A��*B�6`
�9i���p׼ 0U�݅IK��c�-���#�4'>�PA(��
ɒ]�B>�� X1"C��q� �/Ɉ]���r�E�;�óaߐ��e=,	@��@���s6��["&�)�\+��U.v�I��!j��Ғ�A7&�L���@�w<��J��JQ���5�r` U�T,=�ʘ"7ˀ�h�v{ m�Q�N����M�w���+0�,Exŭ�.�u�J�/����A`�U`孕�:���b녺6k��6OĈ	����L�/�R�s����Q�g�gXr�H��M�C��0a�S�z�����v��7hS4r~�P��	N�gbj-��*F�~�(i�'HM��a��W��`����4px�|��I�bop�g��3`q�H��n��B�ta���	�au�T�$n��F��Q7�	�}tl0&��%H�x	D!vf�Ȩ��0�vi�W��Iô �B�Y��ѩ��W�}y,)��LK�*]eJ���bM��g҃Lʤ<��]����pjք48�0C%[3@qB4���.,�g��31�P�E��%A*��Ab�}2��#']0�O7$�c-,Až��#A������1?���R���<}8"aH��*td)��M\�GȨʓ8���5��5w�Љ�#�^i��Ol� ͨ!a\*$B�qi҈�Cl�8��LQ�Աj"� �H,!&h�ݐ�\�!O�{���62�8sΚ�~�"�ڣC��1�,%(C�H���$O�k����D M'�Ι��Ɵ'
�����̼u�����x`FF8`2؁C!;SwN�Q`�"kz��fÞ?��#EGŘPF�8n(Թ���ߵ�f���j�����)*|Ĉ�"a~����&��;��P�N�S^,�[�-�l��U�c��N]�CF��\�S'[�H �0��
�O%��0%ˁ�������p�d∌V� (�gKZ�K��a
L!��(eA{���oN
��&�Y <����@�*oN��Ġ-l��1��H�=n��"�K��궯x�<$Y5gA/sW����	Av�? �!�$��Fk���A��&���kq��J�v�Q�F��P�TIRl8��5�T+_~�Ę3s"Ra3��/PL��ѫ�H�Q�)�0�^�R$�'T�B@���Z�B�?�"�T�N+�����n�:"'ǐ{p1ǣKl	�)�{�x��� �r>��'��RO�)�hT���,b�"�ȠO��'�8h�gD�r<�p�U���L�ּ���{J�h�H�^�$��M��=a@u�wDQs;�\��h K����#F��M;sk�-v��	�d�=y�<:sJ���z�O��$DV��� 1�T�b�˃�s��!�$Ľy�6z�
�5�2��u��Ef|eN�8GB0x���[�j�8�&�#W촔S4�/:�Q�ň�IyBnQ�u�S�L��W�L=��zgȆ�jF�܈@��%n�h��$È-s�hD�6�
4Q���ֺI6��
�(ǗoL����#q�4�ןW"�Э
I	2�&L	/S����(Z��:�hR����شi	�rF}X,�;6,�
�
~�2!�B@�)o�Y���Z
TͳiR�.���0��4t뎗 V��uj�O�.y>b�	�f�*a����ا'�r����*)@�0 ���}��UZ��S �jV+�3�V|2���k>|k����d�R�3
�eWB��V�B����Y,h
I<�)� �d��f�ծrZ������ly�c��T��I�R�/]��YgI�9�Qq�'(/v��U]�qWj��4�La!�W�a�xK�n�3&9�X��V�j�[���R��d�p�:���iF
T�,�ʖ�"~Fd�3W���M�v�x�,�*o����$��r�4��T)�P�*���n���k&z�萑���E���	�	�)��}�I�*�$M�s��l/|�dƇ�N2l��c@F�?���Fba���  ɇ�Wv��O&��� ��Z���';�~ey��]�zO6��C#$=Nz�D~�K�N���bIa.�Y�k�p��|��	�5f���R�78RI�*��Y��uK���(*���A��W�x�O^n-ӳ�'}"��f�6�͇��1�U(6�	�)k0�h�O�V�Ap��g Đ�J|j� V3��1XpƯ��@P�'�#�(7ʛ����u�����T!�V$7�xBa��f��}��kb�֝�A��1"XSޚ�$T0�݋�,[�'f��q���E�'�*̓�Z�6��Ug�������2�O��2��>34fy����$��� hY�b��W%e�r�x�6��-q�T˧@K&���L�)��h�H�6"����b�]#���@3����Ђp�hU��0�w�δb�V������T
8P%�8�R�RW�Ůk�^q�A�W�~���.�H��I 99RX���صo�,���d@(L[xʓbԶa�T*���$]���O��(*f��Ѭsu��ө.`����Ri��wrG�2���B����.�p��剸/6�`f��
��$b��k���[1�B�a�N�x�+N� �vك��,�'r$V`��D�;~���Sc����hԧf��hS
��mH"��h����x��OѾ0C�ej��Äb�\-�.�m��KC�_�w}<X̧��@�.O��� 1�"��W�\윅 �.],"������'Wt�k&��;w�����B	L6�AX#�U�e�&@K���Ayx�rVj 7\�Iv�4u�|$�O,�����O��l]4b�l�P��
<$�6`���|��ʼ&�&D�@�n��ac&W���'>����O#g�:<��\7���u�0b�(��Oe�t�E�QQx�� �	�`h��jM%;^�@C��e�d�ШG��t��M�D�n���\��%5F�`�(��ǘvL)TN_����2�K'g�@���',�%�'h�)C[&]	 �Mz@�B\3�ҬZD����� &��'�M�GW8�	�9(q��?J�DT:�H	!�Dl�&�%A���	K'8d��$�&T`|"��LF$�`oI3	���PR�е�%�N�!-
L���Q�P ���Q"�� R�A���g}�@�Z�P�hҨ-v%���`B���'$�ԁ�bV���T ���Zb�\��q�B�JÏZ�]�8��V-�K�6)Ta�y3p똅t֦qxf�'#��B�LβpVlxFFX�s���q@��/a��['�ah�% I�������X�v���1��گg��ДB	����Yv
 �RS���׉L���D�)~NI�˓,-x��.�	jt ���ya���¢�<�¸��ǅu����&�*"`%�s.M�	|THG,P*|j����!(+�Qӌ�:w�t��)P����"YU8��Y��Ԫ`�N���,��b^�9T��!��( 6 � �,��f�_�C�� B ( fx�)�Қl%�at���{��X ����D>3�&y�7��0C���J��̶ @2U p�#�I�M��)!r���++0߆���y2�nj�rrDȫ��A bE r�����-E*!K��
�I� \��#�xk��'�t2waHD}b�\N�N�� �ܑC��);�l� �ȹ��i��
J�=y��1�b�H|*B��;am��r@��2����
�C��4�-�4,e������#�oM�B�2m���Z0;��D~ң��"�Zx.'g� �#Ut�����',>�"G�M�8XY�K�0!�f��*wn�4�Cu�ܣqѓ,�Tl�e,_��R�TI���`�דI��B�&y�EY��ozB����]+V�F9�wP� b͡g�+�ʑ"��t��� �:��c��?�jt�)�ʹ�%�W.g�l�0@ڋ�.�k����^�|�j���ӘO��9t�R� �|���
,0tz�IZr?�#��=�x a�Rٺc&H�l����ލ9BT��'���q�շNT�86DھSK"��*O\<Aţ��鸧�A�H�y��p�5%0x �Q.�	R��wL���ظtʆ�R=�e)z�|�RPk�O�f4����J4*��|�rJ�;q�4��V��Q��O�YR�aի/ڰ�CS���[�ҵ�Ďz�6�b�[sϺ5�sg_�A���I�d(WÜ`3E�Z8r�m��	���H/{@Jtz�a̺J�h`		PD�YH���Bހ���$��xUۅWK^P:��:�j"9�nuy2ͳ��@
b�)�N� �"O<ICO30�Ы�Ԗ �`|I  S�6���8�c��k�BmyB�Ǖ �dlO07���v�$�tT�'( �Y�� 6�����f\X�Y|FYC��..��k�k�D ņШP��A�5*?z�b݉&��Qo �2�)6[�|�Wk6�S�? PH�A�(b&�p�B�Q11������<4��"�S�B�d%"c`D5�郃	.6�8��
�e�hm@Ѐ?-�*ؠN�1	�hQ�%��uȲ� !�8��L�ѧD�Z�|��� ��xp�}K���I�B?Jh1`�?���D\����D��r���LP�{C!�dÖ,v0@����3�n�2V��72h�I^\�	9#��c�,E8PS>y��L�����'�>@���1�5Ja��?vH)��'"sw)F,?��0S`d�"(Ƞs�8���<Q�5b���2t��@�&��"!X��Z�eRW1!�Ă�XIŀ0g�-"Hl� ��F�!�V�K,�hk��@2��r�?�!��H7�z	�bH��,ب��D]�x�!�AG�8pcC@I�#�2�UIj�!�8'`�0�g���b)��H�o@?5�!�č�CN	�%�u�$;F�G8 !�D�<Bi䌣�nV��|�v'D�Q!!��*b�9D
�,��)s4��vs!��� _nH'����Q�%��%A!��&^��t:���6�
a��n�8?!�PҘ�2&�A*ξ�B/7;L!�$ʎc&�����Y!��r�#!�$ �Z��aa��({j�-ZTj��]�!򤓄`��e��nIzF�H^�!�d]%�.tJ�KI&VFZH�aصp�!�Ė;D���	^�d}����!�$�w{Еta[�^�~,���"�!�D��������ivn���Z�^2!�Ă$C��k'��AR2�{�ϑ�%�!�_$3FF��UlH�xة��A�D����&	�3��1���ø2�(T�sq�h3s�\��Q�ҭ�;�#.D�t�6LH.b�C��7s,ᰕ
g��:7r.帅&*�'aC Q�'(ۨfQ��YD$$~�T�U#R{����	EE�E�KA\4?��v���nS�v�/x4����v���N^�S�t�����ףǗW�0lի�/ad�])�&�p<xxq�4���
��0|���^)D1�d�K�����Ca�7�<���͏`��𩄔{1�Ȧ��E�v��&��p9JL�'��U�V����Ӡ8(!q�$y�t����E���0�%<��!�M�,�g�/k���Ł%}�veC�J
Frm���_1Opm���*�[�[J��9�TQ�cl���f���+��9/Ԩ��aUŦ�ZF��ly�f͌�0|rP
��vY����/# j�$��Ħ����<Y�O��y��)M�#���Ad�Vnd�B1g��'of�Fy���O. |@�!	& ������$E�(OQ>ɀ4,�|���3Ë�]$9�1��O x���S�e!���,�
!Jj�ò��)AY0�P��$#��!��
�c.��b[xl
�ccНr�'m�o:�'rm.��-��,+��
�1�U�7-C�O
�E%,�)�vm�9P��=o��F	Ɲ6� ʓ<���9����ء����EA��0b��O�b�b�߈]P�'�������5F���fƛd|�)�ԄO'_�h�@�xB��O����+A�=j���>Ր-c�dʑ$ĉ'	��d��#H���I
�RڤAg&F05��ⅣI�w��I��?�%�U�����6h���McM|��`I�������Y1D=�hvE=�0��x��=#�OR��ᓚLɞ<i /J�����Xܬ���OB�pAʅ��R��O8X�a�Ƞ+ ���H� N:0a�'�иZ�"��k�v�S"��|B�P�'܈	�
"Ko�����/xf� �'�fL�O��Oz�����q/Ұ�
�'m�Y���" �DsW�K7b۠р	�'<贺ae�cd� G�:$�D�P	�'��Q��MM�85�`����|��'� �y��J>N��c�NT1����'G`ɫ�=t��q��]�L�c�'4���g��f�n)�䍞���B�'4(Cv"�`~�p,�(�p
�'��[���'�ֱ����	�x���� �t�$F��j\���ao�H�t�C"O>��
]���Y.U ��K�"O6��!�
8���1�P*o;ԅ#�"O�i����r|`U���SK6��P"OP�xG�9��0Q�؝>p�y4"O:I�!$�n6L��A�,A$��%"O�E�8	� ��9��Q�/Q��y�01���D1/:`��)܌�y2��`�L]�j��"b<����T��y"�Ơ>2`��e��M^6}�7oԞ�y"$�WҊ��D�@8�ۗ��yB��.&P��'j�:65"��v@1�y"�A�ڒ��)U	���J掛 �yB�4g���X�����}su��)�y�N�W������Ļt��S�<�� B���x�IΊYl5�o�C�<���@lL�R����UDP�i�n^@�<��$ ˮ�I�� 5�lصEe�<	�6�XI��Ѐ�Zy ���E�<��B%8�$�3g<&\�ykՄ�K�<��P�o�ƘC��������R�<�ڒ,fly�cɪ!ip�#a��t�<�E�)pY�7j# w�{�ECw�<y�_�5_�p�V	�{�����(�p�<�G�
�+��9@��MB/b�sN�p�<�/䬀Rӡ�:7����i�i�<�1��! �)��۫
�H�!FEd�<)q(�'�`��զf⍉�&�_�<yQ�H���1�p$�<��=1�CX�<��0$"�cDS�*x�3�#�W�<1�H�/���[�%_�8Y�9���]�<y7�@k0a���0y���`�<1�@�Z�p]+I=�"@�p��g�<A�ł.���'	Bb4�p�(^�<���;o�:aR���Gl�ȓ L�Y�<Y��Ni�ݫw�^�\�*eC�OX�<i��B  5Ԡr*�;~�н1���Z�<��,ʠH:���.��d�͑V��<�S���M���+BH�=��I��Mz�<���Z"`�h�
��0����y�<qC�T6{��%����s���ې��n�<��aH�A���`�hD�m
�S��Pl�<����y>��pUl9td����\~�<�e����]���2:iF�'�x�<�B�J<��1:$�'Quj�n�<ٗ"_�a��d�>H���@�In�<�2k�rҨ��g�X=�ʩc"�j�<ad�(^�X����9d )6�K�<9�,�F`!X�����@���P�<�1aƀ^j���U�Y_� �w�<�*�%-pr�j��X�Tn�+)DL�<1�K�J ��JY�P�
&�AR�<��oE�32D(#�&U�;�l�A�fv�<U�	��)َ֤cMT-���Vt�<Y$C;f-���D��k��˒r�<I���`:�Ͱ���v�6i8M�l�<A����2I�8��^�f>�
�&j�<���E2K�ne���.��NBd�<y�(P�Б���~�=˳��y�<�0��%^�^dk2f݂]&Ԋ#�]�<�`�7U�Z-� E�>B#��JӠ�T�<1OD��a�O��Љ�(zc!���N��W�L
*�5� ��z^!�Nd]��
�l�es1µGM�-F!�� �M2���'A:\�� ls�P��"O"$�� G�C�# gӖj��"OJ��e�0!��hB��;l� ���"O�M����c��C�n ��
��"O��r&ސ
Y:�YE9����"O�}�#.4�T�S$�!(7R,[s"OLL�í�5I�DԵ!u�"O �iX�$�F(I�dP"He͋�"O2�������-T�#OB)"�"OL�:��3� R�F�H:��P�"O����E�Ej����͛$~�Z�"O�q�g$ӾYj�b�K����c"O6�S�+�<R�f�铯 �?
5I"O��3�#@���0P��eb�"O������_#�@ƄòA�6�s0"O�P�Q�b�j f.cԾz�"O^`�H
�f�� �@P�@u�A"O,�9��˙5hH� ��#c�FHA"O~ѱ�"��7����,|���s�"O�*v&�k-��#tcY8A�t��"O�@
����JӾT"1Ë8�!�$"O���-\L�hzuj�T1��R�"Oڕ{$��e����d*�4+N��f"O�)zs���,���7j�3V�Qj�"OvL�S�,\�4܋�� j����"O� ťF`�F���S��]�"O�١U,� ���R��?�Ĥp�"O���F
K�v���pvDI�"O���t�I�Y���`�Enu��d"O\1pF��I��|��ފ9s��c�"O�ă��	(��d�e��$A�"O^1�r����1��I�P�\�3�"OД�ѭ��d��D�E�
+k�~$�4"O��	��l����� 8pȩ�"O`)��X-n���� fԒ��qp�"Ob\��bN�?� �Q���mK�I@�"O}�Ԩ�-�:���BR��|�"ON�1)L y�����{B�dZ"O؍	��g����1�J�e>z�k�"Ol��0Or���l�U
rX�7"O ��
F�F�-��ױx� �V"O��`��@S��PW��9A2� "O,x(��.z�b���"W�v��"O���tK�=b� �Ņ@�m���"O����'׽E��)��ۛ ��E�U"O�Kd��!�$ը���>�MAG"O� �DC\[�T�d)T��Ң"O`��s�U�v��Qh�b� ~���"O�w���{U����"֓N�"0��"O"@�&�vh0Xp6뙯A�
1�"O2ibs$܅?B�Xd,��n�N�:�"O��`�K�8a{Z`�Hȇ��Y*K�!�" ���6���]$�X�f�3L!�DM���Qvι>M`!GȰ9!�D�j��s���$7�ǥݼl.!�V�d&mpa�Z��ÓX3a%!��$�x���-��%Y��� @;!�D�^PƉ���z�~� �	1!�DV~�:��"��}� �c�W�*�!�dS"Վ��&� /~\�h]`h!�N�N��T( B��#5��c�!�$A�!�X�ِMs5LԊ��=�!�$������|�Ī�j�#�!���4D��}Pb�ݽXp������!�� �Yr�؄PV臅])hX�
"O�5*7���vu�U>v{v\�#"OH�@ �	#À$�3�	]:UC�"O�m�"�ڪi�LQH�/-_Xi8�"Oz%*ܚOF�����:0�PX��"O<�+�OB3[$-ag�6�e�"OQ����4t̖x�eǉ�I[1"O�:�!üyXH��M]�^pY"�"O6R9���R@�K�,���"Ȏ�ƨ=�2峰�r�N�Q�"O2p�M��h�j�엪^��q0�"O�tZq��6�J��A-I07 �a`u"O��:��M����A��b*Ab"O��aP���W'���v!Ңv~�UQ�"O���� �^��x�D�4y�X�u"OF�bRh].cs���gqT�#�"O����*/h�d�ƌǟ[}��i�"O�Br��)�0,�s&_�K{��A"O� ���޾wE|1{2���&V<�"Ov�s��1���� i���"O�, �i�|�܊��j�R�Xq"OdH�!D�O\�1"r���h���"OBdcR	̕V��PZD�_!T�tA��"O@�C���9ᒰ�� S(f$`"O�h�թ��RZu!�i޻��q"Op�8��_%31
0 �g�DYXD"OdeA�� P1�%kV�G9#и��"O���% +/m*=X⢔ U�by��"O ��S� f(ׁ�`���jQ"O=�5/�l�>�R�o���"O�U۴���p[�<��{ݖI��"OP��s�Z/h�C�O*�r�""O���SMM���A gM.F�(5�s"O��	Q�VD��"d�
٢"Oְ�@��.W��5��^�<r�I�"O�Ę��V �02
\#{2���$"O�4D�H�� �&?����"O�� �"�  ������F�rx�Q�a"O�,C�,�fD�R̔kw��"O@�"�� ��y�q�bpz��"O���v�ڙBcL�@�B �tջ0"O(��ɸ5��98�ȕ�/����""O�Y�T@N�:<��p@
e&u��"O\���/f�tz��Ռv��� �"Oĉ{�C(X������]�R��$S�"O����P�4jrc9x��T{B"O|Js�T�x���;W�D������"OR�c�NȿPgVPq��͘|��"O�a�'ڪc�`pq���"nB�h�@"O:��dE��5a��s�oO�$�� "O���[Ț|i�NW��X��"O���sE�[��x�S.G�h<<��"O�)3׈�x���lŪҼ�"OHY8rN�0���*��/�l��"O�,y��Ș׈h��^�S6:ѓ�"O��c��,+^�I��b{[!Zlr"Oșj��G��\R�"��-��
�"OJ�T 
  ��   J  �  n     c+  V7  pB  /N  �V  c  �m  �s  9z  ��  ͆  �  S�  ��  ٟ  �  a�  ��  �  *�  m�  ��  ��  ��  ��  ��  P�  � � m �( �3 �: 'A jG �I  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P���OH�=�r�2�z�L�"S��1%�_S�<y��B�&�VM���"w��2�L}��i)�d'�d5ʓuƔk��^�|2 uIfm׊N	�)��CQܑ�G�1�&��F��ԤO����J�l��0��,��Ip�ւj.!�$(�`tp��ɚ]��,S���$��.�HOQ>����2�Px�M�7LF�9Ԃ$�O
���Ϯv�=�wI��1�H���e�pXFXcق$c��-�i�'�1OX�}B�)�2HPV	�۴�ڠ)ے^p`�ȓ(֢�"4@�%O���4��?�.�O�c��F�t	�,(�p���!`h�+
��xR�i�*JfH��R�p���$hn�����V}�� 2uD7	���+7�P6�вb�.O �;�� Q *�;�H��eR�+G\P�p@�|��'2�����G�B%�J�mg�4�J>�'a� �ON('>��'7�~�����iY�5����&�^���,�	$�>���D��$up�lD������gF*
r���;n�����ź�yr �+w���gҾP�R���?A�4�~�x��I�~�R-Z��Cs*B�(a�I�`��b�X0���~��t�? �UP�b�+Oè�s���3'�mJ�"ODt��N���ְ@��3v>b����|"�O���<	�y�M�<Bݼ���M	�=��gV��?a >O��!RN�:�d\'+�E���"OQ�we��Q�t�밈�r��X��"Ov0��J�8(��ʔHK�h��䫕"O��k�Z( q�'ԂA��!#"O�+��U�|3��6bP����'Mў"~B0 ^�Uz�p�Z@zI�a,��y2�V�I4ޤ� �E�QD������~�$�^��o��/48$�b�S)6v8 �
1��'�&#=�O�����#�zf`労�E;F�Qy��Ofu���}||ssH>' �2�"O�3!��zAJTiMW����$"O���R���b�zx�N��%��� "O��)�d]�i��-�1'����"O�� (�z����'�Z�"Ob��HK�#�6�����}9�����M��0=�䮞�*o�5�c/è� ܠ��
F�<��'�" �h�H�9�FH��LA̓��=	Eet�+C��%�@J����G{��$^\������h�n��?�y2l�LU� e� ��:�cC�]1G�.�S>�i>�Fz�U��ݻ�T��8�Ӊ��y�B
�i��TQ�D<Qg���C ���$��j���0�#֯��V�X�qW` -P<��ȓ`D�`�h�7n���7�T�)����ȓ'�V���G�06��Yi��\�=��0���a�!���$���џ�Z8�ȓX�Z$�`�)RM�7"M)����'��$Ē��'R�Ol-��g���yz��$Ղ(Pp"OxLi`I�-��{��X�ң"OzPs�aʝ5e9�?B��E��"O��[b��xnUȒ��P�m�&"O���/�&����B�����G"OH(k4�N�ic���Qɟ�N���!"O�Yv&P	P���
�I܄XEl��w"O� �����0���@�W<��y�"O\x�3hȄ�f9�gG�`6��1"O���w��y�d�g�A# ���"O̹��)�IX���q��$�:�"O6���������V�;b��]�C"O�m*ז ��0��Н#M��1�"O����
%������(=��{�"O�Y���8-�;���2�A�"O��*V��&��c�b�� K��y��'	\c���flٗ&Ƭ]h���4]�JU("D���\&Ad,����Q#w��`�#<��
�HO�O�Lu��(�.y�\�9�N��6�:m����b��E�d��r�Hb���r;x�K��W��(O2��$�5%q>pkW��ty�4�Ԙk���hO�܀a7&ϛ#f�U���|�8�D"Ouyt�ٗL�\A���e>,IS�Mn��ħ��'n��(�� ������Ԃ7x���'P9�(�-M�Pl�C&�T�5��'���R�A�_u�Is�3v,A�'���↯'w�&l���2�l��'G�� c���>��W9p>$�@�'�����f~ ����iMv���'�ԕ�&����	�e�?f,R�2�'���S�H��e�n�AoBKY�+�'mJ��f�G��!���ޅF�4`
�'�$1�דN�6L�ɟ�B�>���';�i��L��x�Ѫ�9?$8��� X,i�A1Â�d K;e�"O��ǂD#n�&���$�3vc.�0$"O�c��ԊtTp ��"��L\��3"O��h�Ţ0�<C���4Y��#"O>-�d�Ñj*��6a�7SL�!��"O�����b���3@��~^r�i&"OP-�"�8A������*jQ���"O*��Q	V-ή�Y���$5X�ە"O�8 -E &>�0c�"#���"OJi{SDQ� �Q�La�,9��|��'3�3"�$>���@� )i�>u��'eX�z��s�,�R�`5W�Tb�"Oz9���<:�S�O�B;j0JB"O~�(���^��ᄌ&(r���"O�x�s"�@�jͣCaM/]��p�a���)J�����n2b�T���Q�p�!��W�h	��DyKB���K*^�qOz���� Ԉ���)2_F�$HE�ݤ ֡��~�6]�����P�+�#��X5�fS}�'��>�I�(���CO�	�I�c�TR��C�	y,Ͳf��(N��B�O�[��C�I�<�ԙ+�E�~x���ϛ�uL��Ox⟤F��+!R�J+�j`>8Y���L;�y"�5Z���3��T\��}��CD���'�����I>I��Cd�V�'�<����WHn���J�x� %�e_�n9����X:�ۇ�Hkh<��-ծ~y�8C�� ���6$P�x�ǣ5�yq��7���=��Ɖ"#ljH��A�pP�Ao� ox(8f"��c�:�O��(�)�S3&4c#�Ѱ$��%h @��F�JC�Ɍhh�X6hֽd���A��(oBC䉚M豀q!ȉ"P�ѡ��1?�jB䉞
,�Tq$�WQn�1#���L� B�`�<1���!|Jd���`�j6�C�ɘit�%�RL����-@"�[)}��C�	N͊�B�@ˏ
H$9�����x��C�ɯ4��d��OW�tmB����GX�C�	�HAv���]�=�Pe"v+H��C��q"P(�vE��u��A��¬p3�C�	2C|t�a�(0�i�!Ɩ0��B��;e�LИ)X2*�8D�<K��B䉃+M�P�"�D�sA%Y6��=�"O���̆�C�5K���.�8�q�"O����
�%�M��LI�e�t8�"O��"G3�x�3����|���F"OԔcRʓ�C#��+5!�hyJTqP"OhR��,� X����
ab Qp"Oʄ/y�NY�Qn!X��R�
��y�H�q�tQ��o��Q�C���y�D��X<I��C�$Rl��Kˣ�y�b�M�����̃v�z#N��y�cʱ_�,�cʆl����3�ȥ�y��گdg6�{��1|w�`R@!�2�y��6�	PF��%z"d�1�yr-H({�~�rw)Q�onn�j��yR�9W�h%��0o����ʋ��y���[��m��m=n��C򋘶�y뎫m�����c�.f��`�ƚ#�yr��|�ʼ	q���+34	��꘦�y�ߊz�"���Щ�H��%��y��V�^랕�@IT P�	Xp����y��J,:��TV�/2�\�'�
*�yB`
^cn�ㆭN. B�"W��yrBܶJ2�k��5J�������y
� �ݫU A�2\މbr�׫��aJb"O,�ڴ�T6�^�QW�>����"OZX��d����B�C�
w�F=��"O�̳Q��oU�r��δh�� s�"ODu
��2K�XE�&��s���'���'}b�'Z��'���'eB�'�f=�d)�*K�T!���S�>Asw�'���'$"�'a��'���'���'�@�x��wĶ�#E�O6v���'���'`��'���'���'
��'�F�� l���IqH�]Ң����'x��'���'1��'���'���'Q�1P�
�(u�P����7P���9��'�r�'��'y�'���'�b�'��L�QKN$Z�Lh���V�euD0���'���'�b�'L�'�B�'�'� ��$����1��iE+x�0�P��'��'H��'���'"�'�b�'~�-8'�	(������	
f�h��R�'�b�'���'L��'��'���'��4� ��$b@��É��1ó�'�R�'���'B�'|R�'���'��vD	c N1�Oм;r�mX��'�r�'GB�'d��'���'�B�'IX�	8s� �$n� Wb����'�R�'�B�'�2�'�B�'b�'�j���H�+<1�i�k�A ��"�'���'�B�'Ub�''��'K��'��xC��M�}&�G�H�C�᪔�'v��'���'�2�'���hӰ��Oh���.��X�"�X��3�~MSsǋNy��'��)�3?9��i72�w��]t���!&��b�^��u 1���զ]�?��<9��i7�i���[pA�ì%n�4��u�~�8�d�8p-J6�&?���:��	P��8��d�'^ш"�NY*0*@�SaʹӘ'+BQ�@G�ģ��~�~Ē1�M�"=>��҂ȫQ ,7�ݏe01Oz�?�����Ȭ�͸��S5v���X�Fаxϛ�`�D��b}����I#ᛆ2O�q[ӽr"��a5l2&r�!d:Od�+���S�Z�a7��|��n��̡��Տz�J`��\`p�ϓ��d*�$�����E3�I=c���`L�C���F �sA���?Q'Z��	ݴ��v6O@�7)d�B&�z@<8sV�Y�Ul� �'ހ�
��� GFԸX��$�X{@�n�۟����ٖQ�J����/O��er�XKyR^�`�)��<qA�������rc��sfg]�<��i�<���O�Pm�E��|2e���R��J��Pٖ�Ԁ�x牍�M�T�iA�b-nJ�F���ٖ՞�������%'%���A�ټl�l�0w	ފ������"�zq��I�y����Qn=Dd�H�-�A�ܘq�ۀѮa��ST���:�c�1B|�xh2&׭o����N��yH��B!��,wZ��k\`�L��Ff�'n$
�(�$ҧ{��Ea�M� "��3��� Djæ.n�"��I<D�`q�C�<x\	"gY%(��t#����B�*B�ǘ:F����ιqZ�����P�`�Va��M���Pl�dBE҅i��3qȼ���ǣE2�@!�[�L���FO��� �:�AB�u� u2�}��31��uYJ��$9j��*�H͕Ј6M�O����O��	�Q~��N�K���q��D>qظ�����M���?��F��?����?y��ZK?�����9.ј�	6��s���#p�̌�3���5��������?ubN<ͧI2�I�a�2 �$Y�XZ�q��i�faRV�$�	����3�I�tȐb�)iS����dN���r��;�M#���?	�x;"`8�x�O�R�'����醕FiY3/B�&��M�O�>9���?�@b ]��?����?�tC�+Yp�
1�_�f�z ;�a�:rɛf�'��U">�4�����OLʓY�T;��@7�H[D��p�<�X��i�2�ɘ'�R�'�^�L`�'Y�hkF�1��X�f�91GG4N�u�N<i��?�����O"��%*�q��?#�����&�7l�����$�OR���O�˓;���{�:�Ё�W��Z��ˢ	��o�>�X�Z�H�	Ɵt��Jy2�'�ݖ����k�d���%'���I�K;[��I՟�����ܖ'��l�dJ3񉚀c�p�9C��Bh�Rh�-U�49nZޟ��IMy��'xr�����Oz�H�p�=I0�\@��1�8Q�¤u�����OzʓI�Yx�4�''�\cL⹪���	>%j�B�Z����ܴ���O��H��>��s�h	����?��s`�H80��u�i��I4�"h��4D���ß���,���օ/0�:�`)h�:�����"��&�'��/K��)��g��/w&`1+gˑ!�ɑ6��?7�75-�<4n�Ο��	��0��=���|j +ܼ\�`��fQ'`��$�qP+"��m�(_�	͟���?c���I%pw�p�r���,(ڰ�ЩtΟ/�M���?Y� ��ĳ��x�O@R�O��J�ױ0�ȼ!@�&��ȣX���']��p�y��'k��'(�Y
�H8�`��Dk&=Ɣq�bnӆ�5Y���'��Sȟx�	Oy�H t�<]`�^�}(j8��d�4@&�6M�O��"��O����O�ʓ�>$���"%��I�Í�n����c&��_�'���'��T�`�IΟH
�A5zsH�7��5˰Ԉ4d��$�"b�l��� �'���D5V��I�

�Ԛ��'4�U�4h#J0���'7��'��O\�䊺s��<�C�is\ݘ�� ��4($�������O��d�O��?�FO��	�Oh̩�N�u�6��A�ן�)PG��OV�d1���8�+�@�:O&z7��f+t�I���a^��¶i��]��	�l���O`B�'��o�`�a`��G�	�qG�/#`�b���I=�D��s�?�~� ��j�D�k���j!MH,c�DL�$V�X���3�|�����������}yZw"ְRb�^�V(py�r�ȉp麌{�O���R�C�y� ����T���4��L�tP�m
�ӛ�*8z��'�B�'���]��ȟ"EJ�4��!Z�H� �l��B���M�'Ꮱ;��4�<E��'X�Ta2B�aŞC1��;���9Vz�~���O"��ǧy����|���?!�'� ��J?1-k��'к��1�?�ɎLMiQN|R���?!�'�ʉ�dB3J�J�Q��������4�?Ib��*���OF��O��<�BiӔ+�2�#B�3i�L��w�>y��o�b��'�r�'����I��!*<tH*���-au��!�M�נX�'���'Qb��O���rL�5ÐI"�n�*F@J�J��J�9��Ǔ�(��ǟ��'z�(��yT��E� ��0��|�����W7���'���'��O2�d�*o� �&�i�64�ю�2Bƈ��b)+L|][�O����O��?9ʲ����O�ظvܷ$.Ixt��M��!�bDǦ��a��?�$еy��D%�`	��)
^a�&��O�~�6-�O\��?)�Ǚ���i�O��$����[�!T>�&U���f�`P �X{쓘?��F/�I�<�O���8��
	l8��
�P_E�'W"`!s�'c��'N�$V��'�,�h�
`���L<<��?!�[0��<�~#e �jC��!�,ٽU���������0�������ӟ�	�?)���d�'-Pe1� S���EK#�>a�v�a�jӄ`ñB��1O>a�I�Lt���ƶO2ĥX��A@���I�4�?���?I%8��4�P��O��	�_W�Dk����fK���0D߃j��m�ybfD�]kh���D�O��ɭ�:5��� Ϩ�z֎.�6m�O&5��Ļ<��?���'�f��B�B�y�<5�h��91ڱ��OT��FN�?��៰��Wy��'MѲ@E����lZR%˱3���4F��E�	ן����T�?�'}ڸP��C 7�pT��+^/G�dMsڴhUƅ�'���'��	��d���t
m�e�Z9���uH5���EȦ��I���	m����$�7//��N��+�m�_"�j�)F!��$�O(��<�������.���^�V,`��U�T$�Z�*@/�L 4�oZԟ��?�*O�Iѷ�x��ЪmL�mL=�r���e�;@��f�'N��� ��c�j�4�'���O����T E�J��щ���E�0*.�I�Ҥ��>k��c��'(��mӳ&J P'�Q�+��M|P��'P��XJ��'�2�'M��U��]�BX��D႗ve�\1A�Y<��꓊?���Ɵe3�<�~J�lU�tl����h��B~ @H&��¦��gLџ��Il�	�?Q�����'�j�3���R=A���'}敺��b�f�$b�X�1O>�	�^���#j�_3�*D	��~y�4�?9��?!�
���4����O��	�Y`����m�#i�@����PJ�`�y���������O4�	�aS�E�UbټE��y� �V�P�f7��O�L)C��<���?A��'&�=["��A
���G�
R�8��O�}{�сM��	����	ly��'��!au��PdȜ'�@�v�,1avj��Q6����@����?9�K)����11l�k�!Dru��[oӔ ����'���'y�	�� B�Şb�D��p%#�!�Hb�i�B���]�����	{���?I@"ɛF)��nڅ��a��.\HAЅ���j들?����D�O���4��|r��	bq( L��xt��gðuD��÷id����O��XU� r<�'h�����M�s�m��BTq�=	۴�?�-O���	5Lx�'�?Q��jaMǫbB��a��������� +�O��Ē �t���T?y�%P�dr�m��t��pA�>���n��x���?���?��'����Zc��_{fLS `ƕ<P��җP����s,z�+�)��8�t��tJS:ik.�hsj��f�@6w�����O\���O���<�'�?饫+I�$��O�n�p*vG	���l���y����O�m��! *WcY-�(��,����I���	�`6�������'y��O��q0+��}�f0�	L0(�k�BCa�#���s����'��O�Iؑ)Զq�c&7)��a �i3r�Z;d��Iʟ�����4�=��e�R尡{���'dmj���w}� ��x��O����O���?9%A[�b���Z�OK�|��ba��X՘��.O����O���8�I��(�Bo
h|�ͱ0�m��9#�"+f�]{1�%?A��?�,O��d�42��� 	~(�� I0cqʤr̎A�p6�O��O��D�����8��wӄ��a�~nDdIPoҒ2Mb�KgQ�L��ϟ��'�m-+���p�@�F�F�65P�jܷ;��iW���M�����'�"k��U eAL<)��/\ƚ��ɋ�}��b����!��`y2�'Ǻ�PS>]�	��,��_�P��eKL;�l��?^���}��'��i��)Ҙ��霒h�z�a�"ܛʀ�;�
�*�I����c��˟h�	����	�?���u��O� �b�(�[)D[?����O6t�".��='1O�i��]�h
�ZV ��.��G%�zx�oړ7]���П �	��,��oy�O���ב ��ꂀ�#^�N���� �6͒�!��3�4���X��Wr�? �x)��8kXhµ��gh�� �iq��'�"��=�i>����|��;����!��\;p�{RHY!i��A����mf*4&>Q��՟�`�Xp���-B��	�ҫ|؊nZʟ�kլ	Wy��'-2�'LqO@ ��-J� g�QvIKcZ�
�V�x�r�4���?����O�5�G�ی��B¥Wc��c��6;���?)���?���'���K�,�*j�܄����F�đQ��H a4�PY�O(���O�ʓ�?�C^����0~�R4���Ư�:%��^6�M[��?�����'����z&���ܴ:�T�Ave�xF��U��dzbq�'�2�'���ʟ\Qs��H���'/�i��ѧt[�)��)��q����Ԩ}�2�d)�	Ɵ �6"_{�8O�aSd�R�A��=��n �t��2��i��]����)C�-�O��'����D�f� �*��0��r�]/;�b��	;!�<a&m#�~B2mB)�x�1 �\
P�#�I�I � ��Mk���?������'�?aW�U�N��)�aF^�VƉ�RK[_#�I̟@��͔Uy�Y��3?�;&: �I��ԏpv>\���Ǩ/q*al�>
��ٴ�?���?��������?���]p����8�����W���1�i}0Y���'�Z��J��ƟpI ��l����Jܩ>$����I��M����?y��*T���iT��'���'�Zwŀ��)�"&�|ʲ�ղh�	�ٴ���O.4��<O���$������nD��A� �")��u�7EF�M#��h�2ݛ�ir�'-�'c��'�~�ѵ&��)b��	X�J��y�'��$��'���'���'x�Z>M�!��(,89X5�ڻR�8�ۖb��uBm�ش�?����?���%��yy��'a�9c�À98����@�Ҭqd�F�����O��D�O���O����~���l�5��Բ�C��P�T��Cp�R�4�?��?����?�-Oj��_r��)��b����H s[�"�'�a`tlZ����ğ��I����P�8T`n���	3]`�[�d];S�R���/�Vh[�4�?����?*O�dȃ2��➤c4����J�c�WXVЗ�z�R���Op�$�O��3h�æ�	̟D�	�?�c -�Z�NH9�HY��*� ��(�M������O�)�4�R�O�i��:��G0�P�R��./��k޴�?�%����i���'���O��d�'N�p�![}�eQ&H �P�C%��>���V�.O<��|�uB@)6�.�j"��2�^$S�e��M��!�N�V�'�2�'����O�r�'�≍#�,@�%��:$��0�^�2�"6�M�9�����O���|K~���ij�P�
�4Th$bB�2��]3��iK"�'DbJ�l~�6M�O����O����O�F3�FA�af?L�܈B�Ā�Fg���'0�'hmh���)�O����Oθ�5�G�%� ��AhC�7�t*�٦��	�a���O�˓�?�/O����B�hf��( ծ�ri���z��PX����+u����ş��Iԟ���˟\�I	^�t�@�kM��OD�7l~Ax�O)�MK���?���?�%Q?��'pb,ǝ�(P':D��<k7��?.�0�'v�'�2�'�r�'�r@�)7�7m�"LX�|(A�K}�(�w�X��p0o����	��\�IΟP�'�%���Ù@t���çZ��S�iP �6��O"���OZ���O���
��l��<�	��1�d̄ =c2�z����A�"<�ߴ�?���?)*O����?W ��O��I�h?�,�����>�X\)�(�0�*6m�O\���O�DEYޮYm�ǟ�	�8�Ӌ*�v!����Ts�F܅-|JI�4�?�-O,��Y����O���|n�q�j�s�(T[����|܆6�O�Ĕ�I1j�o�������S�?����Z����C�zĽ�bH�&r$��j�O��$F��6�d�Ot�D�|�L?!`�)ӕsl��a��"t��ir�ʴ��[ͦM��⟤�I�?���ԟ��	ȟ��t�
���щ�K�,7t�	��M[�.ݨ�?�M>ͧ�䧴?�Q�%2���q�J#c<� ��(+�f�'7��'d��h�J`ӎ�$�O����O|���l(B�h��i_�r/�c�@dÿiA�'Ҧ�+�yʟ��D�O��$�"|� ���;�>0X7�^���oƟ0��߹�M��?����?��P?m���*ݩLǾ�Υ�w��D%L��'�DR�'�B�'���'��\�d�T,�R5�(k&�@�HG�5]Pp1M<���?iJ>	��?y%Ө^�bI�a�	9b��c��9��QΓ��$�O��=�	�-먵Χs�,��^6���(Q�ͭv��'�2�'|�'�"�'N5�?!��!p�T1q a5qC*���
?��������4�'��ڦ (��ܴ��Y�GÅ<A��yI�#��-���n���$�\��쟬�F�s�X�O���I�<.?��C�d� �>D[P�iM�'	剠?DHU�L|2��j�)�m�U)D!.�-�P�ڙ��'7B�'�����T?�;���1Q�e�U���_����`p���.������iP�'�?��'U{��&� �:��R+T*�%;��!	�D6��Ot��+_��7��Ɂ;y T����.DX��R�<{��G%m��7m�O��D�O.�)�~�	ޟ�d��39�`8FfY?ܶ�q���M�4
׀�?�O>E�t�'3��{�CYH��<Jg`��J<�E��{����O
�b��t'��I����l��U
�:6a<y��D�r�|mZ\�i��>O����	̟�)�.�/HxX��de�5�b�qbGZ0�M��%|�񢅖x��'+B�|Zc�3�6��aӢ���I�O�-Yq<O��?)��?I(O�q� e�41� l؄�ѭcڈs�ă��'���'7�'���'U�xj�+M�j ō=s�"�h�%�>5��T����ٟ���Sy2�].A�t�<H�:��lݞ3� ��Z4����?������?���fT�ِ�VF�26��'%�X�f�9�ڠЄY�0�	�\��fyb傰t��9C�m�"CK�Ta�O�-@fn��$$���I�����+x�|�OL�9d��ԛ��0o���fAF	�M#���?.O~��u�Mu�S����%k��40���a�J��c-[:��K<y���?iUG��?�O>�O� 1�E}P3 ��<H3|���4��d[�Z�VLn�:��I�ON�id~"&������H�u���*g���M[��?���H��?AN>�~�F̑�!hLi�g/�;\}nЫ5�զ�S팟�M���?����2��x��'���bĥwm��Q�l�n�r!�6�j�@\�P��O��O>������Ai���	�d�NT(OM�Q�4�?���?�k� D�'XB�'���sC���q�<g�C����jq�v�|�m�-<���
���O���lj�[Ԋ�l�fx�FF~�6-�Or(�vL��ڟ`�	Z�i�%��U�w[�HiEa l������>�a�أ���?����?i+O�p�wbR�BP�;�#]OD����5(�X&����[�'n�C��1�c�����yԍ�(��.�?!��?����?Y����	ܻj_��d�3�l�E�Зx"�i��.m����	��&��I�����h	:\�v6�݃"��0:�U�O~�ň2����	Ɵ��	ҟ�'��s�/��H�j$&�Jb�ߍit-�A炀l�ܟ���n�;^��~�3���P �2����d��-�Iޟ����X��������	Ky��O���XP�}c�4ss���N�I2�1���O���Цse�ŸW�T?���&>0�D���B�h"b�#�i��˓"	~y�'�i��꧙?��'���9v��]�ņ�4_'��.�\c�6��O��dU(��b?�+�[�V���!K��!n���&i�Z;%��ئ��	ȟ��I�?� K<Q�H�Zh�ǂYo�:�����m��!���itԸъ��S�0cA)ș%-~�؄/[>F<�PshZ��M����?���>v"p��x��'��O�����W]=�}�"f��<���g��r1O(�$�O��R�[�������
E��F_�oܟ0Q������?i������)~$v��W��bH �a
�o}Ҭ
�'�R�'ARP�C�?�h9	�a	"
�.��2�^	&I�K<A��?L>I���?y�ß~��,9 m������\0h��0�<���?	����,9�pt�'!V�8�6ƀ����0)Q�B���'b�'��'r�'��0��O���í�\��	e�V�r!W����ҟ\��KyRA.T���bĂp���g�ͫ!����겯���q�	ӟ��I��!�}�.���������j3\�����M���?�,O>�c@�K�ݟ����.���m�6]�e´C�\P��)M<���?�RHV�����l&΀���,b�
�a+� W���]��B4���M�UY?A�	�?)��O�a b�N�Q��)�
C�.�d��F�iE��'*�1����C'}*z��+K�-�*ܨ�	D%ݛf�ƪF�|7��Oh�$�O���Oo��ҟ�R!J�Es�avNƥCQ$�Ċ�	�M�\������ƢR� %�;i����D��,�h�l�������PP�����?���~�M���	39b�,���ә��'Ӳ4s�y��'�r�'A4I��ɍ$��@'�-���R�n�:�S6i%�|�I��p&���g׾�S&l�"bQ�,���$yz�N���<���?a���?���-�����u��p�BZ�x����,�,d���O��$�O��"��O���ڤ@��`h��YCH$�7��:;�h��E��O �D�O����O@���O�w�$���-R*v�8�!ř���������D�����	FMĈ� }���a��~R̅k�
�jvI�$^��	⟤��fy�MwET�x�o/TT!`��P4�4��KF����D�?!��G�^�����x4��F��^��lm؟��	��$�� ���O���?Y�Ǝ�lϢ��+�+eA4D��K����?�.Oj����iݵ�Ĉ	I�p�h����F>
�C� fӞʓK9@	�g�i;`��?Y�'�	<���j��|{(Xa�*�r9\6��OB�䟅#��b?�L��:l1gI߹H�4�ťc�x��f��Ǧ��	�|�	�?5�H<���@r|j��*�4㍯v�(��Q���� ���)��˟(�S��3"v�`H¤��\LBfcS��M����?���g�@Qʧ�x��'���O%(&�CUW��Y���:�L������'F�1O����O�����UT��@ʌ�w|^tZ�F�#�Hm���h�gNϟ,�	���i�OZ�OV�i1D}"R	Yr���[=ra�M≶2�H��?���?,O��k7�*�SU�ыy��I��/��|�'���'���'��OV|ku�ӽNt�q��Y&�9&��ʦQ&�$��ӟd���<�	�jU:��'(�(���I���P.FA���mdyB�'!�'MR[�<"��oӚ�B��(8>�aA�c�i]v٪`P�$�2�Ť"��z��X><�#� ����+��2��Ż�΅@���"O�q���,�� ��`c�RHQ��O�@&�H'�<�&���M���ϩ��`	$�m�l�Y�E-|Dt�O -b�XFɗj��i��BD�JҴ3��_@x�H�葻!_�����@>9U�`�č^�6	{3GO�fKj%�k���((�/W�Y&�|;�"U'U����o�����<.P��B(ܵhh^@���G�@�R�'��M�3~	���6�PM�sa�)u�ܽr��	��L�տy���L�Nl!x���w����C2S�����6Ҹ`'o%W[N�˲��6+5�( Ɓ�O�u���k����s+ӹ��2�	�4��T��j�7�2��	Ο�����'����C'S;3�܀��F�-�
]��'ar�'~>i*�K��n�%���O�&�щ��[�'����'�R���i�%��}�ϗ�z,�%���'�r������'���'WR�wݵ�	矸!É��
�h��!Xݨ�G� �a�	T:��� ��}@:�{w���󤗔i��2�M3b$��A�+6���5��P� ;f���B��aџ.� *��'\��'�]�j�b!(��M�0��'P����v�cӮ⟈᨟tTƩP�|�Q��&r$��Y�"O�Qy �C	cܘ� �O�)cD��F�j�����'��I�8��l�޴c����G�4B8���ȉ�M������?	���?���
�?������-�'k��!@u�M0�$�5���E�*t�0��\��h �M�oD� '�/5ʖ�Dy���h�,�pC�	!i�Dh4���p��=s��đMT1�v�A�q�Mq�
�+d��葃X�Yp�'c������?	��Ө\&�t+�J��ƍX&�\��hO�?y�OH�Y ���R��x�lJz�XF{�o�Z�����8ʄ}谋ʀ�y�@a�v�d�<�@�,���'��Y>A�p�H
h���	��@�;�,DA��?A����ݟ��I�M�<A"F�Z��� sM>	���h%�� .Jx)��=����4�L��H#�"����H� �M���*7�fa`�f����Lx�+��xD*��l���!��ˎ�!"�|2���?����?����J>~�����R��urv%L���$.�)��<����=T\����Ƭe�q�uGCZ~R�i>�pH<i�
C
b�ԔG�32���f���<�P�S�uu���'��Y>]�ql�����I�8�V��5�zV�m� ψ���p۠a�f�Zy�vᖭ=���b!ٟ�b>�NS�:���3Q*�=%JX�N�L�4šN�25�p��%1c:HZ�,]����a���4���"�Z4 DRa׈=b�DS�;?~��æA�)O����O������Y4�%�V!*n��4ON�D&�O`͛"��o�̓'*�/�d�!��!�HO�)�On!�BGK4~��۷o���p0X��O6�D�:-�8]��O�D�O4��P���'�JIB�g�T$zel�=1��Ù'zP�b�\(~��2���EG��&��bb�<IHi�c�Nԁ�G�:i*�I
P!�0������$%��T;��̼a���q�P�j�.�d
5MN�d�O�o�?��?�,OV��ǢJ<j��|�%A1��d���4�S��y�P�]�H����E����M�3�27m�릭&�0�O��U�2X	�4�La��`�<}+���R��!}
����?���?��l ��?�������,i��0��3h��0[���X��9���I?"�4D�Eh��ڐ��-݋@`DLFy�b���Ā&n�AH��A0{�(�u �-c��b'G�0�dк�gϊ`n�eGy��[��?!��Jb�i*e́[~���k�,j������?�-O���/�)��K�&7RE�&������Q�<1bٕ"�������S�����W�<Q��i�BR�Бr�����O��')����bg��B@$X���p�t}r�E��?���?��ʚ�{6ZI�agȱ1,�6Mq�5��O��V�zp���#����V�$`��3B��/E����D#��L�ߴ�M;�	E�$5rD	���/
�:� ՗e��P���K�'�ڼ �N�VaӔ�ĸ|R���#OG\͐���Q|0,)@!^��?э��9O����X�3r։)��tO��+��'�O��k#m#y��4;H�V[T��?O:�3Js}R�'��S��y����p��Pv�:%o+g*�r� D<}ƪY ǇK0a��e[�@� ���
�bs�Hs֩Pk���1�W�Y�Aph�H���:I��v�[$P�0'�F���ЃB�^'D���Uu���@�����w5t�
AYJR.��6���	VcǪr�'���'1?��ظ��u@֜GJ9*��.�d�OD��$K�B4&ux'�P:W��\�pˑ�1O��$NN�����'��yD
�x�2	����V�\�ss�'�M����8e�'�B�'��x������\����/�詁w� 3$�չEa�!K�}{��ޞL���r1��`z��Әe���G�D� b��e�s����j#�'|$��U��g~ȸ�d�ς=R�՟(t �d��51�
�>��h�&>�l3v��C�2U!�O��?��˶�?q��?�gy��'��	3�b�*g�¶J�r`�ŋ�%�BC���t!�	�43�	S-?�` *���HO����O��-~�ݨR�i�Y�(
X�b�%$jԩE�' ��'N���<\���'/�T��8\R��#9�X��ۧ;�������0h�u�dŃ�/9n�PH��?�:�y��$7 �g�	�|*'��%2@��R�o�8��=#n��b�����E��Q�)S�F���O�Y��Ȧ�j�t�? 4�e���0,9�Nݔ;��:��V@�	����Ie�S�d���s��T�@���c�ȱ%��0<1��d�6Kq� čX�y�����ݔAU�Ă����^y�cF��7�O��$�|b�B�@m�1!B�=-D�C��l�X\a���?��\\RаeO�V>$��ABJ:JDPrF�	V����$ɕ�C��W�߱�r� Gb�C�'i��X�S�j��T.��)�rp��ݛt��р2
?Jj�g���
�v���(��T2Ғ|��?Qòi�7��O��'t���p��ד��8KSM�/;d�%#�������T���Y�.�f�T,(b+�(r������T�>�DP��X�;�@04�J�WjW�.�O�e`xo�0�	g����;U�"�'��2��qv��qt���"!�I��g���p�k��c��"qET(M�(@� 
P�1�7GË0`��R���gj"����os�0����*?��	2D� A��!�Ł�D��Q.3S����}�
�������Q��}XP��'�-���MCZ�����ɢ<��䀪:�}!č_�,�Z=S�%s�<9`�J;΂14F�	�����+k̓�?	3鉧�M3��IM6�if�	zͬp����9D�����?Q#뒏sw ,����?i��?ٕ������OH�J��bDQ�!�!��h �DI�HB Iv W�R��Þ+%���)3�P�y2�,".�C� :"p�SE�9-.�`A%�+^ ����6}켬��OD�,�b�U̓8��	q�n>};��P�B"7x�1�t8���������^����G,):�ȇ]�\ 0Dx�!�$�F��(Bm��w�	!I�\Fz-l��D-���YJF�T�'�B�s��X���!�"O#�
�,�bT�&� .f�nQ�D"O�܁��T5m1����[rd��G"OT�ґ��/ht�e+#�ܒw>����"OT<�*����5rf�� 0�p1"O��z"��|t%;�NƝ)ą��"O(���b��B\�E�ک,m��"Oj@B��+S�|0J���Jxr�"O0�f�M�a���V����"��1"O(:p"��z��aPƊB��pYR"OZd��c/Ɩ�*CJ<tȊq�"O��qe�,BF�Z���\�Q�u"Oz��#�#��hE`RS�-��"OtM�so��:����lĻU��1"O�M�uA͡
��1���Gz~��g"O��9��ь_떔��f_�da�<�s"O����ܞjL2)I�d�!C����"O�A2�o3�Ԋ(G>b���"Od�磀= �~e;��"1ޱ��"O��5�֐x�	��,H*�s�"O8Y �K�ypn)���y� �"O ј�N��$ź'��I�6i�2"OXm�Ġ�}W(A�f����I"OVYP�A_�z��؁/G�b�
�ˠ"OXD�ز%9�Ɂ�\�o�͹6"O���OI�Q�x�C��LR���J:D��hT�GV��a�2G���i��7D��j1iѨ0r����d��)�+!�4	��
EƝ&�0ɉ�G͈E�!��-T,���B�̎]9&�A�!�$�.�t���K?K�hXJ2g��z�!򄓛.(P;6 �R��P�2u"X��'�H`K�Ɇ	% ��D�0~?Ft �'cʡR �.N��A䨉�{�����'�� �(�24����M! �<��'&���Gg�u2H�4��~�\�Dz�9SZ�١�ɐ�@�$d��A_�$H&@ʚ�d�T�W�J�+7j���y�NL��Yr�O��P���|l��8�бe�PH�i,%j����s�)�K5�&�!���`���<\O�4À/����"���'�Y��%�	2����D��b�8 ��'AL�#�ĕ���	ُSV������7y��
��P:��*�F*1O�(�<�z�y��ϊ 9�A����2xh�pm<m�t��7�A]NP:%��&HW���$A7Mi���@��#Cތ<��LX�PuuѐNK?I�80���3lO�$P	���ġ�V�$Y���KG�R�@~,�rB�\7%�� �'�%;T,��ςg��rW�+lO� 8 
�Q�|�f�E���ѐ?O�pZա̅+if�4�O���"ʧ@���dbG�p�Q�&I�K�
�R�	�HѠÛ�(�l�oIR�|[UeQ!��!1`dN J�����j
���'{p�7N�|�I`���Kā�Y$`��	D�4[<(�$!��`��R�F���'`��֌W�?P�7͒�
�r���y2*��8��@�  ;zHr�)[�0���P�'��D��Y��[�ϖ"$�p�x��ēr�@�9s"ռL�Z���ϋh*�h��w�B� ��~��F}����E��52�8)#���sm,M3ӫU/�lAZ'��rr(x;����p=ɵ �]�<�BE�e��(KR* j�'���8U-͡+\���	�p�D"���h�Z7{P��� �O�azR��M�l\�%鬼:�a�(�P��;��Rt����~BI�� P��t�������~�oá>�Pv��^�8E�&%�	5��i�iݖs��l[��dͶ3d�M6�B�-��W&��,1O$���/ �T\h�g�H����@C)	��`�B�<A$�B"M%$щ��$��jMh�h!e�_�N0�(K�[��H�R��R�f@���� S
Q����0�|�8@�G�"\ ��@�c�����CT|E)�-1�O�v��ܴs`��"���w�	�!W�\��L9#	6�h�k�9���dǔC=�$2Q���r�&H)&��M�azR�_� ��5�P萄%��=�E�?�4UBdn6Ul������~��3k�b��?�l�����%$H��g�0,o�1����ʀ+����'�ʁ)`��e� �v�	�O�^Qk�'�8Pf�l^1)	O��tE�n�ҡ1M�$B5��n]��Ag��f�!a&�?u�Ot��SfBv���P�ÀND�x�H�-|�6�#��J�8�@<Ot��WnR>6c��T�O=xX�M#!��s�VJ�#ZF�lbdRR�=3�f),%�=�a������I;Βe��U�A p�I��Ghz�$X�U�JuZ���0���.'A���i��dV�T�B
�2�B��7�_�H���H
�<JD-q&Π?�"���5i�tp �Y�&�Z%�􉉇L;�y�G0�$i6O�X�4�m�T0��X�?%�������x���Q'9���UU&5<�	��@�*vX���<��H�
6ز� ��ۺ�PdP�� ��\�z���B��A@,�2��A�F��8%u�&@�-"wh�k짨�	-U;@���%1*]��[�DS4*�2�P�ď/�R��͏�u�4D��!3§�M���nx8��E?�r%�P�O����ᗥ7�J�qu$FK��x�`((O �S�a�Hvd0�E�&x���E�6Qy�lW&S�!X�c�']_ ��O.P  4H�2�a�'��p���24���1S��l�S�'�.��g��'rY���<�UddC��fhJ�UF\Q4�Z�EF�B2�Q9.�5���7�4X�d��>�;��݈ME*U`0+�"���@=r�!s���Q�U��hF6~D�O��Ē4ќ7���+֢
*��-�]{ �;GLM��?�6�� �����>EZU�L��C��=_���c��G�z�Asd�T�������x6p�{��G;t�f6�Y��]Lc��%vyp�ǳm��EL�2���K�j�%Cij=i��'̔'T�g���#I(X��r�\��?y�α~d�0��9���OO�h҅��Rl�<r�n��G�*Xi�G��֟!^W�`[f�K���a��5wX����*}��95i\0i��Q���Ӑ3
n6��Uy"�
����c�:��ڴ��tk���^g��@k��5z�@�T�'�(��� =��[É�1�j�
�S�"Ak^}IS�X�yj�tU�
i� ��fEе0-�E�I�E.��;D��xS�%]�#��+O������\ڑ�����P�>4�'�S�k�a�Q�;�x)Hq�S�=�:�~ZGK@�#���ZTJ�PC��+\�|�i3瓡!h,i���E-q�8��a�V�r�.��'�
��˅2&n�� �f,@���7����yb�)V��Bt@?���q�Dކ�VMy�+{���@$ˑ2��,R�˴W;�z��ԁm�����ĬLQ�� S�	!��(�%�+�Es�E��I,w�:<�f��h���ҟ̉�OQ\e�Ë\ ?0�j�$�0E~��Y��
�,\#<�퐋n�nA@QDX$%��÷ƅ�<�����,҈�P�ҭڇ�07�|Th�@� $�X�Bu-��q'�V�� X"@|I�b���I�I�(,�U ���PP �74+�D�0��0��x�'6�yA�j|�,�'$�(��p����čB>h6Ti�T#C�x��f
\(偒iS�aJ40 ��.��x���)d���Q�w`���*xZ�8z�'Yd8�	(�R1�K��t.N?��]�N�9c��V�KS�T
V���1�4\O��2����.I-!��̫4�{`n=��gZ�B�>y�Iߔ�~*�쀻�O��$�!�°^��`�#%�d��Q�e�N�"<)̷!=���"OZ�QH$���N}?�S%O电0q�E
c�|�AA�<9�6팒V���_�qOR)4�#���d"�°S�+�P�"�!P4���E.�L�0����� A�O����, �`�0҃Ò�B�!�ŀ�4��'��G�!��<I�.߭dG�T��D܏BlrS�؍$l����db~�T���M�Bm�'K�� cNܼz��u%K	'h����'��I:E#��%rf��!*V%�axŢ��z_`��P򉮺?a��p��US�d����ՈgmF�3����	�'�2Q��ɘZq��jun��`4�s�L�a�\���#x^��� O�t�+�k�:��5}"�'}�/2 <��U�|2�7퀍�@ў]��Ѡ�K��y��8K����!�;M���X3�wm�x��O� �u-���T��-G.C�|;`�??��/K�\܆��
�o�aҡJZ�E�i��A�bZ��Rk ]*��9P�:��(���p����Dk���T�� ���͇�$X�Z���/VY�?�O�xZć� ,�q @
H�"�T�$m�!�"� 4�R�A3�,��	����ɛ#����K�2p	B���lʜ�� 7O����C �F�hdQ�DO(F8���i�:�����,���CwY�R���ײi�5���1>h�jz>=i$�'��#?���/!��ȱ�������3��p�g���i�@(o����b'Yvb��0��ˤa>���+ɩP�p�J����������$\O�U�Z�� �y;���ABw*E/{uD���=�\������"�?�rR�|%��77`"����;��c�B(�Px�勻v$��A/�(��I�A_B� +�D�=�¸��4v����L/���� 
�6�$�ZJes昊�
K�U7�qZd�~X�����/<+B�W���Sw0���nD26>��Z�a_)ž�y�
�H��$b��K��4ZX�K�{r3n�
0��_
8�ۄM��hO�������L���#��CUj�ɦq���R����ѬŮQ�H��EKN~��I�#r$��	�H��{$�[�sB����Ѐd3�Y]�̚�=yN�طEIv<�M?J2k�J��Ƈ�,��I��e7�e�p� D��r�f�!�BD��&�2n�TR�!w�fqG#\�zkb(�b Y�ґp�n�Wt�>ͻ�ZI�0B�7U	8�XW(З��ē6R��l�"6��J@��2En\���بL &(c�j����'���B1HOr�@�T3��^�z�I�D���H��Ы^�e� baM ���L�-�j�Z$�16��I�H�qYf��/�p��� Z�	;���p�';� b� \�<�`F��ru����aF@	�Q�	F��Y UC:N��矐bB��5��iH(�����s引R�MJ�6r���䋴`��EK�� ��̈u�J#6P �J�-YLp���ܦ]k��<�!��0���V�w�ܭ�r�;������:Fd�3�	�9n�Q{���be�p
�C�����ŲHQ��1+�P=�ի�'j!d[U$S�4�>��%�I�Q>�/T�i��֘YN�y��0h8�6m�c���X��؃u��Q��3V�Ӹ��{�T>ט1B�����.��g�(�k�A[c �}OJP�Ӏ3\O<3�
�8�����b2?Q��
�G�Ьщ� �<�v�����S|?��^�����t���S-R&E�0iBk���!���
��4F�}�xcJ���'d;��A֎�52�tO���0T���T��a���Γ6ܬ�ò� t�0��X�U���J)/�p	Ez�C�E���\�#-�`U��7�y����x	7�/<~��E�D�H!4�<�R�"a"1�'����o������͠K�`�b���!F L�mڿz~�p!�dĸy@ ��s��Oب1s�`}�B�i�44Ф�ۗ�8Ec��V,�=��5O�|;ՁC�0=�qi,=̪�z�i�fz�K�D�]v��ǔx��\�.�O��O�<	�`°P���Je�E�*�P�#<�O��F�O�0ς)'�^�]D�x���#!tJ��(^>uJ���Ŕ| N^���7��`c�'j��I�h؁j�\�sNH�2�eJ����HO��H0�P�-���K�,\ ]r2$b�Q��4���b�ͻ,J�^��sDŁ�:�'=B��&���?�U�@�9��DkH>9�F�	���j�p��}+����J2iG !uZ� ���+��8 q*<��|)�W��b�(��w�� �.�&]�����v�)�	 a"h�aQx��+B!��)�>�iQ���x�V:�"�f���N<Y�JD>��'qd��'8�Y�jY�mx��	D�w�8�ˁ�'��p�p&���u�*=��������E����O(ʓZp��'Q����?���!��=@R���"�	3��1I�Fz�/��#n!�׎K�'̅��ሩd��	���[��,��X3�W+� �$�Qy�kݰ-��Ok>ԣ�-b�x�:Eˢ�ֲLŔ2���j�d6�C�(�T�X������� Q�,;q<�����8�G�
�&��U*�=�Nly��Z�!c�%�؁�'�Z𦏚� ���E�<iB��!/z�{(8\��qt�!}��ʟ�[��R��ruc� �t��8Q;�O�1ku��#�Y!�'k��yX�Γ�b��B��5"��	~������j�'TQL�����A���j��=a�CA�<�/.@����v��u��9�@C�<Q�.8B�N�ЭP�cOJ=Sw�R@�<�Y+q	������r��%�BT�<iF�U������G��U�ԉS�<I�,�7�]���'N$����dH�<���
S�^)+I	K�L`�-B�<a#@-4�rH��GZ�y��'�v�<af&��?6V�`5�T�#ʢ��+�[�<yS"��w�R��@Dͩaz�|�c��T�<Yuǋ88ƶM"Q�HAjz�z�%�O�<�A��M��q�V�C�!��:3��t�<�D��NP��H���O`Z�p��Br�<� �d�Ż�p8�ɝE��9��"O�]9�J��&"��h�a� =��=��"O.�2ũB;Q�xғ�^�r���"O|M�a���CD@�K���=m�j�"ORp����<�H�k`(R�&��0�"O��ڡ�U�Hx���I�� c���"O���A&�+G�[�Ac���2"O�����/PC8�B���={Lh��"O����4K�I����:v:t�C"O"��`�ђ}s�$�, [�eB"Oy Ǎ/ +� �RMсR��L��"O\�B6�Fh���,G�}
əq"O�|B�$L��L$���͡E�&�8P"O�58�gۚm�f�H�L��#�"Oj���h�2� ��=E᠉�'"O��z4%B�h����%J-Xq`�"Oz҆���J�xD�e�"`6���"O�4��#�~lL4�R%��N����"Oȅb��Z6GT|c�B�YrB��y�,��j�@�٦�F��u�t��1�y�˟�(m�`֞4*�t���yr��J�x�!#KҖ1M����h��yrF�J"�\y��^�v�ƈ���^%�y2����A*�칰g�G�yҫ	e��`�V�N� a��YwlH��y� Ś�t�QWU#(y4����׍�y��ִeJ�$a� �7�zh#���>�y2�@��l�� M;5��"i�W�<�`��Y�b(z���f�����k�<� �B��Aa��^�� jFh�<�t��;f���K�G+/���aC�k�<I'W� �D%sFJ�(T��D!�g�<��	�k����f��e?���
�f�<�0G'0���-V���b�i�<��ʚn�������5	�f�M�<�.-�\��NB +gx����A�<17B�%.�h`į�"��	 rR�<�BY#wM.��7̎�sl¡��'N�<����]f^��v�ǟi��A3�]Q�<ɰ��D6��*�Nȡ���SM�R�<�á��i�8Â�R	C@���lGK�<��D�*r���k�#L,>HH�!�R�<a��J�ecp��l���L�	с�L�<�g(�y��1��$R�N�����D�<����(@�K�a�j���Y�<�#E��*p���C9E����O�<��#\<)�]��0�����L�<Q �٥o���S���",����b�<�7N¸eÊLP�'��3��9#G Qe�<Q�c��g�|(�Z����kr��a�<	�h�Pn��Q�	��{�T��D�`�<�!dӣA���ٸUw�U��_�<���^&UA�&
����Q#�	\�<��6zt�LrU��3��c0�U�<Yw!"A,T8 �iE�H� �j�R�<�E�T������!�d�"��[R�<�#oKE�z�Q1�P5=����K�Q�<ҤU���z恅w���/�F�<�3AU2,�*�3�N�l+@=��@�K�<iD��3 �Q�V�� >Z,�S
ZC�<�`���>8�"�V�.IicM�~�<A���h���U&ϊ9?���+�r�<�C�<N}��ip̖�/�N�@q��E�<A�%P]uX��2��$�y�4n�J�<� �e�-��h��: OÛDd(�"O2:�L׈_�����@�j�2��"O�-z񋒖4�μ���2�vd$"O��I �яM�$A4�Y�r����"O�������5zcDԝI�p��G�Ii��ۂ�4;��@2��-���aDh2D�8v�QAVy��@_(r�A�f/�$0�O���C�	׆����d�z,1�"ON݂�R	/Q�A���MX�"O��G̒�r����%����"O:���c�0p�e�a����"O0�X�4b����a��-�z�["O�p��bπ(hvz�@��h���!�d�4R���'���t��HA�g�E��'�a|2�Y�tՆ����_g��k�J��yd�*@x�l�T>dAX$ے�7�y�mH�z�^ ����YX9hB��HO��=�Ou`�'�������$iF�P2h���'#zu!�"h&�P C�W�H���'=0{@5BR��3EG�K'P��'�܄����K
��2r�P�<>`�y�'ѾD��+Dy��I�i�5�>e��'���ZG�'�� ���W�)�h�(�'&>	At��!@:�݁�&����{�'ں4K�<�v�
�0��'~T�����k� 2��5Z�%cK>��S��]���dP�tc�K��f�u�ȓX�^ ��&�[�(c� <ua��ȓ#�*lp!&�5�6۷c�6
-�Ʉ�Y!<a�EA���0`I9t`ȓk��e���'j�`�T鋶X�ԉ��s^�G�'sv,@BV�q%�,�ȓ~�=�F)��_�6��E��������.1�0&�I�:T��˞���A��_�b�#:�HQ��J�>1m��ȓ�m�┩U��$�!O,PLF|b�ӱ���ӆ/���b�o C�ɼ>�C��fwt��G�Y�f�B�ILAnHP�(7�D,2�[�?�B�ɭ,N8*U���~�`8[1S��C�	'[�6�ӄ�"t�(���(OzB�	!e����Ā��jNXd�6@38�IB��8z��W+Q��A�H�����B3�O��0���9�J]��b�5��6"����ȓm��ts���q���r�&�,TJ½�ȓ)��� bи_�|�R$iG+S8��ȓ" �`���Ҩ����r'�Du\��.������L/�<r�&L$��(��w�H)�NF�f9�����a��o�L(<I1�*��-@��ٟU�R܀0Ny�<���Ђu�4���&� ]P� �K�L�<1G��'1j��&TT
x�d�<�s��+s��1�p��S���Pb�<�v�g�H����
i�$��UG�<��F)G�xDd�+ڱ�C��I�<�s��(4�vdp�)	� F�5!�EJ�<���T�$h���o\ �qKBO�<��Q������M���K�<!5N����pO�Q_h@Pi_�<)A�	$|���i��wj4��vNo�<q7���{���S�\�?�J�S�Bk�<���NL���DE�4r,���*�n�<��l�	kz�ZU@�jM���i�`�<�4�9V�2���H.k�y���^�'��?� 
���I���F��ȅ�#�d�a"O��B��r�0Tr�8D�j"Ov�� ٷ|����b\`�"Or��!�'Y�^U��
�n���"O|�g�J!'!]�W,v�ڈw"O�:�A)Q��U�5H��r��"OV����U�p��=X��[=OI�L�"O�4��O�=T��ݐ��8�lj�"O|�W�ڋRL�E޼���"O>y�B5c�Ub���)���j�<� #��O���#��C���p~��)§
T0�C�J�������%kh�ȓ��|�g٘QS�E���r"@Մ�1Р���m�6
D���
6�Ԅ�n+��ۇ�T�h,�P�=4�����qq���wΖ�0/��@$w����-D��ӷ�πE�dA��,%�v,�E.!D��3�#?NH��rdV�I��?D�4��jS$P���P��[,h`(��#D���Y�c�4����dحj�l#D��Y�iB, ��m�C�P j�e�'6D��7�� ���۳,�[� ���>D�˥���ʅҖ��n{���a=D�Ա&b��oJ�qR,�7R@#�'D���e$V��Y�'�;��(0$D����_�)��!�B�ԃ{�. ��' D���Y�buۄ.�ns�ݻ�.?D��C�[/!b���6���B�&1D����Bxs
��b+�'E�pN!D��H4�	�6LpY��L�l��&�>D�D����"
�LرG�UV>��XuL=D�0��[�7�Z�� �S�:,4yq'D�t���F]: @�_
�2UD#D���ן�Xє��!Ce�E��I-D��12aĆl�`��@�#(������)D���&�C?_��˅�I!��:�+D�(ˤԐHy���p��C���1`)D�Ȓ�e˰c2B�&�E�PԌ]I�*D�0�E�ѽ\?��`7�İv�U"��)����p����#���Bq�+G"O��:RN��5��b�͚(�`�;b"O
%�Ƌ�%�t(��;�Z�B5"O�t�ԡ�>T���&�0��"O��R��?� pkW�̡"�T00V�'V�I�V����0-ŏT��|@w&ǈ�C�Io7$ɸ����N�9�dJ)*5�C�0D"���
(3��0d�B?[�C�I<x`����@��k+�Lc�C6���0?铣,@�x�A�o@j�q�K�k�<�	Ze$�H����V�2�Mj�<Q�)�N��ѥ����ʡf�<	�.$H��,��F
�B�
��V^�<�/+ %���!��hl:��Z�<Q�-�qS�%��ą%�fƏ�T�<I&�ղZ�Fd"���.��pe�Ez�<a�K��H�&< �F�.�x1b�@u�<��A��V��uC�9w8�
L[�<��Ŝ�`&�0�r�O82v�a�U _m�<� g_�0�bq*QO
i��5QDAe�<gA�0>�^m2�$�d`ɗɎ_�<I���)j>%��6�� 9 �Z�<�A�<���:w
�N�3��MW�<� ��2
]KQ!���yI ��P�<�A�X�{�V`ㄚt��IaG��L�<� h@!��:,��;2G�4U�`��"O�0aB��3P���s����)�"Ox����1ola%�0p�f��A"O6�;�%8Y�U+��)?xH�W"O0����v"��a" uʨ ""O������/�^Y��01����P"O)� ���v�.��U"M"�DB"O�!8痃y��P�����1)�Q"O*�C��U6	�����'|��XT"O $㳋'JX@�� �C�08�"OF1ò+�_�� "�-P�K&B]!�"O�H���!���i��*[�(09"O�и#ߌ��S������1B"O�1ꇀK:����E��3��!�"O`ŋ�b�fh.�cE�Q:�8�&"O`���-(�`(�+���a"O�YE�Ρ/�VD�SԎ��"ON�`7�pؑ2�o<{�"z"Ot4���eG�X�n�'$��F"O�E��k"Gc&!���L�>xf\qq"OD`K#(�##��P�ÊN.^,�"O�p!eο<��cI\�k�t�"O 0�!����8`9���"OХ�v ��>�P��:"���"O�\�A��P8�Pl���8�"O�h�AѤvb"�%��*	�$`��"O؁B�!Y�2d���#�C0��%+c"OX��E�!sr�a�ߨj�dhr"O4b�K�z�Sw$��ML�B�"O�!�ӧ$�u$�(y?��
�"O��
�
S�!#�{�<��"OZ��N�qvrb'R�8��i�"O��u.�q�A��|2��"O��1E����w.�6*h<E�"O8tȢ	��M�@ԙE�
aba "OV�kn&�84�6�G�rNn��"O|�����}�h�alʿZk����"O�i�)$�H���̈́(Qx��"O<����U�4?�T�Jr����"O�)x����{ф|�U��
_�T��q"O�x��x ᱅��	���"OD��E��e[dk���6��M1�"O���eh�?2pH�����f��(�"O��C�~���ؐL��ލ�G"O^�g��:�0�c�1��tB"O�q��-6V�K��N�/����"O<����$}R���b¾"���d"O֡�0聰K%��B�#vʜA3"O4}ʳO�#J��AR���[m���g"Oΰ;�M��D���Q��ju���"Ot� ��x�h&�˴!i�c""Oʸ��
K'U��uHц<f,@�r"O̩�$+�Eښ�:U�4O,���"ObH��
�n~8�j!Z�Y�%�r"O�9�Ñ�[��k�a�i�<��"OZySa��+zK�D��̤{L!�DN�0i^� &��f��b�-Ԇ�!�d�;(Y� �d ��tH� am�@J!��%e�REsQ�
~G�D���Ӏ_!��G�I!����66dr�Θ2w�!�$��<�`ݣ����-�(��$�!������A�P$M�ވW&!���(�t�;EB\Ը ��� 2!��G�BYİ�c@"1 �!EM)(�!�� ��d(�.M��Y��΂`N�H�"O����m�UN^Q:��& 3�`y�"O:�HW��4*|Rv	P/��j"O�%�P�H+H��e�A��-f��y"O���a\�KT�Ҳ��B�V��"O��%iD�B���#"ɘT��`�D"Ox|J�#ӳ�� D!�*f}�("OХ�4��d7n�b@��hb�͘u"O�}`GeC�Ǩ���������"OR�3-Vj�H����
i�I��"O�p �N��*g��6�ZTj�"O*��%�eF1*���f�x��&"Oi24�C��hAc1��p��"O&��B�Y�j�X��������"O� �e��
SP)��?w�	�"O%CW�A�}�h�A�ʒ>j�pR�"OT	 �Kө�t���*��""O@�jfk��M�H$�T�<�xHi�"O�p�#��6M���F��?6n�1[�"O��IdM�#:����\�H�"O�b.Y.K�2I�AT[F2)"O(�W ]�n�DS��:�Ti�"Oܩ:�ҧ�l�J�jֆ;H�"O��p'ږτUCc�N &0h�(3*O
x�%CK�[]:����� �>�	�'7�e{1.:M�ĬʆL35�	�''��Qq��(4�re�2~́��'�*��b�_�Z�@�tJ��<�S�'t�8AU����sq)�t ����'�f�6�ʵ(�Na 6��9Q@ ��Y�P+����i
�i�ǯE+����R�rX7Σ�����-~l���44m��GB�X|���"k*�@���@��iU+�4�G*Z�N�n�ȓ��Ѹ4#�A���Pv�ZJ'Մȓ}G�W���/�E��s\����~�qSn��1���J-^E�����it�@s�R�[�\���c �T��i����M�L݁�M��Lv��=�����B]�����G�^x���{yP][�� T t�SA$no�<�ȓP
,H+dM!�ŀê[�:�F��ȓ���bAD�|���&�f�P}�ȓ<vh�g@�o�,;�o����ȓ|0����9u6����/G�[���ȓ�,p��P,y��A�FY�2�ȓ!{�-JTK�0@5`w
^�x�ȓV`�AXVN��\���#��]"�ȓa�&<�5�N�HK(u"䭉�}L���#��!z- �Q�
�sfn���o�څ0���-�P(�d��97+b��h�`�KFO� �����(J���mBT#Y-j
T<�ӧ�4y�L�ȓ2<4@`"큪8
����AOo-*���P6�tX�
��Ia\]Z�CQ�>C�`���Pzt�L�����N@�E�Vm�ȓN�&d���У8��XBG�bfʵ��䂰�ѫ�-耰2b��L(�ȓu�8�(f0v�P�NZ��0�ȓj`9p<�"LZw�p��\�ȓ)v� �����'I9u��x�ȓAq0oҼj��1s��Tg�Ԇȓ����<_��¶$�WȲ1��"|�M�Յ�r�b���+Ie��ԅ�S�? �YBS�>/�)���N�e+�EB�"O6EJ�`Z�4����H*�ј�"O� Xc���W�B�ć1&|�`* "O>y���J"K���矑vܙ"�"O���)]A�2QH@-�^ܫb"O�uB�%��ф��+.�d�#�"O"ۅg֨g^ �� ��m��<C"OF����6N�S����ap"O�t��Ԟ�`Z�4}��3�"O����Y\B��8nӢ9 2"Ob����Hq@�����˸�>�C"OШ3���D
��΢���"O�%�J�n��K��N�֝��"O��+�Ǥpƒ�1�C�a�Ԅ:W"O�I:0��
c ������$���ے"O�0k����>�>��sN��#�2Ր�"O�uJT�J��]b�m��5���{�"O�i
C؅8Z����N`��"OPh��^�r`���!��=@f4� "O��d�=EJ>`(B��GҔ�!r"O��8��]XM���gj%m����0"Ox����A�,�d���=�jD��"OL�� �[�E�V �G�&4����"O�d�(��L-j�&�"Ƶ2�"O:р6���`�VE	 E�9�.�qR"O6�)����V�j ��?2��"O��kT�A�=&0�wMX�z ��U"O�50ƨ�����J�LUt
�A�"O>I�v��!�Z0F�D.,3�"O��*b���ŘFO�d�\��"O��Ȇ(T������a1"OV����1Q0e�f�"��qu"O�x�$�B,+\�DE��3b�`"OXTrr*�pU�	��V.{��"O�a����\V�`�Fzf��;�"Or����H% �%�[:I\`c"O
aP%+vu�l	��R19�e��"O~����m����w�{�"O� ���L%,8m##�[�Ի"O.�b m��Gh܌�C'U0I<P�#D"O��h���`����S��t"O����n��8/Hy���!a�j}�V"O@�9��a�D���F�	��P""O��� ��<�|p���ƥx���"Ov�{�
U1\�8�s�Z� w�-�"Ot}�`IPX)@�Ǜ8�%ZQ"OL$�ѭՉ�>%�!��I ����"O��cT�f���o �L>Lă�"O�`�t.�"Qq�m;T�	L*ր��"O�� �.��d�x���/�<��"O�d�ˈ�!�h!��LJ��H9�"O��0GD��]��hQ%��!'��F"OD{CD]� �l{�˂��z�"O��R#��i	�) ��3)( y	1"O��k��6-C�z�>U��S�"O�e�aϱ	F	���R>Y?`t�0"O����ˍI�;�LǉG(��"O>��$*Մ6%r@Д��DD`	�"O��Qa�T/]ބ<1Ν.aΞp�u"O �h���#춝KTmơ�9	F"O�����Ŋ!0�<Ƌ�	}�(3"O�|Sᮏ2(k0X+���5耬#�"O�,Т��_K��	�g@�4z`�"O�%R*˷,y
e
�%�|�P�"O� r	)A��@�)��..�\��F"O�DY�gXjO�zy�ÅȶbD����)c�搵;�N�A��)�@)��&��z��T}�8��*�n�^=�ȓ8N9K� H�r��(�q��_�`�� E9�x=���ZHӒԅ�!�	y�T7~���T`ȉ=TQ��z��1DC�@+4X�vaQwf�Ņ�*��a�� 68�q���O�2��؅�zB�����I":��,���4&��i�ȓ��YHWl�#;�Y���t=Մȓ=ؙ���g�6e��dE-p�"��ȓ
�Α��hY4qB	�1��,q�P��\'�h+��,q+rP7�èF�HL��3����	ڭ$�f�ZtJ�go����"%(��S�J�R��)^1��L��0�򑑣�͖En&X���&�@!�ȓC�v�{�mɎT����D^�)h+"O�q'�F�$n @��+�
r���!�"O��2�m�:Z�Ȩ�u���!���"O���uA��A2��Q�{��4"O�(7��i��$s�,���#d"OT�vJ�5��iB�NZ9zli�"O�Xh%��$��[��^u��P�"O��s�Ȉf��b�N��� �"O�����L�G��)B	T��X��"O*]+tIH��|("��'dt|,[�"O��
�B�([����� KlL��"O�5�k¾8� ���FN  ����"OJ����,=�J�1SE��+��""ON�0��p���{�D��YФR"OH�#s�?g'D�%Ɉ.�Dԡ�"OԱ[�CX�1��ypdS�a�jR�"O��3�0 ̦T�-F3LTF�j�"OZ�ӏ]a��t�Z.:�p�"O �E�A
:$�8b�]/}�(��"O�yrD$T�S����!�?<��"Ot���� &|��D��/�=Z�(��"O� {UR/y�T\�S��} H�q"O��qB��5�p�g�)o�(�"O,� b�BEl�g���"�L,2"O*=�5`2c�<�g�\�U�~)�"O~=ST/�J!C� ��/s:��5"O$i��+%V�����5�`��"O���4�U8M�$����k���e"O��\${�:Y��&����u"O�i��Vb�-�sbWxKd�Kf"O��
�ش>4D�@b�q=�5B�"OVt�E.R�m�8����4.��0X�"O�Q����
.�Qs�FX"ek���F"Oހ��I�Y^�4c��V[\�� �"Ov܋V�R+TF$��L3� ��"O�e#w�ЩQE��۵+U3=�� �"O<���G]kl\��
�+M����"O���F'�kq���t�Ή0�\��A"O)�P��5%��!ш��I=�y�"O�A�7Q�� �!]b�8�9""Ojp@�Ϡ&p������"X��X4"OVu���yn���a��W���"O�XRFE�e��@xp����ekQ"O�m	�cѨV�����U+��u;p"O�B5d�<j�����)� =�@X�D"O���G3D�Z �㇀Yj��$"O����� �����ȍgM
�� "O� �x�Ì^% ��}H�ԽH�!��"O�� ��J�<� x��ɼ?ʈ�!`"ON�`�ȕ$Vw>���-q���"O�e+2nV���"�I06���R�"ON���A��Q2t@B @:N��d2�"O8xr�̷m�&Ph@J���A{�"Oh5Cdl���H{���+�� h'"O64�����0i����
Z|J8!&"O -!��}��R"�́w���v"O����Ʉ$\�� �"
Q\1�"OƥǢ�
tK�(aO-;u��1@"O�ݒ�a���HI
�@V(�@�"O�ex��f�2,�H�v* aK"O>�sI�Gax=�,�D�"�b�"O�\z��Ѫ^�b�`���'K�,�"O���r.��&RVd���Ի�fh��"ODe*�-�) G"��P�(t��"�"O���	X�y\X�R���0U,4��"ON-)�JͿR�"�&�޲�4m��"O���
KPB��H��B���"OLI��2}A����L׹
�N<�`"O X�,�]��Y��lƅʂ��e"Oz��g��mc|i �&/[�}�"OrH���\��Ӏ�'J���t"O�M���V�Bo�Y�ꊢ2�l �&"O�$`Aaܦ4wRٙ�茉E�TAK�"O�飀��?j�������*t�'"OF��I�L9t̠�)
$�"O�1�&!y�� I�h���V"Oy��c�o���{1"
<
�D��"O��K2�>.���!�6_ &�x�"OhA�V��'Ar�h@�/#��mHF"O��beM@�2�
�I�ڡ�b���"O	iA�Ӻ~)>L���J%��a�"Oe���5�d� ��Z����"On��SJϽC�4q)ƾs՜+�"Oh���� p���#�A"t%��r4"O����1DQt�z��
93v�ʐ"O��2�
8"jh����ں*��"O��(YԘ[���$�Ĝ��"O�m�;E�1���"�R"Oxq��5(2@�T�èl[�"O�ѱ4����>���.��5��u�R"O�}	���� >A�do�7�H��"O<X8 �ń}7h`�$���1T"O
 HuM�/9���7�}��M�A"O����)u�x�K��[;����"O�ʢ���|�x)YVH�?�Rp"c"O�$g�ל+��8��e�;W���"Ox$��@��W�2(��N��L�,�yүR+ssh뇁=��� g��y��d�lLA�GF���u[5,ٕ�y��H;3�VqJ��\�a��#��yRG�
޸41���3IL|p����y���	eZ�b���@���Jܭ�y2�ԙe�ΡCPKL(�	�"J�y"d�>>���SE
M*��4����y"i��K��Y��!I�|�F ��ހ�y�(�8��(p`"�{X����^�y��C�c�ʽ��a��ql.�"��$�y)�<�,�ɘ�o�T]30ȕ��yr��0���Y�n��i 0L�
�y��R�r���*�l�/mB�`g/��yFФ>�ؐ�!ʐ t�$H�ƃ��y
� d�����|n*�+V2M�(�r"O��c��t�X��º%"�ٹ�"ONPp��<S ����
�L!2��"O~ْ a�vjX��*˹I��s�"O�}!��^�a�:y��"_�KLX�y"O��zǣ_����g='g���"O�DZ�C�:z>�s��-EPr�� "Op�e�xkr��S�G)�Ҙ�s"O|!+ %��5�l���D jC�"O\Kf�w9��;�A��%����"O�yJ4D� ����SA]�lᐉ�0"O��r���x�S��O9@���4"O�
�l�X&�aՍՔ{�!�"OT4��PE��4bR��|.L�cV"O�D��k�
.�@����1+��1�"OAY�OL4-�P<�U�Y*��"�"O"d�n5 �F'>z-�,�"O��$�ؼwx�mJ����k>P�*�"O2EI��\]6��UF�8?4��C"O�D�+�	�Ґ��Z4�Y��"OA�㢟*���:B�4/ &���"Oj�2�ǳ;{�iS�d�)[�^�w"O9�h�3<�����3QxF)��"O�������4��	�<�"Jt"O5�pKjGȱ�tH^�dкU"O�q�G)L�=q�FDz5!�"O�����0j���s�l��
š���yR'�E�ХPV��&[�F�q'��yb��0yy�I�cX0N�bq�vBΰ�yrM��~�!�׎A�X\�F$K��y�Y
wx�H�`֟p��Z&n�#�y"[d3<M[��T�44�6���y".�8AL&4*#�X2x��[vI�yr�7{�<*Ǆ�u���R��]��y�e�H��画eH��VQ�y�,V�'2.�Aw��S�Y�v��3�y�+ڙ)b����ɶ|�@�	��yrEO5����dD+o�ĈUŜ
�yB�{
iC�`H�b�N\���_%�y���_��\� �`x��	DE©�y�$u��I��?�R�S��C#�y2ID��`)`)G�	Mvp[�F��yrC��?-�<h���{S�i;RF���y�@S���K��Ůu�q����y�O�%'�H�UŔqK�B
L��yrK�� �4!�"�V��iغ�yB(.'�(����'F�1qD��yB�Jzf�0��)�&D� �x#i�'�y��N�B������7�܈���%�y�ʃ ���`գ,2� E"l2�y����W�>49���U� �� ��y��N�v�T���ǛZ���G+��y�JJ�T��� �|
�P�f�y��(\�:�i�v�:]�DJ�y��=zl�h�eĖ e������	��y2��Amp����U�h�`�P��yB.Ҙ\�ҀC��a���^��y⧌�F�u��똍ifR�A�,O �yb��?mB�!��v�R�����y��'�1��Bk�f
�dW��y"�L;f�8X�	O�6�@t@�"�y��"0�4�x�垻d5�)	Pŗ��y�ܷ�H�I��Y�op��1�H��y���-}�5��)\�m��q�QB��y
� x-���;�h]�n�
/���"OΜ���K���۷��\@�"O��@'B���i@�K�IV�"�"O�3��s}�xV���,��ɕ"O�l2D$�j6\��$cG�^���"O4\; �4�ltC����� �"O���IH� ����@�~���8�"O�%̊��*	�
����%+�"O�ġ4.B�2~�X *�9u���#"O@��DiE�	���2q�$��"Os/��k�=�gB�wW��;"O�]�wE���d`ተL��"O�|c#oƕ3$���aOX�3�����"O,x;�ϐ�:��;i�$Jh��Hc"Od��1�	*�XE��	�d$æ"O ��5�Ȫ6�"����Ղ6�"O�,i�r�Pxz`&ٗo^���"OR�Q��8jƖ�SC�S
zG��+�"O^��r�Y:c��,0��S�v��E"O˒.�l��˘��h��`"O��E�%5��ك-ԿK��9�1"Oܑg�U�]���$�ɈT{8���"O�,�w� A"��#p�Z��"OfI"֢�A��xcm^�5a|��c"O���u�ִ&�Lh� �wrQ�'"O��+�EF�R�N<�R�Ғ)�\��"O���g�> �A��3]����"Op��u�\�O52Q�u��nڄ""O��R��җAJ��4K��o��`�"O�0s$�
V�T����u�Es�"O����,�v�Z�@�!<�� �V"Oj��r+D�O$�E��O;��$)w"O}��'BM����ύ"k���$"O��� ���A���8��D�Q�R��"O���G�6GX�!�MN�5t�B�"Ox0�(յ붸��b2[ �"O �K0'ɍJ�p��bѪ:%�5y�"O���&*��=(��"A�&��x�"O�%@c䓵v��ѐ@&&:�u"O� ��[�Q
^�� ���X{�"O������U&��0�I�*I[�H#V"O�����#U&т�g<R1"0�p"O\ ґ��|^��jf���}̺	+�"O��)�������,��@}��"O�M��_�0s���L�V��@"OMXIR�T,(-���ɵ >�KQ"OF�����~�]�u)���dP#W"O89�d\(5��(���?^G�)[A"O}�p������O�`� P"O���Q�V	��V��"t�T	�"O�5zw��#m�Rmj��(|��3�"O:4��B��o�|��G��Q&�3"O�e[%��%&J�\� �	�$��i#�"Od���у2Q2x"��O��&��"O�a��4{s��aL�-QȲ8�"OHq��K�3TCf�ڣ�
{�x���"O�y��^�fv�pQ�J��0�f"OBL①]�(�w']0�jу"O���a��.�6d��ݐH�����"Of�$O3#�BC�
�Pzl-{t"OZ1I�GM$^}j!Чl�4j@�а"O�cd��/�I8�)�T�u��"Ov��.�*'�^ �6��l�5��"Op�����(��E��4^,Z "O� |t���N��J0��cT�t
���"O�y�a� @0p�p�B�0���"O\����
h�ca�)+���{7"Of�p�
�'�D`��K�H�h���"O�}JD �/o�8�vL�?p�1)�"Oppze�۴{�*��`�A�fxf"O�R�$JGh��qb�e��L��"O�m��� -�ʁc�b�v]��$"O���3*E+L[vua���"PL2I��"OV5zP��%��@�����d<>���"O�!� %k7�p��M=<,��kR"OV�9�a�Ix���$��K�q"OhdY��ioH0�(M�!�a@"O
���%ՊD������(��}��"O~�С�М	��I�s�:A��
�'G���v�;��L�"c��z�*�h
�'!$K�|��11˟DԆ-�	�'B���f�Y$k�����<h&���Ug)S&�pM��	�!ú��q�+D� `�&P!f+N�[b�Zy�l顫)D����!3#��� ����?U���G)D�T���Hպ�y6��vdv��k:D��8�kM�9�U1f��������8D�xӥd�<X�Ai��?B�T[�(8D�T���*)
Z�2W�F&0N�lB�;D�l(�#F�Nz��C�Ȓ~��3PA9D���λ"D1xU���$-�0���5D�����_<'�b�� Ę%���q�2D�1�n�'����}猰���+D�9�T�*O�P�o	�2�~,a��*D�(C�3�x�Kg���@� 
-D�$[3�(;�P������x�P!� 5D� �� �EÜ�0S����aB2"3D��(Sg��R\�Ф�e|\}*"1D���7��e���1�XM�v�i��"D��&��#���C��q�d�2UO"D��Z�Kڷb����'���\P�֠>D��+c�\�]�^lIGl,e<��PK=D��أ��Nq,����� �i2`=D��S�i�XT�C6E������'D�$�Qo�aLxs�F�i@ժ%#&D�,�G ��O��Bも4K��@d�(D��k�����T�C��e��H���$D�t���-L1���P��;mb�1�L0D�袅%@�d���gC���X!8U�-D��5Β+C���0�����*D�\�2 ̚�Z���I�eF'T���#	0A���Su�G��29c�"Oz���cgP�*�I�!�ƐzA"O��S]F��P:�%V�&�d��"O�5R��������?�b�z�"OАr#��)}��	��%{���r"O�0�� ��:Ɋp�Ưf�0�"O�����X"-L���\ d"O�<+��#��B��$X6�A'"O`P�A"E�r��lh��U
��C"O��`�M�).��Pq	�;H$���"OrHj�c΄C� �#
"���"O��ʦ��EC'*���R3��[�<��+A<Zz�
 ߬_���q�YQ�<1�#��[�P�˴��$&�� ���K�<��AO�xS2���^�@X17	J�<�4ퟑ�t�B�D5Ճ�b�^�<���?�t(2AF�Mv�5�6�_W�<� ��4�d��m��'M&�"O�W��� �#MМ8��)f"O������9q1"\�1���h���r"O�T��*¼N��RIV�&�V\��"OD�Y�R�~�T�k��^j.1�"O�ᩄ�QwY��I_�����"O�1@�3<T��j)I�v��1"ON�����p3�j2�"�z�"O@�q�,&�9���7f�5�&"O��Au��4��<-!�:Ȣ��K3�y�¿#MB�a�n������y2�Z�R*LЁDh��JF�� ��R:�yB/чnA����Ғ�R1����&�y2��_��X��EU�^`f�����yR��b����U ��b���!���yr⋺id���X�l���\9�y�E�&�R�1��a#�i	���y�d���C$�*���Wf��y�dO���uѲ+Y�u����Á�y�(�3(k2����R<,�M�pB�5�yR�C�b$�I���3|a�x CJ�y��A�R�\蛕���)�Iȇ���y"'��~��8�фX  ���*����y��13ǂA �# �zEz2��y�m\��P��]2I�f�hu��9�y2�	��li�afT;�8ŀ���y��͎[2R`r�\�a���.F+�y�Fִ�*}a��o|V,�e���y��F;C���䘆c% !����?�y� Q�H���(��(l:���yR.lZ� ��"]�MO��&� �y�V(d�AtO*F������y���Y�@S�Ĭ? �K���y�	8m�����6a���xQ����y�Fnw�[W
0�h���y���%G��ು:wv�o�y���;���K͓D�|�෮���yr��5)��Z���1���(�8�yҪ �c���P�$I���l����y���KnL�a��9x��ެ�y��&E���0RlS�{u�a�� ���y�X�:��%��#ml�#�%^�y�	�|��t�e�b����ޘ�y��,��-0���0V�\ s��y�IϨk'�$��.��Ld<�7吳�y�(F�	��U�4�h�舠�y�.Nn���Aټ��B�#�y����> ���(�S#�:�y�(W�\���fIп#�V�{���y� 6lb��I��ޙK&���yrC��`��BCQ��։��*�y2�oA�� �� rb��y����K�R���'G���a����y�#�2����D�AE�=�2�yR�E�-8��&K�� �i/�y��/3��ЀG,_'���A��ybl��'{�IK�{�z����y��X��4c4A^�sb�C/���y�X6�D����c��ɋR%�y&�'��qpr���L2nz����y�`���S%dFn���T@�,�y�hĲz��h�-j �Q��(��y��	�y�('��T)�dj����y����n�)�$
��H�\�灈�y
� `��� JOnݓ��րN���1A"O)Ȗ�t��$�'
Եb� �"O�u�/��|Hq+�!(���"O̵�D�HV������E�w�RL�f"O�Tiad�D8����*?pǀ�yT"O�m�p%�..@RSd���ȅB�"O�Qz1�ܥ"��q�ύ�5���+�"O|�r$�M-C�X���-:�sP"O�{t��R�9{��K #a~u�"O�A���YT�~���Gi[����"O�7ǃ{��#%l�/HJ��&"O��vG*t{q�vj!df�a�"O`�	���tЁ�.x`����"OȈ�d��	g��Rv�E�/P�Y9�"OR)���Վ'ϴ��%��8Hv��"O�(�Â=��UY��<02�Ii�"OʱH�mE(d���K�>;�n�cc"O����o�$����ˇ]�ډ@`"O��9AL7G7�h*���!�1P2"O�H4fB�	�����N��l��S"On�q��#J��鍒<�\�9q"O$\��ˑ�0�Q(��F��}�"O<����uA�p��G�(/���Pv"O�Y�� ӭ��d֐3��р�"O��s�*Zj$��Ę�}�U+4"OTA���_�(���>~G�$sW"O`P�F-��lSHĘ��Z7��"3"Ofa�����h�z��)V(�"Oi�V�T�Q.DT�1��7��Ч"OHx�1�˵tΌ���]��(HH%"O�䃆/G Τ�Rr�د=���"O�lks���d�)O������w"O����Cʢ<Z>(CCQ�
�F��B"O*U+S� �b��}�V�\j�(�p�"O�E��h��
Ep@1��p�:-�Q"O�8��],����'�1;j���U"O�ي3%�.x�0I�		MJ�� Q"O��́�$�`X҉I,u��"O p
�@Ҭ]L���(3�xhb"O�Q� ���D@IxfJ:M���s�"O��10	�N܁�4j��A�E�"O�(	0��4oC��A2Iz?hY�"O|�I�B(�.�sH�!�\ɨ�"O|h�q/Ͻaf |q
�b7��"O��Q��P�p�A�iX,N��T
"O�	a�F�L��B�H�--�0IP`"O���O�9�ִR�&D=X�)x�"Or����*)���
�+P�I�٣v"OP�����l��)Bʄ<?42��C"O�Y[�I��
��X�i@-D:d� �"O���g%�"UX��QhB	/*> �"Oޘ)/Ċ����1A�*>H� �"O�a��0T���g�0��"O�<�w�p6lʑ�Ϳ~�l�R"On�*�X$ `����p�^��"O��� �y@��G�W��b`�"OZ�x���wl���^1J�n�G"O�u�R/(���(�/�%"p5�"O��7�J�-�LY$iG� q
�"O8X"�YjK6�x!��� y��"O>���$	�~���mA�)��"O�0NFmҘ������`��e�e"O��8�Ƙ�_��R%�]u�H��"OΔ��%ʛS���Y����iED���"O� V��c�R� �eN�+0V\E*O��:`�QZ6�� ��[bD�`	�'�0T�-��!y�:!k�!E�lDy�'nQ�4�L!Ba0��K�/7tS
�'��l�Ъ<#�L�w�M04o��	�'V�X����0|�@�,�̥��'o&\p�FM
-�֘�6 �4z	�H �'��a�,�}����H����'�!H�Y%CתYhE%M�q!���'�5� E>��*B.��@*�'�lu�CȘR<`������'��7]�!����R���'�pPړe�mX����[�(m*�Y�'��D���R�g��(�� !RnD��'6�(0��-~�$��"ל2���'�rXh��;@�\`2�5~c0�X
�'�TY�a��:K������y]�0
�'el�����m�b����G�t��9�	�'�`�	v/�Z{�l@VJR/B��`�'G~H�pL��a���A� 1����'�.�@�Z{���ʡ���)�l�H�'�� �\"Ř����Ų�e[h�<������B#D�� ���b�<�����) Z���ʓ=k�Y���i�<iԹT�Ux3�G�:����b�<扭\"� �D�8Pa�c��S�<a������'�7"t�E)J�<�2��>o�MB��6��t+��F�<Q4�G��A��CW+W�N���A�<��GZ�n�����"s�.�x_h�<�$f(c��Ȃ������ F�|�<ɢ)�-#�`Pcf,??��(��̛~�<�"$I�v�<���8q�QGF�q�<�$+'!�tx 	�fW<%�E[G�<��+̨nź����X)F�N�<!�J M'��a�F�|M�iF�J�<��`�s��p�T���U�eZD�<qEU+3aR]��� �~zT����J�<����6x�*y�جk�R �W�E�<���<e�0y)�K$W��ۧg@{�<I�D�D54�ԦI
�ћ��N�<�揕�k�X�ʆ+Ы%D:9���H�<��	� yx)�@+3}R�FUE�<q�#�(9� �ܮn<��'�EB�<�ɞ�mRZ0����d����N�u�<�7�@�r'��c�F+�v��&k�j�<�g�a��R�� � �#j�h�<Y��\�'�U�uO�;B�e%h�<) �H�T�T�j$�b|`0�҆�c�<A4jݔ0SXQ�gE1�*xuȀf�<Yu�Um�H�[r ׄ`2�3�!j�<����
E�Q Ꮑ�s#��[B��c�<!Á�&��l0G-܈Q\�"L^�<�w
���)��JP��3b�Y�<�A��=�&h��*�T�2�EM�<YWe�dh5��/�<B�ᛁ�Pa�<��^+6Y|ڦJG�M�l��S��x�<�Qa�9ƾŪ���+ �q��Us�<��DE0	��A@'H�Iy]�!��q�<I�.[�c��E�:+N�8�rk�m�<�6!^�|	"�E^!?��ӳf
T�<���	�bĄ�"�3lb�ZHG�<�Q�*:��Z��Tx�B�*�E�<�/_5 �8U���WvDRF��{�<� m�,�:\W�D��͈�G�f0�G"O,]RfI��oTR
K�V~ �C"OЖ��6M�r\	c� �]�����"O�0����:�~�Ł�:;�a!�"O����a�D���	��Q�BZyP�"O:ŢD�1+�a
e�ٹrLfQs�"O>6X8[QBD���A:NtB�˖�)D��I��1L����	�j8y��%D�����*�|�����(Q�U��$'D���A$
$?ʉؔ��h�	���7D��@Oq�p�$MR�N��3��2D�|(����qD�3�No����O+D��JǨH<NX���� tdH�R�)D�\c��J($�&��ӆSP'@�� 	$D�L��� `�.i0��
D8��D�=D�0�$*�Ơ�G�,HlmZJ;D��ҕ�&w�|�{n�&�8D��Zt�ϫR�R��+�)X�����y"���=����('�PiŇ	�y�@��d֥	�N_!�@�@��y�+�8q�Py!��K8�4���Ы�y�.�	he$��0�z�8�Qk�
�y�)#��xr$	�q��̃�Γ)�yb.�&M��Swd�)4�
�+9�yr`\/ΗO���	�'R�R����ȓr���zҦϪ(�� a��=-j�ȓ/4�r�+S�c���@Ɇ
ްɇȓ��А@H%l����G��x��8�U�V�
A{�!ڶ`N�-�j�ȓ\rV��f.���y֌֮S����� ����c�XW���"O��S��@33�e��㊁I���h�"O�-�A��8BFř�S��P"O�����5����c�<���@�"OT�x�/��B牰A�̈�#��fO!�D̓R��;��+nq�:Si��N@!�d�k�ZM8���3q����艉p�!�D^�OTp��A�֐_���h؁F�!��..�@R�����Ĉ���y!�d@�@W���VJ�Zמ���r!���L׸	���.z�$�YB��1k!��o5�Ġ�#�:-�x��%�߃F!���7 q�8p�)M�&1�G�F�>:!�$[>`4�4s�V�%k��#Z�/-!�N%C�RM;A���ue�����Ў;&!�F6��{p�֑'��4񏕨B!򤚲[��D %g}�Y'�N�a�!�$�R��	� C�a `c�ȇ�!��V���y�� �9Ib%Zp�,�!��2t)�=T×3 �����߇�!�DM�zt���1~���"'�P�v�!�$k��@B!h�|xp�L R�!�LGI S��3���#��J2�!��V�e%2�#DbP�4�ФQ3�Ԟ	�!�S����FGC/4ؐD�RI�.q�!�;�H�DE�,/ϘՒTg�1�!�Đ�ARt%hV	��6�d4	#���!�$ &�t����!M8��\q�!��ӂ�@G�ڠt&bI �h���!�$�Y8]��C�{@1ړ��mn!�dD%:��}�4�۝G��Kq&
7D>!�U�,�H�E~�<`��e�R(!�$I"[Ŵ@���s�f���y!�]9C���a�Pz�V
3��K!�� �X�kQ�/N�[s��-YN\��"O�
� Ov�����(@�"O����	�=���ġE�/�Ԣ'"O���T@֓3IL�{�`�{�*�"Ox�Q!yd⥂�"n8��"O���W�		��Xk� Y6�`�"O@ �U�=��R7`*@��rb"O��ض�V<:��`NT{5(�"O����
�{�鑖���x��b"O^uzbS��t��5GP�/�L�P�"O�TAS�L��I�ec�B��Ѓ "Ovr2��Hp�\A��V�'|رZ�"O����B�)Hb��[7nW�\�"O쁃Z8����9Ū��$�<rh!���9�&������x�ѦInd!�F�w��u�M[�x;�Z�]b!��0�A��I�� �Ƙ�B]�'_!���:H�S䞂gq&�����4�!�D��\�J��R�R�o��V�3O�!��7</ƌ5)�4{���Vi�L�!�D����H6❚*?6ly@�]
�!�������+
48Z����B�nZ!���+o(b�a�m֌BаX���*|�!���ꀤ@�U��$��UKָe�!�DF
k��J��M�e�V�RT�?y!�ͺ�pt�&��0Z����%\9!򄝇w�\��	+��@qѪ� 4!��Z��%3�d��k�4Y���R�Y�!�$·�DD�%̔�8�` ��_Y�!�Ċ9�-��a).mЀ�D�@!�MxJ�+6���ɰ����g&!��Y9 a�P�4G�7' s��!�d��.~]��+m�%Q'�5�!�ΐ|k�q�u��3��)��2L�!���?�v�suD�6Ge`J� �K!�䈸DS4�@``��bFB	�c�(M�!�DW*n�HS6��BA����^�!�d�+F�"r����@�ؐV��	�!򤞅RPP���U&e,��#G@'6�!�d��)r`!#��d'*1J,I;u!!��	L�>�BB�34�H[BL�!�M�ck��x�f��?�0a4�ɨ'!�$ZO�!;B搞K�นĪ�Q�!�ۊeX�ŸK�;����J�!��֠d�9!��/}�r��k�!�D�;6.��BHں#$
(# -�w�!�F�$�+q��V�Źvl5�!�$� �("��[�L����"*K�!�DI�(���ԉ��=��c�)�:l!�D)@Yf�����9�T8`�BU�P�!�^ '2���௄�@�^�!�Q z�!�՜a�ޱ�s��Ovq��.ޤg!���U���E�-��K.�?k!�DQ&��0jƧ6�<=ڡ��)\!�ȫPҎ�	r��#�ʤAvl�B\!�s:j�w�J/�d*ъӱS!�$į<�8tR��o�T�@�o��d!��B6x����iT�����>�!��1!�ͻ�鎽+��8fM�6�!��GK<�	 �B�KI|i�U��X�!�d�-��y��M
>+f�	�)��{!�d�v?��+�M��m#he��-1Jq!�ď�5�i�ϟ�\(:���v�ȓua�\��B¾pt$40f�	@��,��S�? �{�6S�
M3�?���&"O�I���:JF�Mk���#����"O���)ַ��h`5P�>���"O���b��n�Ph�bч�R�J�"O �� �طn
9;fB'��h�P"O*�r�9#`�`B�e��"OpLA�^�F@\tZq�W��@�9"O��Cs`�������e�xh��"O
�����q� �`g�_�vDX��"O�I@I�00��9��B�?jh9r"O���%7�b�1Ĥ=��U(�"OV� p�EL�Q���֒l�<��4"O�8��Sl:$���A�||t��$"O�ArAB��a�"'Œ_�ް�"OV����L�.˸�����"]��"O0PQ���NW�[&&�)v�� ��'BLy�OFa4+X'FB�)W%XZ���"O��j	� 暝����O��Yic"O��K��+�@��������T�'%��<��`�iP�T�D�
XZ�*��{�<�$d���`q�+K640�_x�<q�nV7;��J�i��t����cF�Y�<١�1}:)ᒀ��=�2tCr �U�<�b�Q49���ׁez,cR��N}��'���@��"��Ũ��-_��c�'NP-Dy��ɋ�M�d��#)���y��L�AB!�䛫���Q,�m�n��w�/������7�"�U+��t�Rq1���=iw�C�	ʟ�*Q ȇ7W��jw�4<)4�Z�Ow�6B�IDUrA�U�R����_�t����ͥ��';r��݌I�tC���W
h9��&D� �m�x�"p���S8-�fMh����P�~�|© §<ǎA�����I�<�d����E�ȓ3�(�@��L�}Bư���^�Q�{�֟b?���<ygC@�n.�k3��H����Y؟�!��'���:2B�,� ��d���^ h:���4ON��H*�&�� ��	,\�=��'�O�h2(�'_1�u�uY�0�0�a�� �!�$�=H�ԑBg�طcA�qUQ�H��z"�Ѐ��'_�|B���.8�	ZT��&W��ȓ:pؚ��}��<2$��k�0��>	+OܒO�pu���*��h�㏘8G�D
�'��P@��E�s(���T�)_�b����'Zh�q��;YE�W��;JT ���,�S�� ��wE���QC�Y���J�7%Q�$��Ig\83�I�z5�!ar��0� B��0[{�Q��郙I DX���`��D�U�8�+鑐^8q��")%�����DPd�Id���O����+�s
��)W�,�I��'1x�jGȘd����
v]�[�'P�����̯/��M ��Υjz�s���n�#>��	t!��X58�Q%�L7@����TϸP��,�7���w.6R��ȓ#j�P�ĤQ�zP17԰Z����ȓ@�Z��� C�#�Y�e�f��%��F{���,X2L�����1�Jd+�	 �hO� F�ԫB�KhZq�Tf�|7���G!�y��H1C�G��<�*��-��M�`b!�S�O=��fm�8T�z�: �X���gQj�<�S���J��Êٴ� I�sK�h�'��x����
}���c���k��y2�	N`D���ş�W��lgK٘��$#�OBԛfb�<e%����W1��ӗ"O������D�����>�,=�"O� $ukU�}��鰐�
�B1��'u�d�<I�L�0s�H��΋^�  �F�MM�<1�E�90�K�,ĉ0�T(R$�M�9�v����)���1
l�f�3�"}A�=�ynP�s�P���,
$���ʰ ���FyZ��O�2�3pW�D��$��"��17��Ӧ��>�����b�Пl �M9�I�&̸��0O~��d%P�"�1DN����ً�lZa{��DQ�oV(J��k����t+�s4!�ۑ.E1.R��D����ժ5<az����|�ɁcG�gi �x`�^�;(!��ԹG���� �=;w
�� �7���'�ў,Gy�� ����X�Zp��ƨD��yB�Ea�n]��Ȥ}���(�CB,�y����dM��LүLE�h�e�9�y2��<�*�M�I�(��Ξ)���y��'

P�c��[H0�1��B�'in�@�腹[��4��A�j|��k��?��h�-~��A��ɒ;0 X�F*��q�V
�i�����Q��
�<���KY�/� �X"OvXj�Ȍ����"�d�nA�v"O�\2v�ѐ'&�Q&�I8^��r��IU�D2�S<n��M�2C,��`km�(��B��,0�d�`�ޅJ�lA��7	U����l���p��J�|�F�]���((D��0�&�9\����\X8�5�!D����õF��×C_G+,p��)D���h�|.�DSh�:�� �&?)	�/��lXQ/*u�(�vd
�g:��Ez"�~*�I���:�8�"��B����^�<�!�G�P������&P�(xb�C[�<� #ٲ��X�
�v.�S5�~�<1��W�b�&��.��L�^�kg�Nu��p=1��D,Y���B�G	�wn ��f�G�<)�Eͼ0��`ْj���2OF�<)��K1xu&H��㇓6�>\����G�<Ѷo��;U�u�G�y��	`�F�B�<��b��%��@Z�ع�D	���E�<9�f̣6g�i���2�8RE�X�<	*e��B��/o���	��l�'��+ҧ*Xx��E��JC�oPY�ȓk��9�j�>e���%P1J�ȓG+z9����R!�dK�Jj�u��`ܓ2̬`چ�Y��l�'+@�D@���'��}�F+-���Ȥ�@�rR�8���_,�y�
͔#��x #�qgd�`��Σ�y�9RV��B)f���\��y�<'��y���V�g�~	�`���y�"*$��;�/^1	���KP���y"��/ $H��NM�u-FY�\��y�:<��� �����XD*��yB��$%���i��J?���^'�y��$_��(���0�J,��#��f�^�!"��SNjC�.�z�w/Z�h�40�'�1����Q��䉨�?�tW?�����B]0$����o�����@��?E"Y��Pn���̄�4L��)Q�*��ȓeֵ: G�"�|�0�P6R���7oܥ��@��
�b��]{���ȓm8"@J�F��[��i��̓8(ԁ%�<Ӕ�)�ӅF�UȀ��+a=��W��[ϠB�	
�Z������x���h�Ԑ���OL�"~jA�]�S�ҡ$_?Wz�S�`�y2�T�@����W,еl#����O�<�'&���f�A
|}��9?M�ܴ�(O�~n:� �-�V P;v�p��J�%��e�'K�'haz��؞_��%�%lν{��9���yR�׆�bi#�C�
#dT�r ݟ�y�a���5��h��_z�Q�n����hO���e���i|D�C��p=���Q"O�D�u�ř)¼���SO��"Ot�f��Ѩ�:fX���Ȇ�i�ўb>�O��9P��:.ll���0"����A������4��أ$�J��p`�-N"<�	�I%���)U�p��d���S~ �ȓ"�)�f�B#y&v�ؤ�؜nN�͆ȓa�@]q�l˱n�X��@�3&`%��*Z e�6�0�Q3�F�4UӐL��B�|"���pt��.J41o$�ȓo�"�0�(��D[`�tQ'q:����3`����R�J��hSںBF�x��@�
��ǃ�s��{��.i_<��E���8֏Dc������+m���ȓR���:�	�T�Z�*�c��`����4M�y�.����d��k�#T��z��<q���4��X��d��I������l؆d��8|b�Ew&����q��l�f�� 2��6 �0�ȓ.����Ǡ�0�6����qk�=����#W6P�'"I�z(�a�f�c�<���;�:�L�	Z(�tae�F�<AR�N-l�	s�_ s:��!b}�<�f�&'��� D�0��T���M�<IB&�G^0���C�(R��)�F�<�R�X2��� ���^4�K�~�<��� ���Q�����D�<���<���sA�ڊZ�]��m�B�<��#�"i+r��,ֻr�}�S��}�<A��A�J��{Qb4CuZ�{2kSq�<�"�\��ꆃ�,T�[d��b�<�T��<b�0��0A�(q��C�<	H�?eƀ `�	�M���q�J�<ـ� �=(]�G�E���d�q�<��n�
LN.t���m�t��A KY�<ɲ�ϸ$��a�m��4�,����~�<ɒE��}��0�`�[�id�u�\y�<q����:l��KR�i[�aA�w�<Q��[��.��J�v�z ٧	�q�<�'U�q��VhT5;� �rG�i�<agF�~[�ͳ�G��e&��P�'"T�����n#�dA�+Υ;�\�U�$D�P���8c״�@�o�B?>t��%D��3�ľ)v�x ��V�p���!�O&ؑ@�V(B`�Ι%u:lj�Ï	u㸼�R"Oa�V�ǻ)2R�Ð"�x�U�"O �3�]����@��d�p�"O"X{���+G�,ɱ�V8Kh��"O��a���/Cmt��¦J��L�zU"O�E�b��4���e�(Ŭ���"O��j���X�2!c��F���r�"OpŒ���/�T�ps�ĶS��A�S"O��E�>�f�
���<oOhS�"OSj��Y���W�U!�"O��:�Hƛ")僅�0e|:A�'"O��@�#rx09ӎ_��2s"O�ĹeI~>u-t�4×K	�re!򤟾��d݌��Ix��45l!��	Z)�A�f/�'P�¹'	 K!�����	��|Q$I��4J!�� �"DZ3y�(��,R3/j�5�%"Ov��P�ٜ�:���m:tR�ջp"OR�7D���<���!Hm�L��"ObE�Q�ݡBm�����y�����"O��Ƀ�V�5���Q)�:�2d��"O�YpgN(d|��yp�7{��L�@�'xj��^�>�	H?$�(�0�hQ�Q�QȦC�I)3⸙�e���@SVH�	E���O�HCf(�D���"�;�'21�ܳv�^>&���Crɖ����	�&���Kb���Γ��
���	%�4ySN��>���qH� "	x�X�'���)�0�3��F 'fn��fg�9�(DsN^�@��s��]�4�\�O��ЄL-��O ���W��E�xMp@OU�g�>e��-C ��`�k�\�j��'�D=�D_�����,s��%�7˔�LN�������^8��'
�����Վ<��Ղ�%�:Uה���ie��q����Ԙ�����%��֜p�g�/\O��I���]*�h#$G]`q:5� D��b�E�	4D|�E �'V*)b�X/].�PSć ^nm:%�� F�瓩.��a� O�Tu48
�N� �N�?I�M?mB��`�\�?E��D�t��`��EU�Ĺ��OY�����[U��a/�������2�̭��˫|za" �(�f�ϻ֨�YǊٟrưiJ�Ҝ{���'����M�p���+� ]n���K��y�S�j��	@E�#�,�"4��i�u���Xp��	ӭGB��FAۗ���Y�嗠�6�r�}�ɽE��8��H�"
I�P(���'���
�-�(9���	fF}2"�I�D��,�2�!C�L�$��!�6mE;C7��I�#��=L�;��,DP�#�p3���{�(���"� �,L�|�%�G!�����iȑ>�8��	I_�n�xKY���(����p��\���F ����Ai	<�>�0gHQ91d�xR�ڤ8Byj��2��O΅	�GA�d�8���J�
���p�\8t��C`J� f�t [����yV���'غ�>r���t[�%�GN	<}��cp��e�zc��}_����;v4HH�OV�lq��s���'�v����
Uњ�k�lW8
0���n��?��Y��x�����	�8��
4i�'��.1I��1�˃L��aX��x5��*d��D�_qO���Ǘ�9�,�+�0<T��" (N{d%ʃ�ӻ �H�Ӆ�+����G":� �c��3<UŸ�@X(OxV!ig(�f�lYB�H�t����soԓr�y�NA�!c��Z���O�SJ�B���"|�ԩ��f����v@�a/�� ���i_�y���l �;�4E���c�K�8�LU�C��R�A1��Gy����2N����͜���O�@���(- ���5w�RD�9*����c"	]XxH�@��o���!B�*5�8��e�X��˚�"����#!Q@H��l����6� ���;q	^����8a���b��5P���"5䎝BvFͿh� �O�H(*�٪bj�6�>B��:ddW(q� w䙄(��;M��DKp�B7���tJ�a�a�F��r䄗)u1O�"2���C�&	it��8�p5H��Ϩ �P�F�ِ���d��BLA�6-9�a]<�j= F���%΢�����V�`�&A�L�4�P%n�P0�(��5�Y:$NI$L!Q��D�
�|\����Cތ��ЈLiD�jԎ�|0�� M	H���D��C�tp�!��D̤�DL	OoJ�R��>���w�B5L�xt��L�h�j��~eԕG|B�)�,ph�I�-\�~�q�ֆr��5����Y�,X|]H�
�^hhEq�@"~l�B!%��v�6�̮���A&v|�rQ%���®�&>�jF��;U��Y	�@\V�'X����F	N��Y��?�:f��C��U�&�e��a_�]�| �rF�8P�kr�P>��5��.o��+C��#�y�!�[�f���'f��e*	{�ѢS��}v<#�4�J5�0o��Xq����OgE�锒��)��'��*;��@&����!b�Aǈ'*��5� �Z_�A���� 2d�����/Y��u�&�C&��9i��\x��,�����)B�_gx�Ȓ�U9wnvI��X>�&L��F�*&D�[��W�)���CIÖYjf��Ժsefm8DL��9 �E%M�j�YI�씩F��s�[P�1O �3 �R�ɸ&���G�^�*d����@U�C��%��*/#�0�=\^-z��^-։������`�!F��ȅB��-%�5p �<;��jQn��$ԛ�A!uK�Q�ry�4PFA���C2/WV�x�	�c�]Ѱ]?��"��&���Y �G�JJH���6%TQ2��� Xf��d��m���89 DDL�*8�Mj2��5E�I�sӠ�a�Β�'���"�Ɵ:��Z�D�<M(҉\�e1xĩ��#E���J�d	/U}ph��hP%l}��5ET�Jȶ�Q��d�Շ�XPR-�4l���lP!	�Wrڅŕ�O��'��*��)"&� �5��CpH
�jɕb����΂]D���DF�6��dYƫ�q+� ��$h��c�TN� ����{�:f`­LT�0)Ĭv���2eAE;e<�*A�ŊB��'�l�բ�	�0��UΟ�T�8� W�@�X]��`A�țw֬Z��W2@	+6%ۋ�����L(a���9��T1`Y����	�|΀
�U1@;E���P0��jE��L[E�N#K�����'�P`�q 6S9����i�D���lc��c�I|����%|y
��bj�#{}^D�c���:"Iҗgњ)�x!��ivj��[w�*��ӈ͖U���s��y7���9lf���슝E�,��cdG�h����CF��z¾�9��>LjP�.��=��Q�j���+,6��
`�0��K���(,ܠ��[. �V�!3kQ;f����2��~)��2 U_�(,��b���B���!ΜJ��$����с`�}���.�L���qNL��'�O�J���4�mӂ�1A+_��IB��39���"�,=���!&�*5�H>�偟"�>� ��;,X|�#ޚX���f@�8.�����۞s��07�M?i��{Q"���a猀s��6�Y�/����.�q��g �k���6JS�1�P������
\���<s���[G�1Q���S*V��f��92�^����Y�����5P��) �i�% �`�T�G,O��K�a_@��D*�֩D�j�d��1��OL-�eC�!���'H���Z�w���xA��`�⩃� �n����:AWb��e��(�*���O~�{������ςT�����!s�ʄxԭ������I�U��*gZ���'��&��܉����P~������ �&DS�/[)9�.��0���?j�=ூ�����cOS:X���&�0�4d3�/ۨ:�&�� 5�� �0�2`)+U�I�Cp�D�U�	� �@M� �y̴�C�-yn�x!����p/�4��,CԶ���K�'q@2Y'BLO;J�r���-(��MJ�p.�<��E�BѺ��+�d?�N�7Bz��p������AK�qy��B!7gH��F-����3��['8Jc�'�j�BQ��8���6
8钲+J�i�}��Bd�41 r)��Z�T�,�Xq��2ȨO���g�`�( yV#�Zfʄ���'��QV�a9�(�F�	.	����i��a(G�`�ҠqQŀ�8����!�؝vVBaG8�άB5)�T��qG'st����L�T��xboŔD�t�p�g�8u۱k�i�XPq����M��,\�o:x�Ѣm�	,����@�I��Q�VC�*�ꡀ�螇8���F���D��ѺqM��
��u��,!lO�=)�!����,�"b�� ^,`���S~ʤq1�J�'L��"V�w*��'l[$o��"�՜]$r��1'�yǼ٢�$<ٖ9`�G�w�Z5sӆ1�6�dI	"C��i��#�9]���Q�h�Ԧ�����aX�i�N�FCJMSw@�)֮�H&%�5W�\�D�qlī2MJ	gU�ACN	$BI\}��O��J�m�2mN<���]b/��!�悙�#��4��BV>O���B�T�n.�I#")��+n��T_*B�L	����&\=��. �c�Ly��
��5fH��!U�px͕�O��dj# d�'����s���Q�-?�Ur��ɾ���O<��x;$���nP�7��M��ӜdP��F�5���
剕��P'g��1�~\�
�R�Z���YdF���&T�x�T��.��}��A���&�A��G�DN��b0�^mr��a��p� $Ȯ��A��!���>� �F���{EN��+`���˝'���Ez"Nxv��J��5̜Ѐ5nL�I������ه����)��kon1B.T7bx�P`�*=�tp�v�"�DYC�A�������Ƶijb$y�NU�p�ɢ�tD�P)	Ac"���.x�7mT*:�s��0���q�ΰ@"T�Ba�=��d��Y�_�4c4b^�D�2$
R5*n�s3o�J�V�����@�0}�2�<1����4-[�V�F|�K!�ҍ� KS��6јpc��\��<�.�	�0yi��
5,щ�ˋ!�ܥ�ЫR�"Š�OW��UT9kzI�`�={�@)��f��X�T����TX��J`��$���W���$��vp�t:pHD(��m`0�� ]�Py''ˤ�^��2�݇ ��V�)[���b�A�u��+7A�cR]Q�� ��9#�.ѧ!k�#=I�- �5����`��⊹"�(���~RcS
<���sR�ׅ`0bA�p`W
m:&���i��!�h}H��W�t�����:���K�W�a3jU� ��y�#c"��(��*f�6`��(�%�MkT����3ulJZ ��D����MKw�ݰz��U� ��#5��a�4%�J�qp�B�<�=Z��C��(�kR�Ԛ�$��A�ܡa,4�k��$�L�>���u\,!�(�!w|�,Z�Y�%"�Tz祂�b�lb�'	�$Δ;��m�u�;a�~<*W!"Ê#�bͥAՀD�w`J'U�T���T�4� #4�H���d��j��1�֤11G��(���;�riZ��D��[�@{���_�>����Œ�Q�1$mЭЕ�ۦ}R� 35O�k�	fe^�!�E� K�djc�hO �$"�wi�V(���ܐ33f�C!��ٱ�Bi����`�ӑO�n�{']�2<�����:᤮F���{#F �\5[���g��''�ɺf��7�:�gM�,ZiN�ڞ'��tQ#S�r��؊�f�l&�V�T,iU���]�܈��'׮�9a�M�p�h�	�H�VIH��i&���F.]�7Dj��	a�\��$M�:�AӷcC�dw��IA;,��\�#�':2�r6�	)��b)�8 ��';@��(� ]�Ln��)���%v�A�b�ؠF�,d2fJ�*N�&�@r�'�REp��]�/�ԍ8�吅zu�h$�ÂK}�y�bn\	Z
���E� ���܆*�Ʃx�xv�@T�B Np�M�®�']�LY��@K��2�V�Z�#!��F�_�|���٠`Z\��%`��qxp	�/�*,ז"��;Z�E1�gW�C�l���-��fPL�� ��r�'m�,�wa�t���&#+
��Ó
�Z����ɷ��p��P��?�r��Q�V��P
I9<�(	e�6-e%P,�9����C	T�t�B���E�N�(�	]6g���7�I�ID�l�|S�.͑8�0�P�(��?��4c*С	�S�o�c5��T�H�O�>5�hd�J�9@\�05�Oj�"���%�
A��f�3(�42��׮f��,h�O�E���Ѹ�x!;& �P���P#�B
���u
�X���.*4�#S	/�
|�ד��X�󫄻��%��%l،�ȉ���TWV�2�g��oҘ�'HH%�܌3��|�H
@�̊x��`Zp�L�5TP�*�ONy�e��Z�K�&٢�HG�x��ͲD0
t!�.�(�F���b�v��8cT� 묐��
T�xyB��� w��R�,@;C��`5h�%1��5���)��CQ�ˋ��O��PA�@�#k��0�%
,@�����I�� �fH�`_��"�/�>��@qN�� ��eW"y�t�1��vlp @B&T�J�kBB�b�<�W!F`&�����F$�@�~%JUXã�s���s1��1i	�̸�b�>��p(�A;�O�(����;\y�XG6�b9i�o';a�r�A�y���9�|�4I��Hڕf�ˤ'O�z���!���F�1CF 
�(��#C�K�����#%H����˕(-"p��"b�P	ě}n�IA�,D4!;ɨ�(P$�&+�� t���M�1Ǚ�	�Ա�%���~u��<�}���	IP 8)��kW5{�F�y�Р7@�|�d��%�h�ڇ�y���'q�dӅĂM�����R���@`�V5[G2��P�3] ��Re��dE��dBJ?1�שu�| �׫�$���N09:�k�E�,]@��"�8��?�TΉ�GR�`)Q�9?�`� �,��BW�I	9-�P1�	�q�I�r	K"�~�g�	oDPt�S��JX��Rdşs2���>�0�s���%��T3�! S��J��#���R��r�	þu��TpR��7-ZE���$�w
�5�((��/���*��±J}��1#�1}�"%��ϯD�:$�t�ޝ0�2˧��,���z)�2Lv��F�D��YP�O\�G��d2��_��~��)_6���R��'7!�	+Q��A��u0s�B��Hb��3�~��W*G�n�!t�Y�+\�P`&�Bq�h�2TA!�y��%bz:)��(�hO
���gS����Ab!�,�N�iv�U-q,�; ���%xĨ�Ea�F�������ʻp��{��ܺ#s��j<<�Cą��2�*7������c�'e��C=��`Qv�՚K�� �	
�ʍ*�jaFk��xK�TŪ��G�����h�O䀓�
�P��
D��+�lU	F��;}B�HCE���C���/��!�Y� ��i�����xaT�a�>��a�6��e$ �)J	FMR��!Б��$'04e���fJN7(�B��`£�O`6$Uv�µ[��N�%6:y��l��dNH8G(�:G��扥'�\	AAK�:��x8��ۍq��hri��Z���KI`[��g�̤%�Vi�;�M���5㪑���sq1�ɺw��� n�.(�
���'�����4�v�R"��6Cp$Q�o(ғ@z�@U�W,��$b���=P(�qV��Qj��g���G(��0C�)�r�k�Q�u��b��3e2v���8t�~��P�� p��qj���w`h��I��HO�I�!oQ:S� 	t�N�3�©Kd�C04��q���pL��b��DW6+�(�%����(7~$�@{t�03��$!��X�rD��bζA\.$/A7J�.�ѥ_ F�$k5Dr��?E�4f�ɹbJ��^�:6��=H� Q�ڟx����i΀�	��E\�JB�./�����̈�� Ta�/"��͢��*lÚ�QP��GV�
Ҭ��<��f��dS"=�#��*D��)vIE,(c�<+�%?��*��d�NV�?Mb2���P�TY�L�
^Y$b4��ct	+_�@��잷)��s�<B���* ��M��Yۂ� 83��G{"��
%� �p�'9���0&��N��P�.��]���;g����O�#��i��$?��D&�N��Q0.����c�0")긑Ѯ��P�ӢH�9:ў� `LH>dr��� � (Πz�X��h�'�gS2й�f����}��Kȥz�ycv�Ia�
hX�Y��h�W�6fQ0ԡ���#��M���;v��0��,L|�Y�f]���Y�$�3(L�+A(��'������.9����:7&��3A����l���� e;n�9A�S8=d�j��L>R���3,������p��� d9剛v[��zG�D�Hԉ��dH�)7��.t�DH���şM��I� �[�T�Z#�d*� ϲ'ڼo6Qx �vj�r_
�W�_�.`>d��B�c���hwE |�����',�R��(�"�	pmR�HL���MҫV���Ҝ�.U�D��Ms�� �?�s Z�)���S�G$T�(��M��b��q�&�X�=�l �í"LO�|6��X3
��f��o8��D�%4v�����1<�"�Ig�CKT<LJSg���i4Iϻ�?���Қ��	�u6�b�6��� S8]�:�r��Q�iV8�=a���(HR��L4����AV�g��X���M�|��c�H(P��[��
����qy�/E*��h�W`��'�Q��BV/AYS��r���sRΙ�9-d�@P�Tn!1��{�ӵUl!)/O�m���*�<1�M�[�5а�O��@���!�0>!�a&[�L�k��2r��D(Х�oܓHk&�B�7Ob�Xe$�5a��t�C�_m�	y�"O���T�W�T���ݑyZ�IA�"O��q�̕�3��t��U(!��"O���Iͽ#EXɺ�)�P%L�I"O,���9 �&L0g$b����"O�̪ ��59M�P ���kl��	P"O$h��a��	����ަ:D��Jv"O�aJ��@�gL��x���h9^���"OF��֦IX��A���3I�J�"O�;�GL)
�B-�G�3Cd�ș�"O ��i#6��Q�;i�Xd#@"O�Չ�eB5R�V�Ѐ�":���!�"Om�7�"Fd�h��C��P1 ͈�"O�E��+Zk�h�s��S�1�"O�`!�.] �����K�H�(���"O���nM-N�^�� $�w��}1�"O:I!�^�ִɔ��+6�Qp�"OҸY��N2�p)b���joa��"Ov�{ E�W�L�k�0`�=�t"O�M�3�N@ ŧDW��IA"O�; L(yk�!Y��K6{����"OPDy�nP�@����b�՗>�:���"O�`�7jQ NQdk�e�<db"ON����_�_��PR�R*]ϔ�8�"O�	�L�WJ=�6'�(1��m�W"O8Ae�~^iS��E�R��=��"O�q&+�!��\� �Ey��A�"Oд ��$i�\-*T��8a��"O�D����']�&�H�x����"O��B��:�x�,C4��Ȣ%"O�(t#�lB�Z���.-���;"O�|IVɟG����#B�Ad�k�"O^���A���`\�#��8���E"O�8��5ӄx��@�?E7L	#"O��c#�1iɤM�p/U5& ���"O�;񄋦}k^ ���I�W�͢�"OJ�	���ms��i���o���3"O� J���<�� �@|�X(:�"O�ǣ*�L�;c������"O*5z��E�J����D�l��)ZF"Od��E�*��`�擻܆X1�"OTxq�$�9���7��-�ؚ"O���36���[Co�;����"O6m��i�$f�2hH���n6RiA"O.ԣbI�6� 8SG
#$<�y�"O^mAF�_��^pq�	L(�"O�ȳ##ݝC������%-QP�`6�'�|!T	˔T?�	/z� *��܌�9<�C���@{FbR_B9P�k��$h�O@1@�G#'n��q(4�'z|� �$H�e�1��4E�\��	e�9 ���5G�X�o8H c��M��Bp���c�J���#D����'�(��?�3��T0�Spmώ�%+��f��1$lSfl^	1�lyz�Ê���Ov\��I.��膅�:O����2({�����Ћm]�����'��6k��'�:�[��]?!: ����b�l\XB�Ӹu>��3�C��#H�ԍ�qΞ@{d�i�d�U��	\9ZI�B2H���PĜ�Ѕ�%\O�Ȋ!��Hu�=sD$
(�4 �!k��(��h�$�\�EB��J�Jà���ٲ��Ou�5K4��)�:�1+H�)��擌4("=!�%�1Ͷ��0!�%UB��?������Æ�D)�B�͊I"![!d��I���Qǚ��&����@"CP%K�v7���>u�ѲC��j�v�0�t�E!Tƌ�M=�9�BGh(���>�A ��S���	�BB�8b㦕�����F$@j�)('A&X����'o�'�Xub&� vFM�5�Έ}�Rt�XxiZt��tBI�>qu.��b0p&.¹t�8���OV9R����`Gc�*�k��ҹJ�~�cUn�h,0��C�q�6�ˤ�V�U�f Y�v��m�%H�4:��p�� �-S��ޔY�jU���,O� �l�X��X���1r�Z�a1Ã�"[:������e�=c�o> `QbX��4(0�^�v�B�i�#�'S4����e�L-����3w��Ѻg�"�F~B
I?7�����&I��[�I��`����U�V�V��U��#	�sS�œ�O;_	x)0�,ߕ9�H;��<(����� VV��I���ɵpV��ۢ�N���"�!�6:�%G�>l�yyA#�>��!�,3��	s�J�tf%�0bC�������Q#�J	sh1��B$(�bC$�Wv4���b��a����b��9�J���4]�1H�'(���=) �(5�9���90ݨ���;�2c��!WB�!���~G�dI�C+3�-�`�E�70ٸW��:���%��Jp�l�5i�)�XRa�p�V�w�6�m�q�'6����
$�Т F4/r1���`_p|8�aJ�	�j\c�֣�80��g�y�B�� �\��h��5�]��!Ȇ,t�z�^�\3`���L����E',v�2�́h�����D�Z��P	 ��:,ҕ�7��mb��ڟ� �W�C�^�ph�
�%`�������|�.�U��2��uZ�{�y�ъǶ���p/&v�Jtm�<�6 z�2��%�Q4*�p�����%���K�Y�u�B�fӆD!G],��� Ɂ�[���s��ɔcq�}�B����
���K>3�di�܅(�����$S�8h^��F��3���Bm�88���F�9"m� 0h ,�.=�#��9;oP�#�Fς6����͓>*��SƖ7ft�14L�5vhE�- ��vQ#�GGk��k3'V5<��j I7�j���q2�P-d�H���aɬl����/�&� �z�N��.�䒆�˝�f�Q��Q�c�T��R!��o������$�����*-��#v��o=� �q�Կ]�V���q�
1��!1��ꗫW�[�p5�T-c�d4�s-X �a�U��1MBR�rƉ�;ߜm b��$_�`oډY�$�P�皱	H��dw���g s�����K6���f/ړ<*�h�ܺ7}j|�ʟT��nQ;@t�e#��0�iE���H��cǟ�R��l A\�Poj�$LйEy�Q{5�̄3�91�f�6�''�8灗�`�`��ɴ*�`}��4�:��AQ�	,�Vŝ,O���ï��q  l^��녻같�`B�2\��P���N�҂Z�.��P�Hc��9�n
#)p����+�I�j�,�P[0�J�c�;d*r�"�4�Y��M�5;´kv� &.y��A7�ԘC�`<)@�
��*Qd�=�&���@l ;5E�0rl��A��1iurY��$�hqxM1�a1RQ"��Pf�9�&���,Q�7#خc� �2U�ϛl�2a��m�$:��Z��+VH���Γ��>y��CY,g�*�5�Ιh�"}i�**+J�#mL&��h@ l?Qq��je<�0��D��j)�I�����F��A��ӪI�����#,r�1���מ_-�D���F����g�0sh�����eњ� ���\2xrͱu�7fԜ�l��*���` ��8F���"hՋ4V���R+
���+�j�2,�J��~�� �"Rm�Qyt*�+�Lu���:m(�b�V-P4�����QD���{1�.26|�b�#[�E �)Č�8f<�&��(ٔu!ؤ���:�T�Ü(P����ϔ^z*���LC�I>"�-?�@T�G�̭8r�0&�@���-�Tp��J�-9D�����S����'�X�a֐`!���jye-�j≫9�,���[P�6<�e,)H.�꣭��<�Dk)=�.|irÛ4H��0	� M�С���Õ"?�i�D�����+�+;�:X)c[4H��8@!M!vI��q��A�A[�	�4MW�nx�	�v��J��H�`Ua�fW#sB��WJ��DS���~��.K8#z�CR�4)�ҋ��y���<"%P0�QҦhu/}�Ƀ����  �q�]R�]�`�,ݩ�Xv�� �O�-J��3v�+nH��ދ!�r���̰|��%V�|'���kR�E���Ħ��I��P��H�B�HH���:c����N���D�@� t<m�CF K��'v:y����M��=KFF�Ih]���VSÉ[�al�Y�'T�(M���04��=s�Ghez嫒��M+�f��`�N�瓭x��I�� ':��eĮ(~4ɒ�)�$.*x$�§`H�a��h)0b�._^P��b^GEF��E�G%OBA!�G��s\��ht��@�'DTmy�G�qX��P4D[qv@ʠ�T�"y�,��DA��SU���3���s l��<!cA�{1:U`s�J��n��G�@1BI��2����<Q�� ���@I?�:��mJ�V�x��w�9�h�!jÞ*Ҷe�F?z�����'�\�� �j7���u�li%o-u�MSu�J@D�a��IW�<�
!'��TD��H�A�?���,�}#��Ԙ �
���H�CC'��<���K��Uq�e>�I�~(�G�I�@����/0��@хh�d iRk]�)�l�aHΔ\�����Q&��m�R�G���x�EH	�f q!�ݤ(��ŕmV�,x�)I��	�=ڑ�h���:O��\/�L2���
�(���+���xu��@�.c����船'u,����	 *ѓ���,]���#��Szq �?*i��������K�Z Bӏ޻6�� "tN�<a!H��{�ܬ
"��9X= �éӳ���� ����#p��*�.�?B'2��� "�x=�5���d�{���D��(p2�ցY��B��D�(mC�����(�Z}��^m���*5���R�T63������{@��FP�^������>=��Z%m	�"a�!Ce�[ |L6Y�v�r��U���T0aє�!�'ht��Geļ8�PM�!�W$l1����+xRL܃۴H1������!>���Տ�}{����c��N�p$��kM�U�6�Gሌ6t��bAK��2���(p���D'v�Pb�N� |x�ԩG	Q�m�AY嫖�G���7GL{��6�ЗS�h
�o
#}{������l�]ae� B��$���/.Lm�4h��5�<4�DK��#=���"�"yJ���Ml�� �y�rmmڜb�$�&q��}�LE�Ua��qFO��%VpPrw	$j�JX�&d�>�`�$t��]��,D%Pk���GO�5�%�݆E��U��B� B��I�e�6��p�Y=n�N�� 	�"���S�8����&��0	��3BH��8�h�`�\T<�y9U�61����c�ǈ5v�� E#��W�XAS��>>�Q�XA�G�et���A�_⩠LZ�v�Q�G0�DX4//��L�2^0��T�=�M��%Dd잝W�Ǖ������u����f�ػr@vT�	�1�>��M�2p�^�˗A#J�^A�Ó�j��:�!Ÿ|2�Dn�P0,52�FZ�aR�뇁�"H�PAU�S!b��Za��x���ΐ�"<�p/_�PRh���ɇ�T�#�h���h�'�/�U�?s���sǕ?pA����#�"e_;uV�+��|��<a�4$��5���T>xU�W�N��4MS�'�lC��ɃL�@PrC̖
;ʌ��4m�� 9 �BAz���!��w8|��ꋒ�*�� �G�.~�9g��i��a�N)�,�6���P����Cp��́iNb(0�T|�)$��`;4��B��X�aq樘�dSN�Q��(=�ᙖd��!c���a8<�q"�0_�U!�H�?-�q�,�x}���Jʦ�p�_�	":���o�&�ay�R>{PD��Ş�u�0x:��L|viA�U�&Lv�ywk�%W��d`���FI�$�v�<`:�L��sne	���%#@`�1���?=�����HZ�\�a�O*{�d"=�C_z��`�MI�K�n�p���<�~�
4�<c ʘ�E!�@�D���<�h��O� ���bL�AI����mS�2�[P��D"�T#��Ͽ�yr�޼,��e9&"�=�"ɻ�Gޕ�M��Eӳ(�P����&|����FL<�Ms��5�ۤN�xUܔ�ߴH0~�cN�IYA��"$϶�×���pfĝ��	r�[I3x�>�1�P7:��
�2�Lᩗ囃�a��a�Q�^�0S*ԟ{Y���p�m�;R�L�x�
�}T��QL�6A��K�F�?q4��� ��+��0%i���D�	��5
G��D�Ή�&L�PH"C2�a@�*݋;f���d�A�W��z�#�B�Խ�#��O�Lp�4A�|t�(Իt@V�
f
ަ��roE�LF{"iݐW����ǩ�#��Ȼ7�.��a�JڻO��i��#dsX����#����a�ޚ��8R�E�1�6Ӷr;��C���F�����[��,	IvU!Ӭ�>gO��b-s�̂���0���[�dؘ#�6�o��X���¦X�yɒ+T?C�Ʋ+� ��h+dz� ��q���@��ő":yI��[�%��Hv��b�ɜ5�P��%4��%�D��O��I���\��q�K���S
%�t!Æױ&��$*'��qѰ��6���
��B�1pv���b��X�� J�t�E�ƿx�N��q��/UJDn�n}B�'z�:uĕ"O�f�R5g�>y�J��!@ǮWOL	��h8%xhAG	��c�/L��Px"�Ŝu�!��M�:X�X@�ՄL�z��[0G�4�#���CV]��Y t�-���Q���>���X!"VȊ��S<y�����GTx�̂��Ӽy��'��i����<�iWH��z��h��އX��Y�Ҙs�,���mA$��#?��A�E�L�:���_�^4�pf���clƭx$ hP4g/'�� I!j���Um�A+������
�e�� �ƂR��hC��5Au��C���m.,����'m�!������Z�M���R�5"��q��w�E��o�?4P`2U��W�H`*��'�H`��վ���A$	W?BօҠ�V�ܱ ��FX���d�+
Te�h�	�fl�Ŋ��@Љʐ��W�ܵ����Y��I5<���'��2\�2���GO� E �	2�(�Ƈ�"�N�)&�Q�Q�P�H#�?��*�=4�ڶ�W?Ef�y���8��A���,j&`��f�:�l����;j�Ґ��n���B蓋>�����a@���`�櫟1)�8����k���_��uid�D^��y���\a��4�JH�Lժu;�cK�܉96�CX��#�'O��m��o܉1�u*b�v 2M��^�L�ޥ�'�0���$a��	���.5q��:�6eB6�����b�汰��ѣ)}ax2OI��<;��x�i�sǊT��#�Kޤ*�� ȱn~61ʢ���Y�#�;�z *��0u�j��ԥ�<�ͩc��<y�$ �;#���7�Pܰ5�SgMذ#�i��:��`�BPZR�Ȃ{P��O]##*�I#��E'#�ҍдK��&�G5�����B,�e�d�	eht��ш
(��
Ób� �Wˁ-��<@b$΁<�(II���#yܠ$�"�ɀ I� �shҕf���'I!G��F��+� ж)���3��?S��i��]T�`��k��'�H���;tth\q��J�8��1��Va,d���c�R��aj.~=A��O�D��V�HI�뉲=1����L���He��]�V�A@B",X��Ŏ�n��E$����K�m��Y��> (r`�T+[���v[�L�;���>z��iF�V.QʨE�"D�\�Cg`�l��e�(V^�P`2d�48w�R�i�|A����+.A�� yե�\s�S0�i|� �F��TU��u�ܱ5��v�_
We][e%Zx�1�c�lw��8�F�O���N��W�@a�CM.Vm�i��Y.
�D�@U��t9��"UƟ���鲈���8	"��B"m^ 4D��p�M��<X���]-$��ZcDʈa�B�Y`��"��2*O�QA� :�<��;LN(���S?�i�#!�4՚`�t�� s\�)Dz�.���&��P�nE�\"�!��Z�N��0_�Y�0)S��_�"Ղt�u��
��M��2d���@B-�Z�P�� ��7_�0;6�^!ݒT��	
��a[��y�����u��OL��aɖ��"��a��n��q/ԙ�rmq�NӒ+�����1htp)әz�(a�Đ)@�-�ɔt�"�1Ag�� u\0�ڰozlG���1���<���U�E��	����	5&ʲ?ED�:��_L_�y��J�Pa���-G����i 
l�j̗bp����gVr^�)��&�N�i��%Srt�I7E dE�M2�nE�6xrU���HO����DZ�s�Nũ�e�
���;�*$MN�1x�)՟nW@L��Y?S��t�$��t�Zѡ��E����+�
�'KA�	 0�Wp��H��+]�hs��]�hl�9�j
T�'R�Ա�C+`��*wn�0��P	�A�uL,�;��@,ώQ��J ��9DR�^��b��-��H�a�rC0�c�A�/ΊE�j��%�<��A���0;2_�+1DЀ.,�$�>XPr�Bp�b�.Z��X=`Lr���F(���!)B?���C�9~��pb��J��X=7j����ڏ!�0�� @O�A7����W;v��P2�(���X�K$ϳ���� O+�����-ԼI�����:���2�M�G����Y`��GjfL���C�0'Z�r�o?.�b�DFZ�}/:�X�*q�8Ń�-<Ml�%�"C��hOְ��h� e��ç��,<���5.���(Jпy�.ݪ�jMY� ]�!h�#b��gN���5���8ꤠrX��tØ.)���`1$M����%�u4�p6��2?L(I�@��e)r�9D&��'Ni��댜}&H����G@e��� TX����7"��[p�1t&ڨ'	@}����}%B��E��Fn�D�B�Ҥk��<K0�Ԇ��S�x� (&`�b��,]Dy���b4���t�b�"��M�f�D,����k�2'��$Q�
݄itT�b���P%SIO�!��e�ƧE�/����+�<���@�P�@Qp�O�<s����(<�K��T�$��c���3�ޔ���,4�Ǡ��}��ɯ6��0oZ&�a�aǍ�aM�y`� 0V"6a" ���~�8ZV�T$k5�'���3�A+v�B�i4'TƩ���ɿ9*�N�Id�&Rڕ��4t*$X��2�hi�d* �2^5�'��A)l�h1G�	S����_�t���@(�jX���ʎ;��z�(�t)�C�R�����T��9��>��	���r��@��ɟ�P��ؒ-H�u`ɱ����C�9|1���^�y�vj�H�����_�!�ɥ�ֈ�C�&��E�7K�WQz`X�)Mq>�|��ɦ5c���1��<}S�O��c��2mw�BG
ʮ$]\����;'^�(�f'[�u���R�ծ��O���Z��<!AK��:v(1r._�<�6*�U?�S�q����Y�64�U���:s�{!��.BqO�� �.׀�0<�7H�7	���P ���
�
52��C��BT��p�i=]�f}���P��C�ɋe��s�jN+w��S�A)i6�C䉔o��!�	��K���p ��0e�B�I�N�6d�'�٪��������zC��x�ȰI�,Ǚd��e 1+�%x�8C�I�G&���E�G� )P��%��B�ɵP�T$z ���%	�8� �9n�B�ɛ.�V�D��P`�p��OSF�B䉦U/�`��`5^��X<,Y�"OЁQ
Ѧb�6�bFF�+Gi��"O.t9rm - Q�$V�ORв�"Oq��@�5��L�΁1��c�"OF��#��A�Չ�\Al��"O���bD/~��H�*>HFP�C"O�0��č<Č���(�:�� p"O��i3w��,��͝�w[�ti�"Op#�$K(���iW,I�B.���1"O���,��jR�aJ��ݫV�~\�w"O���m� �D(�+I�&� �#"O�D�BN/�t�)�I�)X�5��"O�p�b)�s�=����A��@�"O�\aM�0b���OXl8��"O��Pi���Ǻs5��!w��I�<I@)�1/\���I�d���'s��H�ca��M&��B�+FgRD	4�Ɩ1�HpÀ�6O�1@��Z�l+�]�� )$\�sv��t� T��J�>�p�IQⅼg��nWjX-�ᓁ^X�uS� �1H~��nE' C���E�5�6�x
çf������b��E1���!k��`fHp�O�����O�f��1�#�(R�S�aW�A{�I6�\'`¬���O���t��'$Y��٘hҝ(M<��#�3�MC�y���M�R��"���#U:�x�HS����V)Ud6�#�)�'{\�y�c�=uϺaz؁z��mZ�oz.]�=���i>� ���	k��5����x��$������'	mzӥ�7-P��RJɟjM��K��]\qO�%��MK>�����\�>�	3X�7�H��0�'�D
00n,�h�{�����'7��Ec��GL=�ë\��#�.<��{��)ї*�ڥcg��:�Z#$��F�;t��=%>q��X�x�;⸘��I�%���Q��ɤ>���y� ��?Q��>%ŭ?���iݪ>&��u��eb��!r΄$AYԩ�c"����Ls'&��>t�He��N�FJ݊��
�6�K��Or1b@�>�.T@��O�>���ưI��<��9x	��Q�sӺ�&i4��*�'2���� �p?aOҐ{��ͣ��߱p�	�B���&�&	��O��*+��s?%>�3��d�	5�\�!!
\�OQ���.]��T�p�Ŝ����it��S�.���)�bȨy�0ՊƦ��#}|��J<���F���|�M~zb'�QT�老j��s��Y���FR�$��-�>���3���A*$F:���g�p��չn�}�4BD103�����S�O�8=��R$/��ɍ�q��,�b���J`*A�" ,��s�"}R�@�%<[J��T!�1\.�E;�L�Ѧ���G+��y��)P�(�;��1hF�	*�~	�A��'P5r�V/^^B�43�!�b�ه0x.I���
�$B�I �J���"^���'�_�B�ɛ"r܉#JN�N48�nɽ$l�B�I K@����ɮA��p���0K>!�D�<p��za�	�P����4t3!��3i�A�$��z���a�
��y�!���.z��ʣ��z��	�h�0I�!�d�6]Ǽ5Ѳ��$�(|�'��
�!��Z

1L��̦wa6����!����f%�bL	�M��6�@�6�!�D!Aꂜ�A��5(.D�UFn}!��%c�`fȓ?G��$�&�	w!�dXNQZ(�?nwN�3�dН,e!򤛂��\�`�gN��qdь9@���K�}WV����4u��Mz�T��yBi���aP�іfA�8Y�%��y"�W�7��Ah%�֭^s��Q���y�Oӝ,k�Q�A-�:W�l��Яˣ�yBj�<@1(�0�8��Œ��E��y�)L�FC�@	��٘�2����yb%_34�H���#v���B��҂�y"Ǔ�l�d)sA��-vH���y"��;-@|��w$]��=�� ���y"l��ɑ�E�1N�*�����y"�
�r��GD)8�H��4���yrBͮo�!C�BC�2���P��F�yb*��a�ZX�a������q���y�*.2�9�%��#p���eg���yҮ;P����č�
��Z��5�ye�wN�P�A&n��,p� ��y"G�=4��YR��:��"�L+�y�H�3mt�U)� �b}��ȕ�yr�� 8 �Ya��H6���/�y���-��E��NW�J1BM#P�C��13�(��Ա)`��ӅIu�C�ɥZy[�^�����Ο4Z�C�I�,i�Xs3�#_��)��#I��C�I*��d"�Γ�[ǌ�!�^&��C�ɴ?���B�
*E�.�c�-�vC�I�#�n�I6/ף&���F��lC�I�qB�I͝����*b�C�	�B��U�c,G�B�|a1�D]��C�I3���å)a���re�M�a��C䉇I|�+1�ڭ4�ft�T�W���C�	�d��Q҈f\��2�B7I�PC�i�h*�3� IS��	�v@�'qn��]�)�����b��y���@��� n�tN�Qgh�s�&C�?٬I��"O�<�GjtLj6�Jp�2��"Of��'k�Q%ڵ+��9	t��G"O��������Xm����c"O\����F#�:`�v�˧f� ��"O�Dyg��%S�HP	�-A�z�`�õ"O�I��7KG<m���9]ʘ��"OQ	G@��O�tU�̻6Kȼ��"O���5�Շs��k,��{;:,�F"OƬ��!�E���{�ҏZ�b�{�"O8�{a�[;JD��d�D�r֕:"O��ʓ�zl�����)^H s�"On1JTl��d�����>�����"O�BF��
�j��#�=s8��2"Op|�g��+e�$BC�0��%�P!�$��iJ޸b��#b4�!�ߘa��D �g��Bp0�B�N!򄕦 �|��U���D��['ٍ/ !��||0-x1�2�����G�)�!���TM(�@#��@,(�;�D	+z�!���sVt��M*KB��!�֏]�!�d��Y���)�\��@��Ʒ�!�ʨ ~PSg�&2��`��Gh!�D�P��W�W9��3"�I�y�!�$ߠWyؼS ��Ь��ǂ��!���Nt���Soؔ`<�Q�E�i !�$ )[��XR�P�nA���Aܗj"!�d�!�%)`�V<�	��A�z!�\�c���P��,(K@��6��K!��'hɜx�@�=9�\�t��k!��K�kj��3LI w ���ǽu�!�d�*ИjD�^�o��p1���9�!�d�e� ����"�-!u��U�!�q�x�C�-Y��b�2�!�Ĉ�A^ ���]!
g,�LY�!�$��A�$q� �S�QBJ� r���-�!�đ�'[�!�瀗�<���e
�!�$Z�Hw����E�c�dI��=Zp!�Ę�d�(�	-� ��33�
�b@!��&:܁G�V��.�*��K�}6!�v�V̰A�>��a&-�x�!�D� FO�E�%�nd�Z�M��!�9L�F%Y���1fr���O�!��O�<�4ȱe�H��l�"b��(�!�D��@Tz�91
M'k⑪r���b�!���d����G��O8�`�q��� �!�$�5�ॲ�-B=�`�>!�dGr�ځ�(�qq� �@�B�!��J�x�4ؠ3�6TZi;�HO�!�DK�A�|���I�#?B��D�N2h�!�G}�2�s	."ȡ��D�]�!򤕙w��2���n�@�`��<Z�!�D�6k����QT�<%���7�!�d��t؆ s���8r˜�H�Ǟ,�!����TA�A�P�ԁ���\w!���LƂwIۉt��eV��
^!��=Ot-���0��3s0Y!�ƎV����]4c�TU��

(Y!�"uލ� =�>ظB���E�!��!v�U��[�t��Ύ.z!�ަ���n�]���e�
�'q!�(L�\���t�ؐ�7dK�`!���d����Z(\τ���BXkM!��+9�z���"�	K���AB�4�!�� ��E�Ǘ;$.���˚C��Ж"O�ЊL�w�\��(ג�aS"O�� �:�����ϻD�0�g"O�k��X�>���s�����%�f"O�`�A_r��b��*�D(�3"O�a�#T1��m���^)n:��"O�� ��цo@�U��U�e4E�7"O��J�!�&6R��q&]�(8�e�"OlYI�őʬ�(ԥ�t6hZ�"O[�J��Pd;)��0"O��0�`��Hm�tks�����s`"O H^�� � �P6Ԁ�"O���&�U��H��A�`��1"Or��+	�7�\����ˉ5f��P�"O����S�D Ƚ٠Ĵ�LA"O�Ā�E��C!�	��dÒ\"O�U[b�F�h����Wm�D@XB"O�X T��k2X���9{���t"O��`7��b��x�b+��0�|�a7"Oh$��$�vx��s��d�& �D"Oz�)��Oc�H�C�Z0<��t�E"O\����M�P���l��p�B]Z�"O�q�"H,I8���t%��*j�-P"O��R�(0L4J��� �'Xb�g"O�`Hb��,�*�ңT�6��X�"O�\�Vֽ.7D\�@Ӥ7ҼQ��"O�tQf��-@i@�p[@"O� ��L�����I�?r�q"O�rd��*ԓ �ȆO|���"O��;G�N6ABv���H8A�)�7"OP�b�J�'�P���3ܠ��w"O�l+��-u�f|"���,���"O���cλA}�xhDS W�f�"O��
�C�܀ �W��/��m��"OR�P���1��tC�P�^�d Ѥ"ON�9��N�<�ck� ���{a"OZ�Sg(�N_�(:v жT�F��"Ot `�&�:_#�`�0�֕^�@��3"OD�� 臽h�:4su֦ƺ���"O�l�ע^��/Ѝe�4���"Oh=�b�A B���`�Ι\���Bg"O=�eF��`���1~�8�!"O���n�%F/f�+��>�Q�@"O�=KCC=��	���S����"O���G.�f�;��@"�:�"O�%��P�Y��<���M1=��Y�"O���� ?+��Mх��e��}��"O�L��Տ �]�SI��gtp���"O^uڠō�N��Y5���8��g"O��W��H�H��*R4MX"O�|iv腲 C�`sQ�6=5 �zF"OD)B�KC h�fp;�D��y�"O��+ȼ�0�)#�P�s�<�Q2"O���Wn�>-����a��
����"O�J��U�m�*p��ޚ�I"O�Y�(�{d�B=ldj3"OF\�B��W׎0U* %����"OF��eO#TE���qCQ�k�(c`"OȘ`B�V:HFJ�I�a_5Bh���"O����3'l�� Ɣ�c �:1"O:���삾�$���ɾd�h�"OB-k4�P�t���X�� ���Y7G!��		��ړ�ŬKߜ}����+!��$Ku���(<Rs�1��\��S�? �	��54�X����/�0���"O�U�0�0%���r�B�:d���P"O����:,94!�v���B	�4Ғ"O�!���y*$"#	�=N���"OV���e����Ȥ��(<&�9�"O���%� -ra�5�Q&L� ;.`[u"O��(F�ĉr(� ҇$-�xJq"O>������b�Ղ��x����"Op��1kA��$%rQ��܅8S"O:�gmP�W~�J���
���r�"O�̐�IM,iF�X����"O���؈p��"2��6	����"OyRA9w2��ƈ�KX��P"O�e�SF�
��`'�8I���"O6}x��݉\�e8�^�6HⰡ1"O�Ivo�:1��r#��"[�l �"O�)��d��T�����gdT��"O�s���UB��)��>tN���"O��Q�A%e:��J��V3D3d	��"O�|Re�D�pq�C�M�k#��R�"O�)z�ƛ9(.�eN0��c�"ODH@P   ��     �  �  S   �+  �7  �B  N  ;Y  �a  Cm  �x    g�  ֋  �  [�  ��  ڤ  �  ^�  ��  �  $�  e�  ��  ��  .�  ��  ��  [�  ��  = � :" �1 (< CC �I �O �Q  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��e��G\���,0DB�1U7x�ȓfN����ģ���"'	(|�<�ȓ5z8uBFF�9!0\�4�C)?<�ȓJ&���GF�Mܔ��D-��ȓr���e V���)�I�_�zy��IJ�'\��ؓ�
CYP}��mɸ�x�'%��`�/5Z�}37�͂u���I<ى����VBYQg�����ر�̅�s�!�D�_b�	PT�Ժ�Bh��O��v��O�����O�S5i2p�$> ����H�Gn.C��u�P*5�Y/������(�7-.�S��M[�hQt�Lia�Ā!%���%%�V�<aWn�E�z��uK�(J����(WQ}����ɰ>��IoǨAe�e�v�Y������ RrG�G�0q� BC2b>X\�"O��#N��Of�� �@P�n4�
F�'�ў"~�A[�W�~��14dҥX�f���ybL�2|<����]c����m����dw?y����$�	z��(�;~،�R�����<��m�l1-OH�R��L�=����]m�yK��)D��  =�d̊���\?j�2vBi����S��M�Ҍ�pۂ�AwI���h�:���G�<q����;�T|� �%,G�ҕ@S���o�M�d�>i�y*���b��\h\0�D�/y�x��KO��y�l@�p���+��{䫏���'A��'�d=��"�9q�LA1A�FknT���d2�S��ȟ�;�`$)����.�<1T�����'Aў��
�c�����;\�y�$�i%ў�}*%�G�,��Y��t��-L1�pC�ɕ(�Q�Wf�,2q �kS�O1:C.���(ʓY���8V+��~Dv�W�F�` �ȓLe����!<��Q�'W���|�O��=����Ӽj�,�q��d�z�P�C�Q�<��(ɚ�Tx�"�H<0��b�Kܓtʣ=�����'!��H�T NZ�D�����|B�)�S1%� �8��	W����/��4�"=��E`>� �A�=^�����	MOt�Fy��;OhE��i�N�`�d�w8����V}H<3bA0Y
@��1h�!�*��l�s�<�O� 8v�IP�ߌI8��MY{�<�!�K�����쉅P�@�u-�v�<9dځQ��A���ز��}�<i�K��
� ������c���� v�<�Q��<3�9EH��N�*�F\�<1��S�|�"I0���⢔{��Z�<���7�V�rV���w�|}�զ�S����<iw���Y��
s%��Y�r�����S�<	1�F�T�rq�N��
e�.2��B�4B�ظ;�e���Du�� ߝ*\ZB�?A���"��2a�x�ݷ/�>B�(�^Ig^��:H
� ,-�B�I�Yf�̘�����a���ߐw.�B䉍2��9Ç悸+T6٩�&
�1��B�ɂa4A�S�U�[F��q'�R��C�I����S��%eȄX2B�	 {�	��Ɣ�'>�B%'(�0B�	�5��q���+HL����"B䉚k?��S�#Z��$�F� O��C��۲����}�C�k]�C䉘9�r�Z��N5e� �7�
�:�C�	�vRvd������ �c�+M���d��lnZ�i�B�*U;p��a��,G����&D��E�8�j�٠�T�j��,i�&��*,h�'�>�p'+B91XN��#��8X�:D�ё��A�dȉ���I�  ��6��������u)Ģ!v.t	� �..3����"Ol�3�AW�(̮�� �ظwV��a�O�7m>��?A�?qw�ח:����Bi�"+vx�g�{�<Q ���EIt[�ߠo������O�o�<�|���?#�<���
��%�6f�Kx�,�<��^���1�]$(N���� �<�ϓT�����XX7�]�4�<!�|GR�2"L�*�ɞ�<�Dm� ��c��B�I	A�p�K�EI\�l�'�Z�U����z؟Tڶ��.�N1PK4.��S�)�O��7,V�3�a�eʔ<��K	_V><$����	 n(��3�E�`��r��<��#<��韮�	�F˸=�?ݎ��e�G�C�)� �yB�(ֈ}�Ɂ
�l�r����X�E*Q��D��;~�p)�G��l�ڀ{��	����ȓzb�1`��=�%Sw)�!M=��p���Ĉey�}���@�?N<x��gٖ�!�-��T�}�(����E�-��Dr�����R�K�H���R��T����?�y�kµ&T�|��ω�r 8u�+0�ybv�R1dl��88��DI���?��'ᾜS��E���R*^�D�S�'!t���M#N�ܼ���ߧg��n���
�HĖ��I8G�
�8�@+:D�����pD��,?p����RI7D���7'��%x�4�E�^�D�7<O����$��ҩ*�)ۊ`-�BC+�4�!�D�d0y�a(�"�p�C�B�ў܅ᓰn�f���X�ƕ1��W%-W�B�	�1t�H�tʐ^\X �W����	^�'��<��JM�d���`�M�<p��TPHS�<Iǉ��s��H�e�9	FP0`$숏t��#rQ���=ц#�"� �W�����;�	�m�ў"~�!oN>w0��*`�߂�$8���y�*B�IfI��C�BՌv�"H($���'ԣ<Y�OZ$FxBF�N���Q���/o.E8aT	�y'�x�碑/Ԅ��'��sq:B�;'h,�8��_���B��4}����Dۥ%t�O<qj�)J�FZ ���i
#��@j�����hi�c�����	?K��t0��J �0��F)�+bh��dk�R�ߴ�M30n8m�>թ4!�\��G Og�<!�͐�IXh���5s��!Cc�<�W��nE��f+O2[�l�Ck]�<i�Ӿ(8�XQ�P-gɚpQiRS�<I�j�huP�"�(	���p�M�<��,^`�|��g#S�1]�%y%n[K�<ɕ �~�
�G�Zܘd	KC�<���F�T�=��#݊ �Ʃ �iEA�<Ѧ��!'`�a���^}�)"�U�<ѤE� -"&�nK�vU��6i_G�<���H.v�z�oj�t��GO�<aS`S�-��I��nF����K�<���. A4�s��7y�̬Ȑ(_K�<ٕd��"���{��\�=ːy�@��[�<1C�G^���:d���{�li�C!�\�<A`��L��� ])㍻�Ȯ�y��X3*f��aH�W| 5���y�KF�	*PA5jJNu�C!�y�-�הA�dhǠ����R���yB�S䠌�i%L�����yri��P]����cY ����M#�y�4V���xWC�tV�&�P�y�T���(x�X�K�eaiW�yBO��^� ��G�N0��pÍ_'�y"�nh(�CVFL�Bl��:�٤�y�+W �bĉ� A��p�B�J}�<9�J)s�DZ��ٚ^�"�5`u�<��k�e~�X��W,X��ٛ��E�<�s�M�}a�Y�ć^%a�����L�<! ��B^9J����Z �M;�Or�<IpNԓ7҆�5�7"X����o_W�<ق��-W�u ��5Z 
t��R�<�6�6�~tp@ �16T�a"�y�<�t@ܰ���	3-�.$�	�Sr�<��C�- 8x�펪���!�S�<�gn�"g����F)!�h�*� JO�<�A�T-tN�m��n;-�^q
!�F�<� �u8'���,u!�ƺG�Rт�"O�H��F-L�vԺ�m<Dk�(s"O�=��r��C�,�@<��{�"O �����]cTL�W7��b�"O��R��8Y����2+P� V躢�'��'��'��'���'}��'a��{t��$����rn_hȺU���'~��'��'hr�'���'���'V���n���4H��K�LaЁ�0�'���'���'nr�'���',��'���y�#צ����[=Fr�'?�'!"�'���'���'3�*A)��P���P�>h�#c�Р2���'�2�'Wb�'���'{R�'���l I����U]�D�B*F�C��'���'���'�b�'�"�'N���"a�h�����(A��MO�n*��'�B�'���'���'$��'�2M��.��А��4ItL�Al��'$B�'���'6�'/��'1҇\] K��4��0jr���y��'�r�'�b�'J��'�b�'^2�ۚv=sKH�dE��؁��'���'ob���l�֟x���ɦ;�I��BX��� ��2��I����	ΟL�	ߟ���Ο��	�����82/|�����-?s�UG�64s�'���'tB�'�r�'e��'y�R�t-� ���nx����
.��'mR�'�'���'�z7�O��d�>'��8a� �0k����$�� ��'��[�b>�'��6-M'I~6��F�N�
ִ�
��
�ppBǗ��[ݴ�?�I>QfZ����4udBq⌧S�|�Z7m�'t���R��i=2&D(�m�O.�8�<Z��USJ?�#����	�bU>*��(9�	ҟ��'7�>ͫt��[.�m��	4K!�\�0�W,�M#t�Jr���O��6=�����!��$(cG� "0HA��PȦ=��4�yX�b>]�R�#(��I��=*�
k	}x�=9t ��y�_	gɂx�g��Cў�՟�"�n�Pƺd�D��.l"�9�s�4�'��'$7-�'?�1OL����&J���bEFز+���	!�ɸ����Hݴ�y�_����OO�\_�b�K[�hq���"?i%��gG҄��Z̧[M�d�fσ��?���@�!�\�Ҧ��/�����_���d�<��S��y�-�_<��)aA�#.�Nl��C��y�'l�L�畟,	�4�����-Q<��<) e��t�n��DZ)�y"%k� �m���$Hs�D�`�Jܣ��n���eܠGg:�B@ǿy�D`2b(E�p&,��W�j�L¤�#-�j4�'C�8h9�a�e�)R��r�*@�l\=��>Yg΄"���!�`�{�'߆.�@26aB5$r�R���Ye�H�$u?~��#��5�0;%ڌ2�0�ڐ�@�o��(�6IM� �*|PEd��ID��
�7`��0� +� [X.�i�eB�|�訣w�	��z��f��q~���E�Mp��GN����[bʆ�G �ɐ����K�l���o��+�T��\`x�R��Q�9�틵1�<(1���
�B�r/�,�x0�)-]V����<�S�N�h��nZ��X�Iҟ��S����{���j�K�4Uy[V��G*�f�'��̱Q�"�'���'���~JG-p\0�I�0�V�
��ɦ��ݟ��˟����?��'*�5��p�>s�Ȗ�!Db"�������E��Q6c�"|R�� �� �tQc��~~�a�i��'wҨN*;$�	z���'4��@<9K�t���J�gQ��Yc&t�9�<�6)Z��O�R�'Z2g���f���H��X��␽;[�6��O �+�)�O\���_��'��'�f��ҳuv��r�V(��* I�>a1ItIĽ�'&��'�"�'���S66�Z�Sg��N���գL�(�<��'7R�'8��'��'9��'��Z% 4vМ7�U0��8��n�����O����O����OD��,4Z��|����]7QV5XU��N�mZ{y�'��'��'��-����M�ǋ�,Z�yf [�*�t����V}2�'�R�'n��'(�UI��';��O������y<��GK�{��c#�i�2�|��'�BnF���O<ɑ��%,f	�ܜ�ڝŦ��I˟��'��2�2�)�OV���b�i@V|��QdT��R�9��iA��̟p���<�V"|*��a�$�]�CT
<p�!�a�`���G�&�[T0�2�i_�맫?���Y0��,r�H�3�tE:�X��ĉb��7M�O��ɯ���S�t��ēj�Йꁭ�17����L�&���l��Y��Ϧ���������?2N<ͧa��l���̇kwȹG��hv�m��i��ݓ`]�@�	ğ|�3��Ο��q�)6>�{a�ؐ�U�S���M#���?��e�� �x�OPb�'e��3&��!I#$E��#F�r�����>���?�P�Pj̓�?	��?�@N hf�X�C(lZ�3PeG�&:�F�'�\�xc!�4�\�D�Oʓhn9`���0H��Q����x�Z��P�i�2����'���'U_� y%�]C�n�q����8��!ާ��%*L<i��?Y�����O�����`��Ád��ӷ��V�6 ����O����O*��vp��0��1�c�Ltp슃��K��A2rR�l�	̟T��Qy��'1��Y!����O�ʀj�EI0l32a;���t$���(�I��'�ps&�I�$e|�=��`�$	��5��*� ^�\l���sy��'�b��$��Od�T�\Bf�� R(���Jٴ�?i���H=� &>��	�?�XX����5'�$SE���H�7� 6�<!���?���t�O���t�? J(�6��oݦ	@B�>�����i��ɫ|0��޴)_�������䗥�Hb�`Μ�7-�Ff���'H�@ߍ1��)�g�	�x[���J�	����D��R�6���5�2�mZ����՟��S<���|��R�O������R��T���f��x�I��I�?c���I�BK�i��6`�p6h�#m���9׵i��'|�8:�O���O���55u
��d/�%S@����7�!�'x��'Ȏ�s�yB�'���'z��� i8����%��$)(�hy�����?�l�&��S����ry�8[
�(�w �LyT��&�?�|7�O�����O����<��[>��i��+�H9�i�
TɮMJ�����O\�d�O����)f:v����b��-��"Zn֩��Q'����?�����D�O���Gn�?��A뒪1v�p	/��bQ��{�Bw�z���O �$(�I�ȫbFL�"�7��+#,T���E��}:`�����Iԟ���Byr�'�vP	GP>	�I7t}�d�6- p%��3~@6!�4�?A���'8@d���N~�&#^�$�Q�2ԑ8��n���L�'�� ��8��ay��O�
łU	=�t�w���;oPT��4��۟�������
c��s)Bi)��:)8�Ek�	�&��)�'QbI�.H��'�B�'��P����L:�eV�2���P� z�,��?!u. �-�<�~�tITx��aB��,i�̩b�����sf������H�	�?����D�'��X:2�Z���P�e�Ϫk} (�8Tbw�ȠD1O>��Ij�&%���V�`��xXF�� @��A�ݴ�?A��?�Vn˽��4�>���O"�	't<��D�+�n!���Fa����y���.V�D�����O����Wt b�Zg]f�CB݋7Y 7m�O�Q9��<���?����'Yf�9u���y��l���ҟ]�JQK�O���U��:j��П���SyR�'H�	���� Gn���4nf<)�H�<7������	��4�?i�'-@%8�*�>А{��:HȚ��4{����'���'��I��p��E�x�7E*v�8L�i�9�ʑ�ve�ɦ��IƟ��I}����O����"�66���rƚ,�x�P�@U����O����<��o���P+�0��J�<L��80���#0�9@ѐG&�n�͟�?�)OH�·�x��G�N���̇p_`��1�Mk����D�O��X��|���?A��z��0Q�޵R�pRE�\=2`���$�O>X��B4(1O������ ͱl�B�ǃ�:C���?�$b¼�?	��?���+O�����<;&��5]�4 �5/[�}����!�'�&c�b?�Ұ�V�d�����,���e+3�{ӂ��b�O��$�<�����4�$��V�/�A�f��1�xGF��/)�l�U�Zd@��9�)�'�?9E���	�2�#{p֠	7B%=���'T�'�@"�U�����P��R?�ţ�;�6yz��I�y�]`��"�1O��2 �R`��؟L��i?�Q���,��&�W�x�QƐЦ9�������'���'�����hɎ�#��<ɥ�M�%;�	�G�X�f7?���?�/O����mm��[թB8!������E��`"F�<���?����'���BY�A�CHiD��X�R��f*ċ����F�'�����4P�j4cV7`�\��C	EP<Q8b�Ħ��	ٟ��c��?YsgH���0oړ"�ܵ)3 �5�:Ԋ`lA�Wiꓖ?Y����O��TF�|��o�Q��8iu`����M���-D�V�'��O���ƠSi���$�xmʹH�v��O��sN��cG���M������OP�;�ż|����?���{�,����e�Rܻ3H�_��p.��'�R���i >��y����2G�ؤ�a����/JA˴_�x�I�+Q�X�I럼��şd��AyZw���ѩ�6Rm�0ʫw��O������@���4�Z�I�O~�(Cf�&/%(��D�`���� ��a�L���I�4�	�?y�����'%6ui��K$7Z<L��oʃd�K��f�*鵠T8v�1O>��	/V<�vFϭ,�%��N�b"�^ʦ����4�I:ƚ������'|B�O$e,	󸼒QC�$,@\���ģ[m�c�T��E��'�?���~B
Μ��a��Pmv��)��M��;�$"(O��D�O.��"��*+����VL֤��-�'̋6���H�Ar��C~�'UW�����s�����E�O�,aj �9���� ]y"�';��'d�O�$�4$�<Ҳ���s긹C#�Z4ZJ��g�R�	�����hy��'�\��Bڟ���GF�� r�(
�g��J*���e�i���'�R�$�OBp:�H�Rћ����B��=�@�ss�5���O����O���?�ië���O�X�oߔL	&�j"�ٯ��%(ď��i��@���?i̗֯@��%��I��E2^V�����9QJ�F`s�P�D�<Y�j���+� �D�O����� �����Y�$)���1�ʻDL��>���g�p�3e|�S���
��yP�S����jG�P8����OB)PP��OB�$�O2�����Ӻk�/WPb�ܹp�&�!�!�c}R�'M�q��������D�O���/��ԁ5��nY�{��@��27M��q�����O����O���<�'�?yWFLZ* k���,CȾ�qn��?��v�0IR��k�y�O��OR�I%� hPA,׹_�n=�v�Q� ���iob�'��'��r��i>i��ǟ��p�T�+�H "��K���?H�8����-_kV�%>Y��ş���P�����^�RԬ�0�
�T�&�mZݟ�s5��^y��'}2�'kqO��pWE� a.u��l�!4�&0K�S���4V����?A�����O$�⇉HC|`� �JH/��d 5��ʓ�?!���?)���'���a/ɿP0�T��dC���!�a/��	l��O�D�O�ʓ�?��ۍ��D +��x�ğ9Զ��G�A��MK���?9����'��B��/��sش4cp��� �
΄p ��89O&u�'=R�'r�Is"(�P���'�X�'�@�G/���N�j�����z�F��'���LS�DFTO�A� ' ��zv�Oq�fhp�iJ"U���	$iM>m�O��'L�� N���)&F͚S6�b���a$lc�`�	�K���K'�~�q ׁx:���´pHZ��
l}��'�l}���'�'���Oz�i���hA'ʀa�aB�+@��BB �>Y�Y)��2��m�S�'P4��9ǉ��HM�	�H�cZ,m�#zq&����L��ʟl�Hy�O,��|6"0k",w��;1�	16�@6M�z�9��S���p#�II!r�U�*Vd�	qÃ:�Ms���?Y�?�BE�/O��O>�d��\���os~ܐ�뇹[+�|`+*Ę'�'�O���'��'XT$�v����ݸ�&��M��f�'B-��P�H��ӟ���G�T��ӥ�\����K\@C�h}�58���OR���O�ʓ�?��B�dL�F!$���[��b�y�(O"�D�OJ�d �	� x��b�	M9����b��S�����X�Sd�I؟���gy2�'�l��4ܟ>���P)*{��A �'J�^h���i2�'iB��ORm�4*�<0���I�����]�<Du�&E�����O6���<	�b4��#-�p�dԤ0"�d2�|Ҷy��7���o����?)�"Ǥ`#�D�I�"�X5H`J�L%.-sA�ڛv�',��'/��R_�d7�O&���O���J�p�l%*	ҢsC`L�sL/x)�m�퟼�'a�(����'2�i>7�+�N}ʆH�v���@�tZ�v�'�A��{�6��O���Oh���$�3�ڇ.̻j�]��k�{@���'`�&["�|�O�'ev��)�(�|8R�3�M�x�%oZ!;Ra��4�?1���?	�'�j��?�� x�A%G�V��9��+�G`��r�i��P��'�ɧ�Ě���'��0:r�%��ub A�'y�d v�z�>���O4�D�G�To�ǟ���ğL��ǟ��<7��U��?���!o�b�|r�E�E��O&��'��i��e�4�UJ��X�� j��F:��'ҕʓ�|Ә�$�O��d�O���O~�d�5"��l�4@rQ��Q$��ɥ&���I�����ȟ��IP�ӷ�ԉ����,�1��m�;6SY����M���?1���?Q U?�' RK��e=ֽ�����b��WA��#����'6��'Ӫ4�e�'drS>�آ�V��M��
a��83��5X�̈��Ñ�p=�&�'n�'d�'�	��|ڄ�c>U���G�MvȥWæK��5�MC��
>0�
��?����?A��?��F�'��Q�# 81�%Ta0$}	�͚P�6-�O��$�OD��?����<��'�Ľz&a��t-�Ѓ �/��@��4�?���?I��6W����	ß��I�?�zf��U�|��+�Dڤ���Ò�M�����OT9�;�`���O.+>���/S���#�K6K��y�я�1�M��?!�iA�>�V�'���'����O����<n�����w�j�R��$�\�l��y�b�?�g�	8
�Y�1(Խ bU�Q� �w3�6�^�@=�n�ן���ΟL���?y�����i�<M��&K6%�(�����u�$pش	�p����?!.O�	;���O�݉��=�M�4�]�>�0���N�M���?���>2��w�i�b�'���'�Zw�b�[䄗�P�0��'�_ȅ��4��Sˮ�S�d�'��'�EP#��?��%$��2��w�v��ףs�P�m�Ɵ��I̟p�	.������CgF_xe����>g��
��t�2���T���O��������O��d�OD�sAl�Yj�����ĖM(��v���\��l�ݟD�Iǟt�ɦ��ɥ<���n��p�F�]$TV�`��-K���T �(��<i-O`��O���O����%m�,n�52��i%@��VH�����Z��k�4���O����O����<������۫O�� <*^諆�5QR�8sش�?	���?9��g�7;�@H�޴�?9�S�9��(N�-�u��+
��t�q��i���'s�]���	�AF~���0�^ޭ�#Is�(�J���^�~�m��t�I埼�I��@�4�?���?)��+>�k�N��h!Ej � �T��iL\� �Ia��S񟘖���4/�F=�c��2%�|*ʈq�L�n���I�H����4�?Q���?)�'��.��}RF��>bpD81�(�!^5�Y���"g��I�,���Ē~��K>tKD%�d�U�.�.����ߦ�����M[��?�����'�?I���?�o���x1�N� 8���A7ۛ��,'��'V����t��t�OX%9��0'o j&�]������l���'g��'RD�K�m�Z�$�Of�d�O����4��&��抙T�:T/���b�ЦE���ܩp�2�$�)����?q��'O�H�R=	犘�O������Φ	�I� vB��4�?����?a����Y?�rE��xX����cX5h@����G}r�����'K2�'���'b� � ���}.��2�
.�y�'�5����'PR�'����~z-O(��ޱ~h6)m�f =�G� +?G2��16O>˓�?����?�,O4�X�$��|rEe߆1M�s�ՃKIĐ�0�K@}2�'�"�|"�'���͉>^�o�p��H&�:��	��D���듲?���?�,O�豵G�@�*:���9 �N8U�[q�8Jڴ�?�J>y��?�'G�.�?YJ��	Q���1H /�2%4�r�DfӾ���O�˓+��hĜ�4�'+�T��H��jY~M���R�T7��O����O>�A�3��~�ǃ�n�JTY�*αs��t��Ֆ'h��QG����O#B�O��s�@��TeF<-�P���3ajLnZ�����۴���M�)�S�1	`]�4,S�{�� ��%��u�
7�
A��hn��p�	㟰�Ӥ�ē�?i +���М�ۼ�ʽ����>Zț���Q��|��)�O�j�I�xl�y��K2W��1�c�զ�������$m�b,�J<���?��'ט�� ��&u�4���%�J�bٴ��C�\���$�O<���Ok�E(�q�f"I7n�՚@�ñB�f�'q�F�3�$�O���&��ƞ]#�C��9@H}�8�@�P��-b���'B��';�_���De�`�E���7ym����2�ج�I<!���?�M>)��?B.��?In��J�b:�����d\ġ�K>���?	���dS5@|ͧ��1kA��H�u��
^���'�R�'@�'�B�'��E�'�)�4o�&gK��hU+��
��H�sı>a���?	�����-R��$>�[��(1>�,�7��.����$���M�����?�\<I����I	�|9c���!N?P�� �pӊ��O��uЛ���'$�\clre!�������kY%~���i�}B�'����f�'Pɧ�i��o�����ѹ7Rx�B��ec��]���+��M7V?��	�?�!�O�8�R��@H����M�
�P
4U��I�2~|����\E��V�K����U���۵K���M�Ao3��f�'���'�$o7�4��\B�]�!Sl��Co
C������ٟ��'��#}j��`E�P�!(J�9��
�mʆ�i��'��� J�2�'��S��l��n���Ĉ���v"�<�6���$�F��Q$>�����IVPN���'0Y�̔�2���<���4�?� !B�nY���D�'��>�tP)fr8�c])RD��qF�~}J�-��'���'�2�'k��U�8�p��I(I0vaS�˛����SQ�Д'�R�|��'��b���M2Al� ������W'wn��
b������O����O��	r�3d?�nud*ڮ�����ŀb�ژ�s]����ݟT'����ݟ@{�c�>9�� =�$w��8"���2u�SF}2�' 2�'��ɳ"wp�O|2%@0$�J���L\�#+��Ǐ\8[���'��'3��'{���}��֨���@���1� YR'�΀�Mc���?9.O��k�F�S埌�Ӭib]�2�ٔ��0�v!r4j!��O���[����'B�Y���֯K��y���.`�`opyBG��i�r7M
v�D�'��dC7?YC��3�pq4�,.^2	@�J���������S�,�S��x��4�U!%%���j	 p�m�6x�1�4�?Q���?��'F��'��/�-�x���A!�ؤ)c�PPj6͉%��"|���E�$��O��<�Tͪ�&��/+�՘дig��'p2�b�'x��D��2�Ri��"�P۬!1��Ώ����t���{�&)%>��I��	*�n%��,ҫt���C�	>MlYqٴ�?ٓ�J"`>�����'�r�>1v��b�rmg�@w��� �DG}Bυ���'mr�'8b�'%�<>�гG/��	F��R��d.����'�"�'�R�'�'�B�'�$m`�.���y�+];P�V�q��+5��O����O���<1r.R�󩋲�䱨��̅J�4���R#	�������H�����	���=\bE ���O/f�ţ	X�H�'W�'�2T�l�� Ė��'Y( �vj��h�r��)жE"=)ƶi��|B�'�B����'TV�(�C�&GX�	��I�?s��4�?�����d��`$��$>����?�(a�ټE*v��c���3%�A@�� ��ē�?���u��Fx���%2���{����&e�k́	a�i'�	O�&p �42&��������D��C� �*�!*�"bO4 �f�'DR�>�O���]���^��9��Fţ&$�@�'�i���1bLuӼ���O��$�|�&���	�j�!����� ��
���4Z��]Gx��I�O.�" cǬ+X>M��l�"�h}Ф��������d�	 }j��N<���?��'��59ŗ*\dh��k�Yre�}"nI0�'G�'����+-��m�-���0 ��v�46��O�y� �|�	˟4�	B�i���Q 3m|0���N���'a;�?���?Y,Ox�)����O�����׼u��A#�ę�Y���$�4���0%�0�O\�
��� 	��!4��J�h�$��O�D�O�ʓ`"D��5�~$�2/<�R�J�q�"�k�T���Iʟ�'��Eyb@=|&�q0��8sF�\zu�G�����O���OH���O���
�O,�$��� a0��޷i`�Y#놾rE�A�i��|�'��	�&�
O`��s D0>��2RdZ*Ka"lp�iN2�'G�I&�I"H|����Rs �(���b��պ^�Q�dkX7G����]9.S?7��#-:�,sv�Iy��XZ���6(���'���L��'^��'���P��um>�5/�:pQ�W�+�6��O��MW(eGxJ|�Aƕ�"W�3����
0v�ڦ��M{��?���b՞x��'�܍��2zE�7�:+e�Gj�P�4�)�'�?)U"�.?{��K���F�d�����T���'���'�� y��*��Od�d���ed��G*6���G�>��T��&�ɡ1}�c�����4�ɑAv�(��ͩj�R�ЁfT0Y0�xٴ�?Y�A�	i9�'5��'�ɧ5�`E�����΀�9$UI! �����/~1OB�d�ON���<i���7b�d��0�Ҷ/��єk�mr�A㡜x��'�|��'���O�/4�*�G�%)"px�D3jĸ��y��'Rr�'~� #��
�O�J0�q���2��3zDI:�U� �	̟�%��I̟xZ�+�>�� ��W����pf�:�^5i���V}�'/��'��I�x���KO|��f��{�������u�r�2�ځ &�f�'��' r�'-�젉}�J�N*�0��q$)1�M�I�nh�dɚr�n�T�8�f�9t��7bO�L!�- ^�M��m�K�bDsM�	���)S?c�9���F��y�J^YH�BL�)'�Ds�bL�u��Q���ݓ$�L�0>;JT��KTS�m�MA�8��C� C�a����Wt��	���N��)��͓|����tl���I�f ��Afj\^�Ap�C͓h\t�!o˙h��5�Š 7M��A�Mv��d�윿Rk�BgnR)ti*@�T-pHP� �HǊr���'���'c��]6D�R��%2_�&:G�S�KX�rg(\�40����\�m����	v̧[��a�g�d�lB�b�p�R�	�E
-5<٨D"='6}�XC� 1�eъI%��>)Т�>%��A�"��2���\|��,[�B_��d4?�t�Y���d�'5��`���ˆ 3ƎJ[�p{�'�p���)M���k��P-���Od)Fz�O�RS�hBtɊ�>D H� Z�M�!J\��h���Ɵ��	Ɵ$����u��'l�7���9�Bi�~�3�kŜu���#�F�Z3���t/˴U܊HXǫ��v�<�v���(O��0����6�� �凿g��t��Lo�v�!��0Vl|z�)@�l��0�eJ�&�d�H�#*��ڥ&��t���]�Z��Z�g�9p��{��'���w��m��va�0j���_? A��n�:���q�&�,�ȣ$�,�c�(3ܴ�?9(O:II�I��m��ʟ�j�'U�M�`�R��0Q��4��䟄�ɃD<�	����	�k���y@�In�	^`x!�I�;x�|�tbD,�(��ݿq�Yc�݉nH�I��1��eX�b컰K��n����aA����O��n�䟸B��{a�(��W,衢hjy��'=��|���Ə2�ᡓl��4���U� �]D!���확�2 	��2�[#,l�JgF
3�M*O
С�@:<R����O��',Y�}��/�`�K��b^S �Дt"�����?�P�Y,���(f�����S��^>��c�W�B�4�K+Wnl� f`%}RMދF�l�R��
 ��~��)��D`����)[��X��O�{��ٱS����hnΟ��2�/�&4��0��:/U8�CT_��?�ϓ.���0E�9r H­ ;G����Ó,ˑ����@�A��͒#$ǹ2�J�
�o��M����?��=�4%	'���?����?Q����K#�|����
�e� 
Q�	*$
ui�lD)��O�"�R0CK~R��x��]�:g晒��Cs�ՖRY�e���<F��S�+5>�=�噇+w��3F�xۣ<�H��Ŋ6q| [
?MV*\�7KBy���?�}��ߟ��I1��D��㘃D$�{Wo�
#<��ğ4�')������W�s�&9�p��<
Z���N??�5�iS66�7�D�����<Yqō�|6����B�	ʖ��WHK�h�����?A��?1��t7�.�OJ��u>��QV��b�
�z��p�6�@o1���4v���0��.h���gvQ�4hE�L`�P4�kޫ;�>��qg6tF� f��*p�69#�,��`3t"AV�Q��y�KZli���cg��.�� �=��d�O���#��v��Knn��6�۰U�AJ�@U�6B�=�ȓ4�l-�g����t�8!�� r��<�F�i��P�43�5�M��?yd���m�X�i�ȃ�FE�W���?Y��P�	����?Q�O��d����]Q��A������/�%JE���b6��#a�DZu�#?�rH�0<!���W%K���j�,[�@����	�h�ŀ�d�Zl#��I�o����O��`<��B�"$���1%*�4�ϓ�?��������Wȗ�I�,���׍g���h�OX	m?c����0&m��Ò`�7����Hy�I�%�6��O��d�|Z�����?��ͮp ��@�#̐!�Q$M@��?	�|���dՋ�D,�P�ʧ���*3f2���/�^F�ѱ�Ϊ2R��V�PBgE `���銝r7��b$���<n����M�DB�(2x��ɍ�M{@�i���� ��ٰ�"��M����<Q��1���O���D�.Q]���@J�	G6����Žj�ax�� ғoT<P�AL�.����)!�@V���?a���?	v��be����?����?1F��ty��pP��#�(L���@L�#�Na%�\41b�G�ӻ=�����Wk�!
e���u�Љ�Rh�.��ux��X�Q������"�|sk��>ǖ�Q�-�G��O\��R�`�ＣŅ����5&�6 �:�P��-;]���<��G��>���OH�D��7�j�b#���.p�[`��I������O�9��*�(Ѩ��gKb��H+�7O��d��"�4���|������\���pCj[=uv �J KӪsƚm�kܖt�����Ot���O�鬻�?I����D4-nl`�A��G��@Xt-/+�Zm�f�	2w�X��F�r�B$�m�.X Ey%H
~������<�u���Z!1��#7�U-@:d�s	nX����f'H����Bc���'����&�.!��zfI�	����$e_ �?������?�����'�x	p��_�'=v��K��3L�M�
���p���C}A��
��V��<9c�i��Z�$����MK���?�FCU5j�nL!v��� �"Q�1�@��?!�4Ò�i��?I�O���h0NӅ2����'�����%@!���-6�li Ǔ_|�p�)-��fJ�z�K�}�D(�a��/#Ї�.X��D��9�O������L�8�Q0�11�,�x�>O��O��"|
T�ݬG�-�q�3,�)���Vs<�i����J��)� �g���[��'*�>j�	��4�?�����	�:>� ���7X(��0O�t��u�Ȕ���OD��D��<o��� �E�14!�`��C�*ыU��|Ω��<�sbZ�W�ZШU#Hk��L(	�Ƶ��mJ�r�Īs�U��򰍜-��� &�a�= 7���R����\� f�8}BN���?i���䧮�lt�tkr'�j?����ɇ�V����<	����<�Q 1��!S��0 ��� ��&�hO�_@�'��0A�9Y����fM�`�$|#��a�*���O�����cX���Op���O��4��at!I������Fvxv b���prH��lL0N��Dt
�QY�c>�%��X!E�IfΡ�f��H��HS��7>^��`R2&i\�	��7%�lhY"TD�4-^�\j`yͻ0��P�p�K�j�v��ÃCb�
p)��i�˓ZL�i>!�r�7m���b�	65��������"��ȓF�
UJ���m��� Q��)��?-���$��O��3�l"�&F� ��$�&]�u���CF�)/�nQC��?���?Qն��$�O���5ϒ*7�Zs�8P�7�TQ�(t��@�@3*5����Ȱ=�O��g:�y&�ҩDJ�3��@�T|.E���\�V�:���/c��$c��_9�hOV}9'nL�e� ��! \4@�t��n̸.���'���'��ܟ��?I¢�xB�P��`�l(����j�<	2M�4����τm��P	Ze�	��&�'���B�8�ܴ�?����p!�"�.\*<��4ܻy&Z��?a�	S��?������3��)	O>	��ϛW!�q�âë%�Aav8��9����H2@FM��~r�	�y� ���d��Vqt�S$��p<t�͟���4S���'��(���+}��1!T:'���Z�]�x�IH�S�O*���ҀюO�͂����x�
�'�t7��N����'I1-}L�A�nN��$�<)RA��
ٛ�ϻ?R�SSZ���ɵ8*3�ަRʔR�^�fDi��ɟ,���2G���b�ޯO�%�p������|*sLR/E*��1g�.<j%����`��3�dKEEÑk V�kV.QࡃC�p^�P@��O&h�Ǎ
�P��j�����m�K�8(�.�O2po�'�H�f��K&ZR�)2u�u�H9!���y^�B�I$K��sc�*��!x��*�hE{�O"#=Y�&�:i.�*���;P�0h �_8���'N��''2Q�r*ǝ-z�'�r�'+r֝�ä��h<)0���WTx �J��u�A� d��B2�XF'�_̧��7��=�1$��FH8s��8���y`�֓+c�����Ψ����#(T��T�Xʟڑ�AT��y�IۈL'L%ɲ��-e���;���3e�7m�ky��1�?�}����If��I��D\$v7r���p���Ɠ/�`1�@�ΖUE8���b�)|���'Tt#=A���?�-O��8�N܍V6ε�0�F4	i̡�)��`!Q�C�OJ���O����ͺ3��?y�O���jr�LH�����n��=����EaM5e�3	LD�*�x�U�'��p���F�U�L1t�Q�-�:*VXB�:Y��
���>���0� ��v�|B�J)挳W�K6_�}���X�d(��měF�~�$�H����O� ;��ˣ��1}��H��0>!O>���
b�{àѤM�(�2E&�S�2M�v�'剂G����ڴ�?���E3T$���E;dE.XI���"wU�As��?a"Җ�?���Ƞ �ј��9AuJ�:f�HH�q�1Z�Da�%%��^QRh��I�s���w�`���#/�0Tș����L��d�䜴z|ؗ�'@0E����?����?�k�`|�ժ!&���.�Z��'%���3� 0yRa] ��a�1$�v0�;�O΄og�f�Z�q���nK$#���	Hy��W�;��r�'��Q>��I֟�!�� �:��Ĩ��G�ah���؟p�I�,��8I0b�hI�P��@��
 �ڟ��'�pu南*���1�
+)JѤOzE Rd҅+!Rʓ�ϛ�v��a"�-"����#�~���1L�ڵ���]� mҤ0p��J�$��
g��'��'2�BM@�眹+G.�"�߃DDY$�$�O��dN�|�Uy��;!�v��`V�&�ax�C5�[9 �ńH�Y6Τ�+Gx3dA
�C0�?a���?q�NN�-�85���?��?y���l �Bϧ t��h�HYQ2�9<l6�CG�[�`�%ӏ%�n��T�aӣ���d�5/��I9Ԋ��efQd�.X���"�s���X�@��L�ȓh�(�FՔO J�x�����S�	�;���4&�
Z$��P�6s6��op�
��	2=���Y����#hz�1i��I�E}�RUM�t^l�'M�}�F����x#"�3��x����yr8O7-E���$�T�S�?ٖ'¶XĈ�2$����r�� F,����sh
0)��'Vr�'|©v���֟��I�1%
���ߛ;l� �!لq�ر��	O|��=!�@
�-}�4ı��H�s�Q�s$��p�L�$���+���P@��o�lA�'�}'j���L2��h�UJX�I�Q�����şD� ���cX��QF���(�$�O��m�֟H�'�_��'�����}4��A��)1������]|yh$
9Q�9�����I�M>)q�iG�7-'��O��4�,�:�ߵ)ۜ�sL˛x?�Ax"Oր*zJţ�J�;R��˥"Oȼ!�
�*P�I3
֨B|�<X�"O�DP6� �g���K.r�4�"OΑ��L�V/^��
��3�"O*=(7鈸N�!��,@����(�"O��1�Q<x�@x��M&�z &"Oz�bF�j���AD��tf8�$"O���ĉ/��"� �7l`��"O��9�oC��hx�.�1w? �X"Ov�K��(�H��uHK�t�� �"O¼�DŞ�v%�(h�@T�q�����"O,X�Ӫܟf>�92���6h�i{�"O:�8&#D�h�Tp��41^��s"ODy�,Qh �"�$�;o�"OLI9�d�t7젒fC�?M���!"O� �$ꎙF�kG��J���Bs"O�ęg�J,`\>9��AU�>��Y"O`ၓ����=RF A$ko�d85"O�X����9AT)8��.*D���"O��1��p��)����4[��!�1"O�0삖�h�
��S���w"Or-�'���J��y�BX$�`�V"O@x"�n ���QeKǹ�Ƥ�A"O����"Z9�N�p��b����a"O�)@�Ztrd��W��#V��U�q"O*�h��(ψ}"�ڇn���f"Od�&[l%��]�umz4��"OFœ�ШF�zZ"υ1wl"��"OEjmq�n�s�/7O��8"O�RDG�-�p��N�0BV���"O��K�HF�����&���:�"O橂�K�5��zu!Y�\`9"Op-�e��|��@J!/^�'���$"OF��W�SV2�{�M���	:�"O�, �ݤe���Z �D�xB�`a�O&,���"P�����+�����P���5�a@X�T��%qcә�!�Od*|p��JRȍ[��<�@a�@��'G��4#щ̘ް��t�?Q�?QlW.qm�*��$#�D;�"I��p��� ;rP�@��B��\Rub�1�0Ÿ��5Jt�Y)@������	���,̫y<�b�*RK�V#>!���#A���{1��lRDHd��
�J��Sh6��&.Hk�|�w�c�<�wH	(�٠r�7E�E{T@[�<��-n�)3��J�����s@)�h��=�A���f$zB�V"W�H���*O�$��ϔS6�QࣅqE�I�R�_��M;a��@�J�S�l�6���6�)� ��VA�-3�8E�ZBZ@(�' ���D�Nú���8S�Z��A�&'f@������=�.�qѦ�\T�{I%4A6�rA��G�(�!˙��O"H��.����s�@"�d8q%�X�&��cX� �#ƅo+��Ȁ"Ot��s�]�ew.EF�6uh�ñ1O��Xr�C���"׏WX�t��w�-�'{6F)��
�G�H��"(I�^8}�gk�b<�&(�,c��̊�LZ�0�4�#R*
B�0҇ߌ(I��K��[5�2��|JK>i� �/X�x}rᏃ�l��*�.r�'j� i�(�yx|p凓�<)-ON����E%Q�PIX�R9>8*�&��
-?XU���U�(�ᇫ2�	E��Q�J���4<޶�j�h����Q�D�*H��eK�f�G|%�1ؿS��l|�p!f�1�0�"IY��'�$(��A��'됭��� � �]YQC�p�'Hb�q�l��?H��k�j��;��B,��uw5����/�T�!����<��	��oLT̻���	�h	E.�؃M
m����@I(vI���/[�<<��?a�B��<�E�[ �E{�j�<{bڱ8�Ά{�''��rÃ^?E����9v��'4� �5C�3I>N�Â*��3^RX
��>23�9���l(BY:�%��@��!7�|��O,��2X���Z�GMHѠ�X�[�c'�-��!�Q�ĕÐK�����i>�X�O];Q��ɑSF��dM"%u��u��D�<�r3�ױY?�$PVO9��Ǒ�֣?�B��Op ������;�$ ��͔�o4����xW����Or~�>ф���mV�n��7d��עFs��YS�n%<Od��ӪW%7s�xQF- ��zB5x�\ �����pXў`GC >:�@� �5p�O����3T��l�` RM��9��7wG00��V?# |xۀ�: $��	! ~���nޏ7B�L��b�k�L|bS
�O��z'�߄{���	��XTiK�8����Gy�eT�x:;���b=&�X��
+V�F䉳��'T<h�k�˨�`�'�:9�����'o�IY���(!˚�z�g	*���X񦌴u̌�O����=��Z�l�'P�m��Kw(�:� �1��<�Va]�p�2�Gz�A!0� �� ��x�GF̜��q�GVaA�G�Wx��s�OF>%��@�ON�a�0�k0g�
J(���B�$N��=��k�`��'�"Q
�̹�p�#����Ma�I��cN���F,�]����hVU��8����G�a��v ���2��I��O��u)D)���"''H�d�`�
����e�>�P'O���$Ӆ	8pE��R+�$ ®ԋ'+2\Z�H�!�Hb1�_"blJ�z�:O9rA��&�1O2@�S�"2�  &�C�N���('*�ze(! O���UFDf�'_,9���my��Ņs<�=C�͂��yᐥ9WL8q���	�����
,�Dh���V�K�}��a��\@���Z�9�@���IE�<�'
��\ ��dPI?)��>q@d��-`e�M6��; J���,�5w�(�l�C�he q��6YZ�"<�"C[�w��=�U���Ȝ��Ē><w(��	��0:p�H�O�;_B,�'Y�_�t���C�=��Q0�Y��K�C�[}�dK{�t�kc��<Z��u����W϶峓Aכv�^̡�AL�?I��Om�e�?&�T8����;A���aM�$2��7m�:gxTty#�O�L W���On�س�ؒ��ke�M$<PQT��O�,K��	�I�h�	�hp�`��xpi��.= ET�>ꀴ���S�Gơ.�p<i�O�vP}�;S\��"�ӱV1Xd�7㉮Q�f0�'m��k�y�X�͓~��"���1��,F&&��w�ᢡC��GW�vR�*���(O��xw�2Ea��A��W:���OF����q�����(�m�<�@�j?�yR7O2��$��peF��ŭ��~��	�Ɓ�!�V0��FR�B�'Õ*`����a�1`��	�'i0��7��8� ���/B�
 ;�
:�j�I�uX|P��	N��4+Wj'
��	 )߼T1���A�2C�`V
V0(y椈�'.���2�H?)
	���V�_��̢�J
�ns�u��I;5D�mZ7E8n�CW��J�8��\�@ ��Upj�����q��4��iRe����z8��ф��=��e��
	�}"'�Z5�X�A$ђ`�ᡖl�2r�扸�-�.n�Q��,
�&����BE��x���4&���4�O����:D@hfˀ$t�����$
���b5OI@#%��P*�F;h�Q��E,M�ns�1����n�TT�o�D��2
.��2AU%a}�I�Y�As�SZ�w:Rpa���<MؠҖ�ψY� ۢ+7��̅�ɨ^ٞw̴�U�]=�`aS��؛R�x��D�<��I��-��l�rO����!�^>�a&��Gt4��2K�Y�Ұ�5M6�HO��3��z�|l�-Ҍ�Xј��?��˔e���Pao�2tˮ����`�p�0�dP7S��l��V��4���4K.����OX��ũ�7(�){5(���T��i>84��%/d�䨄�J��8��L�pp� T�u�ܻ�'�[V@9�5��~��Ν���4�)�������
�ի%V:�ⴢ�",�h�{$ J�@�X�Xf�����R�x?�s��]�APj��#~L}���B�~��'�ՖUV�<�s����y"�Ŷ����9Mt\$���[06c"0c��H������D �?a7^��A�NS�����HL�O�Lu9��Q�{H�8�1�]�V�h����=ғGo��`��dߌ��e&X	�f�է� ��@�-�10��  ���9>�rI��覅nj��y�'��"K�#����~r��(֥M�.���u�:\��)��cӺ��ҭ�r<~���|mZ}T4O
0jG�V=48́WV���2/C�.�H�*2j�7��݊��>�B�G��~r#ڒ.��E}��B�Yj���?B��� �eӮ9Y��(�i��c� R&���*}� v?���Z��V�4 �\A @�>]�~x��-�.�`L���p~Y� %�#nh 8I�	ϾU��\�s&A�=
d��� ���'�z��@�c�d���@hR�HS?X�WBʴS������=K4�2 ��M�Ԩi�m�	FE�*_\��7hإ&�>H�c�.ՠ��A�O.4�y����e�i��銵��*P�Ć4�����cW���r��U��+�5U0d-�db�0�>����-�y�C�0H.��I��-���F�[�>�z5�T.y�le�恜Gz�ɋy$r����t��=�G��M�'�Zm���C9C�8=�7���y#3�Ħ<N>O�y��fAK���0�~�n�O�5�֨�Z��e��-̝E���;v�L�(�l���'XT;s�p�Y*��˹=�N�[�O���B1&��vD���K�(a��'m�c���q�<������1UΉ�\F@4;�)�'o��x��b.B��(c�Fg��ː�>���W*�Y�ʚ�a$�-���kʛFmSP�FV���O�BXq6�ԙE�0�s�f���\di�k�D�,��i�ua�˓�l�t�[ �0 �$��O?�vЈ[�1YAG����B���?�a��U�$`ʠ��	T��	�p��?#=�Q�`���P~�1��D�?x�p�U˙����O
�]�D���~y��?�g?ySN-'�p�ber�8���O�we�pF�
�p<�nB!���"Ǹ��O���D��x0�)vT���o�O��3�	���X/R-���$Ոi���SRJK��PXF��VK�X
�b�;��+��|je�ux����
I�]�����J�� ��D�+3h�����:��G7�,��i�����BB�^��a��yN���42�\Ij�C!p���$��	v�&�#�g�'����0X���GB��9S��(�'� 	�aBO�?$��7ۮR���g�'�@A������!��ME�%�^-�3�8k~m�$��K�D��Ԁ��4��\�"�xB���a�����cO�}�r�A��E/!T����]�;�џ�e�W5�q#"fY
XP�)�
Р�����^RE� ��<� �]�^5FyZw�����	("�F��n�A����Ϲ_ܤxDx�4O�Ȭh��� &:, �Eտ3?�iD���@�lZ�	�m����>5�(-�De�t����Р�4^��dQ*�0�	�%ݦF]����c�::�ܴ�R��u��?:p<Р ��^�z ؕ#�WZ���/N��뱡���T�=���ƄZ�fŬ;���u�,Q�B�s1
n����;�.��%D!�@���=_p����	f���[�&̷Z+��`��
�ڜb"`�%��}�1B���s�ϧ�h���^e�Z�I7����DP5Ǡ��qm�%".��pK.m��?�v�֕���lӏPV�%S* �:b�9n��T�TX"���	��c� ���^�Y�F��'�~Z��D�~��q��Η7w��X!&�"�d�E���et �b�+fd�F$\f��̸Sbr�H��D�#�Y�@�Еb�ʍy�.F�0�^�zb��W?K��xfɌ�LD\+�O�� 	PAJ�3����W�G�����@��.l
�Ju�F�WǨ���֟���X�<�n���u�M�<��b%I$O�\��W���'Ϝ]��G�gY�@F}��֊t�<u+R�+R���Ё�	Zh�J�C�b���J]}"�Ǩ0�,�):���8����X!F�2e� /zF�qj[-G��ui�O8��&�E�-=Xz�H�(L7 `�����p����ȑ=��	$L�D�|�ۧ��
��Sf�=��4H�=F��� 㒮b�0FxR�C"��4X`�<N����	�E��i��(Yg���hI�!��O�,a$@A���5v:����x�:���	{�� Na�0�<��Pi΁F$���CG�Nc���g��.u��eLR�t%������'!�Nu�3���b��2eE០�ЈA7��ɪu$���'ߊ$qu�;b�i��*��:Ʋ���X2�ܰ!�*��~��"��zF��۟w_B)A/���C�cvP�E��4e���Cv�L 5hv�=�1iShO"U�����mK�	zt���5 ЊoZLM�4�>Ec�Uߴ���a��դ�z�D��~�ɏE�%g��1��-�Q�
�<ѢЯU�D�!暹'	�0�%�|b ƛv|B�E)P�DmE4z��b�/A 4�P���q�D����	5TV�'_��#r��7[�����ûF-Hɇ�ڸM	�FI^�<����-{&1��˴@�U�I�L��Y��dD�tCL�x�ؒ`A���#�5D��D@����&�� �t�cM�O$q�@�>.�\��$����y34F� N�hq*�%P�!�YSZ��a�J@ ː�U-�!�d�*MN�dX"�U� ޜL��H s�!�䑋l44 z�A�"����&�Ȓv�!�DF)�lEEi��x����Z�!�ĝ{ǒ`��يF�ؽS���?!�ؗl� |�׫X�z���dc�!�D1(�R$��W��[v�K��!������'��=P�mH����z!���B�
S��d�N��Кe!�� �mj�`C�P�6���l��kЩ��"Ob����*^i&�SaA�0b�`�"O4��pd�=R���F��XKL���"O�Ț�%#6�H�b�����r"Of�	vK�I��X��ڍz\����"O��$�#��R �I�?Wѓv"OzI��+Z�U[�G�(\���"O(ɓӥ	:��Ŀ"<<��"OJDS�	C�`J��aI�Z3�"O
�J��*n�EI�`	��>��"O�ċ���&��U�0h��"O���ET�t ���K�5{6��r"OND�G-
\x����h[��y$"O^X�t(F*;؀<!��ٿ]�0�pw"OL�6�3X X|�c��f�Z�G"O}��Z�PDrA����*G"O"���gՒ^̰�H�A����6"O����$�WL��g�t�����"O,5Q 	�j(J��r珹,�@5S�"O
e�y+���!^?X�f��R�!��ֈ�,pSTク4�q���9!��׋Xp��#ѥEF��6��0!�$Y�m^���T�Y�,11⊞
!�䄰sڨ�a�	��#u��� �{U!��4��a�!+�roV$vHߍ7!�M� �&Mr򮬑QEǿ !���
&;D�XE�N���y���'.!�D�7$���b�)Os�*�Ӂ㌅"!��ϒR�D���,T�a��Y���"!�$ �H�6�j�N��f	hE	M�!!�DU(���#HƸ&8�L���< !�$3-��AR����7!�dޛ]����_7f$(��	}�!�d�4B=��av�ڤ}"p��4&��;�!��<mC��	Q�Ū=4�`�s�]�!�Ę M�.LI��S?3XXH6�=�!�Dƾ��e�O�b*G�8�!�M�i)Fؚ���#B���ĳC!�$98E��g�E*՘0�Ϳ	!��%�v��CO��!�ǌY�!�4<f�hFf���|��	�!��O6U�D5��5 LG� !�d�3�H0Ɗ
��j՘�ꕑjp!�dG�ij1c�D)t	�S��Z!�䚹\�,���GO*yB ����$
W!�4v�f1jv�*̘���T	A!�T�w=�
��9�$����"�!��� t�K�.R�M[�%*R�[8c!�$�� NN��eI�v*کٷ ���!��C0������=x�JG�ʭa�!�$� r�hD�w��`�`f�
!�!�ΡV�8<���QJ��� G�!�DH*7�4� ��"[腱�I�Eu!���+7��!��Rv�AT���z�!򄀡p���p�`J��:���`��!�DB��������#�P-�do �!���g/(����rl�$�E.��C�!�d@�T�r�����w"�LV!򤌡\p��1��Q"? �!�9C�����Öc�t�̏� �!�R����3D��V��!��� �x{!�d�(@,:�P`&�� #�#ǆRr!�$�~�`�I6ƈ"\����-b!�D�$)`	9U�[)�������'K!�� �e���/��XR�e�rih�"OZ�05��G����NL 8���` "O.����8F<����7�*�"Orc�[(q������c�"Oj�R櫃7hiNy1��#9���{!"O0��@�Ѧ2�҅k0��/.� k�"O�0jǯ�X���v��4>!Xy*��'��'��8��iG$h\��fL�z$�� 
�'Al�QRl�3]^���DC:l�����'�*%���>��L�vE�c�.!�'��49���5R�=���Dhh�9X�'2*��)���\AvA��]L�u
�'��;'A�T@����$�&�
�'za�W�������T.�
�'>��w�[!
ö��'�Y,Ȃ\J�'�09��`��4
~���MS�\�E����)����9O3��gÀ k�m���S��y��;ĸ<z2����Ig��yR�M�1���Pg�O��V���$؍�yriA/3�<���gL6�F`J�aƱ�y�A�8#�y��N\m[R�k7��y�S]���%�d���Y�$ɒ�yB�H�,xʥ2oR�Z۪�K�	[���'�ў� i�a�d� ������Ɓ��"OBdӐᐖS�t���/Ȉ$j(�!Z�h���+ZM�$I���'_�s���k�0C�ɻ>�����Y-Ѭm��*G�x8*C䉩��"�+��h	b�Q�eBC�	�4Yr��Ԫ7�.5���΄!rH��[؟p���.#��x%�����e&�	Y���O&~1�
? 9���*��=��'̝��f��a��h	!\�m���&D�Lt�-�-���fJ��5#D��#�F:����3/��bu`�eD?D���Hܻr�Z�[�&�� ^:��ǭ7?��OO>yzgN�i}�<��nY;Z��s�G:D�X��
_��<�s�| �I��7D���b�7d1I�t��:��5D�hq�"�L6����  �F�qh D�����?zjaa�A�S&.��;D�XSN�8&d<��'J�!!KFa�wE9D������)���*M3l�(����3D���oúpvŁ&�
(p���Y0�,D�<�)�"�V�!A�۟`���j�%0D��2�V
V�NM���>��` T�*D��iTe]�٠1��?8lt����;D�< 㭋�mK|�*q]8#�r��6�$D�$+cHہ+)�]"���~�\q$"T���a�D�/�`�s-S/$��2�"O�����M� ��L�1��%8C"O�%��MG�nR"�Z��?z�
���"O�)bUII,�i��H����	c"O�4�u+�<���4�Fbt�ȳ""O\eȁ�F�얈�w`V�;��py'"O�P�mE�C���QƂ�R�,�"�"O.��.�=E�M��䊔-��Xk�"OT<hF� �Z���dL+��m�Q"O>��T<aۀ �6- �@�� "OF�:��2�h��E�%!$�C�"O,�
rU�s4>�s����%2JD�w"O�܈�m�F�d�`F
��2"Od�0�@�aDɱPKV5&��P��"O��2�O�F�Rɇ����Q"Op� Cʇ*h��-��H �;���"O� ���g�)@�4��M�S����"O��	���ͦH� &�b���H�"O�����i,U��B��X�̑(�"OZ��!�'�>�{E��"A��yv"O$hbˀ�YM��t�M.P;�"O�����	Q��!�!ؙI�:h� "OlPPN��`�P���+S��s"OxP�n��w���Q䎓 ��O��=E�$�Έ;�VTi�%�< �4P���_��yrӡpΌa3D�B ��(��yS<k@(ȱ@˘3f�H���`��y���6~�0I�B��-�� ������y�BŲTO�|����r;��Sb��yBk�, Mj|Q�M@�b������̶�hO��䙰n� � ����j�43@E^�lv!��Z>ɔd�D��n����O:cc!�d	��U%υ l<ȵZ�9+�y��	�{�k�A�c%�a�\�%��B�	"Y�~����J��:��Y�vC�I��t��@Ҧ4#x��4ş�r!C��$�n�����K}X��!�!�LC�I*c�b����֯MI.��!��#AVC�I�X�Q�j��|����J��}5RC�Izg.�CF�`%ʅ)�
8�xB�	�	����%C"�h���Ş9�<���<Q"G�Gb�$cP�[���f�@��(�Ob�����(w��!AcA$P���"O���N��r��݋ (��f"O6���U��tAĭS0f!�a @"O�4@��*T+(��v"Ռ5�,u1"O�<óG�~W����G�.u�"O ���HI:��Pc@^��Q9��'�O8�(���+C1`�3A)�i�z6"O�Qz�.S�w\*�H��gf4J7�'��'�P�U��<qv(R�-�8�P	�'��p��KV�Aa�I�"yR����i���O�:��A%��R>�ڰ��}8�'��I��J
�$�&y� ��*�Rߴ�hO?7m�h�x�@��^�0�h�����5�!�dǿ
�� ���*)����䆠�!�d�%V	���#
�:]�����ѥ(�!�WI���RS�'y��`�C@�g�qO���Z�P�����8POl�ے�S�O�axB퉮�&�j�*�#+�Ιs'B:"7�B�4Lզd*���m�b�"a�)R�C�	�,O��k�τ
L���`���}$�B�ɀn��iP �ޯt�IXC�[?i��B��W������L�j)��J#AR���D5?�uL�(|M0����n8�R%_T�<	G��@��<al(r>.���"�G�<��CE?'���q�鍠^��`F�KA�<-♈���MJ"��Dn%i��Ňȓy���K$�A�2e��실<��i��F+z5K*�:ff`QG� ����ȓ؝!a�ơ-Z�IIS &lцȓ�����k� ���[PK[�`,���@�MKF�C�%��G�@�@�X��~E>`3�g#5��Ԉǳy0����
X��a-N;	������1ez����!�tl�J�O�]���m3pD��T̹+�^%kc����̇)%����%#M� %�S���1	?���ȓ*�HZ���r�z0j��T�赆ȓ6h�\�M"Tt���F�G?9� t��S�? ~d�֌Q�b�B\�R�Ìa�X0�"O*i�r+XK�8W�@65!́B"O��*��� �.i�d�[�J���%"O0���߁J�\P��f
;l��Y��"O�,�d(	���j&��at��x6"O�!8D
چa.����� L��dҷ"O��C�^C?��VI
 �<mRf"O���;�0"��J(�0A6"O0A��]�!"�ɏD�%r"O�I!���	>v�򨍞~(�i�"Ot��e/k�R](&�u� �"O��Z��J%S��4��3�n�4"O���$Ж3���9���C�J|�"O� �3��*���Cdk�Ê9@�"O
��"놸���;w�1G�xP�"O�i��gʿ��(q���� "O��H�	?�X��F�7�4H�"O��ٳ��P18郢O��;��yV"OZ��
5-�:%������ja"O��A �[p�u0�@�[��Ic"O�p�d�%q�E��I
,a8�A"O���VC��j�٠��g\!x�"O��&lV;"� &���V�U��"Oq2+�<��G	A���t �"O� � ����=�a���+�%
"O��,�
ؑrQ.�:���"O<3�,��*\IQqNE�N�v�Q�"Or�!"��Tj:e9'�S�0� �Y"O6e��eߖ0L4H�RA͹�~�"O�(Հߪ-�q���3R�v�q"O�⇢_�!>��ѯ<K��T
�"OT)�M�=(`��o���ʸ*�"Ovd`"�M5+�j�QՏM}�6t	�"O�(Ic鈬w����,Y���hp�"O9��HF�N����KZ �e"O�]z	F7J,l���:��"OdA;#�t�H�`��7�M!r"O�X��e�%�N9�#j]�.l��p"O6�!��4��}���Ue��6"O��p�2R�܁�ïc8�8�g"O�P+��_5�kҦ\ F2ZD��"O�\�6��	��)iP�c��x�"O�i�fW�\�ee&��97"O���q��ML0)�%��E��"O�-RU��R����ўp�xKu"O���� ,N��C$�4t8D��"O�� a�Ze����$Ôjl��"ODa�	2�Td��Ò�3��"OJ�s����]*�LȀ���ܚ�"Ob�n�Ӿ�s��g���"O�a3�ь[$�h3!�8X�Z�B"O�d��H�&i�)�w�[#{5^A`�"OF���+�"mDԑ$�Q�i�`"O�()�D˥]C�T���&䄙C�"ON����KzB���c�u 7"O�Ta�EV��Ē���=�^���"O���	�c��p`4�Wؠ-�a"O�)ȴ�اg�8q���	�I]b�"O�@*��E� �1/G�y� "O�(����2DY?����d�<�$ㅐ�:8d/ 7�x`Q�f�a�<)g[
`� %!�*K�*�xhy�J�X�<��öv���(��Ȅw� ����{�<���8I:�٫��+Y�(��Wl�<�  �ɲ���h�6U��)�5g�	c�"O�tb�!^�t9��1�F���Ti�"O&�v�A�S!vđ��\�K	�dy"O�A����F���_"$�1�"O�}B� E�mź��Ú�s��0!�"O$=���ؿK�^������}��"ORU���&(�R��̺yA�- w"Ox$s�@�0GD��T.)�Q�"OAq\yܪ��B&75DT��/�D�<I�//H-V!�d�=*,j��SB�<	cC��z4���牀�w��ct�\|�<y@�s^iie��/#^���ǫ�A�<���G9EK�{�V�bDiU�E��C�I�]a�a�lP���$bv#J�
�!�I�8��-��a���T�[�B�8�!���V�L����	�e �Ȱ�!�����`�%��9�&P=�!�$	�2|�h�
Y�X�r%�&&ͣn�!�$��SE� �'��:�Y��x$!��2J2��! a#2�c��b0!�F�o��y�B�Њ@���O�`!�dWu,$0cA)Ξ�\�o�:\!�D70C�ЊV�H�����b�@!�P�E���7HH�(7�@e�+d#!��լ]�acb���\��+�(*!�� �@f���4��_j���p!�S	$ʌ�����:�^�K����s]!��Z#,���C�ᅴy ��4fC�ZB!�I�p����b��z��\�`�PI5!�$���ɗj�M�(,X�@]V5!�*�>@�C�7L��%��o�o2!�$H NB�pr��8#��-Y�@��Zy!�D۟;G��y�Dȯ|!�soX^Y!��:RQ�3 �td�ڳ��,!�$���z���OZ`���	'6 !��&1.=����Dix�ٲ�(\!�đe�0�S�.KBd�93�m�-^*!�dΥi���ʀɓ�>�2`�Ы�;!�$^5]ɲ���[�JU�M�� ɫ!�^~P��C��eP0Ě1N�/P!!��%
��@��3V�����o�H!�4�,�!�
0a"�(776!���I�|(Pg�VHzQ(�#�w�!�d*�̼Z ��j)��"M0N�!�d��V�F�Q!JH�tj�ڔ��o!�K4p�uJr�O�?b�|
�	��w!���Flu��,�3`�Z {��B,XK!�Ći�H�Q'�;t&�)pC�!�!�3.�*�(b'2}d荀�Ҕ\�!���-X]�Lr�DF�V_�P�E�&�!�X�V�� �߬1{z9KФ�@u!�M�K�&�A;uz&�a�	�R!���_~�d�DAڷJe*Xӳf�oK!�ȇ9�hA�#��Ot�%Y���9=�!򄑠^�D�R�ۂn��Y# �m�!���$[���1���0s�&�9d�k��'\8�a�ӛ<rp��'սm���3�'J�����0jf�kJ[5f� �i	�'�"@{���s�x#'�̀c��E��'��A�%�2��g��]:�x�'�q)�Ŀ4�F�[pFB.VuPQ�'J��Z�i��]�⊏�^��P8�'�Y֬�|�Y򯐭Y4:t@�'w���,~Lz�Ö%ܻTn ���� 4�0Ɣ�@��+�eX`LjyA"O��8� T,i���a#�3F58"O� 9��ݙ,���U�P��	 �"O�鉠��>E� �R57" d�%"OV�b1��XP �`a�?J�lؒ"OL���	l|T�p!�M����"OLuy���1����@��I�&�"�"O�a��X�j<	p���?/��R"O�� ���%F(L���ǄO3��a�*O~�C�ꌫSX������B	�'0*�*�,�I�8mc0`Y 4��'�\�"w�A=�l8q4<'P����'#�ɐɝ�I�XH#ψ�����'���iAv�h�K=�LQ�'a Tx��Z('h��;�Ĝ5�01p	�'.�(/Tx	zd�0.4�Y e�9�yD� ~>�U��I+s�be�@N�y¦?Bl]�ł��{4\�:�N��y"-J�!��1۔�Y�)9�4´���yR�ߛKh0}Ї���)<ƌ�cg_��y�N? ��!m9'�]�e  ?�yM�L�"daeV;�~�IRQ.�y2˒+<��%a#bD9�P� ���y�A��_��TK�	̉[��� �y�I���&E��ǋW����ON��y¸԰ ��U"oՠ�EL��I[��ȓfPn�[�h��EU��1�Yb~Z��`�X=�DJ��U��H�WQ�e�ȓz�xL����y��9Z�/y���t��T�F��V�B�U,P�!�䒠	�p@Ƒ�S,08��$�!��_�:��yVB�_b�+��I8s�!�$9^�9(@�rkV�-`�`�*<�!�Y:
񂃠�<6j��G�W0�!�Y�q3��GM��iT�<:�!�ʄ=�r��g�ˈIԘ��q��C� %���J2�4y7Px 0�Al�C�
:�H{�H�>.,\�7(	�YL�C�I4m���P%�6E$|r�� �`C�'k���bQ/S#`��F��J�:C��.�����ˑ�Xg(�x��)	C�	�3\���ϖw��̒%k<��B�%� �� �#ar��|C��ȓV�$s��_�7�<�S�K�vpl���s���nŻR���G�<k�,��r�%8�E��1��D���4��m��AZL��$BC�J?�Xb6�
S�f̆�e�@�%l�-\ �bQ�Lkv��ȓ_��$A�l�"҇��J����ȓ5�2��6�Զ_)���2���a,�݆�/�����4|}�`�H�����PP�󃕉w��$:% ,&"���m3*$x�kǂQ�b=JF�2c�.��ȓ�H��ホ)<�`�)wg\*^��,�ȓ�|��u�P�F��5C��_ j� �ȓB�̳gžZ���j�f����i�ȓEd*�����)D�M��ꜛb@,D��4�yrg�-Wà��F�>�J؇ȓYV����U�y&%�U�\�jt(!��8f� ��%�P�N(��8fi���j�cD�CX���bEЬ\w�ȇȓA����!�^㸱�&ޥ5U��ȓ%��t��M
$!���傕d����ȓc�,��Wᚫj�@r'��X��S�? �iy!%�kh�E���cd����"O���Q�6}�2�(�Hr�"OXȰ�k�@c�ѣv� }B��A�<�.E/I,�xu��Č}�W�RW�<��_,z��9�� 99���J��l�<Y@ δhux�ʕa���5�d @n�<��FKu;.Diր\�`����.�U�<Q��ǭ�
���ȫ,����@�X�<�q��]Ą��%Â&*Y�1f�W�<q�#H� �
Q�B�:�K���S�<I�+�5l�����(ĿqY.T���O�<m��p���#�D�zvl��e���y�J��,��(�6�2kq������yZ2~H)W��W>�z�Ͼ ����M�@9
�KG�&G�UR���5�̴��ZU��c���u9>�j��X�:��5h���g#���@��K�[�P@�ȓ>t*�+�3S��Huh��r��Ąȓh\�S��!1���JFE�=�ȓ|3�p����U��=�g��*z�y�ȓW�RdFO��[d ��&�����%�X\9���JY�$v�U>q�Hх�K��E�2�Ǭ���bP���6	��y~��M!~R
�֎ȕ Sp��	O*��a�3Y��sT��d�l݆�h��Es�&L�JX �ѥO�#?ڜ�ȓG������\ dN^U�#��aU�P�ȓ~��	����t��{V�N9���ȓ":4xE
�_�\ɹ#K׏N�^\��i�  ٢`1H8�۴x����ȓ*3t��1dÿ J��S�E�hx~�ȓ#� + �/��@��g.|,��ȓW����#�E/'��q�&�'.�Ji�ȓF�d{f.Y{�����9;��=��p��j'�D��Ȩ�R(D�m�݄ȓ3����юB �`��P�<��ȓj� u�Ղ
~��Q�	$�l�ȓ �`���2r�x�E�-j�<����&`�GI��,�p5&��!^��ȓ��Y�C��	������&���u����&�<M[��0WB�;z����z0	��S`�٘ �<mKf��ȓmo�D:"���+��D�aG��RL@��ȓ3ƪ�HS���ez<0���D�Q-<(�ȓ#��e	ШԾ����;�J����J
�BL�1젰x��]ara�#"O��+�-7�"�	�$ŔS�Б��"O�����$6�
U㞬'�V�a"OIR�*8w�М��B�
$�X�9�"O��:QC$r�h��A�Ԙ��X8�"O���@",4Ey ��a����"O�9z ��;P�R5�8�>;�"OfU
�b�'Cn��J�{����"O*���IL kHn�أ�J?Ҡm��"O,ݣ�c�K�\0���*֎8K�"O�<��B�h��0�`�ڸpZA��"O0 �樈��\ҥ�ؤ?�43�"O��QP�'�V���Ÿo&B���"ON�Y&�s��H�΄&��3�"O��1&��k���$rł�"O|��D�U�N��v&	�j^��t"O^�j�O�}�|��c	Yw�W�y")������@�O2.�v ��iQ��y�OJ��X�����p�I�Ɇ��y
� �5{Ah_99NA��_�E힐i7"O|$�26:>x�r��q�@1#"O���Ț�7^,= 1d�(-�r��V"O `h0䇢?R�T��J�.�) *O��J4�ǥE���0��j�8�B�'��0����%(�S &F,d�2Y�'(�H�b/�+9�Lq
 ��7VJ(��	�'!�@(���0�>�[� T~��)�'J@�9�
�l6�p����J
�'E
�k!`ۃaJ��� ���	�'u:�
1�RVSb�X��S�b	�'Jc�-��t7r�
�����\��'����͚!2Db����X�t"�'� �y-Ӏ8\I_Uu���yb*æG�Mj�p��8�y"�Y�eyj�7VU�K�y(C.�j4��P*C8�Z�h���y""^-@�4Q���>�����y�ȑ�<�ݱ6U <Pr��r�5�yB�
-KJA	��.�H�s�ď��yr�_tf	�����&�r�y��#�yB��A����p��*t'�	�����y�Â==V	q5��5j�r�C����yRG���P�B� R���Th��X��y����V��̣t�ŏB�4���-�yr��7 B�� �Ǘc,�17C���y�`p �`��$��JV�I���>�y�#Q�p�m���op�z��I0�y��sD ct��d�<u�G/���y2Ƒ	_"�pa'@\%�Th'B�9�y	T�\ "��DEfgJL �	��y�F̔j���@�ŲLH���yRgς.N��	�*>�,0��T��y�)M�W���j_�C���&CP:�y�cO�@0�(���1� �X�E^��yr��1�\�`a0S'��s�dÍ�yr�L�8���C�&�p��À�y��M9Up�D��T�9,�y 7���yRj�+nM3�M<5@�)�jǠ�y�@'0Rn�Iu�_az�Bp���yR@A6u��y���Y�J�Z���"�y�
�h��Q�TY��+�,�4�y���y���ï�D��v(���y�̓v4�2���4��]	�$��y�l|Z|�)B�/�>�*a��yRb	>nz��١K5%{ĕ�5�H�Py��-^��wMS�.<�"snA�<yw�gG�y{"�-<|�#h�}�<9�B�Lt��C�2[
�!"�S�<9�U�ƈ�uD�]i�K��Ue�<��'�5AP�9B�Ƀ�b�ꐂ�j�V�<�$�9j�4�!o�,f�HD@n]O�<q��&��q��<����'�V�<��Ö#�V����-
�x9ԉ�\�<a�j��%���{ O� 3��z�CZ�<ِ倠O��YZ(�f��𚖣�^�<�#[%ff����m�P�:���n�<��c��C�#�`يZ$dr��m�<���3T0zh���/o�` dI
c�<3���9�x��DN.""�D�A��x�<Y�'�b�`(qm��VW Sb�j�<�&�:V�,�[��ٯCn��wJ\_�<��h�c�� ,/�^<UB�X�<!��������Q*dL<�D$DQ�<� �5ɱEW�3����J��i1�"O�����VpU�K0v91�"O@��"�ӱ�ԑ�&~�,p!"O� �t�G2Jy"=2�CS 3"OB)k��(|ن3e�ѹZ52�"O���Q��P���҆��*��Xd"Ot�2�c��A*X��LZSԡar"Ol؂֯È
�z��$�T#g��D�4"O���#,A/��"�V�#�0�"O*UkԬb~���4nU�<�ڢ"O̍�$��:?8��Oh��4�"O�����n�Ј��j�-+��l#D������l�x��DI�hY�?D���g�ߊY6�d0��(�"�T�;D��:��PN^���.U�DQ��"?D��0�M?U$��
�
;aoZ8��!;D�L�̉<��Y�#i�4 �H+�N%D�P�Ԣ[9na��7Jr,�'>D��!��(E����Ў�u$fTҐ=D�,�6C��^��Š׉��/��p�>D�|�G (f�
Ӎ_CⲔ�1"=D��J�I�"_�(�S�O�~N��G�'D����+]3�Y@�EA�.&TUieF&D�`@��؊!vJ�A��_*��xI� #D��C J�`��EP�eK$WN9�6� D��Q���K�)	�ꉚ)aP���?D�8�"��KS������>U(A�3�)D��c�OJ3$D"��%d%%���a(D�$��W�Q���!se �y���8�2D�x�B�7�! QC޲�֍���*D��X� �t(CC(�6(�u��L)D�d�b�Q!e	b�@�	U�&���g'D�X��d>k�$��d��ȣ��0D���筀#<(%P$�P	63����.D�HP� �t�Z0�2��<��$�1�(D���3��13�.d:��)_���a�)D�@�#�7��EB�$�V�� �'=D��:#	u�>�ĂS�6F����	7D��ڐ���Q9����!�=i[̕[��"D������NPr|���ͭ|���B��&D�4Hu�{<踣�*��p�F�(�%"D��Y�$L���à�Z18:�B�,"D����Ƀ*S=�y��ł(�)�G>D�8��j0\ռi�5��HϮ�3f%;D�������
xM -1.�t�:D�<H�ƛ,Q��$ J0|
�Aǫ6D�\���-rh� �t��=OD�U��2D�����o$=�Q��a<F� �m6D����.G*[X2=�����Y�,be�9D���U���<PC���#��h���5D�<�q���lؾ��Ԣ�-ʬ��3D����(�+@�8�h�Z%h��zt 3D���3lQ�vo��%��m v��k+D�d[��ޔ;����T��
}>���tC*D���׏�'�z@Ѳ�PPn<�Rc&D��� ��D}�-�4h�FAX(q��"D�d����u���z�ͳW�L �g,D�P)5�
[�����m���Q�	.D������8��w�Ȩ��=��,D��4��*6N��T�۵K���e*D��KRm#X,^��3e�"<�<��'D�҆#[�r'��4��(���da8D�t�d�G�B��M��MҵF�ԤIU,7D��3���>"�X.P>"]�P�G*O� �����H����!�'[���@e"Oh<�"��=d<�ӧ��w��	R�"Ođ���0Q`r����W�yppq�"OJ䁖�Nu)��� chUW"O�I��S�vc�hiR	}:65+F"O�H��H�s�`[��z[�QY�"O)�1`�jTܙ�0
�>��mx�"O <�!��|�,ᗈ�[ָIJ�"O�9�gGӺ1'�-���
t�Ҡ"O�0��!A )�=㠬�-@��bf"Ob�렢����NV  <�� "OXu+ �J�i�����P�' ��Y'"O�� S˩w��y���2B@̀E"OrT/��L܋��?"��{�"O>����O?�uȗ˒q���#w"OyQf ����z0��?���	�"O�`��)Z�~}�g��?�|8"O�(HF�D���07`�aX��f"OVIP���8j
��2B���Iv"Od��ቜ���#�N]�1��EH""O�d��Z8����-@m�B	�P"O�W䅢/�$X"g�DcL�Q"O`Y��E I��Eۗ7�a��"O8��+S�WRؚ�X�O)d8ce"O�Xp���Q����C[h"a�0"OLԋW(�<KP���#����T�"O ��σ$c�n���K1;�fx�d"OdH{����<�����/E�&���u"O�� ".Y�2���P�eE>�n]k�"Ol��iRs(�؁e��CȪ�2�"O�p��(P���Hq�
[�m�^�S�"O���jB�<�=@��<|��E�v"OZ�җa�.J���jn�'k��U��"O��WE��QJg�Yo"��*"OtQ���>I��.}��E��M�<�K��H�Μ�DI�ܕH���E�<QS�:����c݄p7(�X7gLZ�<��*� ���C� �h<hB��z�<i�i$������94�p@pB�<a�ͅ,���(�M�[$�	R�G�f�<�j %d@:ũqhQ�t"<j��y�<Y�G92M&��@�?-~�y�KAZ�<Ѥ��S��4�����G���c�R@�<!�W�p}�Th�P����i�B~�<1�MQ�_O�	����>�D˲�O{�<QE��h~H,ѥ�/^f��S��z�<ip��'yS���hS.��tY�.Lz�<!w��"kx��p�1�}˖#_x�<9�F\�d�9�BȡZ��u�`�<C��	���B�C{	����x�<��IN@�ph�%� '�l��e�}�<Q��_l���PiZ�`�)�w�Ky�<1�mZ� �"1�n>q�b{�B
x�<ɳ���%j��2�=.�h��K�<��T�sq�0��aW�s���0�9T����٫~V���E7�̑ab$D�x���Ѿ�S�fH�}��qS
#D�`�g��a�PI���1�n��ua<D�d��Т�T��b��<�j��,D�I��M�ḧq�V��F�#�m+D�H���S�G>�}q�$5X�\t���*D� j�.ŰeE I����L�ӆ)D�p�f��;����
]eq�`(D��C_5�@��B�-u�� ���9D�� ~�R�JC8k��{�l Ob�H�"OF]0�*֢k��1(���l�4Ak�"Ot�z�x�I�j[
'�`�J"O(��pg��и��G�/�̓�"O�R�L	����#�0`�"O�P�bo�d�p�'�Ec��q2"O����Hn�z`f7`>��V"O��ӪW9<	�a�DU�*p���2"OB�馨@�P��M�4Ɍ�vi�f"O�Q!ƕ����G�$8 p"O�Hy )0#2Q��oV2-�T"O���H�nq�L*7��*4�D"OhPKY4O`�p�i�V N�9"O0��)zҪX@eT�m�B���"O,e�C�F�fz���@�2�VA{"On\��ē�b�+�aS�|(��"Ojd�R8E�d��W
E�
dRl�"O@
S�<D�h���)Xc��3�"OP�P"D �`���GQ��@"O��[�&�dc�sw�8R{�a1�"O�q�cn[/P>����5hIa0"O숢�]%ye����Д?���B"O���R��{b����S 2�� "O@��«�ˮ���±oJ.`D"ON���f�7F��*AM�*bEp��"ObTiC�	�=��(�m�5:��(�"O��A� �TSb����[�C*�D��"O���#���-@�廔n��5"=K�"OV,�"a�/4D��ٓmɰ$���$"OIH׏������,-���0"On��Z�x�
�-R�`��c"O��7��_=<�p������;�"OND �$Ֆ|$ڀkM*��"O\d�w��Q����"I[&%zjИ"OI�J���(0�ӈ
�p���g"O,���s,8��V,:�\�A"OL9@��0�By�1����.l�"O��qU	�p���
q�L�c�"O���nE�,%���Ӿg���X�"O�K�m�N`�!�ՆH;ƪ�ڕ"O0��q
� {-���'K�	�,��"O�찃�	Wmf �g*ڑl��!�"OJqϖb�r�j*�G���0"OPĉ�
0P��Däz��ؙ""O$��7�]E�q���:�luk2"O�0j��	�� ��\k0UP�"O�����њ5/ 0�@dۍs�X�f"O���d��.L�"CQ�}è0Q"O�2Ro�3)��h4�Ť�b�"O����J��a_B⵫PR�M+g"O\���I��UF��D3��˕"O\Y�碘�Gs�亡���:#:�X�"O���GB�!p�P��#��vs"O^i`�-�:�\�D@���Y"O��Հ�dZ�	�^-p�JG�s����6��̉"�L��x�q��tY�ȓS��9��V����1�gҋ`v��ȓf�l�K�.-�����c:0��&M�1	ҁ�1�G+�:ΆЄ�=���Рִ`�`\a�߳_����4ܨ�M�KiĐDGK]w\@��mr8�2�˸B����Á��ԅȓK	l�04�1*�T�y�Ļx�d�ȓ����6��_69B�%P5C	���S�? � x��2����O�ftX�R�"O�ɻȜ��*�f��"O*i;�����"e���4�(��"O\t��m�?��q�-�'�Q{"O�1P�,�:lŬ��TeܠoS<���"O�U�6,E�x���PFF<LZ�h@"O4��UJ�&A��U�fL32D4�a"O��ҒDP-�D�Aŋl����"O��	��ƨ8�jm��K\1x�윹�"Oh�8E	ϰG��#�ô��qrF"O�KE���A��I��T�
�ы�"ODP�r��.�y#��=�|�b"O�dQ�H�^����Śa���$"O֝$��p�0P�	?� Y��"O���2�ߞ$XT���
�eٔ\��"O,ݒ�AٸK��M�1�˺m�DqB"O~���Ա��{�
��h���"O�ȠWM;KVrmx��ċ���K�"O�zD,�9D�H�c��,B�!�� }"��Q�en��Di�70�!򄐡� I�@]�!��
?%o!��>�^P�P��%�����O�?aB!�Ĝ�Z�	��K6w~��-V(!�d˭aѮ|@D�ݬ	b�Q��^�il!�DL�WiV�i'g?�T�X#��'�!��ī/� ���jz�H8��P�+l!�D� �l9�H]��q1�<XT!�$�ȴe����.X���(y!�G�+��\�P������"d�!�V�*��\sb֞	�d�kPLt!��K]��Ԩ�`�'A�\3���7?!���)O��ǃ[�_�HiJ4k��N!�D
�2�"�����:�dA%^)!���$�6�;p��S+*��1$!�ă�oF��J�+�7;:ֹ��#Z�yR!��)�8���F;P��01�@#!�!�dX�=�h}�C�
�jH;�����!�$�U�j�+��L�0z���� �Q�!��˿:� <X!,�=��ݘt����!�V�E��|�W�	�Qvd�Ϟ*�!��c�~]I��_,hA�x�/�7�!���d��P�-��Y��m��y�!�$  w��c2��*"��}jVM9L�!�$��E? �!՞ ���5�� !��45��l�'dH���� �?
!�DL��>iHV��5��36�3'�!��V,¬{c�.xcΌBG'^�.�!�d-�fT�%K��z1
�x�ƀ�^�!�ċ�
A�C]3�@��Eƹ�!�d^,<���2&lh!a�U*-B8�� "ON=�G��`1Ĭ��ϐ!�Ny�4"O�-zÌ�'"�	!���a��Hр"O^�P7�̬My�L�g�)��"O�u���ޒe!f�($�аM�(���"O����x���N��mrr";D�lx���+�H�Q�N�V��#4�.D��sN՗v;�`Hr�R�dP��� �*D�x�u��\��q��*%2GF'D�xcG��R�;f��7q:jT�v�7D���u�:W$��R�M`��5�"6D�8 �[/����p�/�z��+3D���%g�W^�<�bM�T�z�J��.D����
�>WaF$S$��
�*�۱-0D�hsQ=!�4h�C ������.D�� �T�S!#'��JE�	�G~� ;�"O� s�i_ U≯B��Njy���"OJU0���l��8���,bl� "O� 0�m�	��;F.���z`��"O�E��dY�F2� �&NZ�*���c"OD��c�1��rr�%X"���"Ol�cB�0�����l��!�"O�) 0��,�2pk��_62�0���"O�(%V�3ZZ���B�!�����"O�p0n� qPP�1�R5J��q�"O�9S����)�LA�b+(=��"O��xF�ƀE�,8��K՞� jC"O����7:�T�'lY4��`p"O~���߅^7�,j���&�9�"O�œ"E
D�I�P0|k���"O�V�VP���D"t���:�B�e�<aa�G�w���뇍�!��XB�Ky�<i�aY�#;b���j�41�f�W�w�<��7IдAJ�N�3\�� �D!Jz�<��(�'/�d�B�v�^A�4#RM�<A��t�L�����n��5C�u�<!U��}:��F�:a�d��@k�<��J�����p"^�]�%���g�<�e ��/��4Z��']�IYpKFJ�<���2:�2�{���IK���!��H�<a���O��a�+��>OLtC�p�<��-ԵP@�Y�V._3�bA�p�o�<A�ꋐ�Z�����Eg(�cь�C�<��G�q,l�c�� �I;���f�<i��g�������5 ��_�<	���!<�ROވ=��b�L�u�<���E�����4!O^���zfGj�<qq�C���I�i�k�f��j�h�<�R��j8ȡ��H��`[qQo�<a7dڹ0_�Mi�,Y4r����u�<���@�8 ���	be���(�]�<�5cW L� ��+�:^^2`���b�<�q#U�|;�v�tW��ҹH�"O^ҕO�7w�	��ʭt�^���"O1�B�R��6�Ts�*y6"O�!�1D��\$cU�6i��d��"OB ����?ɸ\�e	�g�d��"O���b/*E�(P���HR0"O��q�"�L�DC"a���P!{�"O��
-�%b�<����ڸ��"O�`��Niv�uළ�2_t��S"O��3)R<Z%$���#d�go��|!��9Lyp��'�Ń)Y�p7,��;�!�diF�aCB"H�9��öd�!��U�j�\���GQT����B, �!��oǦ(2�M\��`�Ұj�T�!���r��с懙�\1��
Gi�$�!��ҍ�����KX�Er��_!�o�����k9�̑���!�dM)B�	YA	���͸S��7!��:uW(!��cV9XK�i�!�Ȇ�!�ѩI�ݡD!]�<K�k%ʏ>&4!���s�!�"� c�ɨEB�.{.!�$��+覠+�ŃpY"��b��!򤀫`5�䢣 �9g���bD����!��_#��$�rcD/dˠ��b��-�!�d�t�� K�&�8UcE$U5!��9<�����׏9�8���Q0!�$�>H�y���.ܒ�p�C�<� ���ϊ�t�f�ؕA�~�8%{2"O��ۓ&H�L־ͣ��=&�blp�"O���g�TD|<���שO��q�"O�ԫ��:J���J7	S�$�T"O������k����ˌ=�V4
"O*�#rC��'a����Ӟ��2"O�1����(}���Y
� �e"O����0 �T���k�,�9bg"OV|xC"FA2<4�U�J7����"O�D1w╏l¸ݢС�'{֪��v"O��*Ei\�#�$񲠎5N��l�T"O�q�'��,� l��IX���K"Oȥ�E� H\P)���9t�Z�8�"O�����/]����f��w^�2�"O `KJ���G%5au�$�y�kh���It�ʸD��+Q ��y2H�=�0Wf��93$���L%�yb�L�?�@و!o�.[R8Z�,�yrn 5I�h�Ƃ�G
���bb^��y�*��r<����0g.��bٚ�y"m�=��1��!~���s��>�y�I�U0Yz���|U��D̵�yR�S(g�JU��n�,y\ �y�._)uݬ ��]�&h�q�y����&����E�5���s�[��y���1>6��Hv�� -���6k:�y�gJ�7,`A2��6�f��
/�y���^�mY2Ĉ*{��DI�a�e�<q�/K�N4�YZ�-Zo�\p�ҎZ�<�u38��d��ޥ@Y� �c�|�<�T.�*_8"a�,�"�BLFp�<����-U3���V&�o  ���Vk�<A��ѫvfFL�c�V�l� �mV|�<9��G!°��%C�YJ�jR
w�<�E�3�蕒�iŷ
PZMRsK�<Imc�!�5&629��I�<��E�:/\�@P�4sޜ�Yi�C�<�&앧8�B83q��0C�x9ֆ�Y�<�gM�4An��5l��C��{rn�P�<�"FA�	�dݗI�8����Pq�<q� 5z�ʅ��ۛ"�*m��
D�<�� ����@T��?+6�l#� �X�<�An|�X���?k�@'�U�<���c��&�9N��A��Q�<fO��T� �J�7�6L�BfK�<�цE0C��Q�⃀�`���P�Hn�<1�F����`�e�9�rA��g�<qGo]�Z�z&FT$��3���<	"���2�0�Ё�тm����B�<�D�G>M���EFP�E*���m�~�<s�P0w�����Ӿ��ݻ�EP�<��/��>p� h�)��օ��&G�<�3H�<d�����Ғk�q��|�<�@LЛ1����	^�|P�,�B�<���  (\�y�oS�Y<����T�<sS�1
�@�D�	x�n-�&HFi�<� �$*P�s*�[^V��ʔc�<�7�µŨ�;�I�<?z�[u"�`�<��$�B�q�㗻P�<��V �P�<���+Q��Y�S��UՔ����AI�<��,��'w���
��)���_l�<��+;��<Ѣi�+M����CB�<OR �)��V&N�B�#�@�<�"!R;�b��E+Pk�x8��~�<� �q�f�ʠ2�`�Z����rC��Ӗ"O��Rf�^�X�~I����)�x"�"O�gp(� �J�P�4Y�"O��y��"�V,2 (Q�+���"�"O���@׀tY���ڔv��D�"O��مN@�d��b礙�{� ar�"O��8��C+Y���b��O�_(>�I�"Oܸ@7��4	�4ɋT"��"Vy:P"O&�#HH�[j�q{Ҧ�7p��w"Opx��M	J���2�c�3FԈ�"O:\n�M��!V�X���G"O��B㖻 �n=	Ta�8V~L�#�"OZ�j'���p�� �9S�ပ"O,�BW�p,
��eT��@6"OTāP�0�,�Q����,��"Ox]�RN�Co�1�&�\1Er��+�"O���lĪ\g�ЄL�EC�Ur�"O�aJ�nO*37LѠ#k�!nJB��"O~�.
*e*�a��lĞ3�ZE"O���W�łn�8@�$�ף]���"O����2�Ezd�UM��p"O�i�H�2�C�@<`ac"ORqQ�F�,/ä���Ǐf��"Ol� ��|�PQҦ
,!�N��s"O��{���r�l��7�"���f"O�\�DiY�jz����b÷g�Bk'"O� ����mF��"\��LH��"O�����OR�b�|�L\�"OZ�)�/��22��Νs��]�"O��#Ӭ��1��w�]*�T�ɵ"O���F�ԹK���֤S�3����"O�ٸwGPD]���%Lw�=P�"O���fK�;5(�3v��&kW�-�"OR�	�D�Ɩ=���\ H!�"O(U�ծ�.Nb�Гh�K��kU"O�h� �B֔��H�#X����"O`H� �צt+z�A�d��5� ��"OzBUN�Y�2	x�Wh�"�U"OP��a�J����dB��Ģ5"O�	1���)C�`��.<�z���"O��K�臓m�2�)���=Ҕ�`�"O�,�7.�7v_������`�P7"O^��ܸN���дj�4@��@go D��R�B�#-ql��3d/GR�V�)D���b�tr� �e�Z/��0g(D���R��v�3��!|R��gO:D���7�I�W)Ҭ8���*�n���D7D����Y L{�����JF1ɡ�4D�@16��{hb]Pb#Ǣ^!:i�
1D�����m3�-pb��ؕ�3�+D��Qejؾ)JB��$�Ĕ1�pd��6D��s��{ �t��'B�xj@�`c3D��q/ւ����AI�'�Pk5�#D�ċ�g_	�\=�#�@�>�F�Ѕ!D��y�_�p.��&#(x�:�4�>D�8���=F*��ӂOr~����)D�<�ѧ�"	xB~�B�(r�>C䉗�N(�mY�oBA�C�G9�2C�ɣ �\��%S�H`,9r��$�B�I`"����ʐ>v:�3���h��B�3i�T���Ԁ+�t4��LN,#k�B�ɛ�Դ�f�N =�J�"��L=xB��W9�Q��GO��pa�V;�lB�	�"���Yb+ �J���J	X�cVB�)� �RŪ� �@t�4I80��I2!"O��h�B�f� ������"O6���ĳ,�h�X���x���"O�Ai� \�2?6�����+�b8"O@�G�1�Y���S)��Ss"O�lѐ!ZV�\!�#�̟y	��"O����9"2:dHS���d���"O�h�+�#�-� L�#[�aW"On����#8�F��Q��:R�̹Q�"O����&��H��R�([?g8=:e"O�MI+�1�9c��WVN2��"OJ��������h�&?I��"O�@�n �\.D�0�@,DH�1s"O�]�#�چhJ\�@� L!OCF�cQ"O�5j�B�#�VaHf!G��ƙxR"O�ps�d�t�r��t���v�Ҽ�"OR`�ᨁ�H䒉��,}}��b�"O�Q�Q��$?
�����\E��#U"O������ }pG(ٕ}����"O�-{���&=B`RfᏰ8�F��b"O���-<C<10�L��R�R"O����iY=@�aB%�7ư�ӗ"O�1j�j��!1����b�҈{�"O�T��뜝0�;1��$��P�"O����a���1�D7+(lM��"O�93� 8^^�x��ס(j�{d"O��A1�(�
S��?����T"Oze�!͐-,�,�y�L��8R!R�"O��%֐CGn�4e��J�u�V"O@��!�^�D��P�_��X�a"ON�B"��
2�5�R��ݐ��"O���쎥ya�5aQ(�
�r� "O�x�f��4}
,�s��=g����`"OFaI��DD �2g�"�eQR"OZ-EH�.UU����R��c"O���!Lɸ( ��ff]��v��E"ON=�b�\�Y�jC|4 ��a"O �+��/�V��R
�9'z�!�"O2yg�'3i���§V�\�0e"O�@*7$B%1���,2uPJ"O����Su�t����lݘ�"OZ@�ܧ'4�Eᱤ��x|
���"O&L���"eB�\�d�i��PR"O�Q�Dh��B ��@OW*S���f"Od1#�K��
,y���L�03d�"Opq
���w�DJ�nN�Rv�Y�"Ox4�� ��EQ�A���R�g�6�"O��KFVp.`լ�/�̭J�"O,p�2f�&I��؀�M8���R"OT��(u^��	�3nz�3"O��BqB��sT~,"��	5�
t"Oj4�P-̋3�r�2�L#�� "O(E���Wy�>�P��ÖY�2�"O��D�V?]	(���.���+�"O0�hE�Cbn,��*VV)6]��"OI�ߏF����Y�H�&)	�"O��,�u��؁Μ�!����"O������b�1�5b
���
`"O�I3cL�G*�����CJ����"O	aҁS��%���X3f_�] �"Oe�#��-�l�"umE�xb @�"Ox�a$N�0���- �m���0"O$�ivJ��}�x��v���B�PQ"O$e{��E�������q��H�"O� P���J�0eA���%ײ|�&��p"O�р�,�34���'�	��-��"Oz������<K�Q�&W�S����"Oa�rj�?C��Fު,|�X��"O�tؠ-;F����e�$��|�V"O����(F�]gΈ�E��(a��]�%"O%03�^#�~%���R���"O�`�u�ՆMU�3��8*-���"OH�i���|�y���Ծ@�	"OHU�^1mN�-:�B����G"Om��D�%: @�Vb��XL�Yb"O��+�9x�Z�YO;:�	�"O�8��]�\�Dr���1 I��"O�=�un��R.I�a��	x 8Cc"O�a��.�zz���j�-�לx2�)��2Co\��@յ;S�Xؔ	�X"�B䉳Z6
����� \��L0&V5`�`B�,6�%xL͓g�Dy�Ψx JB�	:?"t-�c�����+KA�C��RB���?L#�P"a$��^�C�	�~����&G@��.�B�J��:D�H�.��
�
P`���@�)�<D����D�m������X2#%�tK(D�,A�N:��@ug�j�����;�ɲa�az�IF������ʘD��HS��]��yr��9?tp�2�R);�:�RF�ǽ_'�7�-�O�1Â�.jf<;��ղTOX*�'�Il��߅Y�	�0���f[P�!�d��i/�ܰBC�l�H�;�ɷ|�qO����R��_K@�r���%i����iա�e}�!��^f���A�ͦd�!��� 7����9}�lQ����!%�azr��§S5L �R�Un5�$N!OK�7�)�����!9���zݶ��S�5D�*B�g�����ޞY����5D��AS�_�<m�Q�te��_4���01D���d��le�"�i����ke�0D�8zw, �Y�@�(�&�Hڈ��B�+D��Jҋ��;�Lp�'J}�P�k�O)D�(����Kd9��ǧW
4�q i&�}���O<��c-ZF�����"xy�!	��Mc�{�̇Y�4𔨆�3 9J���=�yb���,s�i�0Ɣ?
�xTJ6GS�yD��2}�d��b+Tv��I@�.(
C≂O���c�OX Fo�J�,�$$��b������%�ӓH����`S�v>\!(�kì!˂��d�<��g��ԩ��%Q�J�;���@̓�M#ݴU/�O��_	�Qs�F�>fn�т)ٮahf�����Y©W(^���m���hɇȓu�H{�m����1�'�Y�:DxR�'����O|ӧ���ޓH�V��E枚17�0�"�
fn��Ɛ¶H�"�'�x��ݫ5Z!�κ&70q�ӏ��!x8���ŲiNa~�T��� ��BF�e�,ͬ����)?�����=95���V��2!-{��P؇k�t�<ɕ��$`dd��ceW�S�ޤK2l�t�<Q���ڬ ��R`�]3W��K��%��'�`��y�A�H�	�d��Z�C�Iچq�B s��=����\��B�Ɋ]���4j��u#t\:w�u��B��,1~�S�C9_�@�Q�o�.��6�/�D�<E��4PƲ�X4�Fv���E��MԬd�ȓ{�6�a���w�P�Ь�0/j]��#[���疲rCj��n�
I�Π��Iz��1}
� ,�A�咵l������W(ѷ"O��i"��f}�ɒ� *r�+cl&�S��yR����p��p�F�!+���,R�y򥇩,ƭ��en"�B�lҵ�M��4���&}���i)BH!d��Y��*'H��g58���'v�48U� C@��3"�2����'��hRV]/���a��3$,�����'�I��v��6�Q6���2�Ɔ�%�C�	$d)�d	ϣ:�h���t�4B�I29R�I��
[����I�}H�C�ɌO.$���"��|�� �5�Y�o��B�	q���g��|�thQ�-�>~�B�	s����"V�X߂EQC�
N5�B�I	c��ku+�>�he��D�.��ͥO�ӧ��<�H��4�ߍ'���Ӈ
U�~�����_h<4NF4~.�dq���{F���SV�<)��6 p��mU�]6�m���H�<���A}Y��A��M&H}s�&Ʀq�O�ӧ������o��5i�M��� �D9�yR��[^d cI"I	�U�cА�y"�cL����q��<3�Iѡ�y��)�'s�p���L�e;�KE��(����?A�J *C����"ѩ�2���#0�.���
�|��%L�jz�iQ��DUJy�ȓR�F��w��s� y�L��&�<u��y Ur@lD���D����p��?ɞ'�Q>E�'u��Ǫ�%T.R���)h����$�@Ph	��X��qĨ(���G|�����~�vg�.Q(6��c����Y��~�<ia�Z�Z�B=kĨH���i�#���&��5�5���n�gh@�b��݅�I{�	�Z��i"-�>NY��JL�Z�	A����S�ΞfE�e������ZB"0D��襢�5���l$4Q��1�	/D�8c�6�@q��:aI�`X&m�ܢ=�O��O��A��Vf0�@�:c�ܠ!%$4���Љ��)~��5ꃕ2�lU1AL�O�ON���E�-�蝆V��BAV6!��>lqz�cq�;]��8�-�d�!��2_P��FEFn��e�4m��D{ʟ�2�(=
� T��o�%g�vx`F"Or�q��ZD�Xc�πd�Zu!3O֣=E��k=�R{� G2ad�@�mO�y��O�=;`�h�b� "�	��yB���A��d �K�fHQ�tHS��HO@�=�O�����1S2�(p	ƴ8�(1*��;,O�˂f��
��NZ�����"O��a�%M�6�\��MH�Y�� ��"O:��3iO������+��=KR"OV ��ds�|js̚��51�"Ov`)��H����f�4
��QH'�'�)�>��)�:�Њ7@_Z!�IX�J�'��{M�7+JpJ�K;�A-���1 _��:����M����O�>��f%ζ(�I��Cӗ��<���5��2�HVfO�-+�R�|���v�Cpi��#���O2���[�V�F�㇃E/u,ɐ��8�ў0oڪ]��>e�PB��y�(pC���W�@�A�D�O^��$ū���c��ADD�4�$dE�c}8ȉ������4Ϡa��Lܛ9���hW�5Q��X�c-��B����Ќ6lJPQGk�%����'�4 �2��z�S�%-�d�Ѥ�c��p�c˜V~��l���y������|rO�,7��Шr���2����<a�@#=E��'F��b�`K�F�2a1�o��zm��'H�}�'��9&+2lxL��*m`r銚'��
� ���M+$�<�q%K<Q�p�q�"O0��4�G {R���V�-��$"O��A�aеq�����O�v|�̡��MX�P��Z�8E`9h��j�(�
�H7D��#K�52й@7e�quJ�e*D��٥,�>4���ā3`����H5⓫���$7h�`t �����2�'I�|�0�y	ǣ.4��K���I؜��I�i���F�S�Of�4�#`R�R����Hn��!�"O^:$�ٯ�&��m� {f`XQ�	@���I��@l�<�fi��3�ܒ��	<!��rQ"XrB�F!�V��u@�'e(�Ҧ��*v;����C��F��y��'�T�	��NG�<%�29��Y��'9Z�*�j�]���4#�%|f]�
�'@�"�4
�� �]�hk�'�Qۥ����x�# /X�
�')�����UG�["$�%���'�
�8@F> @i���	[6���'�q�Sܠ$�����R�����']~yj&��'���I���"# DH��'�
q���^�k��C�c��22:�@�'�"�`
U��
6M�Vg�E��'�Rd��M�eK�JL$R���'�����F3{��1Ҁo]�G�Vm@�'9*)�cHǈ;���p#Z�9�H�'B���dCJ�w?.���&ַ%�^�B�'HJ��#e��)��� $W��'�B���@�/ .b\��l,+��y	�'�@q�� �%!���W�W�
��TJ�'q�H# �͕K#*���c�#:[jŻ�'��p�M[7y
����,d�$P�':��i�
@d%"���[Pԥ��',jM[���~��U�Lh{Фb�'�Q���Ao�\�rŕ�1��ի�'�Ab�B�z�͒����*��X�'ht������,Ć�����5����'C�p*Ѯ�2���8!m��8rBU�
�')�`2@oM�d��s/��0��H��'��%`w(Mo�=q�!Z�z�R0�
�'�,��f���L4;�@?l�Ȭ�	�'���k�I��m�TxU�j�����'i�tH�)Կy(|H�G�m*���s8�q`�^Bb��
���>���n���87�Ԙ�� {$���6�Ňȓ6ۜ��u&K�/V✢TM:s�6���c�@����(&づY�`����͸"mA/Z?B$���9"�<�:E��Z�x}A�fؑ[�HB��/U�hj�EY�I�⤁�L�� B�I�N*xR��'6_����U0S�B�ɠgxNIJ�\�z��Q�vHІ��B�;�9z�`� ZY�U��Α�M߸B������j�2B�����	X<
�B�I���)��'Rv�pM�VC�	<`��H��+,Z��m�T�)k�C�)YUz}jpk%\�f��ь�j5�B�	��f��vD��t]|A�(���B䉡`܄3BC�P}��N~ɨB�\ǂL�R���B6�Xca�6,r�B��?�����߽[���C䆚$��C�I+XQ�5;��?@<Q��e��5�@C�I�c��{ugݖ	Y��C�V�
�PC�I:K���a�$H��(���@B䉉�BXsȕ�Ir ���׍!DB�)� �(�F�~uh����՘Q����"Oн��@�r$�<B@��5G�b�`%"O� �V�! t@Xr�U�C��k�"O�4�ǥR�C���H[nB�h�"O���`iQ*e�4��g�]d��w_��$�9�qOQ>]�DL�Y���)�\R��(D����iNw�l���óxZ!�0�'}BK�f��Z!LO��c��^R���ߔ)�8�ʶ�"�ONm��^J��1Sb��G�j|)VG
3q���e�̐2'������!|^Y�EO9d'�#>ў�x��H�T�z��΄ �O��ݨS��*7�4=xM�+����''r`L��-;�5�N��yB9�M�<��2�\!z��0�g`��"~�F�,��@�g�k�Z���l���y�H@��H��'M`�Ν"�E6� %��$	�X@��]+WV�]I�����SR%f��C��#@Q4���+�O�d���rA��Iq�A����M.l���iF�>P90T�:�OE��_ �
 �D��Q�Ĉ'�ɼ���;P��\�(Xr�ON��R� .P0*P/�=4���NU(&!��]�u��x�hV�
$
�PT��)����ՙ,��"�!E���Iz��M�\#}�1;=dl�aj��$|�ˇgG,]ɌE�ȓ~���M�D������.vn���M�0+�P�!�9l�T�:G��m��Ƃ���'�~�j�i�`�<$���P����-Q���`xӌ�JE�/x4r��>�:�Q-�V�T:��3xYP�K���g��x%�!\O�\c" ����!QE�D���:�[��S愅"�z��/1Җ(��� <!kF@`A�+u���C�� n���S�>l��8@#۞Pц��b�BCN�T�ơ��#�A��l�F� 1��+5ȝ	7֌	�+��r�##�����C6f���1�,Рӭ�&�����َ����'bl(�C�6"μphV��5��@�P�L7P��#,ʄa�y{&
J�H3���!ɰdHf�5��h�H>�n��m.59ᮉ#sfuK�H{�'�pI���S��$�vi(䜄r��┪Q�[d�Q��̪H��I�aF�"K������ք���D��Ҍ��8?Ab&��E}V �@(��zD�TFC�<Q��E1� Y��F&O`<�R"攝@wB(���Ӗ{�lp��&�, aH�YC��U���˗vH�T%�J�5�/� �*�Si�ϸ'mVDҲ�ɳ�dhG�ʓ@h�hT��,��(;(�p��iT�ƈDbLt�2i�2�pX��KE~�0���/̌X�T��-_&���E	2#\L��l�M�L̈́뉗R��K��0}>A�#lK�#w��z��ȿW���'S8̤�	gX(U,��+e�3{,q��� s��J�⩟��P�Ӊ��Yy&�
,!��9u���}[�|""=.�~�8Ae�>?�(]ѥ/˧�M����=�:���P8 4�ˁ�Ȯ.v0�c���M0����:\���z��u�����O ���S�B
&�x����vP����'G.@���N"�:�%�;x���4�@�@�9-t��;��V�"��*��M�5IUa^�D��R�)�?QS��R�����:��������Ǉ�#��hf�H �䨁
��l#��co�,a�i������6#��(��	�����
N�[.�\;�D�,��Y:�91���EBȷP�H���I90������c��+�% +.���,ЭVr�0@V/_�[�
�B�;��r%G�g��Sa��%���CLP-Vp� h6��L;�X31�P7e��e�P�N�£>ф#	�[UV@��]E
]�D|>���G?obx�V&X+��fiƽ���lb|%��Y�,��ᩕ���t��v&W l`�����Yl��x�B��E��1,�|��n��C �O�ia�F	6H�h�\x-&J�/cw���4K�h�\����+�!:Ǩݳ��86����W�~d!�Sڼy�6�{s �x�jq���9���G{���.�\z&���.r�*U�_�]��u�bn��e����g� RF�!�E�4-�DB��ڼ+y�"5d_1\��Q�b��VY��#A�4�"�cbND�~	��0EA\2a{�o���08�3X���d���v��@Ɂv�k���:o@,-I�m�/
�0G��L��&��p����r����@u�4h�E��'Ӛ��'+�]�;���.����`	�����"A�T�dN5;�$"�[3�2�IB��T�#�H�%��-��� G�@�A7>�S��E�MJ�f5z����4�	���l�<�#I:|��D�a�&Wh.X�7iO9����,M�A�e��H+¨y0��Sc̩��Q�8������[�PXv|q�ƀlc
��C�	��hO&p��H_�k�́�'�R�CUfy 5dC����fʝzA.�$EׅTH8D�!H^�o�Ե��$ӍG]tUh%d���,��U�Mz%�6C�L*)�e-�-ZU���7�O����B��1|�� �AH���
��'�e[Z�`���	&B�L�&ď��O��(CBg�
~��lAAN�g�¬�©l~v1��I3hdXX�!͵9��уE3�{êX�K(	 F�#?Tq�C:7��y���O��!�J"�ȕ�̂&	 �(@3�Ў����17r�A�,��&�ru�u#�$h�1Ovy�#T�m�z)+����F�<A-�5\:Hy�'�R��%-�Z���E�
�jL�����:_�&��U Z[��<�d�=�F���	�b��8s$B3m��d@��͊J�`��6M0�6(K�V҈��g��P�dC1i��DUgL�M���x޴�L����`���Ȓn�	#rTRaNխ~�<�-�ҥ�Q�H�[�6Z@�KQn��b�������.!���h��++�̙�I�t�a*¯P[�cf@C1D����!04��Sc��1�`	,�9a!� zx����a�H
�X�57��F'h M֐>	�H�K�V¦�@�M�J!��G�S���I<�й��N�}.��֦F��t{c� 
�d���N�:q2��Iߵ3<=ȠG}�Q�U�a ��b��� ːQ�^-4�x�bZ(�\�A�2aq��b3ړus���G�-&���a��O��@w��3|~�r�i_�r�f��oK�qy��hC�V/"���	'�� I��&N�0�*���� �r1�RD�+tg�d`a��+L�0R�'�Z�#�FËZ�Ze��dW(=�&���	N�J�bI1�=Dh��cl=��T�$	�7�ZQ�C�V���䓧X�Rd��N\�z5rF
��O�*�����Zc�е�I��>�B�,T%!��Y !�J�o�Ό�K�/G�Fu# �Z��i!�gE=y���D�F����1,�����@¡����� �6F-��,�|<4�0+���?����<�E��MGw�)���=�`<Q�Û��]P$��q�@���ƒ?�]�p�A|�i7�վ
�~ � ʆ"
��a��F>c�����۞
�x`Qr�K�0v�c��m����*��hOl��0K�}��}p���c(�؂��������^q��1If��MC����9� �Ӱ.Q�'�@���ta�%(�w��K�.ӛw<���]�`�HA�}�'�6�Q�c��e�Dt���V���y��2�,��^�q�F��2E��;�d�A��u��qbw�B���z5��*m�YSF��{�����U6�P�+o�p�W  ��3�5@��ʁDe�cX,yh�Q`C �$�񭋙\)ȉ�"l�q ��B-1Ѧ��U�ݫ,��I��|�"旋q��(�!��"�t���6,`|�3wE�-@eN���<�F�R���p_ �j�F��Ed�s!��3"�'%A-@dJ�(�V��L���:v^8���uf^��?r��5-��)f���#z�<�s�P�Z�����	skD9�?��	��%�X�[��
s*�I{���~��)l��b�ܸh7�6cVh���L� �V�[f��S1��-0R�	2�F$|�b��d��Dq1��X&O|d��)�,L�uEy�d��P]Y`&�#Gr���KQ��kT䔡V�H��T$��z���a�H�FFBR���II|���/�;�ĕ�S�Z���-{��j����v�lj�,|��`��3uʱO0T��L�0V��ؠG��I���k�l�'^��%;�'/��	5�ɨn����uG��}�}A �ۘV)����i9[�4*`'ۗ'��%�I(o����%��!z�U�;A�	�&T�LZ����-���y14��<kV}�$勜
�F�	0��B��K|�`S�/�$�#�JS+HtZб���!� @���Ml� ��T�?��!BH�6y��X���S)M@��3�1��5��p5��8������c�i3�W�&��s�M�\׎X[6`����`%(��ܑ��	7a�y+�+�Cm�d���K�������Q\hit��H��d(�(O����&�RRpAF�&ذ1��	� #������^�B�d>�$)��	�j�.�2 �D>%Ӥ	V�$+������-�T�Zw	����� )֎�RN�O� 	��$�� eH�a�BX�-k�$(�z
0F5�T��a&M�R��Uf%��m�|��C�o�x�ޤe[~�';Ĩ��'Jæ�&P�wx�����4(a�!�e"��V.�@�f�:I�2�ۂ[%�eJ�b_qf�aA�*e�5�5�ߧT-��'0Uò�ڴ9Nur��ët[����D�q]�P��ԧp
>�j�%�.I�p(W%�7?X]2�`C*��'��=!�g��p�v���^�:�"�,�&r�+7��N�����#��a��1	�g@:v�l)���8�
V��� Ŏ�*�����\0:W���B,X����@�+̈́2RazlVq;B���[>�bѰ��%-qz�"��ĚLתِ���� T��W撚P��i0�ܚQ�1�����˜Ϻ���9�����޺H%>��v#�q��t�j)vEu�|٧#�?q�\Lw�G�g_B�R��|����G�"l_h<B&��MS����M��H�����e�N�=2��>��e�aHX�Y_�q�Ġ��-�$�"('����I�a&d�R l9��i��� 6	g 8D��`͐-D�:�)O`���'�M�q�Sy{j��AL,f��]R$�.(M��'�u�\�@h&M���}|`�<���
xu@h�6��1O�6E�$Ǉh1V�ȧ�E�iZD �4/R�zEfT���ċxvD\���D3L�:E�g$f�p�8��I8)��eӯt
�����@� ����bAJ� _�� �i;�l��6 � ZD�U��.s�c���e���s�'qٔ�j� A>b@fl 8��d2�y�8�_w �F�M�^|6��	4���W��;E�ʌ�����O>9�H7)*��ZG�7~��Qq���!6i�\�"O�tg�\�GC�;� �P/�6*~ȳ�
=8L�l�Ц�[�&�x\Pq��q��I8n\�畟�y����$��T
]����n���=���H���I���I�b�90.�2����J�]��¤��M�D���R2��8j��a�M��0�(err���,v���'܂�C��-�(�Ґ�&`��ʂ��=6Xl:K��@�Q�*d��[�@'�o��
S<���O�Y��s�$�0e�m��aS-N���@�Ο��<!���8:J5qQ�=��`b���a�` �Q�^�n�$��B��(�F!'�]�A�;/]X��O���6O�!!���~6-¶'X^qI����o}#W�_�H����F��x��!ڑ/���{���5����X�,��i����4�ާ_^U
'�>7K�8bg�^O��uJ�i��t���A�X�ӳ)�����D�Nxb���'9�qS�Ǌ;Ω�����z�f�&˓1.n�����;hl�t���Wm3�(I�9ƽ��N4y�l1���2�ȍ�񈟱_�!�$�M�t4��	fn;��S��H��Hq7#�b�ҹۉ��0�𕱃��)� ���� iR1K�i�;y���L#ܴLsp�T00��ѳG����!mK4aDcI�!,�����T�$�!���6�Br�8M�NMA���T&�i��+�8�bB�9!���#&a0%���[(���`�H7�%!�F ���Q*_($�����%e2-�;l�t��WJ��|gbIJU�E$$����(}`z�@��x�kʖS����f@�J�ⱐ�`[��\qu��bغ�
��R���XTb�N1�ϟ;�(�HUk��!h^EQ�핐���� 	��V���8�F��`�H!�aϞ9�8�xݴf���%+�0���ȟ�vYF(Rv.Y��P�1�ءx��!# `�ݚuK��:�=�7�3wYN<rFA\.j�>	�%#=�!�#��-Z'�q�&�`\�<B�C�#;9����ۅi�0!�E+�	�G����C&3o���R�3��F��{.8l:��(.v�x��k��7��$5m���" 0�ܙv@�{)x `+�'�����7v�h5K�ƒ��91��J�'Ҙq %I�(���;7Y3n1�,���ܽK���B. ��n�&�5X��ѫ�@θ.�������o6h����IW�LX9y���.U��utEG(? ��cŬ�r�;A'AW~"Ƈ�Z#��p��� *������ qet��5[�v/�8�B�
�/���� ��^�5��:Aְ�H� �<�p��	V莈;�!+	�����N�[�uNI;EƐ����!�� �lI`��x��%a#*�t�Q� ��|�G)7��)AG_# �ta ��0x��5Isʛ�w�)!" 
� ���iF��1���A�G�6hV�R��Y�g�& "�ʈ�a�b1S���9���"��'��S�e��_ʈ�ВK
x�XaP��ٌ)�(8���I0�����2̇]
p�c$J��@��HA.i:��ʔl�(�s��;#@\�Ë�I��ɹ1�"�I�a�����a�{+� abZ�^f ��)9����#T^������`EF��`�j�ѴG��}c�
�\bi�	F��u
zݙԮ�{Mz�R�	�j�����$j�I�+\��'L"��I�T��� U�V�A�BRJ�D` �}�{�k�%2�R!(�㐠H�`'2��U2CoP0)�d��4�Y7E,u���E �E���&��cPI1G����c��l�Iñ9�Lzs�Q�pm4�&�Nt�'7�%[�G��?�cG�M!�H�y�4�D/^�b�֑kv&�L!>��G	��D���]�dd�(�?��U+&�����Hp.@Y�����ia5"��i첵ۄBd=��#�l�S((�ΧKs4p�C�= ��I!�g�r�EF\�s�U����Z��Y���[g�aGxr�̸n�>�˶��26���L�-�� �Țr�T�PC�$[�T�B��1d��mXǨ3�4i�%A�/��;��p�R�HcN��|�;fE$�C�k�h� �;Eq�&��9���r���u�&~-&TG����1qB��k�$�4�p�y��-H(7DK�WD�AS��`���O@��SdZ�2�j���>�GG\ r�<Yr�[�O'Q ���{�)r��B'����Ѕ@�E�|�DBP�Dv�i��',k��Qs"J@�Г�O�`@K��haތ���R�Q2�(���{�@��(��dK�E۱c3�HRQ \[�ƭ��δ!V�v#�$�5��h�)����H+
�C@+Q8YDErV�ѕg&��C��c7�hA��'$��sr��g?�tq�+��U1BE��B�)���	B�kT iѤ[-`�"(�W�^ U�F�~�	=h�����4k,���I�1^2��O�	Ö�@�]5����fX�H��P�^h\����,A)�M�m��T���A\�hpp*�!�@��۟ўt���A�W�.���a8�R���)^�Z���xyb
�
��O�b��s>�j�+7�Nи֍�^����V���fŅ�ɬBۢ�2��ʘ{E�U c��|�^�"�mʩˮ��wD�<qː6����,�w��q�Ta�n�U�|��'�t�AE,�w}���u7x��E#4�`��I?�~����-����|���H+"h��d�	4s_�s�P �!��XK�9�<,�|,��C`�!�d�V+и��[*{,�hFi	8@�!�D�,4A��n��� �B�O�L�!�Вy�m�*��L����^�N�!�Q2
���.�H�������2�!򤒾T�����r)y���M�!�� U��	@�&B:�Ĺ�RN�T�!�ov������~�еj�E�d�!���=�22�J'vj��Ӎ�>�!���NQ� �2�Ǐ[o�6l 7Kq!�Ȟw=��b�2|ob<����0d�!�D�-/�P���D��PGn�9z!�d�rP�=��ś=X���R�$b!�$�=&�n�a�4@r��<.��
�'r�rǯ��&�F�HѪ�?���	�'�p��E�a@�ŨeM�1�.Ɂ�'����P!ݔ2K�$j%���)��[	�'�@:W���� ���	[��9��'�8�Q�K�+��Ƞ�"��c�l��'�\�i�&\�I��t1���e��T�'�"���fK�[�2��a��f��"O�|2ϖ�}�=�gi@-����"O�0;�)��n��\۠葮m:`��R"O,�*��V� H�s�&��//�9��"O1r",>\� �[�FA�3B��2"O��⋱2��R�L7�Xi�"O~�k�R�-���1�"«y��9�"O���v��6��$�#�[%@�<q�A"O������؃����E��"O��aQ�Wj���#�[�~��t[�"O�����&U���%n��r`^0*p"OJ8h6�� �ण��Ҕg(XJ6"O�s kV	��Y��g��QG: �u"O����a��\b�� �8�t��6*O�����c��Œ�	ǀE��()�'ȴ�C�ێ.�t�8q��aY�;�' ��쁒2y����.A3[� ���� �Q��&�=N�Bh���R�.B�"Oj��5jO3>�T�aՏ�0.�v|��"OB�2j�JL6y�U�KVw���"OL�)fH �U9��b,�?zi> �B"O�G=^���u�>��y�"O�r�	#t�J  G?D�8�W"O���'�2��ZfO^&6L�w"O�53�X2{��\�RȎ.pֽ9t"O8	s��<�I�!��D�:)��]����G�qOQ>�)�%� Sٌ�W��
���GB7D��`R��]\n��$N�D�ڀ#� }�	����@A�Ԉ ���g�0�b�>Oi����e"�O���r�j�^pm_L(j�� n��4
,)B���	b&�0&�K /)B��%^�[��=Q �~'��r`Kb��"���I��	���3�9Jx
t"O�{�h%+K��VH#q���'��A�¤I�h��,"� _N?E��h�rhX|d�P� ����L!�DE	0��cP��q��E�R�Ƅi�\�����D!��܆*�~l��]?#=��b+7�\�`�S�l[5A�NX�t�檂�H�8�Qe����Ĝ�gH��A6��)%K�` F�j���C��ð7��Pa`D�#9�<2��'ғ?νd��PD�pRLQ��� QM�D˕�	<;�L9#b8G6B�	6���Sqؒ ��`��	�#j�6m�6w-�(;��jX$Rt-n0aG�\c��6-�5(���ϬP�z@@�"O�q� /	��Xك�޾\������7	��Qj<l��٣e�M-��S�S��c� I-(1!D��T�H%64
���<Oƀ o��M�a��%4��׿(!T
���x:Z�H�/�*�h��r� "�i���	�p=��e�0Q����D�b���2C,�tybꆓH<��J"�L1l�da���-�~��~1�f�7k����! ���7�N���͙��<�y�j>@m��-����[��;N��e���|�
\�j޺%o:��dj�=Ha�_w[X����IM�0�];��p��Ɛ� �(0��
�A���DP�G��Z����Εb��֪
J�����;;F(Ν��j��pdY<'2��<XG�T\�X}0J>1%��d�a�-��w*�Y��)@Y�'p,�Q0��Ӓ�J��k��Q�'ßD q�-K.n®�R�ӭ@�Z�+���SզȂ��*Pt0��y���*Qv2��'���KR����m��	H�J��	��'4n	H 蜴y��@�$��1k�������u�WI�4L��%�6��<%,~�!!i�&�Ĭ3.��z�
����7}rlܠX�N���%��d��X������X�^�`1�\���ѡꏺy��y��L�_���G�۟^�켛竘X�<0��?z��١uj;SIA�_�V�hY����=�5�s���p=yp�O+G�h��`G� ׍��?[��Q��#=��Y���w�֔��e[�Gx$�C@YA���(?]����������#d�FQۇ�R~��q� �>[�\1$���m�H�3jϕ5N �E��ֺIH˄�.�{ �AZ.%�P� �^��bMQ��z� ��B?�ŢU�h���W�`�T��3���wE����=�gH
*�yN^�}_0��)!~���*w\>Y0D�%z��1�ʝ���6�1w��"w�\���t�1ͅ�c'���*sS�Y��O˅�L��O���2�=
@�O��J�)s%�X�+�|����~��T Q��1V#���B/�	?
D�Wo��A�	բ�9,�h\@%��qW�I��!�=I�l0 QK92Ge=<O�d8`��UAm*F(���\Eǹi7�H8% %e����WO�!Rr��F�H�S IJ���>x��hP�E8k4�L(�Q$f�jsƘEZ��$14�����I�ve�u$��2tf\
cc�8O[��. M��bF��6M���W� &����$�)fv�U�4Z�}h���ڮ OƑJ'ڷO���@@��k�iט�A7b_�@��eA���U
F5��'�~	�u�˛gXܹr �I4jOި��O㶬a�����\��M;3�u;�� )XΤ	A'Y�;Ov��0c\�1��b�E��~�q�#;4�i����b��ظ��PYSfAyբ�'9z�QV��y[͑��T,,q�c��f��Ȉ��Q�]YpMa�b&9y�iJֈH��̦�ZL��o �60�f	6k��p�a�%lO�$�Vm�`��0�r��,jȡ����# M�HYʋ,��̢�&]9s�R�DI`�� ���O.g֑���Z#I�T��
�p���ɗ��>!���K�=����+<��X�b-e��Ц�ܧ3s�acU��E�|�p*ŨQ=4D��X5Vh�04�?	�H����ds�uS�Ɛ@�j�����*U7"tS&�'�
��G-ǎZڞq8��J�4���y�H�$�ɵ鑭z�x����Y y����R�\�ݺ�#�4j�^�[�H�}$^<*��E=mӦ�T=V��(�Ǣ!DQDH�P���l�ў��6M�=�U�G�T�� ��[8jْو3�^':u��P�箙���9�e����Q���X0�[�kߞ%��)V�x6*]�3 t.��[EϏ��vų7�REx����LzZd���p`�D{��N��`��G��sL�Y��	6SW��D�-�+/s�X�u�H�Rxz�z�L�.4��$!A�:_�az+W�Af��H����bNT��#�Fw��y2�h
8|�,'���]�|�7i&1��X� ��
vF�O�$�1��8[���``,�?�� �{f*���B��o����
Q̓n���ujN�V��B�+~�6)]3_���(j��@Ѐ����B׉"2���V�ζ�����.q������*o��dG{
� r�!������@�_�.��X')"٠�x��Ow��K��Kr�j)��mڏ	�����޿#���)��ň����Q��ݢ/�=N��Ja��bL�#�/_mx�d@�%�~�T���i��s��a;D$1R\��Ŭ���)�K�5EGU8�@E��W8n�� f5b耇�,g��2$l 0a'tI��Ɇ~� [�L�YU�<�% N�Y��q�p��0��AZ���(��oZ�F�'&��	��7K�X+�FֻM!���3�ݟ�8Q-�k�q��K��2ȫ�:��s���s-�i�nTp��J>XQ�pA�:�V��jk,��Đ�*@� J3���7���F��,C���$"0	(�2�o�o:�=A�Ά�'�FP0�nI&<��S6��E�f\Q�D"�p�ӎ��c���TN� �^|x�.H�:��3�i����b�Z�eD�ө� G����V��Bڸ� цD�0�ax"m6{v��D�
���T�/���բ	,P�pt�p�,K��ɲ�/3\)��U,G7�ŢL�4��
h �eɘ�g�bx�%ЫR�B [5���O��ylҰU����6+!U���h�
ؙ�([��}}��S%
�@��4+�'P�H�4\KWllӮ\�4�ߘef�2ڴ��!c#-��{c,��EL21�Э�O�a( ��*H�����N�z'���؆ �"����i��@�Q,<̂m8��J��0�+��.�CYʢ�r%U?(��[�		�`
��iX���1�2t�*Ip�c@�J�jeХ�h�'t�QDՠL�ۿs��!��Gru@p(�Mˇ;��Kǩ_⦁���O�	-�}��G�z�6�kT��8���2n���3l���uZà �*� ��+�1�nt��lݥ0���Q����9䎚7�.��+v��11N�B�)	s�ӏ9S�r�N����9�.[�1�"���%A�r��qA�+c�̬ѷ�C�2|�I�R�5�O��tg�����b#F^�
���	�f�Lw� p���/v�$����؁v�RQˤ�x-u#0I�-n�[��=}���_��q,@9N��U�֌B�m4��E�L�0ލ#�"�V��	����%�񁀣� X}8u)�?�0h�q�Q5؅#�bԅT����
$���� \�"|Bᗑu,He�T
�� 5���C�p`1	g�U�L�ʬ��AS�_�6P*�AVS�x��y�'Nqs�!:��M�I�I�ߕ6{�@a�'�D#�4���&{��UiC'ty�=:�b͠I�]�w1�V�ð�\�V_����X7�f j��:�܅S����(O����ٜ2�|423�E�8�\1�aɖ�Ը!WL��v���C�v�(0/�q�tA���N9�Z��V��Ȝa�ׄ{p���s�TPB� e��P��RcI��m�<1�>�R�[)K�T}h1B�+7�d���L'(����(��xH�� }$���O#N
�B0�`Ͻi8�ɀ*�<x�*��h����6#���j���(�<� d�;2^q�&N�t���隺�� 0p�h����lλ;�������7Vy�N|Z�a�� l����v;�D���U4_�P��(:n�c�#ɖ_7Je�q�ͧw�-�rC�s0�p�E�4�	'.V$�(��IU^���}��@���B��D���優R?X�׬	�.T&�8
��\�r5㔜ŖP��e��<��]�Ϗ��q&�&=�3*����� q�9�(O�1��'%:�Cj^�� 25�_�nR�@�q"ՠh�5C!�ӣV6�ˆE�6�%i�1�����	��Qӂ�[�Qxcϙʺk`k�"/�Y�7�SCEI�e@�z�'��r�`��GT��D�Ϥ(��(��K@(tjAH��=?z}9���:�x�
J?�$$�sCW�Q:����>9��?}Cw�R+TٺÑ� {B}�e��Sf�)�C�2 ll$��?[P�o�5�`@p�F�i��Җ����� PcL��|�&���kw��
�\!+�^���D	AD HYt����w(�+>� ␐U�A��ٙu���BQ�#�I�j�R4Ȃ�
H�^��K�IZ0���.D/��̨dM�>#��=���S�k�X(�"k�N�B�[�+�H^:��6��s�\ɓ�<VNtA��	&
����@�ϗ8���Sŀ�W��D����&w�(��T�EO��`e���bVTuJG�S<5V\24䛏T5��!v�i�j}nU�9�Fct}�AA����ܚ#�һv���S�%�ԛ��d��{Q����'� �a�ѓ;F"T�J�^y0��	�K~�h�7SЄY��k� ��R��Od��V�˙7�DI��?-��kFm&��Qs��6;,� O���|㵃�i�`��_��xQ����9:a-� g`��B*���fK!�*(̧U'6��H�d��D�x4��!K̳[u���>H���'c�ղ�NȦ}:�EFy��R;	�ux�kY�4�h��)n�4�� �@�ty�e��������
�}$��\�8�h�
�럸��lK�u��) 0b	Tzx�x@��'�M#�Δ7D"=! �V|v�@ +��`ʴJ���T2d��q�Y�D��� N�#d�$	��ש��q(DN���j�+����X�A������g��hF�!f  Q�m��H%T�GC���I&\��C�m�h,9RF@�$ޚ)��"�|>ֽ�F�'|�(�TH�oAb�˃�́&g,q�G��H��9�I<=L� (���Xw���I�2��r5FP�w|��2�RZّE�1�L�9T�]B��T��D�X��k��ԛD������4DR��Ilӆ �6dC�g`Ja�& �qy�*��kJ&HSF�Q�XK��2b�*�()�=!��IPC���B�t(+�-
C���sbH�6cToF0d�,� �X��ThC@����ٓ0�������k9F�yd"ђ�ay�A�t�f��#h�� )c�bF4$�δYw���g�`�ׇ�u��X{��w�iJ��I7|x�U(Gﭟ��'�S�0F�իC�C�yj�5m`]���լH_P=+7��#P`�O��R&n��A�ވ���
�:��e1s�
�c��:��L-Ǵ�k��dc�����$*�|�û ��qI6����M����H��U��ݺ,�����KS���ɻ>7OI6Y/t�0�hR(fS0a.N묡�w�Z��bXt�Բ-�"	��Z:}B��R�k� F�H%����D಑�D��i�y�%"�_c���]&g���`f�Y%8=�]"�P��S2~�q ��I�l�6����J���)�$u�G�¡[�ʄ���A�=�xEZ7)�|�><�5�L8J��I�t�����I�!X��y�̕�q�Hic �dP�@7�5i�T��	�q�B)�`PaY��hw�]�j�Xa!阔7p��l��\y�E9�H����[?x�3��Zw�yI$H���Q	�A�uW�W�h[�%D2f"����Η6��a[��ґ.�OD)��FW�'U�A	��ăy�Ĺr�U�kfbeR�g�B8���s�r�2�i�cPP�&�B�q�~L@�
/c�|Kvĥi2�8n�u�j�
�)Ƴa^pڦ�Cr�F	�!��Y�r�MD�L�t����<!2J��(���yĭE�G�:��a��%��U��L�C�P�@D��?�4)�c��tĺ-��ؿ3���D0��SWl{	x",� f(���I�d��9��}��@ʳY��H4���vXZ�[3�K>�4����D��!'%�6��[�O�_��xD��uZF�K`>�� �t8C���G��d9FKI�2ca� ��5�]9�͏�'���G�3_@�YC��`q(�QAG#z���bl�_��c��kp8�a狻+�L)��!�8go�0ɮ��a	�J-
L�={3G	�2�xe��>9\�mbWmGވJF�x~��V='Ҝ�IU��t� ��7��O�d�"��U�8�3���-|�$E�Eo|?`U)�Y�<��U3�O�$[�:Ĩg#��4�U�cI_�t�.Q�5��:dY1�Ù�8��us���%X|� ��S7�!��AG:����G���)U���yx(���Zm{� �銜S5�5�ׁG�;����G[�F�(E0Ŭ	� ���ꔩ18�p�ŋ�T���� AA+n�T�rS�J4[�<mxELIIܓZ�<�#�;{���9��ɰd'�ъ��X�z7���7���Fl� SF�-H�-�wc9���!&�2a.���T�Y�?��� �	:�`���M�� �"ҍ]�м��؆�����i��$X��m�:TH���-��ݩ��Q*S0�!�WG�6z�څl�79Q��
�?"��d�ƿ6RH�t-�1�@����<9����^wX8i���s|��3�K�&FqrpeLp~���E ��$�K�e��D�4.�ﺓ�eƓ�<1�"֟�צA�\�� �ʛ#�lM"𩐙rk��!E� 1��)�h֦���;kvdqG.e���)��K����	�X��*bJ�qXE 0�!C���u�+!��<�}"G��[S��ӯ���BN��S�6pYTIы.��Z p���ze.��@��@���,������8^�pP����!�����oV"�&D���M�&u@��Z>�b%R!ςY�vL��O�����#�6d�UG�"��CV��}@6���f�)Q�8�o��f��ҏ�ֱB��L�'O;^�\Ib�_a�d5��ȀZ�|��ٙbE.�Q+	%�<�P�����a�ҋ�n-���H^�p	��Y���wPzA��	�s�0��/3�L<YQ`,Tp�[�h�-q4 ���r:��T�L��:��$.�$f�
�CްM�Јh�oR,H�`��6���$��	� ͒�NAf}R�T�-�paɩuv|���ˊ8)o^��R������	<���ۊ�t�W?������OP��͏L>N�Ro�>�X�P%!S��4�ģ��T�p ��5Oꐂ�`�=��<���W�qjՙ�� 
h�+P/N�n�r�;��Q9�H�@����i�#:s��d�A�-H�XE��.î��V��m�b��ϓ/�������i�l����d���J�-�1c�����̘�l�@��V�,eݾsvO�Ü��FlT�jUQ?��E&m� 8�d�<(�����X���'����̘|�Rp�N�S�O�*`�e��'̬���;[<�A趎�O|��0bLJ'Р��#��������t���D�E��h��3�JM�A.L��N�sr��~bĠ�0���2<�б���ؽrj|�R'�T���1۳/=�O=�v���~���3D�!F��Q����l����']?8B�ɲG���F�T��!�` ���+"d�i�`���=)R&��g��h�f- ��Zۘ��`���7��a��Un����̈́��S�OM�
��	9~� E���w%���'��%3 NL�1������k��MR�'%Z��&��к���K�`�jP��'d�4(�(T�j �b�؀[���3�'�
���l����	��«{�hb�'D4`X�꙱}4M��p�Н��'�>��%���SN��P@
;r�t�K�'?>�Y��N�_�������s�� �'~P��M	�rZ��P�r�@k
�'▭8�ǔ�=��P�����-B	�'	�WF�:���դK>B`�*u�%D���G�H�NT �`ږ1��Y�u�!D�X� ,�M��=��C��-�yj�A=D�(31iƛ]�R�1�� ��ӆH$D��yC��W��]AD�����J#"D�и6��S��J�M$x�����&D�`��"Β��4Q�fU[�H�de)D�D�A��6AP���Ϫ[q���F'D�(�dˇ*�A  �5F�$ta�l"D�|���/;!N� Ԍ�����E:D��a�f�0;�%�r�Kk|�0x7<D���mJ�`TxI�KI�x�U�'D�xbd'1GWʜ�`�ҩ}�r #��"D�d��Ú6@6 ���׌1X��x��!D� i�o
v����u���ufB�# �>LOr�B���4.�-x��zl3��1�^Ĩ�l� �r��$��V�2="vNE %cQ>%RiAZ�}x@���:��sE���	�7�p����Z>�
D��+�r-��Cө��堣-�<���V�M�4��v~��i��G�xtpbK�z�0��B��ɭM_�ū�4A��R'�c�OҒW�0��P���ۿ��0���O�+�OME}r�	ma��͜?N�5�#W�5'n ���������T��1ac`��$?��|ڒ��4eP 8��"�
Q� N�$�����yReC�=�a��JQ��m��/е!����eL��y���<r`�^�)�AVA*Qh�<5(r�H`M�d5ln��<��&��S�π z�0�eTr��L�y�8O��PV7}"�1�'F��O	�O�*�!gL (��YJ�k�����>� *�Oa�4i� A
�iE��NY��Tֿ�� �V���%��yZ����O�ɟ�|���
r:�P@"¤$��Ex}��'$7��!��)�'G0�ش��\�~4����!0<%o�ß�s�4�`<��ܴ\籟�a�4�S�Ǣ��\#�P11O>3aJa�S�O�F-�q+�9�U��
�%
ɰ�Z�L��`b�"~b�'P(`�DW7c�����L*���dŰ�0|Q�F����^�z 
��k�Ve��x���Jk��|�'�V��Q�N��
D8Tn
�{j�,�M��`�<�S����La��NL(�u-ТRBP;�'IB���y��霺ZJ,�z���q�DI�ơ88�έ���2�I���O␍&?5
�	�.��1 ��}�}�p�c?a֯i�����0|2@�hÄ���;Q��;�0�M;��<��'��韆 ���)Ҁ[X�9p��_�ry����l��?f 	����C?���<g��c����<��#W�^�+T"��r���#S�
'ʤ8z��U<B$�~�M_�%n~,c��]Z0
Q��$�ybl�7|h��PHVDh�؋0
���y��YfT���c�=��5B�	F��yB&3dV@0�"���ȗo���y�@� ꨕ;�n[�x�^�a�
�ygnII�,ӷB�PUK�<'^.�ȓ6��� �d�"6Nܚ�*�O[Ɇ�^ d�9�ȥK�>��_�Rvj4�ȓ���G�8B��q0�	���28��FTi��Ň�VH��bG�Ǯ�*͆�)�����.�;���Ңo�<��h�ȓK�)�e��*��6��Ą�R���KF�\w�峵O�,u��h�ȓC�(���鏝A��i3�i(R<�ȓ'�"�E\��!��J��H��6�"��c@V/^���R&J�:�2`�ȓ
�R�h��_y�؍�5^��FT�ȓT}�p�Sk��@K�����NG����w,�8���V2H�|M���6)4�ȓ}$�,+���;��]�3M�6Ui�D��40�+�iӡq��<�e��)6{lɄȓ
"`��bL��t��ѝ$�.�ȓv7> ���j�5��	�51jՅȓ�t�3턓o��ce��7]�����x��-�1 a8Ec�/�(F*�ȓU�HMj�	X�=�	w`W"U����ȓg�<[�N֚(�X09���Y�4����K4��/O��Z�M͉E���ȓLȀ�����Bq��8fG�8w�<�ȓD��XAM
�_!:`��Ǆ$Qn���fDy26�R
��d�g��L.݇ȓB�z &�>ڂx����w��,��l?��0�-�wC\U�%h�2
 D�ȓglMsf��>y�4�a��[���x��a��̐Rtq�(I� h��&������V�]��5��d>0���b�ZHY惛8]������ ��|�ȓV���1���*jnܒ�dO�q�E�ȓ�^��Q-rt*D��K�t��+0��X��=
$6��h^%��ȓz�H��@l�	jϚ�R �Ф,\Ʉȓi�ɑe��UҠ�a�ըZo�t��}y�,���K�w�z�p�@ƥ<� Q��x낰��J@�bSx��땻?���l)�d�5�ή	O�aB�0nj}��3�p�Za�0F�ش�7k�e�攆ȓ-q�a-�1�������y���ȓq&z� ���}!:�{�H��u�t��S�? D��&��:#�I�.�9Ϣ��"O����ū2�6�;1��<�.�q�"O��ѡX��&YY �ƶ$�R�Z�"O��"�@�|ST	H�M�9&�޼h�"O8���G��y&�`mN�l��E�p"O��JWE�/��ʖ�C�
�@�b"O���e��:=���4,�M��%C "O��	A�N�sz�h� �?I��i3"O�̩���6P2��l[	h(��c"ONX(�T%!o��A�IJ�7��T"OhDҵ,�!S���3�L(z���"Ov�e�V����uŞ\ilxx!"Oh�R�UqE"�wV�Kgh�"O���CkU�g4\Ucݴ<�Y�`"O|����
o-98䁅)}��
�"Oư��j�D�v�Rp \�+~�q��"O��*��Q�Qv��]T��"O�5�B��:4�֌ARW[~��r"O|$�� #b���s�Yx���"O<ٶaЩn/ �	�kƃ]�z8�T"O(��CؠŰ,G ���xP6"O�<���������E�v�0"O@������F�ɓnƣM��)�"OԈ�T�F�pn����D�J��8�s"OJ��ԖKXȹ�U�&�B"O��#S,�/$>�b���/C��=�E"Oބ!0dġ[�ڤ1�i�{t�{W"OPD`���~�%�B9C���G"O�C�P�`^̲���W���d"O	jB ��j�U����N�iS�"O�6-OW7RݹBk�#Um��RR�+D�0sɔ5�^t�G�o�t��+D�t����#`Jq�d�jОH��G*D�8H�)҄R^lٖ�ʚ@�X3w�&D��V"څLchD���Hp�1�w�7D��JAJZ�Ix䣐�Ć�N��:D��󂉃U[��˄�"A
W�7D�<�C놁}�i	��J�&��"��7D��{R�*;�h�V�G�B�ï9D�B!��1})V܊d�+¸��4�6D�Ԭ]$%���q��C�h��3D��*	>NJX����d�*�e1D����;*��"�k�:�(�s�1D���$��YAf!��+-	�Uʠ�<D�`:��)[��س�ʙ1T�m$H&D�ȩrN�,Q���Ȍ`�X�q�#D��XmN�D`���/Y� `�d D�x#��|8X�a���>�ȥy��8D����y��5k�%� cv�u�gd2D�����w��T����3��"7<D�4k#�)�����Y-k���"�8D��[���8tB4Ыr�W�c|X��$4D��p.�!L��bB/���yz��6D�l����)��2H�r��eX��?D�`!4�¦��yrDʓ�YuT]s�C=D�H4��9#
|��"������k<D�\����l��³EC�Ŋ�� �8D�( �፠D!��W�(	ghH�E�4D�d�!�ҐL���@�J�u���K�j1D�����=4JV����		K��Ic�-D�x�UΗ=_*\��p�I�[Sz���,D���d�]!*�>|Yg��vI��*D���fI��JE��8o`E�aH+T��di��g9
�QF%��i��z�"O� ������;o��3���3�fH��"OH�r�I.bԉ���@�~�Xd��"O24ۢD�����9���>Z��%�v"O4�SM�hH��9a�5,}ҕQs"OlwĊ�\zX�AE& ���&"O00�%;E�	��� 2�V��C"O�M�z�Má���v�`7"O�U*6@�_�d���N��6|"�"OZp�S%Ǣ2�P�ϊ�A�vpP�"O�D����'��i�P�J(uf ��"O.e� =;2���E�Q����"Ot�2���Q��uŉ. >��!"O�!�2� �8%��s g�* >`�&"O�L0c����q�� ���QF"O�1��n��a4h��/�![
D0P�"Ov��6_󘥈�M�6$q@e"OH����lM0!p���T�Bg"Oz�4[3}�X�X�(��]a���"O�x��-<�C�❸HxtՉ"O�%9�a��>���k�a%0�ڭ�t"O\d����5O��!�� ۊi��("O*��īW
�%h��á[�&P��"OPt�3���QK<�pe�_u�P�S�"O�,�t�ηFT��X���m�hĺ�"O~)��iBxuR���I��k���"E"O� p��֎Av,}�H��O��l�"O.m+��Ĩ.Z
��h�V��x�2"O�UGᄰD2J�bdhX���i�"Oִr&�h��	 G�%Ш%"O�THפ��K~�r$�Z2g�"5"O葙�EF�O�&��E�3�� "O ��Q%�0bH�A���B�"�t6"O8�0f̎
Uh�<Zc��#D����"O���f�5c~H�҅��$x�\935"O��C6�TT� "��i�H�$R�yF�4z6}�[xBn@B��^�yRCS=vP^!ތh(2����yb��4Cֺ�
T��)Y>1
1���y"���X1x��H׽3�x�P��y�JY�bb� � U9X0h #Af��yB�Ǵ&r\a�J�&]Qfq{�$ɓ�y�o�,~�t��P���Glؼ�yB��D��h����8|8Գ����y���6V�`�''�@���P��y"�݇i���Y�c��l�A0�����y¢�;`0��a
�w̄���HG$�yR���\l��2��l5~e:`ǌ9�y�e�3,�l��� P*_�� �t$Ѻ�yZa	� ��D�QPi�L�y����$��t�׫H9HCD4)>�yBO4J���3%��v8V}�Rj�0�y���� OҜr}�4�Ō�0�y�L�
B򂄨�Ïm�E�d��y2FDS\����rLI�OG��yb'�1xT^���E��8��!�� V�y��0c~��	<C�n�K��C��y���%3ǜQ+ R9qT�P�1�,�yR��35��H��E�$By������y���,���)磏�Y�e��y��Ӝl
�H�(�����A!Q�y���Sd9bFҳn�å����y2 J�Y2~�!�W;v@[�����yR(��`���p���>��1	L��yb��;��F/�3iƕ�pG�y
� ���&��.��h��E�J�BC"O�a�-#F��ףʃB�&��"O�ܒ������0dJ<=�F�;@"O�	qCL@NR ��>�40�"O.�Sa.�*�ڬ�e���Z���Y'"O�QO
hz���0  �/���b�"O٫s۱j6n��C.�/�Ƶ �"O�T��ъU�
��73p�"O���@4v�H!;�퓾j"��5"OԠ`��*H�0p�M�.
g2u��"O��p�,�gC\�^a��+��U�y-�Y�P�i���\�ҼBf���y�ޤN38H�7鐫`K����Ҽ�y�I*� � ?]�f���j��yR睨�:`,I�[��	���yՓ;������1[�*�Ջ
%�y2��R� 8iaFY�<�T���a�!�yBi�$�Z�	R�H�`�`#�Ĳ�y�B �PU�8�0 ގM���q�G�3�yrA�y�zH��J4F����ʞ�y�F�8) `  �