MPQ    2*    h�  h                                                                                 V�E=���,��B�݈��'��`f^�X����b��zʄ�u�?��]M�q:���J,9��;�d�؟תD:���r��S<���/�kv'� 9)��v5kQck���p���t��0Jzc��A|gE�ϸ,�}x<%� �%6��r$@���ͨ�)5<Y��π�`�����
��}����s4�t��u&�>�x�?J"r̢A'T��;���gh��LZ�Э�8�� ,a&��[r��NpG�#�� Ә SEc�X��"T0q�L<|�~q�T�u�D�s/af�-ΩYc��D&�e�8�\� ���[��L��G�㖦�����I��:f���:k:�ax���<�|�����x4o`��:�5�H�P#\#��T�w�Y;�n������%��'�r�+�J~T���iԐb1�R� -��H�q�b�Ğ��� �]~YX�����6'����9�4W!�����J%�犻��L"��S�muW��|��_�	zA6��B��������T=4t�.2��L=��c�d���.;�HGK*��H8x�V;�X�`a��:��Fz~��"B�os�L�6m֫��x��Mw��F�%�ǁ��\x^�K����R��J�<��:җ�R����B5�| �c*3#�=�np�t�H�_�J�������j�&Yzd�".�4�k󫞶OG�����\�ST��6Vȶi�d���F~����*���lh],_]�;&�&����Hߑg m'�"�����qi�������A��Xތ|ː1�'ǆ@�rh64k"��v�k�^A+-]��살��y�(\Y�D�0&7FL�*��b3 9xP�ٙ���N�AM�I��X�3�\�n�60��w�}6D�N)���[�I�d�l�v{ZV�5�D�����Y)�6��� 7C]�5��:�|{���tОG�2L��t��!"m�0-&�lsF��J�b{rE���Ҧ����.�<�V`�q����T����A5��7��	���/���I�fI�"� 
�CZ��rN�]�%�����~���Y����l�So�ͯv�~��m+YjӖ5a��ϐ����Dti��r1������O�Z�0ˆ�eTW���&�vэ��Y���CG5���Ue���^L�R�|"���+t�?�33V��~� ��	|�n�c�ҭ�8_L�A+J)&b�D������9��s�6N�~�����X���Z
�g=N5��8ָ7a�6�3X�s����3��x_���.Q��lȾ��#�F�G�yeKn�1�.$+J�");b:���|���oJkNK���%�VXr��0b��2bg��\`��c��O�L�}�r2vh�,�ە�P7n�`�YD�������7Q��mcO���D �0���BTQM?Gc �#�/�r�5@0���'u
��f��Y_��h|�ש�~y>�@c�|����&��ޮ��$W(tL�m���)F�E�,,�ɖ�@�����f,�c���x�$w�J�d �����,��)wĕMe(12,@�~��k�V��jM�<�ױ���׶i��9n�L�r΀>����
���o3�X+���%������he8"J*�'0��Ȏ���m���	��]�|�.�V��>��c�C�����,	��W�T$�~*�t	���@J�(���О�x}�-��ܚ�����J����������2V�3�E+�1ᰆ\�e�n�è����8��;9f��}P�f�h�}3����~pCӱg��z*\���Z���rPN����Q�����߀l�sH�h���j�m9�(<��`��$z�FWjb���:��v�-oU��>��m|��Կ�Vtd;���|�ԛ40l2аyJ{$ꌞ_�W\�[d
���_h%�@w�"B[��(�Бd�࠽��b�c�xDq뺢FG5��:T���.��am�)}6nT�=�
�8"�]�d,��W��Y3Ȅ���&<@ߤJl�����ͳ.iJk�x^ݹ��4�J'�PV��P�t,� �,�)�������9�6�U�9�qv��G����R�<�[�/��x4��Z|m�����h6��@��F��A8�%P\�Ί��f��D(p]�\'��6P�r <e�E\�`7ޯ!��`-�ټa�0��+��`�4J����
2k�M�j��m���E�}�
�.�=(��ӦV��>�_& �ls������ed�ܲ�+4��ٶ�΄�1���a�ӕi���%�v����ߪ5޻#�
b��<��z� ���U���+= q�~*,�ػ3AK�<�[�v`������ֶ��Z���K�b�l��j7�+�Ɋ�ĳ�η�u����`2֠*&x��%z8DX-/�5�1}��1,�V^��uxq��2#��5��Nc�fp����Kf3^@��-!��>DU=�B���Z$`��iG��&�k3��gi�x�A�P��R���b�?�$��2�.�=���T��'�|���WL}&n�d̑��$]>op{q>���)��"�=���2��/t'Ʀg��TC�6ޒv�P��V(шk*�NVݜ-�yU��˗��<4�;1�`i6�|��/46����<:���&Y��)\I�h�eëz��,��nw�
�L�H�?~o�c�Bj��w(�t� �h�x4�_�GQs{8`��,���Tv��-8�\��T��֛���;�lWo��!�!�j�=e�G�ӻ)�����dx�$�0*QE���B�>� ο��2"�G%ލ*�w)��i8�ۊ���oN!J�:L�����{���0��-�'D��`�R����$h�c��$ĢfgҺ߭Y��	�� ˲��7��K��o²�e��K�ȿnꝎ���&����^6�[#��� ����ĳ��I���/T�i.����|���z��b�,�n�E�0�̣foT�eǰٰ=��%.���l=ؐ�����^�zf�N[�&�����i3�q��ϊ^�ɜA$���vu��H k�zL�T��tR~#�j��9�T6��	�{"g��8T�놋`�6b�)��ob�:���W�}>���ֵGW�*�e8�g#hJ6Wu|t�˔�j�hN~Y��/���<�_,�kD*�[B�&�B�ewz��S�ĢwK:`f8V��:�6������ԘX�KS�L��p���J?k��i�LuH�ð &�t�Ytu���,��k�<c\8kDO+ۦ+�cyz��8'�p���FBŘ)`a�\pa���(z���5H�Q��-c�	���I�$2�|$�Y�m_1V�M�;Pܨ�<�]`^��d46)w'�X1��SR��Q����Y�����4�9$�@Hr7C�T�3^�U� ��l��/��Cվ7�b�� BT�����L	ط%������β 0�h[j<t/����a�J*dQ��)��������ju�ә�i� �����[6A�	�!��kH���r7ޖ�.��~�Y,��ɮ}v�:���i�ڻ����c���I���mv��Eg��XP����Ú�x�M��B�畍��[%v�|Z�n�г��C9@��~>n�b�<m�wnQ����)��}�Dd�T�b��uz�
d�__�>F�11��)`���7pv�Sr��>%�-��Ua���fN��{
�M���pwJ��F`㼄�����|^����@��o�8<, ;:M�(R�T}�}����c%������pH�H��J�&��͙�Ug�7&Tģ�}�V��c����&O�f��GM\�����6Q�1i_�B�i��a���*d
�l� _�_�;!�x��mH�\� �I"F&z����qI
�>K2��^�L��X���˫>�'B7��M(S4��A���/A�b�]k��읬
����7�aD��7��g%9Zb�f� �������u뤭cI���X,=�hln#�30K�%����ɺ�����b�d�y�M�s5u����)������u�0o:^��U�vй��ҭsZ�O�}!]_30�S��gx�F��k�{��Y�Y���[���i�<K�?�l���&��'��/!���c����D�*�ʟY�D���Mп���^����V�]�=6���Y|��'��{��ƤyS�F���:�~�/�W���O��0�<�*I�堑�t���r�J����O̊�ȿ���`���:�p�1 ��҂5-�5���ѐ���q��^G���0����a+��u��g+V�b}�M_�줢Yn���qѽ�L�=J���bҳ����R���s�����t����ZX���Z���h��6����]�6��n�Ε��b�-�p�_9�.,��lK(��]��FТ�y������$F"���:�i�|.O�o�=�K�����X-�0}w�2�|�jwӁ�9�;�OG�ʦ�Bah<H۰XA7�c�׺DQ~������wQ�>m���������г�T��xG�i#䶂r/��0��B��
=RE�Ţ�Y�Ph��8����~��[@vO��B��rމ��_�0t�~���T)v�EXt��'�һ���)Q,��8��_�J�K6It��W��䶕(�h1X�o@%>R�f�#V���ȋ�Ơ�`Ȱ�Dݮ�t1L����{���4n��+��o�����c#`�	�GB�c�"�����ĸ�y��b|m���	���ￖ�G.��s���jc}��(D���̒�R$���o���K�M���)����a���������xʘ��<��k۵������ޓ��b�E������.��n�8M�.��5};T�����f�28>�q�?~k�����S�5U�\��ZG�r+���S��h�����:뺐.��h�j~�H��{�ȿ��FR@|�?�>��׌���o��>��s|�7p�Z��Vo]�A�ҥ�g!4Kb32KW)JV���ِ��"[_vp�Kdh�Xw@�ΜB�L��莑�c�X��?d�ny&x�Ro�ջ.G�Y����TTʬK1O.{�a��d}����A�
�*j"���dg�W;G53�QՂ�d@������$f͎3i��xx��v���܎���P?B�"*_��;�b͒,Z%v�D*u��9W��U[G��;���X����<��z/���/��Z�Z�\a����bh�!�IAsJyP���΅�f��(+4k�w¦��4v�M�!�C�\E�ު�C-�DA�9�N�
z����a��<�}�2�:��%?�Ȉ}��[��}�.�i)(S_��Q�E>+�> Mʗs�f�� �@3!��F�4N~4���=�v�Gk����ɒZ&��QK��@a��E���;
�ʠ���C�����enU_�f� �~%�Mz@�v��K9�E��v;���C�;_	���I�3	[��R�l��j��₤|��ev��,���⻢��ѥ�x���z���-
��l^���4Vz��ް�9#�w6���N>�s��\n�wJtf.Ew���4�R��DpB��Z�ۖ���Bk.�y��Z�x�^-PǎRk�����z�~��|@.���/qK��B3��pW��|&I��d����و>j�q�Ω����=jz]�2bf�tb��g��LC�IڒъP���(��O*+g��wU�y�'-�f"��%���`$M�ӗ�t/�p�[�^<u&���N9���IX1Le~��x���%7
�<VL(��?�\^��j�ʑ(��T �)�-׵:��Q���`?����1�v��8n�����v����l�A���+�!��= [����4�aqW�?�$�������j�B�& ����M
����3��)�D�8 荶���N|���X��eF��=
��7�hd�D+K�M\�������@���C���K��-�ː��2��˭<u.�؊�ư��޲�t3e�wOP	8?���&����b;[>�|�&�	���!��J�l����!��y6�{��|��|zi�=x�ԩ+Y�˩S�a��\ۥ����Ϟ��z$q=��j�7v���E�fа���$0�{`�3�xO�^�5^��ќ|֐����v������5��T�3�R�Uj�n,���3�ln�{_lʓK݈�i`�Wbb������uR��>䓳�j`��W��]�g�0�62M�t����6Ny狁��ݝ��,�{�*���B[���}��w��S�ޙ��ú`��8q{t:R�}�H��{����9 &��?�pW�c�,��?�JuB�L�<u�^,W&�c�Yy�Wu�\L���1`����\sj�O���+��zܘ8�
>��9J���sX1a	�Sp�ө�#�m�F=hHё����6��#:$VG|��K�h�61p��M�v��Q���5U�J64qIy'�w��^Rh,e��2`P�I֝ndm9_H��O��^��l S������� �W�T(�`��a�	o�M%m���������C��w�,�?m��\8�*�L)�=������Q�@uq0��' &v����6����ώkc�=���m
�Թ�,��*�x��u���N���G�@zˢ�u�F�� ��@D����w$��|�a[wM|�7�")�Fp.v�$�S��n��C0#��U��n�?��w�O\޹��~�8�Rd*�b �z������k��0��,oڄ]����p�JJryH%�`������oP�N
���u�ң�wſMF;��=��ܒu�^��A��QQ�*�r<G��:�*�Rtݬ��7�7�c Q���}p�HB�J�0���Ly������&O.?��Q_��8���V�O=V��&�\����6L)i�d �$$|��G�*?��l���_�̵;�f�j�HUG ��B"����,�q�销�"��)����dXTXu��k�'���(�4�J��.����A�&]&����t�o�O�D�u7|� ��b�� �o��7����Q����I
ېXE����Cn~m�0�w���E�Dl�Ϋ�M�^�dE���D���50h���v��O���BNm ��+1|:p_���\��t6�(�~�*)+!�q�0c�Z�b:F]��"�{�����Ѧ6���1�<濷�gh)�F~+Bj��J�Ě7���0�����eϭ�?�^���z{��yDM�ho]eu4�-E�����pD)�����S�� �l�.~Ʉ鼒ɣ�UW�+��Ʌ!�[u�t�)r'	e���@��*˿f��[<���Z��>�&�J��65��������^B]5�2_�K� +�#��oVdFL���^�?�pn����dԽ}!XL�YAJE�b�B��D��o��s���4�
�f��Xۑ�Z y�W�qC�mz�6�s!�)E���L�b�_��7.|l�����!F��y�5���$a��"U:��2|i�o�0\K�cٚ���X���0�?$2X�%�E��������B��(s�h�����:7d�r���D�Μ�j��m�Qr+mټ���`�&&��DdTǅfG�G#�]�r�"�0r+]g�
��o���DY���hG����m4~/��@�R�趥�S�d����-t����D�)�ާEܚ�Bg��6��굻K,-�<����gZJAS�g��)���rU���1���@�ža��V>}Ú���_�۠V�����LS�v:i8�eU����ӪN3������{h���L�^�" +��7�����Ёmn�	Y|�A:���.U����c:s���>�����$,vצj�?٦����D�Dr��nfX�㍟��
��>����䳸?)��۪9���E����&�J���n��mt�aȮ�;o�ʗsef�
��]��v�~f�%�Y���\Ѧ�Z�,�r�卧L����
ҕuI���h��vj���\�P���X�Z�TFM6rޚY�8��W�oKp6>���|!~����MVj�z�����JS�4f�2��J10Ì��-�[ZQ�lVVh�Ϫ@�?B^���(���g���k����ɯ/x�T����^G+�4[��TW�J���.v(�a#@�}�gfQ
��"dk<d��CW� �3�>��K�@U����K�X8�iui�Ex�����֎ v�P���=$����=��,����߹��W9�� Uu3� ��=����b�<8b�/'��* Z2h�𞶜�66���)A��@P=C΀�-f?D(�w���}��S��(����\��pޥ�I�-�M�T�Ժ�����&�v���,�2!ɪ����ȣ{�֎V}�r���(��Lo>��7 ��s�r��ټ�"=�(k4���8s��Z�ۑ�	D���p��,�L�{6c����x
�^Ȳ�à�8w�~��U:S���- ���~ �+�X��1~KT����v�Դ~���[����d��n�݃cl���j-!�����)\��I겓�V�3נ�AGx��iz.-�?�ɧ_�g]dV��y�+��c`�#�u_QENzԌ�h����f)L�=��ED��hB��Z�w\��e���k)���l.xn��P�bsR�jY��[��Ͱ0�R.�W9Ɗ����
��5g�Wq&$��dB���3�L>e \q�5���SX��J�2=�t��g3��C�|��,�PXn4(��*���R��y�j�͎���o`ߵ�Ӳz/*���6�P<�t�\ds��YI�be9s��,��d��
�ڎLc��?�P4Y��jC�K(JRQ 4��nG�>�Q�#`کT޿�sv` 8)���7H�Jrn�Q�!&��l�����U�!z�=��$�	���� 0��n$1�=����^�BbG� D�!�h!��=���J�)��8�)��W�Nר�{o���g��q��t���ND��g�H���H�o�%b��ދ�\h������,��͵�˨����+�E�3����P�e�[=�T��؎�w&V��ԭN[Yq���������)��۶�����]�6�|�;,z�b=�$��� �f��\�g�qD�OT\��7!����=���r=+��wf�2 ���@�6M�3����پL^Ңɜ����O�v����f��9TТARt��j�/��Њ��{w���bÈal�`7R!b�D�q�B��:����c>�v`�k�����X��Jg�6E>tM��̠5�Nt����L���&,ͫ�*��B6L���~#w�^hS�Wk�-\�`{��8���:�	�[� ���
��,@�iϮ�pQ�G�G?af>P;�L�P�����&�rY���u|n���t]�cF\���Oa��+��Bzt��8�O���� �N��aD�>p�E���̆���H�a�����>���$�|+|Zh��c�1�UMN������S+��s�74���'�u|�%R����Jk�M���Rh�I�G9�`5H�|��J�^H�Q u��G�:"��N�>��Tî���2�	ʘc%(�ʹ�m�����������U�W�*hk��b��O����BuLUv�!8 �i!�~M�6�V��� k~�h�L�H���zZ,43�sE����A�	�x�u��1���¿��1ף�?�;A4yq��2LY�/,���]�MW"=�]�����v��M��E�)?{CK-�����n�<9��}���t�����R���d5-b{�Zz�:��7̯t;(�'�&��z�t�p�*)r�+�%j����C��
��N�2 �l�`��%� ��w@�F���xMJ�-V�^�����@��P<blF:C��RO�������M�Kc��N�p�Q�H1��J�������AԠ�;e�&J�6�3H�e-����?O�e3�%�\F����$^6Gg�iY��ߞ�����s*>"l��_.Y.;������HR� ��"<QMէ��q��S�t�����X�W��*'8�x�}4���G���edA<-�]���������B0��rDG�K7U�?bD� j��R���k�u���IE�X�}����6n�8M0��m�� ��=ZΆ���z�d�3:�[�k�5�)m�p���o��Q�}6���&F:ˀ���E'��XJң"���!ӣ�0�&��]�WF�W�{�{�R��O΢�����n�<��Ǿb�5����̜�eu���������>=� ��:"�Zr~�5i֨��ݪ��]@͂�h��O�+��#+����<v�S�F���Af~����'*{�&�6����ywt��Kr��I��5�� �a�i�V�����䨧�A,�+`�5�n��bP৫A^=� ���T�d+�t���0 V?J��=���O�n��c�'޷�8ƪL��J��b��_�N�ח
��sz�q���!��X���Z{���� ������6�Cp΄���P��tN_/2.�l�H�ē�\FƸmyv���bL,$|�"���:���|���oC�K�Ɇ�6EX��o0�'�2�ɻ� 
�Z�B�qh�="Y��÷h��)���:7�ލ��.D����TS��iKQͦ�m��9��S���@���TRG4��#�$�r���0-��x
3��{:�Y�3h�W�����~�R}@�O��K��Π�?��՝t�,���<),ۥE�cX�]�Iұ]�mV,h˝UA,���J�z�y��D�����y1κ�@[�\t}V�Yf~8��(Q��V�ȶ�����dL�n!�q����%V������v�£�,։;�}́�Y��"[���X�����
_�mII�	��T�P̖��.�p�o2EcU����Ȏ�����j$�!�e��ܕ�YH�_s=��u��Aa�K%Ϯ�<�����!���}]���G��!�E�Z�aկ�d��n��
�/��iմ;��$���f�&6�.����bS~ac9�x�:ͫ
�\�hZ2
r�͊��5^������0����ɥh�W�j�=7�ҹ7'��a�FHLD��.�k����So��>[��|\�JԐ��Ve�������_�4�H�2A�J懌OS�(Ɲ[U�M�ǁ�hVf�@Ȋ	B�������䃠�o���$�xuv��N�G�2�6��T�B�����.qjya~�{}g��2
y�"?"d��Wq�T3�K炦˵@����Pk��D�%i���x/K���\l�[M2P����X>�,^��,�U��ziP�D�9ޔU��'��%⸉3�y�<s</�̓%�Z��z��V�o�)ޥ�hxA�|P،��{�Qf���(����Xd�}���ʝ��\{�1ޠ����t-C��oS�� mVҼf^�5���2|wy�2Ⱦ���Qc }r����(��q�G	5>� ó�s
5��u�Ğ�0I�c��4��R�ĝ$�B_��j0�$�"�P�����+��{��>P
s	=�m�g�˪�����U�x��݆ B�G~��0����ĂKok��u��v�9��������L[����>��l�$�j�l�Z[��dr"���E�����q㗠G�x��z���-��������V�����#ܓ�}2�N��� 䭑mf$s�������0D��B��Z�3�V��U"�k$��x��x)��P�V;Ra�s7��H��o�.���	�X��PF W�3 &��d}�΢�>`�6qO���Z��s��pX2��t�nBg�ReC������Pl	("Hq*!��-hy�_���>�6��Li<`�>C���/��z���<�⎔������I"�e���GnI��� 
��WL�T�?O�#T>�j��(�� Okj�1��6Q$�`u�<޺]v�`98�#߫R������,�(a��l(���T!զ�=��i�$@��W�t��TM$l�qؕz��s�B��7 ��؃Xڸ�����)JoI8Va\��7rN2��6:ރ߉z���®O�ޤ0Da��C�����S@{Ǥ	웢���p�@�A���h�ˣ��%�� ����в�K_e��x��?3j��F:&�w���[tT~�@�z�%�d�i��ݞ���zp%���|�	z_����'�Ĝ�Q
�W�K�(��
֑���p�^=it٭$q�/�zf��\�7�1��Y�3�D�T��^�����r��R v\��Y��ū�xT�1tR��j~�A�������{��I�Ɉ��`R̒bXfLV���B]�(��>�y���3�[���g�!n6�\t����;�[NocK�@ڌ�mE,���*�$B��0wKDS��8��<`6QH8�ь:H���6��1��)}^�ͷ�]��p�]��b ?�O^+TL&�A����&㡶Y/�_u7�S���'� �'p\���O��+��1z�.U8X���U@e��)�a�p2���i�����HGQ%���,	,�u7�$��b|�d��^�]1&��M	L����b��@G�N�i4��'�/,wI�R���P1�h���?�Ɲ$$r9�˭HCOL�E�_^��� ����Z�媾Ȟ��y#
T^���# 	%��%��%�ɲ~�u��L`���u�+�R��*u�M賽����=�G4qu'�l3�� \}w�y��6R�E�Rwk��.��|��#"��/�,ϱ��n�%�+����vV�+X
�6	ߢ�����j��>�G�6^9�-J���Jk��W��M2�R�=��|�v�Ա	�&��yCfWp�Kgrn�Y���5�HM��ݹ:�fծu;dP4�b�i�zg'����fu�"K�:�'�/k�p�*�ro/o%E&*�fХ[N�{B��T̨~��;Ҹw�<�F�����&\��V^����QXЭ���<}B:�=�R*O�.�����c���ڨpy�MHL�CJ��1�_B�|�{��;�&Eb���� B����O3��dD	\�|��Qfe6B܋ipm܅�>a�n��*�YlT��_�?;�� -�H�|g �o�"�9Ղ�0q��F�2	����]lXʣ~��%('�$��'�4W�X����;�A���]�8u��T�e���ģD�	�7�B,��b�G %��m%2��~�d�I�yXPց��KFn4$J0|V��.��:/��ap5��d{��桒G��5���3�J�E[%ڢ�}��=��!l:&�������
]������U!�0��o�X�F�[6�M{�A��ʠ �����̻<�o�]x������O˜�O�-�������盎~�5�G�4��vM���6�^0�]E!��A�G��Q���F���S���b��~���������!���;23�ќ�t�?�r�:�p��;�����Q�u�K7�b��\������5^���A���B��^8[��N��D�+��ȇ��VnZ���1�u֧n�P��w{���L2��J�bc����x����su
v��a��J2X �Z����u���M ���6�3[�����+��_���.��l�u�.�PF�s�y������$��"}x:^y�|�P�o�u�K�O��L�X^�r0�/�2N�=���́��u�8s���3#hm[��C7Z5�h�@D���[���Q(B�mO�D����I(a�kT=>^G��#�Tr@��0�"��ٔ
����V��YK�ch}6��ñ�~�C�@Ol ��Z���t�����k)���E��x�@�,���k?q,����B�טJ���z�:�_���햕��I1	�s@�<ӾW��V�ˏ9��C�6�ѱ�����%;�L���l��t�m��/�D�#�~|����î�TI~"�|,��E�4�7���m$ǧ	�Ηw�v���.d��*��cp�����~���=�C+�$b�d�`E|�\���i�z��d�ޚ��܆t��I������|WP����������E��6�/	��+n�W#*���$�V;���i��fcPr�iF�BoA~\��w��f��\KZ�W/r��T��b��o����K�&�_ߍh�$�j}o�h��r�IȐD`FC���P$}�&Z���oA�G>6�%|�jf�+nV`���R�ԥ��c4��2�
�J�܌����~[Pzf�"�h�@��B����
�P�"�)�W��Ӷ|�x0�K�&ǗG!χ�fT��Ǭ}�.l�ha�bW}"�:9|
�"��d�jWԘ3�x����@�C;�����YCi6��xʯ>��T���D�PB���sx	�q���,��9R�9h IU�0`��JK�3R>�T�B<��/]M �Z��l���Զ*�,=����7A$�,Ps2��v,rf��(\_���SO���0���3Q�<\�
ޛ���-�-�Q��9X�{�җ?FLއ��X��e2�E�V���ِ*��W�}MZ��X($�V�Bö><�� ~�ss%����89��_Eܞ{4��"R靃kxӔ?r��e��x���@��h����
�X;�(0��<n�t��U�<u�� ��x~��-�ا��K����Fv�����P0a���2.�D������l��Uj#ؐ�56�ğ�&��Г����̳ؠ�xx�R�z$^-�+3�؝mV������#��)�3[Nϻ��R��He>f�����	D�!B�}Z�X�U�ӏ�`k�����x�t�PkkR�yRN�v�+�E�f�.��l�@�E��o�kEDW�&��+d��1�i��>[P�q�d,���Ș�;2��t�3gi҅C�B7��PΉ"(=�*�p���.yAQ��7���t ��fi`U�����/ [��Ǆ<&q�������GIiJe����b��Z�w
^v�L��8?�+O�j�d�(��6 jGdڠ��/�Q_L�`�\޵��v�8�m�m*�@�'� �8�lå,��	;!0Pq=Qy��?�����%��3$�Ys�|��B�� �~d؞�.�3O~��>)�4�8��'��7�N��L�$W����gn!�*D4�uFD�qO�>]���x��p�$t�R逺Km��|�_�-˞��?{�ػ�9�ۿ��g�eiQ������󎵧�&�h�J�[�W��lm�U ğ��=���4����'|�zڥ�κ��Z��ǜ�9�R�k�m����w�� �4��G=D ��+��ʱ�f���������3,e[��-�^����-�Q��v��p��c�fk�T�.Rj��jY�d�@�t�=\�{�ʤ����w`mf�b�߲'��&kW���)>՜��!���aь�gJ6Ô@t�����J�NjQu�����(�|,l�*�,B����.۱w�I�Sҩ���<`�4d8�,%:�pD����l������Q����p���}f�?WY���Laٵ�/_�&��Y��u���1���/�j\$(%O�5�+�}z*�89����p��Ea�h�p͈�N��WjHaɻ2�����PqV$G�|����Y_[1�S�M���ȿ�IvB�)��4"j�'P��r��Ry[�=v;胗��3����9WzH�A��@)|^��; ��*��V�����������T�I��4�	��%�,�)�,���O��2}(9��g�Ml=*����n�Y��k���uWnZu ���t{E6�C/�e�k���^)��]V�jɫ,jP_�i	��?��S�F��� ���p%�5-M���ǳ1��/
����ݘe�ך��JM&x��
t�n�v�ܱd�'П�C��П���na�?�(��,x��t�����i�dki�bqBpzB겼Kމ�������ڕʘ�s�p�J�r�R% �!�A P�@5N��`�"ݷ�9--Vݧw6��F�Մ��cw�^�	�� �[��<�8�:9��R8\�i�\��z�c�p4��Hg��J
���:�^���*�q2j&@,:�����vu�2[�O��?�}\�������6=q�iˡ��U��Ѫ	��*��l��_d��;Bي{��H��A ��"2���]��q5n��i��Jm���PX�y����'.9���g�4�
^�}�Y�1
A�w%]W���	�#��'��DD�OT7MP�}b�'� ��7���l�aEw���4I�n�X�N���qn�/�07�F�}���@��<`	p�d�����!&�5a�N�����'�}	Y���>�E�7�:�#��A?h�%��ҙQt����!Ih<04z��SlFnP/�	�{�P��E���"�UI�<�ͯ�X0#�WD^s���I���(t�`�3�0/ �6��0V�Ы��ʓW�ٸ�]���ޞ��;���5U�#��S��i��ș~Z�CD?`&b�� ɖj	��-t���r�8�K�r�v�J�7�x�L��ꦚ٨���wX��!�59���|�����^3
L�C��|�v+�v�}yV����9�Y�}�n��0��0��o�LMnoJ���b>����B-�@��spO��EF�����X,g	Zq�����"#��>��6�C��:e�N&��z_%=�.���l7�$��i�F�Ny,/B��7$�;K"�]<:9i|<�oQ��K��u��X��0�WG2� ���"�Р��Õ3�צ9�h(�`��T7ի�C/�D=�Ҝ��e���Q��\m
����R��
<<��TxJhGj�F#�r�u90�����f
)ĸ�1R�Y��gh5D澃T~@U@
���9���]��PK��tSe��{�)�3�ED��ԓD�ҧ�1�F1�,������?"JR)O5���z?���9��5J1D�@�|n�R��VO^��Ӟ�^[N�L���<�`~L$���g�Ij�������]��Yo�L>�����OF"e��β#�OfԺ ��m�d	
(o29���.fwG���c����`�s5c�~�S$����[�tٷ8���r������3��t	U���o��dA��$e����p�P�,ϛ�x`�ErxP�שV��n�L��8�����;��p���zf>������ݛ�~W�4�.7��!@�\"M�Z� r��N�?6��׃��Ҧ�u��h7j����ȹ�(��+G�F>�|ޫ9R���Ko���>�|���Ƅ�V[ɼ���*�{ց4���271aJ±��ŕq^Wy[Kf��}8�h��@��B�Ri�o�h��<u����Zƶ��x���A`�G�����T�Ĭ�+�.gN�a4$}��nT�-
o�i"���dS��W��T3���\�@����������piq}�xe4\��ll�\4P��9Î�?�G1��@?,F���({�
9�B=UG�����Y�:�/��<��M/�a�ġZCP�H3�����p���gA_�PP�E�q��fP��(͛�nB�sn�ƹEZ��,\��ޖ5�Z��-�?I��?V��ߧ�r8���QL���224W�f�����Gl8}(�U�q(����=��>��b 90s@��k����1��/�4��Q�������I3�y�Z9��F���r��,v1߱D5�
��
)�Y��x����zU���R>� xb~�-��%�bpXK��;�k]�v���/4 �A��8���^YݴU|l�j�c��1?������S��i��'�����Wxƌz�4�-v�Z�X#��8�V�)R�<�Ѱ���#0�sU(N���M���XGf!��NM�>�D�jNB�q�Zk���$ɏ���k��.`1x��P3�RW1�)e�f-p��Z.��@ƛ"���!7��d�W��&�1\d�l��(>V�q,���ϔ��f�2ΙLtNYgr^C��#�=��P��(X�*	���4Ey|��Ҍ&�ҁ���`�@��+/�>����<a4�-e����IĒ�ej.�}�����
9t�L�A?��KJ�jT�:({� ��K�S<��؛Q�`�,�ްm�vq}�8Z׵���E�_���_��l^\���}!�=n��Z8r�M�B�2�$�3�������Bs�I u�ع&�ڮ��q�n)�C8�Z���W�N���/�.O��,����Te�D�i��9H>�YX���^�?f���*�&m����G�}˙T�����v�Ұ��b���;eD���u�u��(�&g���Q�[�z���0^j���?�$t��kr�0��g�(|,,zUw6���?ԕܰ�7x��M��������9I�;ê�f�|=���#Sy�e��f�x*����gӪ3GIڏJ�^cGR�h�$� &�v��٩^��!CT!�qR�_1j4���{(��@�{	!��h6��4�`� nbNݫ���a���^(!>����|3��NF�1�g���6��t�+��q�Ne_{��T���>,��*}+/B��N�i9�w�ocS͂Ȣ>�`�88ݧ�:>O���?S��`��_~���ܮ�pC[����?҂"��WL�Mޤ�Z�&�_�Y�chu�l#��r�b4\_�/O2��+�E$z��8��[:�6����S�a��phZ��Sц�6H��q�M�x"���+�*$B�|+��T/�1�"pM�k�/��������]4]
�'�^�m_�R�UU���螔��5���c�9K�HyT��;�t^Y�@ ?�ԓ
x:�y���~4y��o)T�Ǒ��eD	�)�%Y�b�D���t�5ʯ8*c����O�Hh *+z��)k��*s�=Ru�j�&� �̞oB�6�����okϸ?���-�ٹ�ԥ��,!�d����%�:P��a`m�,��bw@�p��t��,�����c����I��M%TM�׭��_��Dv�N��H�Z�C�ٟA��n<�
�c�~,���g͹�oO�$�4d���b�:�z򎼆��E������̘���p��6re��%�k��|����TN�m{�}�#���q�w�9wF�xC�)9<����^�c.��ϭ��<�N:��R�@L��N�&�c`�_�Fp�N�H���J���\K����IS&;F�D7C���#�MGrO)T���\�Ч��I�68&�i&���ޮ�o�q�*���l�P_��(;�7��HA2@ Ԁ"��8@�qpjɀE�����ݖ��X@o��2`{'�����ǔ4�e��y��G'AMM�]��$e.�[��~�UD���7�}2^ybU(� ��X�����+
�c�$I�߱X����ꃹn�Z$0�c)��*�0r��R��4d�� �`�||75/�i��;4v�Xw.l����y�:ܤ@�����@���I��DA!��`0�Se�Ny�F���A�{�9���`��fZ��0<R��S�Z.����c�#���;���k�_���/�+� k�f���@�Ta�]єN�R �����a�m��S���X��~5P2�~�� �׏���_�GDOt�rCA�&��̱���Ҏ$�G���D�؉Q�������59ѷ~a�x^v^.����X��7&+(���MzV���t{U�C?n�d��8
��it�Lh
OJ�b�4��,F����sk�� J.�RJ�XG��Z�b�_�]�]��,�6�sΕB�	A0#k_��.sO�lr��dq`F�I�y��ƕ�ݎ$͘O"^�:y�|UG[o�:�K����G7�X�ˤ0�x2DL�ݤ��7�B�.u��tzh�B�7n7PB(�Dx�Q�%���\Q�شm�G�9��{�3T�v&GV�#�9r�{x0^��ˀ
���gY��?h�S#�u~��@@�˳T� ���~��t��$�vx<)=��E���Ԯ#��"E�!C�,S9&�8��GJ��%�qe��	N�舕o�z1c�@,���M�V����~�y.��B綋������L�ni�b��GA_��+P��:)�4���tm�N��J�	"lm.��ƅ�j�x�{�m�"�	E�������.��L�[c�����#o�N�8̹�$��ҦV#�������섰6e�Z���O���r���G��n:�2Jm�+<��G��/�EM7Z�D��5υn�a���/Ț4�;��b�_�f��2�x��~R������
@\=o&Z�~rr�x�z����ك�����j*h,�js�o��:�����i�F9N��o�����x�o7�	>�m"|���aoVV
ˉ^�6B$4ґ�2�wMJ��6� g��O�[Fr���_h���@�YB���Jl���|�_:��1��5��x���\�Gh�s]TC���R��.b�[a��}�چo6G
꯷"��d��bWB'�3�2����0@AS���b-�ռ�i�z}x ����֎l��P��éL��",��K8~v�9�qUl���/�)C��
�<$��/��G�:Z��q=7�
7Y�"���hQA���P����l>�f�e�(��o���=���Ɣ��Ѱ\Ldޑ�+��s-t���e|�qɒ�MQ&�&j���(�2�Bf��?����� �}�o�%_(Z�(�8��>��� ��s[ɵ��f���z[4U���!�S,(��$�u ����Ҫ��h�g���LAB���
�W�Ȟ�,���j�7U����� y~G�A���v)K�B-���v��I�j�f汎�^h��CI�o�hl2�jjL��K�u��� ϓ�Z�₴ڠx�x1YSz+8-Q�ɓ�\��?�V��'��^�O;�#-���!N�}9�����~l�f����ٵ�KD���By�ZF'��˻��&>�k&����GxZ��PN�R��,R��ώ���M.�����숉i���$W�:�&���d.����@M>Q oq`$������6�@�2���t�7�g�1�C��̒��BPD%!(s'�*���ݾ��y��"�m�^�P��]��`˘���]/B���y<��4�����%I��e%����&�Pn�
�LO��? ��E�j�ku(6�� ��xZ����VQ��!`F�EޫL�v�;8aG���6Dֽ���l�2��=!�y=ǂ��u�����Q�$.N�����r�B��� 0���Խ��)$�L��)��8'�����NC�^gZ��0�5�]���#�uD2��4S���q<��Z�|�H꠺����؃�9 �˔*K����1�ϰP���e��)����l&�X@���[Ž=�����d��s}㞐��ы�<�"G�|G4|z�h����S��I��;A�H�_�#@�;ˈV�h���=�w��^�;� �f�z��H+E�"@d3bM����^>�
��1�����v�b��j�_��:PT<�<R`2Zj�ڬ����sEu{�Z ��M��`���b��P�\E�������>�Bm���O��\���g��6yd�t9�y���N`�]�QB䝞�c,9��*��B����w��S�{�����`g\(8�Bn:�M�������g��.J��nP�p�	o�R%?M���^�L�ẤevQ&���Y@�uh=�>�J�3=3�\�FO�"�+��'z�� 8���UM����ź"Ya0�tpL��
x ��iHx��h���(��E$}��|���O+17dM:|��Jr�?A=���4�ʑ'�&�h�R/p�!蹱�갔���3�9��H���6I^�� �w�%����;Y�g�*F�T/e
�Ӷ�	6��%G�_���&(ʊ^g����FX=�C��*����q��&J¸�u��p�� -xʞj)�6c�B��hk�4�T⻖�5���M,��:�_M�<1��lH�|;��O'�=�K�9�P0�'u1�"E�+s����ȧ�Mé��I`�M�Ev�L�;��JKC�����o�np��^L\��z_�K�#��N�d�3fbgS�z�������m���K0/�`�p�r���%�>a��<��v�lN����M���r�S�w,�_F��A�dr
ܙ�^��o�b�?��A1<΄>:/ʘR�i��L��1cLg���5p�8zH���J G���/�-Q���&6 ������Q@��hSSO���`6\2+��"�K63�Bi�jw���[���K�*�%^l��_��;b2�1�cH��b *��"('�q��X��8Y�� 
�nk�X����M-�'$���oG�4�d��[;�} A�B]ͺ��?!��p�Y��D3<-7�˩_�b�H V
������W2��>��I1q,X!����OnE�0���:y���Î��AL�+^dL^�����k5�p�Ą��¶��3Aei�t�>��:7F����9�[)�ҏ ��q�!��y0jM��I��F$��g�){/�1�;�b�}��ˣ�<�v��N ��v�/�ѝ�����_�����l��&n��;z�!`K� ���)�]�l��T%��ث����l��(�ES,�ͯ��}~����@�Q��0��L;6���t&�rr��V�-e��x��m��B���\�N��������F85���r��ڢ^)ȇ��&���+1���sB;V�����z%�F*n�n���$��L�ƖJ�B�b��[�:7S�v'�sf9k��n���.Xb�HZg��:�G��-3�t�}6����𑗐�{>�G_�>.N��l�	!���|F�d�y���N��$�"�~(:�r|�rAo��DK��՚��nX��0�2��L匸��F�Ɛݞ�)&G��Dfh����Rk�7��s��D�%e��5D��DQ9Ԭm�~>�TW�������T�G�)�#ƀBrQ�w0�����
=�����Y�I�hN�Z洇6~��A@����oۛ�lޫ��fkt���qU�)��E��w��"Uҝ'���t",T�����o	JX�1�����J��1��L@�[;H�V�j����B���f,���d�LZY��]0��D��\�Fª�č������c�E�"Ǖ��D�k���%���Rm� �	�:�H���b.���[m�c�!�
}��)'����$3ަQ��m'�E� �˷��\�*Q��7"-�r����k���˸�Ԑb���nE(T�M�����rn��V;�c�U�U;�'ݗ�Iyf􍇤��U�~M�����͗��\X�'Z���rM�Ҵ����S�����\	Ԑ���hGL�j�����#���a��F4�%�a��W�.3��o��L>���|H�q����VQkՉc�W���J4픉2-�EJx�;�;X5�h�[A�Y�3orhBJ@4��Bv���%Mv�7�����(`����xa=�w�G�d����T~�:����.]�_a�+}S����
e�q"�=�dɞ�W݀53��܂�Y@�
)Ķ�Ͱ��i症x��_���܎��Ps����z��:6,�6���g�q/9y'�U�9��.z��k'��9O<_"�/.w���Z�������%���7ۥC4A���PD�u�g��f>u(����A�i�X�oAW�\��&ތ{س-/�%�۫ʺ�ҩ�(��zi��m�w!2�p5��9m�*�N�=��}ޥ�˄ (�&�3�d>M15 �Usv���a��b���O�4��0��q�鮰��Ӕ�'6�<ń�s�W�@���]� >�
���Y�a�7�͢���U������ � ]~�\��؛>K��a>�v]ﴥ*[���ܤ��UI��*��lM��j�ڋ�ƆA�P�P~B��k���䛠3,�xL"z�A�-,}Z��E��n�V����W��
�#HL�i�FN`�����fO��:n���,D]�B���Z!cj�s0���k����>x��PiglRM s���ܑ��7ָ.�H]�Q�@�D�����Wy}�&k5�di��:�	>L�q�ЍF���F\��2��t�Ag:8C�[1���AP��(�\*�:ݙ�by򚶈o��؞�1`����9�w/�ej�} �<�۩�c��h�Iz�Qe�y��ڀ���%
��L�y?���@NAj
P(�� ���զ��\��Q��`�#ަK\v' 8�
���m�Hx֘gfM�l�)���!A�=��e̐��Cn��a�)$XH�D\S���B)\ �]g��t�ڤ���'�B)6D�8������N�E"���KR��ؾE�����ʥ�D͸�/~��Me,�u`�����̀�-�Ԣkˏ �P;���P1�,ȕ�|y�e���d:��a��� &9l�{m[� �`>��i��PRf�j��cC��݄�ݽ|b��zKz�_�u��m�C04�~A����qo�\o�=�cٙ��=�f��h�������3}q�@�^U��ޣ��Vy�v�O��V�ŗR�TW��R�$j�.��k�j�{�Τʵ�#�Z$`���bD8��I��ף~��'8>����2�٘G��"�4g���6T��tt2�̧��N[���Ol�Yh�,T|*s��B}ZI��U�w��SÔH��5@`"��8�:4lx��Z��������r�ɳ p�ؐ����?�5���bL�K� ��&ϝ�Y�`qu#��Y��&w8\��Ohɶ+��z;TO8D��p�n,��ŕ�akg$p�]����h��H3Pλ�_ms���$�f	|a�p�J/�1�!xM�vs�e^�ں�<�4Ӫ�'!7c�R���n������+u9��#=9���H����1��^{k ��T�@���o��4J��e<T�"{��'Y	�*S%ϟ��z���j�&�e�4��B��s�>��*��蟘��AI�3z�u��' ��e0�6��l�>ykkq����8���,;쬮Z���������p�"���F��3�ת��"'@_����C�����CJM��I�2t���v��Zu���М�C�?�7]!n�2��V������t8՚,>d���b⋋z�a7��G��{P��|ڦ��N�p3kr[}D%�1������|N�ߤ�36{�j�[���w��TF]�Є��l�4�@^�k͑��O���C<�ڠ:��ER��<��L�Tݷc����peBH��sJ{�j��#��h�0�B�-&1Jr������,��O�#��z\m�d���36.�"i��U�����zFR*ao�l@�_5�r;�!Ɋ�j�H�g� E�"�l���	�q�j�{Ў�����U~X����h�'����J��4C|f�N^p���AX�]�{'�Z���QL40�Dn�G79�7b� V'��qL��XT�|�Il";X�x���;�n�0h�ڣU'�&5�����!�;d�E�据�2�`5��hğ-h�1����#��8��]�:�.�r�x�v���
7�L�!�~�0g;�D�1F��"{{J>�׶*�X�����<�� �I��h*�����������>��{����!Q�!~���Ҩk�JE]�d���@V3(��I�f�����SG�ۯNR~�uw����1&��bɧӌ�ktA��r	 x��z��'����ě=�U귄��Nǳ��
g���5�
��-���u^$��T���k�+L�Ӈ�VHV�=8�����07n�����K��ݥL��FJ��b�;s�uaT���sa�_�V�@����X}\4Z�9�A��bl���6�3 �Ka���Y�*_��w.)yTl�ImĚ�PF���y=���	�z$��"�P:���|˽{o"��K��Ϛ���XJ�g0:��2:C�g�<��Cʐx��$�x�J5�hY���m޸7F����*D��[���5IQ��Dm;��o�����I�T)/�G;z#��r��60ԩ��=�
������XY7�lh���毹�~QI#@;����#xކ�a�� t$bx�lR�)�Eu�I��Al�*~���},�M�\���6gJc3f� ���q�c+�%�l1�s�@b���C:V`ն%-���E�S��A���lL�c'�X��Zb�З�a�v�0�������(����@-�""�0��Mָ�gںq�m���	��m�s�ߛ�.wq7�L�c��]�������/|�$�[!�L���ȳk� Pل�X�P!}��[�r�Iϵ(]��b���
���}���.E>����k��n��_����;�ߗU��f�7�U�����~H���?5��R l\s�Zx-}r(6]��}����n�ҷS�Kv�hb� jiq�~��^����F/�D޼9��N�o-�{>���|��]ԗ�PVL�ۉ�~.��y�4��2�dJJSSьviu/��[<�⪎:%h�7V@O�WB�f�� N�<1���aQ�?��)x����jG��}��T�Ƴ���f.X��aE(�}Tc�޲
�^�"���d�*Wx�Y3�l��m	�@��mD�d��p͋�Zi"եx6�E��t�"b�P.R.�ߠ���x�_�y,�~@����lS[9�ɚUx'��I5��b����<�u�/�1�� ZTX�yl�@7(�˨�7�A>uP��b��fa6�(H�A�4�L����J�-=�u\�e`އ��k��-�
��A�g�����8�"ߏ��2C���BS��E�ʸi�}����(��[�.�V>��n j��s�!H��vC�=[�܊n4��Զ�v��	U�d���NO���ªN W��մ߂�$���
:�u�I��R�=�`pU\�H��Q I�n~]��V�ؓ�K�i��ރv8��������
��nI��gnlhm jƷ����ċ��������d�85ݠ�xg��zx�-�2�	z�	�V޽'�M�Y���#c
��y�N;���>R���f��_�µoD-�Bow�Z���AJ��\��k*˺?txЧMP��<R�V��t�����.¥�Ƭ����X��ׁ%W���&F�Md�{���I^>G0�qB�����u�{�2_P�t�g�9C�NR�N+�P�@0(��r*��B�t�iy-����lW��Ξ��`A�+�Tz/���X�.<꒔��*���I�+he��d����Fk�
�-�LŒ�?V�;;��je��(�� ֙JP��7��QKf`|�ޡjrv��8�Զ��nf,m+�s~�5�l/@l���m!�5==̫��ʾ�"�<�$��P��5�޼�B�a� �=�
L��y����)q�P8]�F��w�N������f��S�T��W����Dh��*�;�j��������>k�,Y�ho��oe�ˊ6?�ا���G`���eռ��z�F�ˎ�k�&x9�6�[�����F���
ċ����
����A	m�T|}�zƫ��:~��F��#)�>�D�ٗ���>��n�����=�oW�Ԉ<�6��f�ޑ����y�3��Ǐ���^�L�6W��Rxv�\�� ]�R��Tr�jRV7Pj�{��,�:���c{�����ʈ��`��b����Vg�LI�/�W>�h�֍ڣ�ؘ=�g�+�6/�t��f�B�}NVI��}T�A�,ol(*BX��@wR�S���O�A`��8.��:��L�}	��X\��0�_ݡ�$7pt�V��?C��r��LMj����&�lSY��u�Ot5��f��r\�GO�+��Bz�-~8����e���_�p -a�Q�p9��� "3�û�H�߂�����'漘$�[�|�3��E_k1�P�M��-܀���5���l44�;'��^�?R�#)M��K��u��k3�9���HJL��,��^j � p�*�[�V��,����R�Te ��ɸ�	��i%�[������31�@
��L�|���9�*<��Z���\$p®[�unڎZKa c�o�`W�6�V���k t��J��j�$�V�?,�
w�U���D��k	�����t��K2�!v��ECy�Ϙ�������цn���My�������v�<��)mЋ�C�	㟲j;n�ɍ���O� �� ��'��U*)d�}3b]�,z���7�����	�������7pNmr� �%�Da�-��Ь'�N�ȳ�>g�%���I�w"�UF8R��Dc��9^�G� �G_�<Q+:%Rq=�U5Z���uc�)*�prTp llH�I4J�/7��7�O0��L&,���Us�ǉ���MO�b����\�?1�X��6)i7�4�A=�9���`V*<�\l{�q_�D|;����IaHr2 `��"�����q!��|�6��$`�Xq>˃'�';q�%�}4~7���}�I�A^�e]C\�u���G&�)D���7�ƀ���bf� �����T��M����TI���XWq���G9n���0#詣p�����1Ψ�O\��d���戅O�?5MT�ĺ�#¬i*������j�����:��t�-��БQL҅/P�')+!5q�0��Z�?`8F��~ݨ�{eͺ�1��3Ld�A~w<#���DPO��a_�ќr^F�̊L��W碜�T�|��З���6h����]b|���+R�|����fY����SbGү�V~�8B�/�����B���c�x/�t\'7r�������b��� ��8X��hD�	[��0���w5�#L�h���I1�^���#o�hE�+g�J�i��Va��%�A�|W�n���IVo��BQL��^J|!�b��z���I��*Ts\��±ʀ���X�C�Z]b*�K�������6��Φ�J�:Qt��_�\.>�l#���5H�F���y�XԕĎV$p"|E:�h#|)
o�R$K�ͥ�X�DX_0U8}2���B�0���A��]覦�E�h� ۈq�7��/��D)H��f���iQ�*}m����34��PD��Td��G�0�#�ncrO�0��	�
6�YrX�h�o���~���@�����c
y�M�as�7��t�KV�go�)Ne�E02 ���ғL�8�,����\���aJ�j!�4��' �|�~� �-10,�@���>�-V�� ������}�83��y�L�6L��J�S���r�7�|������z�8��o�;v>"}F���ĸ�R���U�mk;	�̕~t4�گL.���J7c���� ���ߘ��j`�$iǜ�G`��#rp���u���c���ܭ�:�P�k����C�)�\萘�%�d^WE�3����4�n~`�����˳�;,6j���f�����:�I��~C}��t��+8\��"Z���r��+�����2��y~��2�,h}�j��Y�s����ȗ�CF*p?��g��]�i o�P�>}nf|���2{�VG�މ?��gE$4#��2#[J.�����I��Q[7V���%xh��@j�BlX���nD�wmɠ0%��v�F�sx��b��G��XwhT��#&].S�{a�i�}��'��
[�*"a�d?#}W��3�9���u�@r��_���yd�f��i]2�xц�����}��P��r��z�p���:��,2�-�'%g�C9/��U35x�d�c�j��	�<��b/d��-Z�E�4���[�k�~b��Y�AK�iPzN��]��f�NM(�p�O`�_�Z�%��x�\�ނ�n�>-�:���ߺ�E\��[s������zu 2�-���#�`���3�9}��NA�(+��)E�>D� %p
s�}-�WVԞ*D��S4&�𶦛{�d�i>�ƕ�2���)�f���������/
����#7�m�U�ې�U7�5�>� �o8~��Rq�NG5K:��W�v�*��7�Ґ2��YݠX�l�uWj��ς|\�Ɨ	����z�;ⓥ����x���z��K-⨚�D��ؤ��V��Q�nǰ��.#~��_N���y>�Og�f�����׵*��DH�B�c@Z�:��|A��y�k�k��e�x���P��uRCO��@$�Rv��mI�.�"j��舺 }�� �Wob-&!��d߈�p�J>Bx$qq����ڐ;�RIB2:��t: �gp0�C�a/��� Pu��(�&�*��O�yh�ڈ>�����n9�`���o{d/���3�1<M�{-��VI0��eV����PM���
���L �-?�T�6>j���(gI, ����yc���Q�a�`�Gޜ��v�6�8F������*�N�eÄ�l�v���� !�~=����ƨ1�9m��n8$�ܿz��ّ�B��n a=��%CuښS����V)��'8��
���NTd���у�������q,��@f�D�(�%4����������f���˺������0�
H#˅l���br �bi�r�e��� )�$.��l|&�YD��?I[GF��L������T�DG�ۄќT��S�|�~]zA�����ԁ�JǣFq�9>��4��l�鈧�S�R�J=��p�0{��:�f�@�Y�9�SF�3��6s�^��ԜT���L�v�U�{����LT�,�R�ij���g]�D�{����k���~�K`�Hb:In�@�MH�ʦ/>�+�������E�X�gv�<6
��t�[��/NQ�,�bʜ��9-,�|�*i�rB3@�U�w�E�S�&����`���8IԘ:*	-�X7���E�� ��x���p/�����?�h�M�.L�^��6��&�[ZYQ�zu����h	���^}\K�O�v�+�mZz�&�8����!l"j�KOa�[`p��P������H��;����h��r$.qU|��=�@�u1H� Mk�ܛbjڰa@�p�4I��'W=�Y,R@��l�
�(�!���Fc97�fH��)�'g�^ť +
e�vX��e�=�����ۈ�T �D��i^	G� %E7��(��`�G��O?��2(�4�%*����F��wb��)]%uI���^ ���[�r6t� ��ݒk;����g.�Ei�ԑ=w,qI��P#<�M���&�?�����<����\�A���Q����7A�O���h�9��MT�%�������v���+��F�bC�-�n���O'��j��s~�\�!�HXd�RFb�\�z�Q �r.��������\ȗ��piˤrQ�%gw��h���G}�N�Ѿ��fӨ�����w��bF0�����j��^��ܑslP�U<��:�v$RL�픐���lc������p۵�H��<Jq�O��k����x�h&'���)��^��7gORE���\����k6$:Wi�����{TE�p��*c�l�q�_k�;�ˊBIH-� {A"�W�դS~q\�?��_"�z���2X,��˞T�'��� �k4�f���b��4A��]�\Y�j�Gc4�%�D��7Tt��!�b�i� �M�X
��ϭ�ǄI��X���s�nVHZ0������x�΃�Y��d-��|��5���տ'�'f��ĄɚE�����:H���ޢЬ9� wՅ`Y!p�|0;��:�F5�R�`*{�|K׬/��.��|�<�dھ?����� ٜ"ޚ<)����W�g�=�3�w��b�Ri��Q�@C�]=�j�_��H���\�YCsS}���Dʾ~�}�j;�g,��%�]d��3�tw��r�|ߊ�v	̝���>�ś3�n�mk/�Ą���v���Z5�\oѣR��y^U$�
R�#?�+�,
���FV<��`8����n�����s�U��LԺ�J��?b�9r��3�G�jsW����S�>�PX�J�Z�L���e�I-�E�e6�s��@T���U�s�_��.�"�l^*����!F�u�y�2Y��v$9M2"��:���|A��oXEXK�X���?X�κ0p O20���	���O-��W��Ц v*h���ۣ$$7<ܟ�l�Dd���/GͦQJ�Um�r���ѐ���4�KT�g(Gqd
#�Nrb��0J-:50�
��y�x=�Y��h�}�~��@��ѳ������<ZsrMhtZU��b��)�A�E����2����d,�w��E��&�J��|l�r6��]~��%1k�@��@�9��V�����$~��9���[�UL+�E�N�z��-�;����&�D sm���$�6��"��3�uU7��]\�g�amFZo	1�Q�o����.-����isc���{Ia���o̥d�$SP�B_��~P5�v�ք���F
����p�������ҫ��(���(�OȐ���߭E�r����'�
ny��L��Ȇsy;G�|�K�f��-��u��ZP~>cձ��V��u(\�7Zn�,r�?�f�ç$��֤��mH��h��oj_��4'����24�F%f�r����G��o#̞>XY]|�/��͈VBN݉t\�"1�4>^�2��wJ	_����er�[2�I�D1khs[@��B�i1���3��ɠ�����	���}x����=G�3cT/u"��t�.N��a���}�M���
֍)"<��dz��W�M3�&l�#�@-�z�Xwl��AGi��xl����Ę�ذ�P�w��u�:���,moO30�y(�2��so���N����@��c�{��~-��I�)��mQivސ�#�f=\�$G�Ѣ���Y���}atlf�&��;]���{��R��k�*G�<�g���@e�fp��K�ox允��(��a�
-���8"p,Ś����	���S4>��50��O/RZn߱
C��z��Z=NR�E_�!�^5�g.�s�����1�:�,� �Ĉt�lw�7ZmgCDl�}��|Zu�y~�A�s<_O�tX�hjZw	�(�c�����/��AC}�������f����Q�(W0F�S�7��Y&�B����$(�ݕ���Y�FĠ Em���,���Ķ�6F�)(&�M�������T�O�c"N��<��]��5H�����v0P��G�O�h�B�|����3ԣ�ܕD��34~��1p�i�n! �`jPC��j	_��O���N�"nz�HM.��63�D�|!�(ȼ�@*N{����o����8��ݪ�6�}��AH�9g~䐧tJ1|f������'�˅㔬�]z�➨�@��狵�?"=W�GP�r�(˲ME]%{"�<b/��o.���7��l��{�Zp�O��������DB�e���7ƌ�<������n��-�_ �#*D�Q����[���<���5����~� VC�8�	8b��s���t6�j�0���9�M�5�i�i�ހu���-�̤pm�%=w/�����şq/{&����DC���q��'RU�3�R��2 X���T�����g��b�� ���R֓��kdvG����)�|R�/ɽ�&Lo�V�0��sy<��:�߬�!�Qg��>���-�Z�g}�yC���_sK�|��X��S�[�T:.��lC�a]��/�7�w`��-5P�S��_ػ�Q��&UdM�o-5�?n��;`�/ۅ}9��E/QD֍�	��#��-��#�я�2/P����TO������o��d��?�k�d-\5�6�	�\-��Y*�d�ۊl�Ԣ��]��H���Y�n�_����nVFϥu�x�s&�-���2u���V/мw�nA��Sr5�
��!�ȝyIi9
����@z5,�EC#�:�a�ov�ȃ�^���.ZY�Ź��"}�}?8���kZS��g�ufͯ�o��R�E#�"����4�b��=��|3[F��oRf�t����mhF �J�IG
h�|��!@p6����G��@N�7>seIR?���!�v&�k#p�$W�M�TQ7����ɦ�0%�_ѭ�\#�4!��!@u}
4�������>�#C0��U\-�B:�!W��`]�kTf������]��q���Y�׆��XD/���n���8��;0�r.^�Y,��܉E<)!�h��d�tq�r����/�T�	vAvU�	>ܓ�Fl<�3l���O���k������z[�7�>؏e#��P�
�os3����9�(����GM�݄�����e��֦$H����.�(��*�&����S�ţ��$e�r�*�(R79j]6ƅ�?�dg��Z\�#(W��p��G��N�L"G�mN�+?5	�D����DO��<Y�P�7YpLL����=~�R����Ɨ� ����^��n�&�jj���2��3���+*�Ch�q.׍gr �����M���2xUX�E`�8ω����'�l "�(%e�0�e4�}��Zwk�;E7�������˟p�����y��(�EEZ�n���?lу�e���AE��ZJ��W��1�מ8=N��<�B���S2 Y���F�9�%�Hc��o��5��\ƁOSf/�F��[\̧\ʴ�/���| ���?��h[l�	�T�[%a.����cl��75��v�w|h��6�{��AY�K�ª� }5��L�����f�?�ߏj���'F���f��s���șs	R�KF�Ǌ�pxC?�ކ�m�$�������D�29쩑�G]��f����qm�O�2ڡ�?|�>jGG�ZB�x���;�_�K��@T�V(uz�;G�7�L.���S���,\b!��IeT�������懎'��3��~�K7$�!2"�fyŻ���r���������������C
�P߯&��"k��������;i�M�'Wl��s��(��-�XD�2�����b�3VCU%�'��f��k����D��z�0�1
b��{�Ug�tjx�Zg�<�(ݶ�I��6��$i���-z�w��'�?!~�/0��+�aO�Y��*	�����?��%�-�9��Ոv�����^�釴�.�����:�+"é�=��t�vv��[Hp�����j���q�PE�Z�H��o�'ԣ�}�Y��o��Є_��!�Xb�w4��C9*��7�4<�DI�b�ίo��onw��w����?W*�j�2#�<ூ�M�N�D�����w�C!|wB��nK�/Q����N�&�)�\��"z��D�s�����S��1O~��'��"@{u�Y^�ZR��Ѥ��Bۣ�"[���#z�2 �^�}�CЎp4�2�(J��u�Y�X�Z�0���mQ弓S�F����K�K�����J��>��}��a��A�̅�5�J�EvW�%V��_)k��7-�MK�w�U$�v�ç�l���+��_�n�d��ϱ���C9#;}�l�,l%�ւ������V�PX�Y�����4 ��{���������1(luZ
�B�X�l����q��Rz�uͧIu���{���8�(/�j�BM
@��lY��FO�%�k���oBv��Ud��g�Sщ��a�a[��j\���jN��x� 鴟?s&hg	��R[����[����l"�M5��v��h���,����Y�oX��<����5���wA�Ӗ��E琺^��%�j'᮸�a��s����=�8S�t��aa�HXI闇J�wף�=J�LK��@ۙ��Kv�5�ךC�.�.�L��0�:�ð��ī�!v=ǌ[��6���m���]�q�g�a��H���!��J*3���n��2J����H�4bÊ����a*��n�>Q�ˇ�bB�-o�̯n�>w�8��x��*�pM����<g�6۴}������|w̄B|^{�ɉ�)�XQ�ALm�mEB)!P��z��J����2�?c��Q��Z�qI�# ���j2*+��F,"�#ހ}�ß����g�w�8�Bٞ�+�����r}�������#��h��͗��r��_~<~��ׇݡS��:ͫΟw��L�����]y���h�
ܭai�aN�-_-������w0��A�o[��j�Mcq�d��6'���j�(���G"�[p�
�W�wcR�����:�t��;=!A�~+�5p�~�E�AT!>a: x��MR��b�=�5\7H�su
;���%���=ʉld/�Z�����{I��$�z`E.x�h�C��i(p����� �FK@$6+u�����6��k�~��ߏ��q6F(�h��B�6�
W��F�V~9�Tcl��T!�L���<�y���C+�P��&/!�O輥�0�=�;�������j-}��@�2��˥�/Yj1�ww�8/vo$���� �H�2E�>���D_�+���"n�7�:F�����ѥ�kƲVY�1�q�M �1�������Q�JG�<�Y�DG��6(+h<��ӝ3�~<4��欠��LB�A�J��@���o3�I��N��kVD��\٥N�ai@��eN���v�1�����{β	��kқW��qq%�tI��Nh
�p����}�­�K~:��c���_MQ�_Vs9�H�xF4��P�߂K����j��v"K���ue�`�N��@���\��!BR�׫`0��m�A��zN�� 3�
`�R�z�\�8I�Ga�v�� MEe�LԬP��u�#5����"L�z��:09��3|�������u�Ё:vJ�G��F(��Ol����<O�g��h�e@�@��\���}���O�a6T���<� �6!�)Nn�����\̪9[ag���Z�Ŷ�[Y�6�)�_n��H���'z�k����;��ܛ]iV�l���k��$�L��R����ΠU�̀�1�V��߇�8�5���Y�*���j�MK0�݁�J����0à���.�}��8f�j��� �|]'3s�����,�ȷ��<�	0_�H�	��rR'Y�3��i���V��5iS����`�Z6�֯^nc[ �8��k���l�����.��0�}�OVx[��Dki ���31|,�E|Ԛ����x�T�#P
�zTi��Y�B�e�PE��4
{&�8��wl��Ѡ�.Ғ~�7�e�R����,��M	�]L�;$�5�q���g����庚 �,���sI5�I����;���K����o�>"�����aJ���*J������t�k.m��W9:��8��u��ArKӊ1�X迃%O���!t�{��):������#�r��z��QH:F�(jH1�%��������dQ���YQ��_��[�`1��k2 ������\5GVL�Y8N>�Fr +v�Ԫ���3��4;�����Y��ZA5��@�	�]�L33��{�D曀�>jNy�@�5e���w�1,p���K{���E�����6�����b�XG�hX���~�7�T~.�Po�K�-�����.��%�@�9�|��Q�\�)��] �nk�u|)��f�A�@M�|ˋ�ZC/"����-���Q(���XXx�k��'M{.�J�[I�O��%�T�oP�q�IP��&_����id�Z)�VP��џ���sq�oh��١��u�A2WJ���+tC��V����0���<�Į�m�[�V������ɂ�-�M�0���1E����V9�;G�4h���=�H�)�<QB�ࣥ�#(]��]!䴂!�}xx��׏�w?��p�vB��5�G
%>�_�}��cBҤ�OvePN���W�#����
-,]o��[#�$��d��*��u�W���\������� ��1Yβ�a�d�9�	�;�e�^Պ��� *���1���v���,�S�j;��~B�a��b��7bЇ�j��4!i��&��Y��ņ]ɫ%[�P��JF&WaD==�Ȫ@7�	��rx��SiX�A��L�g�=�(�Zி�a@g��rh�,�y����#�f�̦]O�boC������o	'P�i���BZ�]��P�:qm1�^w��=�W&,H���ߙt ��Tk���~�0s��th�y&����x�8���W�T����!{Y=s���	\�Ťބ�LMOt�N����ҥy�
paq�E�;"����M�U7��u���'��ըE"���?����5�
�Y��4��0Uo�Q's�,یUy�N͸����a�f,�4X0��a����ʰ�w�?����{���Fv˶Ӛ`VR[H�� zw��o��m}sh�#���Z��K,�_㋉?��I�Q`�q-��3�[�"�MP��Lb�eU�&_�zCj����Bo��#:�p��ٻz�i/���ڰ��B����B/a}��!Tˍ$�,�U����D�|��^��F �
i��>*�&���AƢC.�!~�3���̔WԻ6ix�9���g;�%��=Cڿ�D4�Ə�ۨ�, ��'���P���s��CH��v�򕫛T��6J��^p�)P�g�uB�����KA�W:�|[�J[��;j�[��3!�E���������j6�B����N�X��߮��`m�X�2E���H���C�P�쀊��7߻���:ӊ1�`�p�S����z���J���Ź~y��]�BF6mm��p#�/��)�U����
�m��A����F��+;�X'�dwx�r��p�A��:�:�� ��8Ť1+�m������� �����2l<�X�����X�G�rm\��2�	C?�mj>= .G .��OR����_`���*�/X�T`�VuMm/G�HL��R�F�n��!�?I�\�yTv��_���gW�}3��q���T�!�\�f�V��tN�ry���F��$�Ȯ�����{�č����Z��}!��K�(��.:M�.F���&^��(��c-��ښe���~��b��C����jК!֧Vh`��G�`"0�vby�yǨ#�t�2w����
݉Vc�ޞ����%
��@�j����>JG"$�I��a��HNl�-\���w����
��^�[��zڅVBc|Mcd�Y�q���9&(Ғ�G}��pa�r`5c���|���u��t��=�d~��po��`A�ϓ�a�Y��Jl�x�=�m��0.�VrOS�������t�/aj ����{�M�$o(EE6��qp�vi=;�Pw��ݲ�ؖ$�c��?B��HP��.�~8*��*���
>6����#V�B��˅�i�!�~t��c
��Oqx��o��؊`y�Bz˾�P�	�ac�����G=昔��Ξ����xj��Y��2�D��;��)�j�Ŕwu��v� �XW ��J2�͗�liD$]�{w��=�R�������x���Qa�Y���lVT��
1YV���h�Q��ncG#��Y��9�S�e+#B��Z�3�މ4��������V�<��BŨ@����h�3 �
�)�a���fD��WʬNrN@�,HeiF����1��C�|�{i[n�?e����,~�.��E^kh�ߚ�w��!�b��4�K٠>�=��߆�����:r9�ߑx�C�K5���;��'���v� o�e�'�N�@������ޕv�I���OK:ě�!��C_N�6s38m�`�:�Lb#��eI�q(��&b (b���Q��Ru���E��_͕�5:��x��ǐ<��u�N�:чEGT��FC��O畎г�iG�g*#'Ӯѳ�]}\M7�}�}�Od��T��w~���!�)I�A�P(z\���v78�L�5�$�*@�d��) f!n�F�q
�z-�B�OeW��e��?�ge������a����3J�����U��7�s��QKp���~52GR��SaϢj�"Kݘ�|�ߢDׯ�텮������8�ڻjR�bϢ�|X2��QV�̱��GHշ]ȩ�1�	kzH2�l��H�Rk������i�;Vs�H5D���
~�U�j�
�c�&H�S��kd�l[Bh��)�0��zO��Mxo�Ȯ8k��y�t8��nm�|��"EwW�B�@x�6��>if
n��i�y��}�K��E���
�g��p�{�z����h��Ш7�G��M_�p�,��M$�����$�W�q�s���N��(�����,�)ю#C�Ļm����QG��d�#���>}r�ˀ�J �z�D����X���k�GQ�Rg@�&����\"����X���%�aO�4g��t��RK�;����rw�Z��(:�?��R���r ��j�~ ��k����:�D��R�L�Ր�`!��#�pמ��<���-E١
�C3Ha��$��� �����/�6���7k]`�����SF1�<L���d�VL-�Q�n�_`�Y��k�j�7f�Q��a[�{$-+���I��1M�P7i�Gf��7�SVT�3�k���5!\KaW���%Y�ן�3���H�� �K.y���֦Ơ|���nmt.��^�е�&��k�P��2͏����ۼhZn���S��v�p�������i��=��  @Ҙv�u̝ܦ���X���s����WZ����B�"�8|\���2�Z��Kgr�f%o�:�6�"u����4	׀ӕ�|�E��SJo�F�t�x��ž� �kI�h
k?r|��!�}��V��_
)֘| 7�l8Ivvq�B���s�YK#Ȕ�$���֬Wy�J�����!.q0}m��#ٜT� ��uq[�4�Z���>�0KW�U��zv!Y����k����RTµ;<��؉�i�:�޹iX�R��@��T"ۜN�;��-��(�
���c�*��@�)y��h�����rE��䯉�¤v�>U.��>4�ӟ�uV���P�]���V�݋Qi�e�>0�\#;��P��o�ʁ�tJ�9��J*M�����
��:�e���|���*"��@^*�v��)�����lj�e /*0p]7���6{? ���
���{ƈW��y���m�LzQ'm��?�	�D8����ųДM�j&�ڏPL��$�0k�ު���l���?oZ��^7���~@j�$��J�0�U�#R6�����h���� �}�>�'�+iHx��ME���'Sx�B�X} z�H%��^������ `Z�A6;���]c�,���ս�Bc���(鈷Z'ԿPl)(�մ�_Kղ���&����/%g8����w��BJ$K��$�Y%8F,"%<����o��������.�Sn0�Ҟ[��7\"�1����k�$ F�?p�}h�	B�[}�D�+�ܭr3l߆5��v��h9\�i@h��s6Y<�z�թ�=��5���t�p$e׆�F�7��B�G'�F8Ծ@s�,e)��=/�0�)5u\a3B��]O��#�t�=#e)��fN�^�9��v���W���k�~.�!R�ͅ\:�cÍ���z��5��xX|#p��0qa`�X�Q�T$�U��j0�'B~U}Z�焲���.6�����B?���bj�̞~���c�-���L��vC�uq�y��˛�PG�~PTܧ4T����H��k����|^j�@�ɘ%�2��v9��Q߇j�&|w�vǴ �s O�2��y�FצDu�Gド��;�᭏D&�M�q^\��R���Y��iP���}1Z�,�؋���|����G��Y|��PYw+��(�+��3ܡ 4E:���ˤ������?�,@]H���o3�D���A��ٜ�DpJ��aN4�@;.e�R���͢1\r�0�{&�C������f�k�"��hb)ɚ�����K�E�KּH��}6����D�9Nx����R݂���,���r6����e'�N�/Z�H���w�st~�/)�#�ź��[p�N���3��`�q�I����T�I,Hқ��F ���Vլ���u���
��z/>��{�:�R�����Q�F �u<��:�sG�ęF�7HO�M%�0c�d@�g��0����b\ꠉ}�OA��Tn�K��n���5)���M�s\$`���nBͲ���G�I!�)]��n���zT�PU;�U��;����.������|6��b16��U�U�yQ�ݮ�>m�*v�5o�����`L7�jG�Kׄ~�ٖz��ů��E��v�դ$8o��jo� �_,-|�ޘˉ*�i�Q�s��:[����	�8?H����Rh��ċE�iTVP�/5�9�#�"i�}���h��tc^����ek��l؊��\>�Y0�O�1x�����k�8��񭶽��R|i�E��G�?�MxI�1�{H^
K~�iҚ�L�״�E���
� ��A��GWm��u�ꏔ7H��Ymc�,Y��Ma?���`$+Tmq��ݰ����/d���,c`o�n3��ٷ"0/����p��_�'���W��s��/=(3,I�nU�a�)i�~/�E`�-Tq�P���ͩ�6���r�Sv���������.����:1:�c�æq�a8�v��[%���,���#����^�q0���W��HS�o,)Ԁ�ĝ�+ތ���AZ��~��b���K��*����mk���b���o`8mn��w�Y��.�*'���<]1p�j1��H��aw�;�|]��Y�_n�Q{`���ބ���)W�W��� ���Z�o?��jQ���):�F7���µ���GU�qY(ڞ�+�Ϊ f3qP=4z���١�:_�����@����܅-3��	��'9��I$D�S#��cN�,�@�=|e�L��cL1D�B��m{��,$��Ҩ�B��d�`3z�Ŗh��w�����STg�/K���/�4���L����Y�9潲xO���W`�X�s���ۢ��z�eI��N��ӯ�cZ��R�(��L{}�Z�Z���OpN���3j-U`���V�	�I!���c�> ���y!�%�uזּ�-S��\���Sh:�8�*+���H��guQ��:�@�GFwnFu4�OY���eq�9�g\�Ek��M��\?�A}=�O�UXT�m[�iH��*�)�����\yp�l�D��瘑�ܚ���)r�n��2�cOWzI��?o�_�m}�*l#��W�x����������t�H�	U�Ʊe���"�<��5dN	�FA��>�j�4UKL-��M���hW�ݨ
���շj�^8�CjD����y�|����Aľ>8�ysH��Y�����	]0JHd�(C�Ro��{i�x�V後5�o����ސ���#�ּ��c�W�"�k}��l&p�^�[��0��Oc_$xr��]kV�*�&�s�`��|ޙE�����Ix���pܩ
���iG���o�ٳL;E��
����/�� L�D��R?�ҿ��7�S��{�"@p,�jNMV$9?�$`�3q�j�4�"�M��L�,�X��̏�6�O�tƶ�C�e疀%��
>/��r8J2��Ӷ�U�s��.�k�Ks��񢷽�v��,�����wX�Xu�a%|y`�f}�~Pk�6���-����r�.�}�t:s)�����y�r���\�~RA�ݼ8q�X:�ښ���L%V��4�Ɣ�z�����i�fŖٓ�5u^aS�"�{���f�9���&�H�c<y���vO�+]a�.���3���N�;`1Q<J��z��-� ����e*H�<M�(3�T-���數lds�i�Ub��CSS���4:�r,y�!�d���v��7(0�7bĽS�S��t(d���z��ݴ�O�i�w��[jU�{@[�p��fYJ������a�YN�LA-G��h��wM9��ڇ��y{[_ٰڰ�Ac6Sd�S��E8�AZ9(��*G��p,����cX)��g�����t=qf='�
~� kp:������Z2�a R�G�[�#�=�Yj����1�����p��Ք��Z/�����{�b$:ޗEa���G	�8i�������)��_$����C�Ѷ�̕���~�����U7�M6����A�B-T� ��_�~���c���Z���<أ�y�6�Iz6P� ��W�ܕ!	��z�){ؙ���0|j3r���L2T�d4G��7Yj��xw@ZQv�v��s rD2�I�4�CD#��񅽌ijD�}�LH���C�+D���YɅ.כ�Ӎ&1H���t��Sޯ�ρG��Y�>q��q�+�υ���3�@4��I�2��˒ʹ�GC���W@���ժ�3�|��o��xD^M�b�N�h�@i�#e�Z��|ӫ1}��^-�{6��o5�a����v�Y*��Л�h�r���C�����?�KD��ܰ
���er��%~9?�x��v�V����Z���� ��b�e���N
Ce�6�%���-�]#�vc*�s�L��c�NT�3�3/`����̨�2I���|Ќ =��ͬ���u�M,�x_���ŵ���f:6�K2���Ua�p�˷|�Ado�<��R�= ��Մ�������ȴ�0t�
y5�8:�5S��e�Q�{�>&�T3�gV��y<�־Ή�K�Vʱ��S&��TӼ�W���:�<��7�6T`�8����Sg�!�T U�K1�d&/�-.:Sn���`��I�l#��X�JQ�v��xܛ��s-�$����k��Qٛ�)�P���zA����Ԯ~k�]��>�5"o|��5�w�Y㖜��G��d$��Q����礝�B�n���~���q�4&��ɳ1j�2΄d��D˼�;<n�'�SK�̀4#�������i����F�@�����[�3�ֈ�ȼp]�X�ZҶF��e�"6<�������ZlB@gS�f&U[o. ��ނ("�Ud��m�4�G��Vz|lb����o��t<vp�&dE e�gI@�5
,��|�!��T������7�I	s�����#�Z�#�]$����@���L螽��E�0^([���#�(�A��u�s�4��B��9q>�ˠ0,��U��»��!�cG��	k-�Q����v�XϪ�5�j�\��g�X������Q���}��e�0���(���,*�ۏE`5<S��� N�w8ϥJ��w���|ʘ��u�����QqTc~?քY��)����Ɩ��l���)i?���Q�Q�����#�*@��\�+��,�7��l���h�ߒ/D×8Rf�
�8+G��g��}�G�<O�r�3F�n�8W��]A ��N)H�⒈�s}y6E 1��M�]i��~i�ߔ��`뒘hx���}���CC�W����j�ߡ6���g<1Y��p�����z���뗑Ѿ�~_�]��F����������Ϥ��+e 
ߢ���Ԕt�yF <�+,dX�w��(��Ak8� Fq6g��Tt��W��m�dڮWR/�fE�=��2R쥑�J�����mO�mB��2���?U�X>c�GdeȱA��_�,D�㏫�-T�usD�G�ILg杙�� إ�!�~���\Tx��2�栩��#�n����!�!�f2�1���.r�T������D̮CU���Z���ش�h���5T��J��1x�t9sM`���.(�/�m��-��v�K��$	�b�S�C�0,կ�ݚ�T������v��,0�S�b�B�����t����q�2�ݯ�T��~�]�bpf@���I�J��*����a���NR%}-���Jbw�����g^��#[�Ibګ]!cb9#d�׋��c�(��G#�p�׀�-�c�WU�"����5�t���=��~,`�p��s�������a��/�b� ���#=���8W��d�|�9aߘ>���*|/������W{Jk�$���E\�t�t6�q�i��q�v�!�/�G<$W<l�>$�s�6�P��~��;�Pּ��6Ge�É4qB(��k����~��c-�U�5ׯM_-�>o�y���ˤ��PA\u�
��8>�g`��>�O�4�t���j�ͅ��S�26�5ߕ���Ⱥj2AwۍZv�"��; -��2��a����D�H��,=�	)�x�R��΄����F�~���Y�l^��n�!1C�LQ�$�lA��P�i%�j�P�y*�f�IE�1�.,������?�6��sos$�õ({}�|��.!��@�$E_�_��P')H�{fH~ 9�?ʹ�����U�g������z������ *�yi>+��1i�2ɗU�f�2�A'��:&\3	/������3��G�� �w-�ܰ <��]Ԥ�/y�S4��D]��:�	�G��q��<��(�N�=Ά	���������%�	eR�N	�&ێ��Z����J����ۖ���{!n��X�ǧB��۽c�<�����h��50-��,E�v���0��i���F�iu����3J7��+�����������N� -��m��BDJ���k��\=z��N��i�4ŀ�͗�7�����w&(�5^q{�2�cf�kT^I�>!6�AKm����_5��q���K	�CY��LQ�K ��L"p��ڟ㑍�*f�/���XS D����K������2�\�I;%ܮzfC��X�F!}�|B�BBXI_ֲ
fx�C��%σi�Z���ף�T���. ����:����r��c1���_-����[����QE#��٘�����z1��'Y�9KD}ӆCf~���-����Љ�M��4*9���9���f"w$Kr��x��ld|�:�au|ʳ:�E8�&�wyĽ���`E�������_峓PR�0)�|�N>������1R!7c_�A�^�Jg`Э�O9pfڢ,��,0�˃�t8��)B�gu�_l%*X�.�#�kA&#d���t
�8\P;��b��y�i/�4�Au>=� j���P��:����ɀ������t���v�(�EɹT|c2��!wmBz!,������o6�wk(�����r��$��s#��J��C}z��>A]�����|�慈��ho0��db��,�}��t�:�Ga��d�y�������Lĸ?t�@����hLJ\Qռ��a��Na-�2�R��ww���D��s1�[I����#cqŏd�А�W��b���TqOD?�b�&ebi7�A<�[�u��Ȍ�'a���e��D9K��d��]"��~BC������'���V��;㋓}bn٥�u-7�9%��������Odϫ���`>3�bg����;p���=��#��qšș�9��v�mYT#��T�O�JR�es3us��4Y"���e�=��VQ�djJ ��RXηe.�dx!3�$����>V��1�c�h�����g0]�y>��:𱮬g�Q)��>��0����A�g?��yE�y���KK$��iS��oT|�u Y�#r��x7�`���}S�?Z�����!�d�-7@Gn��7`�W��XC��tQ��}��!	��5-�#�������8��g�V�q�����C�'�h�ݦgk�V��\�5�Vg�}o�)Y��+����U��c�XXй]�Ӧp����n��^�gHB�z̶&ڸ��z�e27��XռR�~nô�S4��O��Χ��wi�z����@����Q��Z͕<�NֱE/�sC��0�Z[o��,/�"�:��啟g�Z���g��Rf��&o�Q����n"�w��Q4�;��|��]�G
!oT�mt�q���� NG�IIW#
U��|��!�E����IM���^7 *I ɗ�,J��x��M#r,�$�3�ց�����v� �0�G��o�#�>���k�u��4p�-���>Ծ�0uhU|b�D&x!C���Q!k�S����������n׈o�X����j����7���;r�����=t������!)��&hn^w�vR9r/�k�6;���vC�U�>^����5/���r	�)����2���^�O+E>Z#���P���o�x�����9T�D��	�c"��4�H0Je�_f�f�:�T����6*�^؉�Z�5q��)�e��
*�^7��6�g�?�~7���/��QWg|��/����TL�Z�m?7D"	d��S��������y&�L�l+�c��T���V|y�i-�7m��?^!�+�]lj,�m��� �u�'�M�H��_�b!��x� ���6(�ՂZx�:�E���]���i�S �����}�&'�L\Ъ���.V��Hg��mS���:��;�LڬK�/J����O��w8�A�qLm+�QB���}���<6�]9y�F<��8�p]��k���)o�<��z�sd)ͫʏ���c��崿��w�`:�#��N���뤏�!C�~��m��-	��EZ�`�1`��p�G���gSz/���7�8�e~�%�]ܮ�F��Q��!���ֿ�v���$�
j����=��\�F'gq+��X��1w� 栯?|A���gZ�]�[���>V�mND���*���Ť��2�WV�%��*Q�T�~m	k�2:)�?�v�>�&�GM&���La�
_�_m�zuq��|t�TM*}u��*GBc�L�(���` ،K�!c��⩬T����5�����J+��޺�s8!�]rf�l��a.Jr��֕���X�J
������q�X�.�GH�
<S�x4怛 �MgZ�{p��V1�!m-Y��@B�K' b7�C�tJ�v�ĚT.M�C���R�.��0�b�<�ǵ6�t�3K�'�����(�����@.ww�@�:�����J�)��6ӎa�aN��Z-)g$�r�w� ~���mΫ�[�Z��c�
^d��'��J����(�G���pNB;��c�T�I�ܵ�>t�܅=ɖ~��p\ޗ����
�a�>��iAȫ���=T��z��!�t��7��e�+�1��/n�܏�{�E�$\*�E���E���Gyi�kh�]���M�8���Q$��ɥ����VM�wn~�w�7ɛ�Lg@6�E���B��i˲�t��S~�Hoc�P��*/��^���c�yc9A��ܓPh������\�.^���iػ��9	`j�V'���2=�^�mD����jٮ�wb��v��A�� T2�����[D��~��aӌ����p��Є����Mݪn[|Yk���9����V1�C,L�z�5�L�0j�G0�YR*9���V+,��{�R3,�x4�Z��T$����������@���7��3M����8�)D��-�NhL�@�P�e��_��1_L��Υ{v�g_��Cj��ٚ޻�k�r�h�9F��8�.'N�j3�K&uu�*@�l�J�g���9al�x�̍�������|"�ϡ�M١ed�RN,ꃯ��	�ǖf��1��1��؛�Ȝ�p�N8�3E!`GP�-g�#I|D��K@ �B���I����uII��Zϑ��1��"��:��T�E"i4�c��u��:MHGAF�ӐOt�ЀS��:�g7���1���\:C}h�O�k�T�: ����ީ�)�&���\tR���@�QӶ��q�)�L�nU?y�^Pgz�0�ok�26���sK�B������K�ȕ�0?W`�j�c��U0XM�2n���
��hzX�5��̢�+��jW�K'Y�)�W�h�N��
��T:�%�(8�lFj�{?ϯP'|��?Ĺk���?����>��?	�b{H?�]�c �R�i����iWp�V���5��s���V��Y�Wɏc�O��D�k8�l(KpO'�6nB0R[VO���x aU]�k��A��۬�|�E$�+��{�x�dʝ�T
��ib|8��.�'i�E7�
#	>�S�I���Sp�m%��:J7��t���؃��k,�Y�M����ص${Tiq;
Z�&�@�B3�,���Ƃ�񯡝��M�����q�[���>�
��m�_J����qdrԎOǆ���k�%l����X��L���>�2��X�V�%�N�A��pr�����(�H(r�G�ј�:�Ih��y����rM"W��~��������:&F��gL`������_���]�́>���O�P0a��"=����Q9P��&�� ~z��y�O�\Xa�f����t3�?ϲ�-;#�<e�0�%�x��� L�#�0H�N�탍;�xi�N��tL:���-V���H(��m4�a��]9?��a�ÃxkD�Q�����>fb�%��x�p�����\7�5�SR5����{��ͣ�@�	��~���v� 5p���ӝM��h�e��G$46���"�.T�� ��EZ{@��;�Mz���[�V�.WB����a���"U�2��Hn,�zP1��b�\��+�"m�R����j�ǧ3�̣<y��X�T��j�b9Ԅ��y"�sfͷ�E��$.$h���� �7rE�.�sg5�#K{u��|MF.e;d�@�s��"�	6��˜��(�5vƸ
��'�wʜ�?琜��$Z���A����ũ����Hr����]��@A�~g:&>����=�s�E�	a��r�=8SNRH�1~�q�8�����ȿ��@9�r��=�^d����#����k����#%���Ĺ�N�SPv�>�{��Z�	����q�z�^|�=n?}&qS��xn��d]��Ukp;��}�s�`�tѪ&�i0}68zW�W'��M�6!��s�߸��<����:���M�a�@�W�k������TqW�Zڀ���~y�Mo %\��:��R'��{����X� ?wI1캞 �~J�4���U�.
'x�{,���y�'�vӑ�h���4��_���~�3���`����F���_DlR��j�c�ܣ J�8��sM��W������$�������Nɶ`-P�-5|X�@�ݵ��n���S�*#���zH��ٽ:B��H#,h�'�z�g���I�x�����9�fBt�a��)�TP����n͜mQ�Pm�����������X� �IIi�H*��f��xgA+�N.��;f���S�W�+�i������;��)���C��gD�m��<ۍj���Y'�Pl�c����C�*��w��.Tieϒ�^�IfPZ�Zu�����V�A�	�Wb�/
�:ǈ�������|�K�U��x�R���((��%�U��[s�'?�%=�����\�VIXl�������jϒP&�|g����:�PZWu�x�^3����]��,0����&"�̼�(�,� n�^O��C>0�pb^����#�Y}i�A�0zu��Kb��!�t	(��1�����3%}J���\k)�� �ǠbJ��W�XV�x�_W���%�u��Yw`]�$�/ Õ��l���5_�dsH�;}J��9QB��Z�lӋ~DcH�!���
�����'�&�9u�~"u��?l��j������	�^�6؏����� K~V���.�.��j	���$��|PD[���V�ٲ7z���a�'��Zx�H���zxj�ߊ��B+��E�z0������Ϫ��a���>X*ʌ��5�b�H�Ԭ�yJ�f��1E��.L�	��wP�_��V��s�ߣ�㥕{�� |/�9.8��A�/@�(�_����)h�{�\� YJ/�Իތ�
,U�����\���iԭ��Y ^_y�������R	|UĪ(R`6'��&|�P/<7���"�SɡG�P��������<��4]��/�*'4���dYf�ZZ�	��hʑ��<��
�nIaΦ�P��&ږ�)���Ţ	��&N)$�ۮψZ��6���!J��׹{A.��Y�Ǌ���	�\�c��hgy5Pnl��p���G�PzI��;��	$��ik�oNJWy�+#J�����܍a��oY�@=���{#��J������\]���n>[��2�Š�Ǘ�k�(C���C(�u3q�[x2�+��� =I��6ȕ�5#z���_U3qq��k��C>Ek�l�IK@XL,c�����%J�/��Xs,w��eK��3�%Ü�;N�\��%�Rfc�X�r.}-��b�`I&���*�~�cD[%�G��֢��$��tz��N�
�6q�Zo���)Ē�&cQ;w��4-����{��:�Q;�]���ٸ�ٚ�x���8&�Y_�}��f�#�M������\�=��*Y�s��m��ҁ�fB3K��qx71w��,��Z�a���Z֘8��������B����e��&���)��XR����ina�s���LRA?�_�M^�g�de�oQ���L$�,8�1ˣ/�tXJ��I��g���lEb(�N������AF���,`t*B�|�[���!��Ι$K/��A�"�@Ң�@Ò�*������9�%����.�������(�ѷ��d�,w2���ymbw,�����6�=(��M .��eC�u�!L`c4-r��J�E��-���!�P>��!�w�T�i�M=a3f���gN��Ex>��8��XP!Ҟ!`|M˩C#j��w�!s��`4�n��SM��F6S�z�O��%;{�f������b�o6y���puHb��g씐y�1��#�m	�!��՝>q���]����:������K�"��,��k?�D��m]w�:"f��/��G.���73�4�|F��,��O͏��ү��~�D�w�e��l72<"�z��ɘ���'���ҵKD�9����֭�ϵ�NB��Nb�և���pVՐ����`b�����?��e�S�<���=!�����h���W���Y�-�p�-[=I���q���ң�&���#����(��韑�R��3�Õń�y� �����~��Ο�lf +`<R����gd��';���fP͎�e���D��4��(��0�;y��r:@�Ϭ`5�Qy>9>�3'M��,��g�*y�㘾G��K�B*�jj�S���T��Op�z�s��M�%7V�L`X�G�GS@�k�M'ԥd7d_�{-�*�nO��`VY�%��1,�Qֆf�ۇ�5��-^��J{����
@�g݈I����Y��-1�kM+�6�s5�~�[ю�YaY��R����/�:������8��t�;�n�.Ϸh�����&*-�����2�捻�� ���Dn[S�Ҁj�۟ ���oiK(��Ѩ�@ ��G`�Wߕ����Z��U)��CZ��|�|�"O�B���'Z�g���f߱�o�����"�l��~�4����TU|֝��o���t5���?�� ���I��
��/|_MO!RV1�F"����S�7P�Ip���|��j�Ú��#�� $�%�&�jL��П[�0�u�ѿ��#�@��:��u��04�w���>$�#0Ŏ�ѝ�b�n}�j�A��/b;Y����y�L�f	���9ĝ�h�f���8E�E��[[�?�,V�cBdR߽�@����E(�r�Gd��p(1\cTq
���P��;6t��s=#��~m�p6�7��-V��a|UV�C+�����=�{�yNv�C��Dڜ����i���/�����-{�C$6�{E�n���R�R�i��Өw����򲈕S$���ɿ�!�0"��~u�Q\�]66�o���B�8U�t�̈R)~�c.�Z�V�z��L؟��y}C`�E*�P�����ƥ��p�6�ؕ}�S��j/^�ɂ��2/{�n���Bjs^�w<S�v1����m �k)2�`�����D�g�m،e�����HT�[���'�;�P$YŇ�S����1�5��
��}��
^�GJ|�Y�|��:o�+�|S���83��,4/5��.RD����C�k):Y@��V�Q�33��ո����WD�3�^�9N�|@eDe��x'i1���ZpW{��M�a4������ם�ժ���+zhLȚ����H~d��m�K��}�y����a>�g�9;�(x���R�X���q�V�Ι8����j�e��vN:����!E�.�q�\�A� �)���fÊ<Y�����[ �;����A�an|	��5N�E��#,3Z���K��J&g��fw{֛\�=�ǜ���p@�q�I��h\�5E"��Q?j��O��%������~o�>�%�t}KJLR�+��ýֆn���7�=���U�"�BXxmaJ���� c\��w�Ct��"0ŵ�<��M�}[���(���q��2�f� ��I�6}\3�����_�U�qO�`�@1jC�vJ�K��L�<���CO�F0h�/�L�X�����K�n�zj)�0�\��.%16�f8YkX^�},@9�l'I{Ê�Y�����%$������M����a�Jr�f�òOKlI��ǁvc&��.�$-�<��0N�TqUQ0�ɐ��w��I��фzJ�����}Hځf�I�����Tl��S1���!*n�ֳnw��'��f7~K'��xl�a�>�ϡ�a�8ó�U8	��k��r�ȍ�κ#^�-N��Rax��X
c�+��������R��_<UZ^.�g5K�� �{����,m���x�Pt��:�^-�gJPl��u�C��� ��A{Wfƣ9t����d��v�pΎ(Y/K��A����N"7l���hX]>W���w�����-�k]('m���n���e��mWd�,��2�K_a6���(m�uM}(�F���<���c����O������cr4�B�8��!!P��M�c0��"5����3;K
���)�ZQm���B�P˙!�[�`�:�x�ejp},ܖ��uR�n��$M�36�4{�#1ꩯ�[�{�K��=��(��ěb6n��8VH�C<g�:��b1�(��"�\v��Ւj$�S�']����د��8�"DuЁ.�T�9^��Y��]�D�";7�/�D.Ǹe7����QZ�!�Ob���w��m,D\�ge�Hl7�� <wO4��d��qІ�7Ҋ�D�FK�Ƀ��b#�#dݞ�`�kFj��V�H��P�wb����zcp�}��Eh�'���8Ŀ�*�:mQ�zq����`�q�-K�����/�j����@��a/�z�A �R�Bʺ>#�p��z:�����N�H�Z�5���B�����ZT�}�7��0@��&�5�������; �z*i��O*iW��pA�h.�:A�_���w�W�җi����ki;��\�� qCuCgD X�!f��c�*;�A'��P���C�6��qh���bT?,e��^��Pp��u}ɑ��A��*�m�]����֡��Y�R9��뉬xM$F�%6�$���[�VP0V1%yd������In����qщ������4���#����Qu6 ^I ݿW���h���2����C"��.��,۬v!I^eǘC�p�Y��lms�9A�YSŧ����0�A�1+����
;v�=�E��0�	�;J����0����� �]<Jq�W��)V���_����{Z-!w6��$a�Z��M*l�1J�o_z��d��e�Qs���*9�W��/Bl霳�������b�6�'�U�9�~/~x��Ԋ˷�x��]#����4&��%/�FL� a�F�g�.y�2��4�e���$��d�_�. �� "EX]�*��8z|q[vY��Z����G���eǾ��)�^�=H��z|J���}�F�+~���~r��;���}l�O���eMX��o���Cb+��԰�(y΍<f�m�E��.PYn�8�A�c^��ڇ�s��D�g�O{��|���.<���f3@�efޫ���c/ur8�j_�gD!�?��$�н��k���>�L-���ٗ��s��U���Hm@s�ZR�^����u�jk�#�^w�t}k�,���eӸ�D�N�D e��������x���E���Pޒ͋����f r%f������
Z؄1;�|jͦ�咃~��QuE���i���~(��YZ0Y¿>�lr��&��"x��[���{X��V`�8Z18�uҁ�S�B�(�4�ZY�٩F�9�%M��ho(�r�O���B�dS�:��Gn�[}]�\jq�"��� �*�?�Ph<�"	�6}[F�O�I8��l�o5Q�:vZ�h�Xk������nY%c�����f�5Tq��w������I��U� X�K�'Ǚ���Psh����y=�t������a<M��.�?�=�����h�2�z��˘�"(v��׀:G�Z.U���Vf�:���V�$��vc?[Ո����,���;Ѓ:�q��<�[H��_��0-T�����<�������.IbiM/��Ύ*��>w�!�q-�b�8Dot�n��5wMA����u*�:Z���<q��gℱp���wr�c|Ğ�ɯ�p(�Q+Px�Ǆ�x�)�H������
�;?I�Q�g��׵�#&�C�PP,+���,��$ަ��Å+����>��8;XGل�:+9Ľ�a�n}��	<��,��F��X8�X�]���ʂ�d)Bjw���:s�M������`�ח�N����Np�`�"��/��'�Ǥ��~C=��� �s!���[��ډ�1���p_2\����z�����Y��K�~��]���F֗;��ﶹ�V��ɍËem�
}�ޓY䒔n��FZ�+�Y�XǴ`w"�b�gA�Ta��^�0��厣Ԥ���mAJ��Q�㠠P�ŷ�/2���'�E����?m���2���?��N>ݮ�G��)ȫ%h�=R�_ ��h����~5T �u�3G���La$�������!V�gfV��?"�������0�4�����c�>�8�0ĆUl�W�R�!tƊpkkd��
k��m)Iρ}4�!:זlPXT\f��]]�z���;@�H�>���ܙ��)1��h�V��T�r�Ai�����dnTvQa�U�_*>�L�V=�C_�������b�y�	v����>��#���P��o���,��9����W��ݔ+~��r�e�뽦4�����&�8��*�A��K������$�eؕ�*譇7I�C6֎+?؏s�����3W�W��������kL2~�m^��?ED�D�)W�T��	z�P��'6|-&[ճ��F2�2��񮕼�Sn���S-S��3�y�	�+�xuit����@usIy>� �t�U��"�&�IŤ쩮>���B:!˽n��Y��~��mc?���Ư��k��y-��E�P�a^����"�~��T2��H���Y��w�j���S��2\�9��,�j�1�w���v�z�L� �Y2��"KDP�u㾟��ֽi��թ���,����xY��Q�2��@��1U#CW�m�������G[�Y݌U����+[]��&��37��4 ��Č�tn�z�@�f���|3Xv<�a�Å���D�%�'�NSv9@ַ�e��)*+1�C�K�{��I�T��.O��d[]�f�~�}O(h�:�㖹�Y���EK[�uݓ���@�rBI9,�7xq������g(���`�ɐt�X��eϯ�N��H��+k�R���w��^:��� �S���N~�3p��`�/r��-�O��I'�J�)�� `Z�����#9Nuԃ�E[d�;���z:�z����%�G�����u�b:	��G�;�F{�gO�-����?gby)���!n\��}0!O��rT):������	0�)�W�ꈤ'\��G��5�����m�%�b��hY)8�n@������zOO�z_T���V�)�0�Tȟ�����}Y����kkH��5NU��̩�݉	�����'5j���-��\j"*�KR˴ݴ�y�S���#�a����00!8*�Oj�om�ڽ|��Qf��M>�J��E�O��	��Hj�M��m�R��Y�&�i�pV��U5|F�><F� ����B��c�1�EkkC�l�"���a̛0�~�O�.�xN2� �kkp��X��9|�u�E�X��z�hx䱭�vK\
��i�ɝҵ)-�R��E��]
+�������ح���)7�=^�샨��,��kM\���Z$��q;�:p��˝��-�@,�����-Ѿ�����Ԇ��:����R�E>�F�˸C�J8���|�����o�M�kf��L۷C���� 灔���=�rX�ʿ%�P�l=߭D�G�s�e��r�5?���:����/�?�=r8����+~X��֋�:�}���L���ϔS҇��y���%��=���!�{1*a�F"(��E#D9���&�.��ڟ�D^qOŃ�a�s���A�3�v�T̿;&}�<�~���Ϣ�+� ��`��H�b���;ϭg���U�M��Le��J�Vo��Hs>�m�i��(�9�%ɢ,ă��L-o�ұ���,8��d�p�AբL��o����RS=��"�He�j�!��b��AF�+�e������a���
Q���j���mG�;Vp���]n��-���3U�����r�?_���0V�p;��|h5TڇH������Q�&�(�]��HA��>}}�>���sk��\�;V�BD����X
B��}�lB��O�oNqN�W�B]؃�
��ob	���/!�dbm%��v�Wۿu\I&��G��K1��l#�d$�	�i���Ƭ�m��6�fT�1CX�v��g��%�ݠN���͘��)����y�2�v��h���i��B�ʐ�6]�-��A��N&$�5��=VN�k=�	G�<rcΪS���WeתWm���>�%荿!@��KrS������.�#��"�ST�-���ğ���.P�y}���Z��f̻�gq8oW^�|=T��&����b�����~k��Ix�s§Ct���&{㾆8��$W�2��1b!FͰs#�����ŏ���bM����&.i�j��D	 5X�q=3(�&���B�M�yBF��4�J��'�t���j���;:?�z��Z��d�d41�U:AX'�ߋ,f0 y�c̸ܨ���y�q��4����,x��#�d��n���$�ƒ��b�F��.�R&�l�+N�܉pM���&s�q��}Β��rb��놉
�l�tz0`&8-�즾ڵ����N(�И]�LW������5CP�M���'����3������� �]�Y=9ԖEY!�H`�������j��ܜx��;�3n7wM[��6 �'��#�5����Ґ{Wq�\�7�)�
�i6t���E�H,lg,�g��/.1i����o����՘����]��U^�"�h�wu"�Vہt��?��>r]2y�"���/��.��7n�q�J��'/O(����ʛ�ךDb��e��R7S�<�-��?�7X�l�7�Џ0Dn�~&��v��i(���[��14P�1�V���V�b�C�� ���ł�$�$����Y��j���J󈗯_�\��g�BaԤݯ6�t�&�������G(�g�q2���߱�I�Jk6̚	$j�f˄_)�&qn�$�?<�C����@tK�_�L �`�"��'��>/��CX�����{KM�&�������?\闧%P�pf7��X=@�}�L�h�I�S
�~�*�7��%C�ꪩ��c��H�q��ux�冏��ګ����d�c%�9�J-�?��Ϩ>�Q�@V��&��)������k7���}Ǘ�f���!�j�s��򸂫���*-��0����*f�ڧKf��x��җ`�����ai(z����8��8�ıhߍ%��ι������R ���pC������,%� A�R��_�T^�^_g�b!�CV��D r�,�ܬ�wB�t��\�
�g�Ĩl����ȷ�_�&A����;t~��P���*������/�/��rA�R���ْ�j����}r�y���������jg�({hɭ8��Ų���m�ID,�TC�j�6��(LO+Mԕ���vW"K�u��c_@�-�w���f�B^���u��P�u&��(R攡�v3:F�ܻ3#���r����-�!&s`P�J���ujo5�ul�4X'n ��M��^6Y��b����A���C{���Ud��P �C+6��w��H�gzg�2=�͵�1b�����=�$���麔���] �#������$O�}C��e: a^�Z��5�[_�#����I��t�n�d�~�β?��$O`�6ǹ�kԸ�H6I~�%F�H5�}U�6?bHÁ�B ���c̿�~�W4c%���-�s�E�`�6�Qy�F�˜��P9���Z�����_���6�D�,���j�7�ɹ��2.���\]��n4j*��wӑ�v����ۇ %��2�.����D�f��$K�����p��&���W�>p�LY�K
���f�U1;U��"��W*�!^KGA�Y��ڞ�/+��֪�"3�\K4fU��Ey���|�����@�ßDY����J�v( �ڎa �ʺ(�����=�"�lq�$eԖ��H���cʂ0/ߝ�� ��{�X�$-��E�UFV�<K�i��4��HE�ވĲ�^$��Iɖ�w�˸1����~���ߨ=���i�6����|�B���������~24�c����.���Aؖ�RyT߬��@tP����R�hO��b[��،���*�j�;o���2�V47�ǥ2��j�fPw3^#v�R@z ���2>K�T�DV��:K�\����9��깄��ў̪�4zY���j3~��p1�mk]G��f���G��@Y�2��Q�#+�g�l�3=��4�e�楕��e�p�z�K@�8@~�*�(��3^UO�'^2�zIDD1MC��N��@\C�e���/��1�i���F{�X'��=������7ެ~��z4h�'̚i�|��e��?�K������]���T2�84u9���x_����炤���M؈�?��^G�e��N} ��	���X�it���P�2ɠ��&���AGN��Z3��`�_�J/���>RImv��/� &~��Ei�if�u�YH��[����[�:���v5��
���=u0 :ϐGѶF��O%�б{ug�r���V\>�}Y\�O�^�T��5���Om)���Nm�\E����4��X��3G2��SQ�-�)>a5n���/��z�G��`KcͿ����vi{ȥ����g���_�!�Xq�����U��s;\ݏùn��KWx5��{�z�͐�j��K�Beݺ9�S��Jy�Et�6#�8��j<� R|��[�,FĊ�����'���N�[	)�mH�=���~Ri�IĬ٫iHlV��5Bf��T*J��w�6Pc�ѡ6kI�lY�	�*j�ۧ0�viO�'x�C�F�k"�H�r�`�,q>|*k�E����@*mxj�=��s�
�(i���;�y����E�"�
����:$.��Ƞ�e�ҋ��7	���t�n�j,z`�M��j��$�5�q������-a��D�,�Z���0����� ��!�X5}>{=�>jJ~O"ӂeBԿr���A�kG�ј�(ӷ	��{F��B�CeX� %H��䲖r�J��x�����N7&M��'Xv�P�g��QC<���c0�T;����^A��P��uSm��>�A@�D��ĵ�۱vfdx�,N}�$:��(S
���*x���+���9���@[��FC�%���&����I����sKl��˒�@P�׃��)��|��uu	i^_^`�-�t���0��E���"u.��T#֬��^{�+Cꇛp��ҏ��OP2Y)���mG0&�!�G�#������AƓs��%]���^�J7aR��\�v�[�@��ňJg�W�4�V���_������'7�wy	$����A�Ll�b��E�_V�du_�g?�� 9}?(��8l��u�`�M���s#;�*�u'f59D�~�x��>����~��H�.>��
a�ػ������ wN��=z�9=����e��9$�M��*+.Vޘ 5 �E܃ܲ�%3=�z �[L���� �|��$0������c�Hp?'z��:�䓇��6@+��Ԕ�/�75�i�̥���u�X�\�JX�b�����y�f��E�\�.fڏi&���0��s����=�X{7bE|	�.R>f�e&@Y?�_��V�) �{ 0� 3�3���k�.p]U;�ᖈ�����H|�+(ycw����ì(U^�r,��'��&ֿ*/��X�~X}�m�SG-*��1����0|<�q�]N�/3��4��q�~�q���$	�ʘ�kx�<��4�����@Y2��U�44�&�	�PN0g��VZJ��гJ�ϊ���[{�5ʨf�ǡ�.�ߑ���㡘h�	�5jl���#�0�s�*���}%�,�#���KJq��+}|�;�邶G��d!���×'���J��<����\�~G�H2����)��2f�l	X��Q�:J(Ueq56�2�Y��	pI]�i6b-c�>�,��_��Eq�E(�EY)CX��Ƈ�KڦlL�	��6q�q��d/̩qX�	}��&K�%�����U(~\o�%��f=�X�d}qg���{�I �.�D�ޓ��%�
�갸N�)����n���nĀ�Z�t=�I;�,�jc+�2�Z-N���z���QU	�e^�R;������p�a����Ҝ}��f��#ǧ��ٹ����`�W>*��w�S�I����f\omK�x��P�f*��t��a塀��=8�YZ��k�7�W�ki%ο�����d�-��RF�v���8��m�c�F�R�y_��u^s+�g���I ������,�l��}ۮtrq`���vg/�lk��h����vCA�y���tD��֨�������γ��/v�A/������[����=�@�ug�?���<���.J�p�(�f7�3�,ƺ렌p[m|��,p����@"6��r(��MZ ���Qk]fK�;X�c��a�s�ĺ��U��Ƈ�ϻB�P�
�;Q���7���3@Ä܁Q����eϸ)M�ս�!�`�P��ݑ�ju*�;�݁�T�nf�M�3�6�y��ͻ�ay{��s�ۆi���p�I��6�x���{H��g����1��)X��Uշ�Д\]fA���e���J����")�P�����^����]9�"@�e/���.��7͖=�V���F�=O'5��l A�r��DW�e��7��z<�ĉߥ�66�K#bҏ�D����D��G찵�ID�����0� j>`V�h`���3b�_A��?ʧ�V�̃-V�9]���������(�pٜ�=c^��0��ŋ���V���]��­��y:�R�+3�����엧3� v
�N\/ C#R���Вdb��ه��!Y�輅��h��Q{�B��0ǖy(�E:��zj1Q�W>� '�xF�jg��y/�!��K��i���S���T��3�w�����祖707�`rC���S�Y��'�?�~]d��-!?�n)��`p���[����Q�����'\����-�lE�$]��(�d 8@3�#�ܺ�s�hF���9G�K�I�m��S��e/x��w�#1��)�{/�R8F��<j4�2؇������7�h+�����Q��}��Ca�K^[�CH���N�`�O�bC9��ux�̦�чV���/��3W�W6����e���N��:�Q5���V���ԓ��+-�n���$ �N�{D3�R�` ���-�*�I�ʋ�w�0 n<퍸����Ou"��S\U��],�[w�:1�������!�O�ue9�:��GZL�F	�_OmS+���MT�g�:0Y����~+\S�q}��O�T7n�}[�����)ϸ��/�\���<(�V��{��0��*��)��ynNp��w��z݃�%��;ܶ$(����l��������!d�i����3���UɕdZ#m�״�������5�iעZϊ�Zj�K�����Ǣa㸯�u�����~@W88�GjX�h�h�z|�&��m�����7��u�]�	q;�H�}��<c�R�'{���i��vV��5��]t�rRb����Pp�cǠ��qk�wyl�ư��𢡊0+PKO�)+x�f��@kj8��E�t �|r:E��P���kx�����
�Ri��
҃+:����E��
k���O�h� �'���#����7Q'��7���,�|M��Mm�$�s1q�&��_�'�;g�,��{�T��J�N���W�-�*:����>�'rˆF}J���ʊ��A��<k�YИر��Q�M��܁"�fӋgX	�?%������������G�A�m��r�����o:�|@QjX��+�rF��piT~�kW��J�:�Z����L9���ȭ��!�ߵ6�ه&�6���٧��	��ag�^"6�;���9���&C�xD���OS��a��P��6i3�1V��<�;t��<�J���ӟ2� ��u �H�I��&�;���Ǿ`��>L�U��:�V}�HA�emm6�v*a9�M���*\�1��{DR��0��Ws�溲#�R0pp��~�}r��֋SKl|�������oL��p7XA�K%���g��ח�'o�#[�ߙ��1��+�p��)�y�F��>���w�ЀmX9o���|�bvm��[��y�[�fd�$EW~:.{o`�ûv�N�y�%r�s>�[�rYM{��|~̬.g�qP��@�m�_��A��W)��B{��� ��+��q��U�OƖ}���I�׭}����0y؇��"�]�a*U��!"'�K(&��/�;p����C�G�N�S֓˘<yؿ]�D�/LW4*9���$�i�,	���`�<�(��������5UT�&"����a	t��N��t�]G�Z6���D/y����{P���[tǖ�u�� ��2!�vshVS�5���H/��������81�Z�0����n:4J���+2�Ͻ�����hʏw�ݎ���'�r��JΉ��� �\LZ��=x��8�"�/��A���w�-�Ɓ�(
��q��2�Ė�:ӚI���67�f����A"ڨ   K  4  x  �  �+  �7  �C  �O  �[  �c  �n  !v  i|  ��  ��  >�  ��  ś  	�  L�  ��  д  G�  ��  {�  ��  �  G�  ��  ��  0�  ��  ��  � 0 t _  R% �+ 0-  İ���	����Zv)C�'ll\�0BL[H<yVCQ��F��e�P(������C�<��	��e��A��+O��$���X@�<�v�C��p�TJ��izsf�a�<�&	�P����w�&H�ؐ���e�<�0i�������^z��B�V�<��(��Fz,Q��!\:�\U�N�R�<yӅ�I~��3��,}��٣�JVy�<a㇊)nt��;G�ʏ���b��Kv�<i�B�r�8��L	�W6�}�=T��zf���R]��0/�6őf?D�haV���  ʔ ݿ���1D��[�
(m����@!\	{�� 7�.D��`ƭ�}`|��a˚t���Q3)-D�[2�ߌ=�v!����ɳ� 8D�t���O�u|D�Z��Y�P�1c��7D�LÐmֱlGfPb��U̮L,�0C�I�[mH=�W�٠d��C�l�&9�dC�IMM^� a!1�>�Ie�?`'�B�	5Jy�]��tn`���JF}��B�	�v�6��V�+#*t�c2H�`��B�ɦr9\�{��*v�h��⡍��vC�I�v��ɐ�ƙ$�P(˅��=EItC�I��9��ǟ l�����&2lC�IO��P��(����'�lZ@C�I�aS����k��p,rI�3%�`B䉅%���Gk�S�X�z'.�#�C䉙U���@
��K�V�j6.����B�I6\�qi��-d@��4�\�Y�B�|�d���a϶l	Ҭ����_��C䉈-�I�����NL�,�ب�E�8D�l�C�*&�n�h��Ώh�YS�j!D�h�$�$!��0*$�b�p��� D��3�X(q~T�אFbv��K!D�ȩrMY>n��ڵ��$V�$�P�5D�l;'N��d�MJ�6[EHS�%D�����£j|)��f�}�� �L?D�,q�
ۨP>&@���S�b��K� !D��`�AJK[�D�!�Y��dZ��Oj4���wyl��p̂
��: GǄ��̇�I\�'؆�Ȣ��{]؈� j]	����Q��/���
���?����&�>6EZD�O��=���bRjI�u�V�R�Ӂ�Ukܓ���H�(���#;���D�ŏv�nqjw�i�ў"~nZ�a��q��e6�-�0�	`"=qǓp5J);tGO3�,e+G��(�ц�s��Hx�V>��RӠ��bʎm��݌���G�9��@�׮T�xDb�S� ߞ,�B�őE�Ψ��f��=�Ó �6�+��^ HZV�2��[���'7ў���I�|]������,��4�Қf�<9&�h���Ϙ'ZLL)�@Khv���$�
D��	�'�ў�}
���'o�����'q���b��K�<ɓ�G;�$K���~G����^�'9ўʧG_�d@Xi�¤0���;���!��	V�O��=B!��.j8�x�Y�6���+*��hO��G;���6'uD4q�g�##�Q��D{*�,�W���P�F�`��	s_Xt���=�S��y�/˽*R�k��M.z��,�΍ �M�O<��O?7�L�R���;U�Z+�|���%ȣ9!���nw ���,k���i�F*Q��F{*��ZbȀ�<b�h����$2=r�ѧ"OH���,��*�~5�M*��B��b>��!�P6�8��`ƕ9��ɋ�"D�� dC�@Cx����䂘?n��j�O���=�Gˍo�hlAGN�10w��)ӎ��<Ɉ��S5}��L��@�d�l�V�ڸ?�C�Ii\�D�ҦR#d�0���C��*�~E�E�	��Q�-�*z�#>���d�~*R��wB�k�-63"ɸD���<I
��[��TR���:�(9#e�y�����Vr�r�#@`��t`�deV]�?�	�q�,�5'�	5ȍj@�Z�������YL��1O��R��'<E{�G3%�89JS"OQ(#�''+�����j�R�r7��l?a�{B�T-L��֝�v}��R��7�Rɛ�Y���B����������GO��m����	٠z�V�>Ɋ��O(чmF��j���-����e��IG�O�؂'	��l���#_�h�~P
�'��=
F+�ٕ�W����O��	f�S�OFXi3'O1��yZЊ�36�����M���E9;��h2	�� �m��CM�<����0~5�h�݂\|i���K�lD{"GW�Yh�A�~��qQ�N�����<ɐ�'Fa�dJ;'Ն4B���T����Š��O�~!�@m�p���ΌgOt]�'�k�'��xBd��tA��y�7eXMb�(O�=�O�*w�5WK�u�1@N���Ұi�!���8xb�1'̎qQ��g���O!�d�R�$Y"閑FY�}ZA �(�!�Ě�R��$�XbR1"���!�D�-B>���ŰQ� ��3~!���Q������b��!k!�����lӢ�EU�ْ�B�ip���E{��th��L���-#U�z�$5C�"O���G��/;oHE��-��Jv�l3�'Cў"~"'d�c��H��!�,/.��2���ybfүt��+e!�TjB�߷�y@�&�<��	ׂ�lqÆ���0>)H>�rC�{ȼ�	���5Y��K�~�<�����i\(����ڡ%SNѸ�gP�'��HD����y��tK�j�Bt�(1�[��y#�QC"&/�B����X990,Fz��9O�۱�ɨBq�%�r�߭�M	�'s�Ms��2+^}����^��h�'aR��>�d�yb����P���y�G��R��@EmX� iz�1���+�y�>1�΁!DK�&ȓT��<��OZ�����R10NO�7/jH@(��b!�D�p�tY����"d���G��v�)��-��Ț/�T-�,�h,��[hC�I�8W*18`c�]b�US�F�!�`�{&���B�U;���`+	�ri�!�b"	�3a}R)0?9u+6_%!�x�L�*K�@�<!D�*yڡ2k�C�θPF�T�'ў�'\���c [:ԙ�v�E�A~H؄ȓ;Ȗ�s�+U����wIC#��ȓ+�>u5������iv�U-(f����<q�.��nu�P;�e�D΄�:�b�<��B�:�[$��eƸ�zvhB[�<Qu@��<�ر����BzqH�Z�<鴀΃%uF��v+�C�$e�Q�@r�'���%�'6���Ѷ� �mU���� ���Y��);DH{����2�"���}t�U��44Y2#<E�$�	�WԾ�W,�M�ŨE䒰3h��q�dI�'���j�2
!NFThE\�����-�^i����"U������ 3�HC�Ɉa���sg;=�����S6��C�)� �ј� 4��,K���`��p�"OsU���&gP��d�x=�h�"O��ra,��S$�[{"�@w"O��T��[�>���:?oЌ"O�J�@k�<tP�@��yp�]�a"O ��W�+�ԍ;F/1���W�'��O6D8���5�ʔI�n�@ٖ�c"O<eGc��QN�(�#��%Ϫ`b"O8���_�a���t;����S"O쩡��+���b��w�P`��"O�XP/ג
Ơ4��C�R��(�"O��aD�0`�تe�2}��"O&<@UI�C'`e#w͑V Z7"OT���W#J&U�"�\;]c��"O�5�Њ3<�A�b�mKF,��"O0� ��xT�`+b��2�4=��"O�P��T
���9 �1$�6i��"O����IΩ[;rq`dIQg�\�f"ORlz��X%JA4TiiN�q\�-��"O��e�%~H%�R&v��q"O$<Z׋�=xn��'fEL� �"O��P�g�.z�gG�g�=�"O�8��^�1�� C�Ȯ���(@"O��)0+�/e6Mz���dM�)�"O��RA��$�2�E�B+��"O��+�#���z'@�%cF�s�"Ox�JŌ<��ap�Ôj��u"O@-Z� (;@���%U(+b�z�"O���AN7�&����ǳfLvLa"OA��#ӭ2o4ݒ%�S�kA� ��"O>�C�_�u��)f#A&U�4"O2��c�?�����Z�x7L�z'"O|�	�	L1���pBZ�5���1"O�8p���J�J$����$J"O A��1*�$�B��U��1��"O�py"fQzh2Q�FU|��m;e"O~X��G�9JV$k'��|�6��"OXM��W=P��I�%�t�@"O4�@CA����rȝ�eʊ�pe"Ol���(�7�>��v�U2_Y�"O�t
cH��PiC�ɴ$�}
�"O4TUY�	�H֟+pБ;�"O���!=U�؈&��>b֌bg"O$Is�:XbAat�Ӳb���"Of`�E�H�n�Z�kW�/Pn i�"OVT���Y+-~v�A7**}Lܜ8�"O� ��b�~����w�Ύ8T�k�"ON�Q��I�:иc�V;-f"OTAт)}X����97Q40@w"O�(�äN(>���@R�yHvx�"OF����2�8}�B,I� `�lx�"O��q��ߖ/�D��v*�Nuū�"Or5��AZ=_��E��/��"O�d��mT�<��!�%��a�(�XC*O:	WM�.X��z�C�[>���'/���Qo��MT�lK�^�[p���'�4,�g�H(�e��O�� i�'�0���c�]�U@��
1Z
  ��'E�tabـK��K�*ޮj�@��ȓ/�%�ݓh�@x*C�U�U����vN���F�&Wdrb��-�Y�ȓ4�|�,�|����I�*(���o��d�m~	�v�O&I<n���^؜�3���'g-� ��#d�����S�? ����ԍy���k�nF<!��hT"O�郤lC�9��pXBlO�=r"O­�䆆�m~�` D$�'j�����"Op�g�H+�,���c 7}"�i1�"O���P8X�Z�v�Ծp�|a�'��Z�`��ݟ0������$��d��[���N���C�i8�5�	ԟ�I��p�����ş���柰�ɷ=�\MUjmH�{Q#�5v^:��I����	���a�����Op�$�O����O��`KC�[� �F��6[	�Vh�O
�$�O���OX��O��d�O��$�Odp�L'��Lj���,N�Y�`�O2�$�O���O����OD�d�O��$�O.,t�* ���C��;k��@���O�D�O��d�O����O����O���O�ٱ�]3rW����n�`,|�%�O����O
���O��d�O����O���O�����:��A95�X�{�4@�օ�O���O����O��D�O��$�O:�d�Oԉ8���6w���7��ne��`1"�O~��O��d�O���O����O����O����c�#{x���B��edH�'M�O��O����OD���O����Ot���O��� �,�|@r��+m���L�O��D�O����Op�D�O���O����OR�Id�~�r`�-P�-�!�d��O����O��OX��O���OF���O��ض�˪|�h��R�J�#�����OB�$�O^�D�O����O�n�:�M���?�R<d^
�qCD�&u��ȳt ������O�O���V�2��O,�n�p���*���+g�)s��q< ��fBl���ٴ�?�J>�g~rLuӌ	�3۶����MZ�F�܉$�O����^��Ih�6O�$�ܶT��TA��J�ɬB��j.^0;�� �e���<1���D8�'9�����δR��/�̴02�i���R�y2�)��4|+�E��A���(��i�/uZ&@�ߴ:��=O��Ş'��z�N�<� ƌ�.�v�P�����V)��<��m�G�:�F��hO�I�O����Z51U�����-r��p�s?O����p��n���'�@a�g��P�9�n&W��i����Lb}b�cӆ�o�<Y�O��c��x��!�����A�Q��XC"��6����TF4��3�r��DC����¦�7D�`9�$ʃ&zq�k5��ny�T���)��<�0%
 �e
W`ҺQ�`���K\�<���i�
�H�O­l�M��|Bb쎍h�`�A���T���GJ��<�`�i(|7��O�9 0DO�;A���HR�b�ʄ`&l�S��6R;��!�� ^�� �����]�&?u�Ug��uN*��FE��B��Y
f�+?��i�
���y��O��OP̠���5-���MZ$.~1���>!A�i�7Mc�H%>	�SΟ��1d	����q�b$J�`k�CD�4㺅��Φ>a�G^�I-J�IW�?_6��'��4��!���=J�P�FR"9�*�H����D�<AK>�u�iB�r�'w���p$j\�E��m� g�d�:�'��6�+�i>��M�0�ibA=����L�"���V��"R���-�yҏ�
lf�l[�F�?7������bZwE ��1L)���o	�/{d�g���Lf���?�*O0�S�O?:���jZiǺ51��en��yҭp�v� ���(�4��|�$�h$iޖ[r8+5-��r�� h�'��I�M��i���
�/��ȝ'%عA �,R�m��O.c�>�@E?��-3�b_u�H�3F�xB���S@y��'�P$s�љ^]�q ����*y۟'��'�Z7�
4L1O��'A �Y��([����߽A]��'@��!\�&�aӼ�	]�S�?��2�H8+��`
Pg�
_����]*S�@8S�*$x�R��W��PI>)t��MeL�2�	S�<�2!��:�?1���?����?�|+Ob=l�8 ^>M�Q�i��J$&�UN���Styb%~Ӛ⟀J�O�m��X��{�㊫i��eqA�I8K�Y[�4WN��jIV�Z�ؙ'�B͉<Tp���E$&��"�JV.Bg�v��MĴ*�n��jy"�'���'���'wY>�-֌L�����D�d�q�� ��M�	�<a���?�K~ΓOV��w�6��@ hr�K�	MmB��W�g�F]mZ��?��O1����M�(��d�#{kP���� /Rh�Q�߬.��+<�
��B �7%�Oʓ�?1�M���2�\=��A���P�������?)���?!.OtloZ%XG$�	�|�	6!�q�r�����PG
�;2*A�?��P�p��4L�&��O�v��x9�ʨR���!�L?��L�'	�Qf^���m#s���)ә2��A��O><�T�ܮ&�
t�w�'�^T��OP�D�O��O��}���)�.!#R�ٳM��x�Ѕ��Rz|)���;=�6��:�������?ͻ����m��-�rY��
�P�H��)���!~�5l}��5�.?�ՀB�(��H+�k C�xr4��.t���1*��bt�O>�)O���O^�$�O���OZ�a���Hv^Ȃd��'	�����<٠�i�<�*��'�b�')��y����N�m�F B��Ig����f�hӆ���Q�O����C%⑈5!��h��2��@P����T����'�<6���F�I�|yK��/r9H2��8m����"B/g���'A��'n�Oy�	��M�a�<QE	�
@����ES$�L�Z�<1��i2�O  �'��6PΦͺܴFu��HgO�<���c5l�j����
��Tm�'"Ԥ*է�
-���c����n�� ��pt#��B��Nz0��t?O��d�O����Oz���OL�?��"Ґb����FAH�>>�(*P�{��	˟�*�4qu�'�D7-7���8TZ8�1,�"l"����䇖fe���	A}�@f��Llz>�+KDت�y����/�� ���n�/��a�@Ŕ������F� ��?�*O��̹߲p���$W���a���ue�+���Q9'�;�I�?���v" �4扑(趡��B�s���X)�I�M�ľi�d%�i���s@H��|&4��G!�B�<т�M<W��)cCěSc���?����	�4�� %�0���>O6DB�f�&�LStNHcy�'b�)�3?��i v�nV�	m���kS攈�.3�ɪ�M����yOw�X��@g"�(��7p8�@�[覥�	�.s̨���n���I9 �Ф��D�4m�y�,� jH�8$� E�=?(���<����d ڧy�v3�I8A�H5*���N���;f�i�4��y"�i��3'��z�B��u�����.�W	r1xڴ5���1Oj��|"�'�?Q��#�8�y�U	@e)	��1[AhԹ=�ةΓT��R����Ӌ�4�����"Yh��&IH3�fӁj\�6,��<�I>�ŵir���y�BW�'&�ы��U���$P�Y�-r�|r�>97�i{Z7�s���'	v�(6�3#�8�R )�q��q�'��)3r���R�D�������:�݂��N��9���WR%:��u�$=�(��4dޕ���D�Oz�d�OB�=�'�?�%�(�j�ࣖ�h}�A�BLS��?��i�| �4]�<H�4���y�fפ\�����"��Pv�!�P�7�y��c���l�M�O�V�&9�'H��;jz�ȕ�X$�HJ�囬J�z��o��'����X�I��	؟��I�A����˚35����Un�L��4�'��6�����!��ɟ,��?��X�ZT��I�búA�D>&`��+\�R�4>"�Ve�O��<�����a�%&�]BN`�A��c1��:rHW-zĥZW�<A��6$�� �jW����dR��B���M��12��G�m \�d�Or���O��4�2�l��)����]�����遬aTk��ג�y��t�:㟰�OB�m�>�MS¾i�lL����j0@!ԬN��xR�6�i��Ov���M�@ITX�1�,����d�rEB=ځ��&rr�q��Q�<)���?��?����?a����+8=�L"�%�0t�
��Cf�F���՟���4*�r=�O�"6�?��^]�rB����*.����(Rf[���Ia}��{%o��d��ī���,�#g� �H���*9:�R�����}fD4Sc��).
<&�0�'��'���'T1Cm�#0�.��荖,"��P�'��]�`Hݴv�͓�?	����� W��`��j��&T�t'X,`�I��$���Rڴ+�B���A=
�B0k�2d�$����30!��?{� <��O�<ͧJ�8�3�ٿ��Yn.�`�M�LY��3၏v3l
���?Q��?	�Ş��Đզ�rE�9ƼK�&ϴ�|L��eOW�h�w�v���C}R�|Ӱ���K�Hv�	�aE,!#��e�ݦ��4���$KU~�G_�H��▄<���\j� U-"+����	 T>x�Iey��'S��'���'�U>QiF�ضL��i��C�+� �r%��M��:�?I���?�J~ΓJ;��wA>�c!�Z�:�sѢ��+�D��hӢulZ(�?a�O1�&tQ��A�6��Շx8u�Hz9�I�#�	6��T�d�t�0%m"<�Op˓�?��W����X�Sk���ҝ[�N�Q��?����?/O��oZ�5R|$�I���	�nr�E��@X&t�b8S��
"@���?��S�D�ش,���l�Or�'$�F���K�n#�,qW���2���
��mP2��	`:��O~����
fp���$�!st��Q�0�V�ۿts�I���?���?����h�>���-QKX�CBC�%=�H����s_��$��I���'?��i��O�M2:��|��gP�`%b�K#o�|��D�Ŧ��4�&�
.q���a�O(�K�j�I��<#�-C�N|��tO�[H��Q.�3-���OJʓ�?!���?i��?I��C�H�CD��%U��u�֫��?�*YX.O<�o�!܆��&����?y�'x��	�1���{E�Q��P��cո�1k�O.�o��M���'o�O����Oo�����V$2G��;�l���F��d��S��`@�%n�H�i�Q�	ey��%��Js�ЫHV�d��*�B�'���'��O��ɋ�M�UE���?�ɇ'�(uIFoU2�(��E��<�&�i��OL��'j�6��Φ��ܴu(�P���9ѪDkSGO:�(��j�zA�'�Tka�>=l�a8g���.e�͢��G?B۪ة�JˑP�^��D*c����]yR�"~J��ԗ<s���ٕT�* �� �N���D�)��$E�u&��)��	�r2�E��(�D/МS�'���0�M��iK�oZ7
m����'HR� !�޸ @�73�H���i]g7z QG�	<R�52��i>q�'����9�!;�L���j��5���y|r�}��3��D�|��AW,��7� �wgzu���v~�`�>�״i�>6�g��%>��ӏU�<H�׬�:y�l�30��7f��X�"�I�ĉ��*(?Q�'!��i"�_���_�D�)��	*$����%"�;�z��-O���<�|�'��7���L�,)����k*
�g�x1n��A�����4�?�I>��<�g�i\��ٳLζXT�H��(�3kv�L�(o�����(̄i{:O8����=�XD��h�7O��)� &�����1��$�6��2kZuHC��OX˓�h��dh���y�uZg-��YֱJ�KȦu�08�	Z��ԛ�w.�@;���!�*���C�&f�=��Nl�z�o�<�O�������G�Nl�{v8OV����E�6el��c�єLB(�=O�h��	�8U��6�ĩ<�'�?�4K�E�Z�cB�޻����
�?����?�����T�5"2��ğl����!��Ź>�.�Ӂi�p>�U��Q����ɉ�M�i>l��>	w��o����jW+wYv�Gm	�<y��9���C樏�S�܍[,O��	�w
B][2�O�%���2z�R]#���� ���l�O���O�$�O&�}���VSLq�)5b �D�c�Ħ:��$+�?����)x�ɪ�MӋ�w�X��g��m`��r�= �'�7m����ڴt>i2"ǚ�<��]��q�.	w�W/u�m����!���S�g�*�䓠�d�O��D�O����O ����y3��@��.G�yq��T���CƛֺX�����?Q�����<�2�8N�РEh�K����T[�	�M�b�i�@�D+�i��v�)��`|a��/BӀ]$�Z�{4P�j�h]���ʓt�~��6��v��(�H>�.Odm�C��9}��=C��:J�-��?���?���?ͧ��ĉ���P��}� R�(i=`x���^<��s `�`Q�4�?qI>q%]���ߴXG���hӬyBפM�D���'ƶ��@iN�H �A�D:O����8/�LxC��W�e��ʓ��ƹ�`���ӈ[<\ C�%��M�|�a>O8��Oh��O��D�O��?�8F�ʄd���Tk�B���ğ��ɼ�M���`~��|���D�<i��S� c�؁��L&Vp�qK"��*V����4�f�O�D}�P���y��'qx��*�\H�E�@i����><��̑"�'>��ȟ���L�I76�!�V���%P�l��Iٟȕ'�07��A����?����:R�ъ&����Hu]���NNN~b$�>�׸i��7��� '>���Ƞ��e��<���U�0vt�A�Q�"��X�cʅ[y�O�^�e� �'�ʰQ!b�Y���ǩ�,a#B���'f2�'�r���$�'TDI�Z����}���	tJ2�	m�%�l�)p�й_ș�Iߟ`[ڴ���|2�T����4&�03*q��7�ܫ��A�&�i9@7�|��@9�=O���,S�i���\!��ʓk�6Ё��0D��H'T�r����$�O��O>�$�O���|��O����,�i�ԉ�a&BB���h��a��'<�O'�s�������l��I����glG&|/B%z#��O��6�}����J}�O����O�x\v#�yb- VP�TIPs|>�ʃĂ��y��2dn���'�<#�'o�ȟ$���y����g�=;,���7�+��y�Iʟ��	ɟx�'�7��E���O����1����MC�F�`��d��h�z��[�Or�m��M���'M�I�Z������I)�+� ��fz�I�T���ec�BFEYdy��O�%�q�e����>:Y .�fS����`��X�b�'���'%�s�en�9��٦���/�4�sJş4Zڴ+�8��'�271�iޑ�7�V�p����2��jh�$C�4w��v`dӸe`���i��D�O�(FL[�e;D�d�D�k�f�2C�,O�2YE)�6,��O0��?a��?9���?	�eH�}+t�L�D�J�*R��$��0*,Oz]oZ�:c ��$��`�s�<�FNՎ(<�=��8<��ڼ�	�O�\l���M�@�'��O��D�O&H�H���n!�p���½�^���Ș*Z�MX�U�hza�B���6dH��_yr��.뒰j�Nl� b,���'�R�'n�O��I�Ms'H��<�eJ�EO0��c�M�\K��^�<�s�iy�O=�'d6-����*�4:ي|�堗�;�n�c�V.M�<�b�%��vz���?��K>B�^������������|�1t,��3��2RעDjŰx�JUnt��Iៀ�I䟔��������7=����V-�� l2t������O�n��sPx�'��֐|,X�2�0�{p���7���q떎\�$�>�!�ii�7���J5�C�	q���O�+����|�`�bI���� ��d�X0Y��r�F�O\��?��?I��C�>u˗�Q�(��,�S�ۺ�t�Q��?�(O>@n�a*�q�	ǟ��IK�tKؗ �xP���̧;�dPGK�	��$�G}B�n��n��?�H|J��!;N$rd��\MpqA�>�����5HM��8�`���М�B$LWd^�O� 
�C!c�lS%偡H�𔂲M�O���O����O1�$ʓ6���lܨ<"��!p�&W1��P6��_��Y�R�<#�4��'9����6�зp���P��8�L劕F֦H��7���x�L��R������4�ɣ_J��!�@y�@^�f�I��*����n��yrV�,����Iџ8�I����Oq����H
!D���s���E���SDz�8M�8O��$�O��d̦�]�Z�౑�"�2~�nh��[-�����4�6��O~��|��'��f�Y�j�=��"ȋ��L�{e]��!��;�ȵ͓vL 3p��8�rH>9(O���O,x�,B��r<��b��xJ&&�On���O�D�<P�i>y{�'/R�'��ѕƄX�t\1��6��j2�'h�'�F�o��hnӴ��IH}��=Vp��ō�����ǯ�yr�'bZ��B�(ZOr��qQ�x��)mȘ%��۟��r��&G���ĭ0Pl�xs�J֟@�	ǟ\�Iǟ�D�4�'H|���`_wո�ÆN֭L�"}�';�7�S7)���_ƛ��'�ɧy����5�Rn�:ua���d���y"p��<o��M�v&��6�8�̓�?����\ &$A�\_� ��j#Ǒ;k����h���"6H&�D�<���?	���?9��?�Cl�$1_�X���|m6`$���$Ԧac��㟈��ڟd&?�I��2X�q@�#q<�8��<�
��O�n�3�M���'P�O]���OG�@A[�Z&R� �ND�Uaѧwq��VV��� \�p.��E�C��{y�ŔN��˕e�#8����ֺ?p�'
��'��O��I?�M�v�K��?ysOU�:�f���Q X&���DK�<Y�iu�|��>�#�i�Z6�����",T4o���z���Cu:����U�H���&c���������%�5l'�\�'6�t@j�5�$�_Z"����V��� �`t���	zyrS�"~���ÎO�-��Q�
�0M�"\�<q��i�����O�<o�۟��'V�����
.�JDHϽYZH)54O��"{�6�e�4�$ؤv	�P�?O���O�!=J��©b�詅'�		�l!�ҩ�)<8,���,��|B*O��d�+�ĉP��[ Zg.U;�R�W��d<�$TǦ-x5i1�	e����Ut�`u-_�0���$����$D`}�|Ӑ�m��<L|2�O��MC�r���(��ҖK�2x���[�:�*�S~��OϬ]`6�P�'��'�����O�\��N[:z&��	�^���Izy���O�9o��.	��f'����">{R
���2?��i��|��y�*f�	�EؘuN� �f�#o�"e`2`��}�ɋ0�j��y�$�I�1K���dB9D�p�$���M �f�X%��*�&�X��<�����&�'N��ӧ��KMqJ��^�M$B�i�tS�y����ަ�C�4��B��� ���#��:ܴ�0O���|
�'�?1W��+ D6�Γ\[>�B��7|��|����\��q8L�������M>,O��O�Tc��(,y��S�.�*Yl�����Or���O:��<i��i?�}s�Q�x�	�0��GK� i�Ȣ�?r�?�U��ܴ!��F �O��*�@�3l8�cRiԼ2�48��?)���&.Rp�W��$󟬽)��A,9���Q.>�"Qi�l�� ���
&����O����O��9ڧ�?�� U��ɢ��	|A�Qk��υ�?��i����_����4�?aL>ͻl;Pdص,���� �/�̓=���~�p�l/P��n�m���	����ɷ�2�i� ɏF���I��/��0ՀG�	Jy��'u�'b��'W�A@u:Ĉe��b�HD����7]��MsW�L�?����?�H~ΓE�\�.A�{b�	cV���sz`�z�S��0�4�Vn�Ox���)��f������İ։����)��Rᄤ�d&�<�ǦI�cxld"�b�����$d��uh��'�y��� �t�(�d�OV���O��4�B˓@�6	�Z�b&P�rI�S(�:4����L���y�.x��pȭO�en�M#�ir��gA�:��P�s��Q2����}zB��'�B&��B����7:��	�?�YZcZ$1z�Ҙ)�"�#�V1:ޔdҟ'��'���'R�'��*pq�Y?n|I
�hU����1��O����O4�l�*_ȼU�'H�7�3�dS�愹0�ԾqO��S����2��{}"�t��lZ�Ȳ�-�2|�p�Iן�
�CW�r�B`CZ%<�(��6 X:p�<}b�(H/���'�x�'��'���'�����̘9 DX=��BE0R���'��P���ٴP�u�'$bQ>�I�n�2@�8MP+���!`.?��Y��P�4`�&m�O2�N��O:uq�$�׋E,lf�"�M��t�ԤS��+Lш�B��<�����"[���JՒ�`�nԮ8�3���3UT ���?*O���	�<վi,FaKm�-+����g�����J���������?��Y��[�4~,ei �B*��9�I�[ŨeJǵi=�7�G(g���B�<Ox�Ű+��U�d�T.���i��:uĀ�j� ��C��I=^�����O����O����Od�d�|bD��|f���Eɲ#LC MO�;~�V�O%�y�'���'�T7=���J���jɘf����S,��b�=o���M��'a�i>�S�?1	��V�N���I7;��A�V�	�EpSǐ�Y�L�	�k��i��G�4%=$�`�'��'B�$ ��|r`L�S���(r��'���'ar[�4�481L���?�p$�2�ŏS3}�ɹt*�y�B�����M�i��Ľ>��E�LX�W��7+N��Ā�<��j��SFB@EF��)O��I�@91P��OpBA�;K���b&�x����U��Op���Ov��O��}��k\l��ڏ�H�*WIȔ4�Z5��VY�ϖ ����Ħ��?ͻGd@`8��>����!b��0��	͓Sٛ�!z��lړ���;�m���	��D��HG"1p0tZd,��o�"P������4By�	^yR�'^��'0��'��k��J������?��U��؝a��	��M�e���<����?!M~�xI�M�$��nrl8rA�� �N�2S�t�QÑ�JV���4C2�O�4�O���%��*B�
�� F+5�`%3eM�v���wX�X�
� .�*��jr�`yRJ�;٦�!���cN�]����=��Iݟ��ɟ�dyc}Ӟ���7O*M��"��v桘`���~�$l�B6O��lZ|��RF���M�"�i� 7MJ�NJι���W�B��-�<3�:�gR�a��d�O��S�FT�{2¡��̱<��'(�k,��$M�U@�"���񓯚�+Ţq̓�?)��?����?�����Ot��cA��}*��ƚ�71=�WQ�l���M�H�T�mӶ�O�eÇ.T;9 ����ny�������'�h6���m�ӯh�h�5#���	�l0n� ��
�*�c�H��V(EP�j�[�,��	�~���)��<q���?���y�g��cWN��3�M{ˮ��A���?	�������Sd������ĔO��d)焓|��f+x(z�O���'k�6M�ͦ]����'���V����	�Dڿ`T3vI�p��1��Jۉ(L!�*O���T:X_�(���%��ɧ�"��!�="\AKs��K���O��D�O`���<�s�i�: �&A��Rpgë�j�C�;����ئ��?ٳQ�|�ڴ/��`��X�LA�N�<<3H!��E�E�ٴd��k�<��I3�(uA�%N�P̰+O��R�۹u�z,��6&I�q8O�˓�?���?����?�����)ۈE�ZE�_05����f�˿R&�mlZ�C��	ޟH�I�?���y��p�󮊷=6�@��N�$h��Nz�*\n��M;��'��i>Y��?��A�����'F���5��T���;�(`�;O��'I˺T�L}s��$��<9���?� ���H���˘0�H"��5�?���?�����$�ɦy�5�ן��ן�,D�h�6��P��!ӂ%����?#T�h��46ś�`�O��1��Y��'к"q�����9J����?����<]Ui�$�0��d����bA2����b@� �0]�����B�{ID�d�O����O��%�'�?@R:CP s��5�dYp*��?���in���V����4���y�ŃH�|��= N���*O��y�mӬ�mZ�Ms�m9|�ϓ�?�'^�+��a����+J�U�k��_s~qJ>�(O��d�O��D�O��$�O^!BT�۹A���+��Կ8�|)�"�<�i��ӄP�X��U�')�ʖ�U��lb�k�<bU҄�Ӣ���d��� ݴQp�����O���l߂L�6\:��:r��!�b�� �v�@�ȃ�	�q��ĉ
"�`�%�̕'h��0`߲x����L
{9h�'��'������T���޴X�v�S�O��|kdD�_2��1l϶j��uϓ9>���'3�'���y��V�r��n�y&��[@�E����W�����'�D"d���̟� Q��L��kFJ�My��OL�ט#Lr���4�P���S@h�dJL���������	���	L��S��<�7�����Ǡ��B��+���?���b4�VNH�z��I��MN>��`R�f�@USu%ȗ	�@�6!��]�Lߴw��O�|�Jw�J�y"�'#l�@��1̀t,��*���]-//,TҰ��@��'.�I�X�	���ɐf�bQFMX�>�z|bB�A8W�\�	�X�'�,7-	3+��d�O&�D�|R�L�n&a��኉�t�VJ~�>���i�7��ǟ��~2���0v1�c$ �zP�G��M��}b���UC�|�*O󩇦k�Z	�A%���"?�~��;l�]ңG�<�8�D�O
���O��ԟ���b�	y��I �M�w� -m8q��mª;�v�%��+`�f	̓�?�S�i�ɧ����>�i����RkA�=�,���4$�B����w��!lڲ;]Z��1�g��	$��0�����'�h�D�:��(ZSj�(�4ݒ�'��	�|��ԟ�	�L��~�͈1x�1,ș����	J���6�E�ad����O,��:�9OРlz�B�؍%�����D�5�j�����M���i#��D�>�'���'J���`�m�<����#s����N[�mp6���JU�<�!"��d�f������OX��C�{6�)(���.K��:�DV��B�d�OR�$�O˓c2�m׈m��') Y�G��D�e���c�`��@ �0@�|"�>��if�7�Q��'�x�wg�6i�`I�g�.�!P�'`2g	$+E:D�FP�>e���?��3@B�8��3��âEZ2���e)��s4���	��P�������C�O4rL�6��hf�E����	����n�N����<���i?b�|�w��}�c��F��-��I^XЁ��'�"6��Ub�4y���ؠ��<!��wL��5Hޛ^�t���jձ{� � >m̑¤W?����d�O��D�O��D�O���/(.Ld����#y[j�q��8���h��V��<r�'.�O4�s�h�f�F':MB0#��
��"��	;�������4�����O0�t��J�a���E�S�D���ʗ/dA�LX��I	(��Pk�N2b�L�&�T�'��1�Q�r�|�e��.�b��g�'���'"���4]�X�ܴ`0�ϓ!�di��
�kq(�
�I�7d��̓S�&�$�J}*z��n��M�	��z��ď�c�z�:�ܹ}BP8��u~��)]���Y�c[P"�O}6��<�v8��Û��R����9
������I؟����(��|�'?C�a�tF_�M������W;Tr ��'�� `�0ɱ���!�4��e � �!�\% N��PJ϶v?��6�'����Mke����.ݛT�� �O쁀ѡJ&<|�1J�,I���&b� V�Hm3BdA7�֒OJ��?���?��j�69���ը$d�p��ꉐL�����?9(OZio��R=���?�,�օه��b9NLdFtbq����D[�O�Ul�*�M���')���!���*�%��j�+i����a�"\�ݢ�'"����|�S�C�;J(d�L>����H�h�b�`ȅx����?!���?Q��?�|�+O�Ln�3w$��ժF� ����hJ֘8#�~y2Edӄ⟔ҪO�l>y�@ ��D�7'��,h H�'&�MB�i���K�IC����A-H�(ԋ�* �˓Q�x�Q�ͤ3�.��.��KV͓��$�O���OR��O���|r�J���Zv!DN5m�AN�}țF����y��'0B���'�87=�Ԡp��<����&G$_��i���ߦ�޴.x2Y����?��?Fop���#u�� U �n�$[:�h�Aҕ]>i��<O~A`���cg(EY��<���<9���?��HZp:A�����P��o���?i��?�����$Ҧ�r�+�͟����$��Ǌ�D�f� k�+?���6�R�������M�w�i����>a�.�9*��@�wρ�rh��TF~2�,,w|)�@ 7f�O��I�@ )7�GE�W��	�~��ہM��,_��'p��'��Sߟ,:Gk�%6��螬de��C�����۴"�~ԃ-O�|n�ϟ%��]�*-X`J��H�W��9�/٨�@�	��M���i&6��)c�Xi�5O������Pmֳ)�X�ѫ+"A�pw �9P.�!/�U�ITyr�'���'NB�'H��D9
�B�a�7����d'ܧ
T剋�M�$&��$�O$�?�C��L�10L�Wb4�
���B��d�A�۴1{��4�OI���6������k�m�������	�Ut����L�j�&���'2X��2.�7TXt���(��=���P�'���'����_���۴,�D���UԕC��L0uJ�KLz���; ���^}r�z�h�nZ�M�4!�B�~�����W�tYgh�7.��4J����<���v��"�g�A�4��)O�����̄E)4!�b˘PtB�a�o��<Q��?����?Q���?q���-Цz��1�0�=$��J�l̡�y"�'��/iӜ�	���T��4�� ���+cT���D�+h����`�'�����M3d�i;�D��:K���'�ң"Y3�1	�D�v ��KD "1�ܚ ��I8�i��|2\�`�Iٟ������#���:��(�R؜�&������IFyl�$�;�����	`��
3O���Q!���QB~���΁����]}��h��eo:�?�K|���y���ZRB�V��C�<.A��Ȃ=�((�@C=������.2#(�W�|be��`�1��@֭ �X�ru��'��'���tR��YڴCͰM@Q!n��I��Ⱥ9X�m{��OD~�oj���<X�Onڋ%l�x+2�չ��I��[8mF�ش~F�v�î �iA�'o���0y�|��摂o��!2 Ntj'`T�&�)5�ƒ%��	gy�'iB�'�r�'B�Q>M;U�&=����K܍JtJ���ٹ�M��d�<����?�N~Γ9��w���)��1�`b����ެ�U�b�poZ��?��O�	Ꟙ�� �VV�Y�<O6�� ��Y�4T�ADî6$1�:O���lݵ)<8��qa=�D�<Q���?Y�Ɉ�+����]
NiHP �*�?����?�����$�����d%?��J4�����(��q��Lpx�����7v�I�M� �i"h���>%��P�d��d���D��A��<���K�]�rA
�j$��.O6��T��a�o�O�����4[����ǎ��dC���O��$�O����O:�}��b4���[(;W�8�[���1C����f�7��D�ئ1�?�;G�B��׮V�C�z�r�m��b5��Γ]����|�`po����q8
p���
n3Nը�"A��xwT�"C
HX㠗`I �s�f�T�_4���d�5�j�ɢ��CT��#�?�!� |�N�apf	^� ��'�H)�gK��w��(g�z������s�iy1ę�M@f�3�8�Z�(F�y!�,ɀ#�E���d����xTEǏ6T�x0���BTn�ʱ!K�My,L&�
i6B �f��7�t�Ն��е�ݲ&PF�('n��"	H�)҅L*�*3
�f�'H��'1�M<?QĆ��_�"��7j�{x�)�R�����	ğ�
�O������� �O�b��5&��2B�μZD"�&�N�
�Ҩ�Mw�����'��'��Do1�D�O���+q���H!�B 5q��:a@��0�d�ٟ4�	���x���j��dx�L)��FFp����@&�m����	ߟ���"����'"�O�y�@K-����.і��U�F�i���'"e͆��ꧬ?��?I�qژ9R�F<q-,I��ks�e���iFb�M�NGzc�\��U�i�����pn����d�'w�2��k�t���3����O�����^��H���i����҈�k���j��Y�.N8�y�
�0j�$ٲfٽg+��V�Ȳ��O�	�֠�.l��+b�g*�h˗��5a0-���ݢWHT�����{Y�Dv��/c���DƗ�BT�XW$N1j#�MS�ִ{�Yʇ���O1:�����1_,l�i��_0a��L�W���A����e �Aw���E�\�^7�Z�)l���� �d���ݎ;"��pv��+9AtAQ���cd@�aB�'wª��qt|�	TFUԧ�i�i� �`��7c��P�	U�)sQ����!�y��Eaa����OC�!1P�)$ RD�?�h|ʏ�Ć�|5�'MB�'���zϚ���Z�&�R�CK����I\�S��yR:<H�f�Or���!e=�0>iD�xmT4s4zd���E
F�������y�`݅gp\6��OB��|��(K��?���?��`Ѣ�x'Ί����%G `8�Ǖ���X?��|�ݱ:���7xK�(���%ziX�"F�Z`Ͳ���[����4Tk\�IR��\�~�h5��~�ݩ*J��f1�����U�:��D��0��P~�'��R�Ư)򔹖�#eB�QK�^�yB�'+�}�)X�)�����D���!�� Ř'��e$��|��r��8�E�R����&��J��I���?��L��yf\���?���?y6��<���OJ�����J)t����- h�{R�O��+��'�
���$K�lcو�Y�9��ݚ�'��:�S�? �0b�H�gDl)Yb�S��R����O�,#"�'H���٣=� @��nM:.��`a1��2�!�dj�Z1����/"�$�	�b�ȬGz����2!�
Ul�*'B�9QbШ$�x�*ݢUY���ԟ���ȟ�� ��|���|:���6<@�iSQ��H���!/�	�Б��\����$�G�(�ay��D^|m��p������&C��"ch�b���d)ƶ�m׌�9�ўܓ���O�]nZ.z��S�=�����ؿX	n���4�?q*O���#�)���^�B|����b��i�$i�B��F{��ĭ3���#ׯ��S�,�y�ī�y�&C7r��Q�:�M �u��'�RS>�J3,:ڲ(����K��5�U�\!r�����џ��I�{(���F��p���fGx�F͓� p>��(���dY��X2 ݒ�	rA;ʓvP5
�4`�(�E��zi@��w>�3FoT�'p�p"���P�\iq��.�FJ���ɔ�M�c�i]�T>�S�-��3�1q��5�"	�T����h�?E��'yxQ�!�DclDҼk�R�	�yk�'� ]'ꉋ-��E��hI�f�^@q�O˓��<��m��|�n�Y�$�,(J\��Q�<����G�HQ��K�%yeZbIZS�<��BS�]d1�¤�$0@lQy��GD�<YΗ��TL!s�(�x�X'�B�<�4�Xd2�1J�dкQ%�` SJt�<�F�?��`��Ь�,p $Ms�<	2Fԇ'&a���*{��<�w�v�<�P�|�h��ˉ�!^P@-�n�<�֥^%T7���	B%F��W�D�<�B�#3b��`᭑"�B@�� R~�<!�፧=I���&��LZc�z�<�&̋3�$d�'�Y�$��a`k�t�<��D��;DŎ�Y�G�x�<��`�??Qti����,��3Їr�<��m7�� I��	��銇nSk�<��A>v}$5�eEφ.#B@�EKf�<���	�n��P���7��{�-V_�<97���yJq�ۻ(��=��-&T�(�̑T � *���"�����o-D�����#6��
�ڲ?Q���E'D�TB��ؑ��%����_a�!�8D�,(�D��W�꽱��R>���6D��(���oJޭiB���o*��q�,!D�DRDb����R�m	 \p�Y�-=D���cR!<�l�r�EU�qؔ�k2�-D�����ע,C�@�BD�:AF�{`j+D��Yd!�m.�}B��@�.�>���;D�X!�]�8hM/E���⦛�&t!�ݤ.�N��/�.S���"L^�ba!������N]P&H(7jɓ\P!��ݰn0v�s��rD���冖�;M!��,�F�����z4f<ۑ��97!���'F\�i�����leSI�o{!�X����`K��f<��Ù=g!�$)=�q�)�|lq��˵pT�y�!�O�ms��ە0����֫��C.X����(���(���p=��	�%!��1'�X�b�S���EuּYf �)T*Z8��H�I(T�
t"γQ��1���޺wKc�`k�d�7l}���B�
����.�	,���{tK�f#�h�d㋌}���O�I�&��c���[�
�8�Ƶ+W��,292e͜E-�,���<%�0@�ȟ/N�B@h�3��Q`���!���܇�i���U��>yt��&ml���.D��8��88�1XjNL����K�l8���h�y�0�a�/�)2�$!GɅ)JI"H/� d(��1��p=I"�%J�n�qD	W&(�(KE�|�|��c�Ůp�����l!��Z�al����"^eb�
�'�}��Oj�1D���9*����A�j���<4(��I�j�H��S���N�P�T�t1����ΗHb����A�A�N4K�HIܓf/����'�"�	'&�&ك�� $2Pɛg�W�}�lp`ve��lB&��9x���i����c�'G6pY:�kTL�x��(�o\\��W�O'Zu(�W:7��c��H.�cu�'i�%t�Y<�0!���ŉ��� ��xB�B���)�f<�(���OB�'4��C�~R�C�x�ha��T�(|�A�Z�S���� .I��1� �]��/�o�HQ�r� 4�qO�����i�df�!%�>����L���	�MS���a?ܼ� �)Ue�;t�'����ԥ��=Q|	H�@�<I���G��j��͇�t�����fCQx?�O�ٛr�ϩ*�RH��^)n,�������i����"��iO����*;OkLL�znL�dO��q"���f�Q���d�R��D̘3E|�bll��tAL�|� ���KB1j���(
�q���@BIE�LA��;[���l�'BN>���Ȁ^dZ81
���C��ɿ���¦� �jЩ0�^�������U\��DAA=I�J�0�|BIQ	J�2��KX�\�T�E
��'
@��l �m xx���X/���'��6��O�a��JM��@�Ѵi[@��p)8�$>'$}Å/��
*�$H��B�hx��q�I�x����*\b�'	�D� ,@Xyir(ѭ�h\��l�=N$����f�(1�ֵyLf���i�A��AϪ<]�Zr�w�F�X��>��~�>Y�����u �h��\�I�Pn��3p�,O��vAJ%�@�3v��9r�`b�D(>󬉪���< ���E�YJ?��'s���	��9�0t�'�H�Tr�
��F�W<X}`ħ�<&�t��h����Z��u��`��"{h�{���'����=��NE�x1�y��+L}HŞb?��u8�ƌ��T��(��FU�8��{[w/|�O���V`�)c	�i��L�4�^��,��0�H��XK�DB�O
@��I��@k�1ɢA	5*��4)�8�.�,��Q�F&@_8��G���x6C�4n(�p��&`H�>q�'ڸ��t�O��'	��` ���o�r���:Z�,��B�� B�2N�i[�Hl�f�@F�B�m���I`Q��z�j��O����O�RZ���^7h�	��n=�@!�8�y��X�E�E'�pB���� ��̍v � �* �I!��8��W�P�@��NZh&�������I$4R�A1�� �8����ģF(7���O �a��u�P ��X20�(���>f008Z�Y��$E2R�x��d[pĠ	5a��fB	���;̶�SH�P���+d.�@8�֘Y�anU������{h2�>a�b�?9��C�3��B��E�6}֭��+�c8����Q�W��[�&��<��Rɜ���ף�dd��~b�8�	���Y�e	���%�M��
2�L����15�@��Qm6ZV�'�L�z��,4��@Eӵ)2�:�}R�B�k�����=��a3��,�(չ2"�O�y��dG���O{���ߏ`���d�Jcw��Q�/���
���:
ƨ�����Y�"���	$	RtJ��YNI�1!ҜఙB�(U�DN���Ɩ��Q�ف9�����^5֠i��"O���L�u,�9�"�Ќ=t0�q�)Oְ��@���2�����g��Ep�Ƀ�B�`M�\�9�8�5�%��?��'�Ȕ��ǘ�\Er����Ȱ�Ŋ��M2DE�!�_�Z-V &���K��D5Z�Bp
	6#XP1�A6�&6Z��b��!/�p�`�9H���{2�8a@�і��5k&x�1�����/׶��B�N�6N�"���H�"0�ve��j4��i�Qb� �_������1��1X#�Z5l�%��ȋ�Z�%zu�	�uB�T�ŎL�8
����IMz�8��Mèq�0�a��P���ƌ��-H�h�ӧH�6p+�ˮt����5*V�(Vܽ��"O�%(�@�:�\���J�/G!F���c(}���?N{��7����l�>m�['�D��aF�(2�aB������*X6c�x0�1D^%e�h!9���+id���5`ސѐhC:e��i�r�X�~�#?񀀞$ �R(��B;�iG�w\�A�G�p�8�x�@��/!�$��J�h��ӒO�zA�AAP:n����X}���<jB�S�O����(�� Sp�hgE��U����'q08(�%�8	#��ԝu�(Ђ�>B�ϙ[+hP����}R��Е�Q�M<w ���VJ�i����Y5M�PTR�A%v��$97��6<ʠ�taB%@��U��I%���!dʵ	�vp�jJ�>��"?�C�<A�.L��;��MK*�I*���S�v�J�$F�_Z!�D]	~">X�w�S�h�HFIZNX���{\��C��X*R�S�O)�@&)�0vryh�G#>�<@�	�'��8�6�ܩ;\TM�G�џ?/��ʨ���b

N��z�,�?6�IC�$�/)nQ��c� VAN)U�F�(�����	�a�X;U�D�ZѢ����[�;��}J�Z��t�(�CJ,J5�����Ň4H�d*UE7�O��s��q�̕s�(��I�y`đ>)�AK<�N@�8���&&J�S��a�>+��-�`ʀMR������yI(	}����ن@
��Z$@G4���ϙ�k:l��>%?��@�
v� G��Mȗ��3���bOA"k���D��#�hR� J)`��A	�+�~��L3�OJ 	�Z������n�!4�4�B�)� f�"�I�m
V���'��xI<�x��'��%'��R����GMֹH�D(3���!_��tpS�E�0���� G��j�	�W��hi�eI�|����SAͱ(��>Qw$ڣo�^������eA����_�ʧ)c�m��V",D��G16ۂ݄�ux�IgjԀ�r��+�R�R�o��4&Fz%	A	w�,����(�R�̻52U n�-fz�r�?-2B�n>赉`�Кz
r�R��M�'mD)��i�LXWGQ������?�i��س@�t�f�v���YǬT�I�a}��I�BF yR�&�Y����[��H�D�Q�p�@�c�%_(�q��	�T���G���xΪ�XD1�#=Y� V
��!GDT'�R-���|*�̏){l�sw'6���� �x�<�Lߕgf}p2G�<7�Q��/C���v�܌O�ઑ�j1�d�R�s���),����T$FA"^�X�"O�%�T�	�`{�:b
Ҭ	��H�M"U��	��ъc& ̘dA��D����7����R���Q0b(X)@ҡ�� %HK�⋣>�01�B
�K��u���L+w2�'
C0#������,�O�}���@�>��� h�(?�$�
&�Ɍ r�|���P�~K��$`�$˧��Ź�n�"I��,�G��!/�J���d��(���6:zps�%	zZ�AV �"_�,`�7ݒ����U>����! U?~ j6x��3��M��y��.
��T�ơ�4��,X��'z��I�*���C�Cޢu�}�����c�K�!���቗t��� �1�O��"�Av8�S��&<5���$�ց|G����(U�a��Dȡ�p
�[s2�*���N:JG{RD12�6� ��ƼL!1��M�Ce�)$�E�TU&@���i�"O8��[2v��%�m�`ɔ��>O�$a�BKoZ�
J�"~RC��"i2�X�[>8�����y�<9��$�Z�V!P�y80Jr�I^ M�t�'ܰ����,Q9�͉�ID�Ked5@	�T\���g�%b�¸zⓡK�*`�����y�lŦ~S,$+���KP~Xr�Ȫ�y��ķB	���Q镩B���� #�y�VN��a���=��x�S	
��yR.���l��4'la��y�g�&�|ᐢ�Χ'5h����D�y��[X:��e�A#�D��A���y��M�R<�JS� j�^ؠ$Ω�y���
1�YE��'f):�a�ag��ȓY��c��P=(�bL���W0עԄȓ~�֐G-�tJ��Y���#��Є�
@�q�悶Rg��)H�lfń�X�*�2�T��P<I�k�%j�}��[��P���b�ޱ�ee�!'�:<��c�*�JV � @Tj���FkC`���%~��S�'ʀ}�~�t�ȧd� �ȓ+���j!������Ʀd^H	�ȓz����"!�H�� Q�)pU��������>�d�p��0c䘘��!_\���!�_U���ĥi�H��~s.y�`�#m�B�ɑcZ'4B(���`��]�ҙ}����!����S5��(WoN��0�c,U6|�ȓe�V�@Łܽ'r�6j�9.C��pD]:S)C[�<��� ʎ{�@B䉒{��=1r��T`�z/�"B��oM��i0��0[D]S��b�C�31��y�aIrpXRgH¿a��C䉆1�-pミ�z+Tt�v�U�C�	�sE��	��*�"��\2|��C�	#rE���1'W�����
͂@�vC�ɚ4�lD���q^��r&�U.�C�I�A@���G�Ɲ�`���5x��B�	]$��(��C�E�m���)	�pB䉴y!$�#���|���I�m�C�)� ,��ҁL�^[v�ROس0w���"OV�q��
*c��[2O�o�( "Oh�����H�/l�v�9�"O�	��n�+L`�FH(�(�A"O������/ь�ˣ�H�-�4�9Q"O�X fK�8� qEi�4�Q "O6�gIK�Q�HHА�ϢT����`"O�S�٩c�[�E,X�b��'����vH�SP���N�1=1�@��'��xKuhW��d�-��Y�
�'��3$ �R����쓧���	�'M�!����}N\�Jr��n|U:	�'W<8q��T6H�T4 �Df%�e��'ڜ�J��6j< ��ޕh�dT��'k
���
SW���!��`�Y��'�8���j@���|�D��U���"�'bΨ�V��3$�����D�Mقq��'�<(I��̽DE.�X�*.C�b���'	�D�J�\��2��J�';j-[B��9M�8X�D ���'mj�Re�Y�ngD�`T��(��ċ�'��`�tAW�l[aIS�ħYz�l��'��a5핾M3���}�����'&��f���j��L��/�+n���3�'I������]>��!��W�Y\�Y@�'�p�� CH�-���1ݶK�r	�'OV���D��|c�HW�B��P�'�J��D��̌7>��'�`!+wALYP"�� [�|e��'8JAqaX�E]�͹W+��fy)�',�A&��x�&�0�4C�mZ�';�-�c�+W���"� >�m��'͂r�#�<Lʖ�h'HJ�5���R�'���a7�J�o&x|���,ݪ��'0,h:�DʃZ��P�*D&`��x�'fƥ�@(���w/k8�'~J4�Wݳd��I���YH�8�' � p�@"7�$��π4^��'AD�!��16��`�!�ȧW=�u��'��S�	3agݭc����sEF�yRg�'|�K�Ş�p���r���ybս ���`�kŌ�Bb����yrKR0�`\[��OcGz��ae֠�y"�U�q.1�@�T�bUi �P-�yR�����N��D
����y���~,�
EP�X�|�6�G8�y"�]N�b�.ņ�f�F���y��z/��`vœ�;Fx��f���yR�ސ9��𐵬�
H8�D�s
P�y�`�e����C(��A�>x!S˪�y2͝e�r�� i�#:�����΁��yB�/��ǧ�2UP]��ED�yr�� y�lmK���%/�8�[@�
4�y��I}�x�a#��:��MxcȻ�yrÊ1ZJ>�14m�eGyZ��J��y�K�,(��1	4 �=W��9Bw�*�yB���y: ����JP΄����y�-� fy��+S(^�7$:��NA��y(��B��R�I�'��0��턾�y"N�(v��y�N�H_�QːES,�M���s�X�c�~|��hC 4	��s"O�x &'	�Ф�h�-p�Д��"O8e��J	#'FP����\�y�=�"O���Մ	$��`X�0?�^�b"O� �	��iX�>��q�7FI	TԊ8ٳ"O.���(t�u`�&�z�*l��"Oµ�1�d��Qa�P<�x���"O@L�1��RD(� �'D�T��	�"O�P�5�P�E����GQ1&��8Z"O��q�I�5	�T"��C1'L�;"O>80*S 1	Z�Ȣ&�s4�[�"O(d1�� &@=����͟$�28�'"O��9�B��6���b�^,N��rB"O��[��";�)�f+x�Mh�"O&)P�EMQ�"+��C�*�|1�"O M:t��$eX���s ��e-�г'"O����j��kN�a��1� �"O���� @�O.4��D��N��"O*5�"�%J�QQ��v�<��"O.��mѝx5��I�!X�lԃ�"O4͸��-h��)Th��~�h�b""O>V����M���_�Du�%�B]�<� ��1:A�$^�}P�Ӳi�W�<�f��?�^�ن�-N+l���U�<�s��h��Ñ�J$U�y�i�h�<QB�+L�80�%�s�h=��l�<�F��&V�.9D� �	��`D@C㉲t�H�9e�
l-�1ЄG�C���ȓ
�r���w"��S�^�^ld���Y5�0��+4C�0�c�
K�	��T9�UZe�U=��J�b����ȓI�QkU��-p��b&͐;�b�ȓ^i�P�V"ABX��d�.7Ў �ȓR� ]0�H���X��n�-\0.9��C4��+�&W79pv�S���w�:��ȓuڌc�m۹YR>��hƿd�:Յȓ�<��GE(H2��2F9&�e��4&*Y�we-��ճ�hƳq�l$��X�Z��6n�~B&	85��( �
M�ȓ VDC4'�,�j �F!�;u��ȓ)7�x`�Y74�������|U����R��Ԡ�,b*��ra��:x���6>8��� U&a�bEj�O�"DA"��<�Jm��)3���qфet��Ij]�!-QQ����A�=.5��ȓ%߆0��!'cR�	Ʈ8;�Je��q��,pևN�Z���P��S\�|��l�V+T.�2�^4sj�<	�C�/��ɃE�n1rYyB��0ILB�	�m��Rq���!:X=�!cǆ\n�C�	 d��S�=IƆ�R!�D1.)�C�q��D�xf���u��B�ɩ]F��I �V�l`V][eF!>]�B�I�EF$���ʘ���nD"y��B�ɋN�^Y�3��,Pu�YA
IJ�B�I2Y�ڈؠჲ6A����©N�bB�I�+4����Ч��٣Q&�"d�C�Ɉim͠$�T�>Ɏ����q=�C�#���Z�I�gC�EQӅ�8n~@B�ɚCI~LBT&�x���1�َ2[B�I:{�h�U��46�[D���
�"O����J�>��l��Ƿj?��c�"O ��&�dלű�@�e:�<�b�>�����H%z�dD[�+Űi8)�D<%�!�Ѱ=&�� �K��Dݤ��ż*qO����D)5Ud�YuA�%��4�����4�!�$�4��Y�$�� TN��OZ�!���5.:V�k���J4̘
���'!�!�� ��a�C��U;���3� ��^�"OTZ��D��9�a^�'/���"O�HI�LՁz� pv��)t���"O�[�)ęS`�PbseE$3^�x�"O��1&�EP�SN>Y"�xY"O"IC��2Yf\�;���/F�p�"OD��ʇS�|�(�Y������-�S��\,�����Z�n�*&)]!򤗂3<t��Bݴ/(�3�� 9U!�� �^,u�șe.T��"ڰJ;!�D5O5���w��o��R��)!�D�`�T����?#���!�9 !��\�>���rvDQ
h��D <;�!�$ɉ眽YaL�<w�p@3`��!���	�p��4H���H �Z�!�$̀:ͮ�I�,��(���J�(H;!��
'qD��bO��
��P1���l�!���k[��fɓ�Jv��B`��!�L�J݈�X��A�"���H $�+G;!��ƕwK\ɴ��IMhC���qX!���ʭ+$g	9,�Æ"N�!��6K���Rѥ�?Gj �D
�!�@\��-��,@"�1���"o>!���vH�1+�mĤ D5����"!�M4�E
�d^�r�T`@+Fk !򄕽(s>���.��S� ]��gǥM!�$Ŋ5$�rgQ+�4@$�
�!�$�vr��I�!K�y��`k�)ڨ<�!��6pت��Ҿ|aܤ��(ƛ=!�d�"Y��d�C1�p)�5�8fk!�;eBX�A�Ə�.2p�s��T!�DW|��2j��5�T��D�n�!���;At�p"?J.-kSfȞ�!�ΌP`d�KP��������5k&!���7�F�8���>���q�n[-�!�LS�Z�z�*C�ppǢ5�!�D��
��#��k�H�+��V��!�D�"w�n���#ļ}q\��R� �!�N*����l��mYn�ÉO"!���(�1��� �U;^Ԋ��A�3�!��ղY�
����72�)��bQ��!�A�}3�� ��-X!�St!��α[��8�GH�H���dAM.�!�dU�+�V-0Ug>�%k��n�!��>e$�d���F"���I#m�!�D�B�^83��̖C�!+J�mR!��V��� �.���TJ!�Zd�؛'��M~ �[h9��"O����Ir�L ��ޔG��D�$"O�3�kS�dW�h�3��"QR"Ozb��X�2���� �*&%a�"O�y��a�1�`)y��9L �!b"O�x����|�V�c¢PF�䥊"O��T�Ö��Q�`Q�bd:�"O0��!�.�ܸbo�B��Iȇ"O�� � �
� �{��,Fz�Cw"O��94�ʁ{DJ*6딻�j<�V"OXMKPa�o=+�~�d����y�i�8[8ĉWȝr8��ЪZ�y�Hr���X�G��ng��Z�d�=�y��ƴ'
<!�㮕���DGf-�yA�dSF�C�Q�_����[��y�GG�.K�,2�iO�@R�%O6�yBeL��:5��&.�6�s���y
� �D�p �3/"��%gق8k4��F"O`�R��..e��fƅWn�@r"O.9b��T�X��0gZ�� G"O�-�g��!��Y��J0[O��J�"O̥�@�!�6#��@�}��P�3"Oj ��fңlw���Z�ǜ�j�"O�HiU!1UTP2En]�ӨAb7"O�E�2k��nE��J��Z,r��"Of0�,U���/ğn6����"O��U/B<��!:r� \r���"O&� b���j���+�D����"O�L1���U�bo�P�T(y�"O���9� ]@�N�&H�TSR"OŎ;5���{@�ō(@`�"O\Xc�ě�X��@2�ޙ8���+v"O�|�ʊ�FB���NHJ;Ҵʕ"O���$�V���c+�>'��҇"O�i�2oԼY�n1
�I�!���"OV���2��H�Ɏ��1"O MC`AM�rk0lAb.٣{��p��"O�����y�:A�L����{"OF����.gI���|��D�"ON�R��0(vȄ�BM�� ���V"O&$j1�ӕO� MC��X�, ��PD"O�d���K�gR�dB2�7�X� "O��*K�-��t�pl� ��#�"O�\�7��hZ=i�jo���""Of�%+[�-��E-Ł�"O�p�r��5�P�s#��y�B+G"O�%�*�41��%I���HF0Y�b"OP����^-�r����XX��W"Oj'��nɎ�q��&zG�8P�"O�e6���n͚����0o��Y�w"O(��X�O �xP��4^��8�"Ov`r"#K�P��M�u%�/M���� "Od�Q�l��`���@�8EAp"O�͉���I����b��d���K1"O�i�5(��1����<u��\8 "O��* 9&d�A�!Ѓ@�X0�"OR�kVhġ�d͋Q@�x<XcS"O�%��l�;����Do�:@�@�2"O"x
qㅵ
X�uC'nئ��=��"O�y���Z�wKb!�7K')������T�W��5(�إ�0g�u��Y��gId��$�-٬iz��ҧC�l���NS������QEH�����.b��,��,��9���R E`$߾p]&��ȓ~��iv#��7 �yE�PZy�ȓj��! P��h*�u!6 :!�ȓRF H�UIQ�L��<��n�4I�"ل�]����ɝ�+�0� J��>���ZM�Uk�̸_|�;.Ê)(����%ྔX�N�9 $���Y˶ͅȓ\D����&0����F̅=^�܆ȓ"�=�hKld���W�����^�Ld�"����({�~M�ȓdN�}�')ƫwI��iH�b�P���G�F(#����lj��%tJpq�ȓXKڜ��ϑ�,��r#��*,�&�����1[&kL
.�IB�DM1P7���ȓjW��b���5�Ќ��� d���J�@;�H��İ!�:\h��ȓt��="�k߽�N���^-Q��%�ȓ_�M9���>|(	�FmG&����S�? �0D�-V@8�3 }�Jy��"O�)���I�KH:@�0-k�D�"Ov�R�ׇ�t�r�T�|q���#"O������`	&��_����"O�H�f��УP�V���q "O��1C
7\���� � �aa"O �JaJ�%j��j�H8
��u"Op�A�תU1�����x(��w"O��TH0��d#��zL|� "OVe
�B��$�T�d���p�t�c�"O�DiV@�(�*qi�<,x���"O�;�Ą&I�Ha��>K@00�"O�X�Vh��*򄴒GG'C\���"Ob�+F�V�jԤ9�Ň�oR��
""O�ኡ�U�v��0���3:RI"O�E�2D��%5ܫ��_�2A��"Odt�'��.x�x1U�w�@@J�"Oj%�B/�{�hRe�,wG�q�"O@|���
rq���X����"O��*�%°!���%��)2F�ʄ"O~]��$m�ec����2��"O^ܙՌ�:;�)��Kӟ(��{�"O��1���
�Ò˝s�.��F"O&|!r�Z�z>dy�@M�C�v��w"O��5�H���c!�2��\;4"O��g M1	��`pv��jK"O��k�*��ٖ�!��T�:���*�"OD����D]r��C�X>�%���y����,�%�`P�:@j���
��y���eȦ�p�oϛ;�رc3�3�y�M�g�B@ �$�bFf��r@��y���v�f`��护dG��A[��y�-�8��{f���_�1�bdL0�y��u^�=��I
-E���3�W��y��X�IP�tATsߖ�X7BH��y�ӛd �@�Y�vH��w���y2l�h��Y�dn��ZqV� ��y�-˗m�.�r���5�4M+MC�yb�C�ia ��A�=|��I��y�O��h�|�{T�Y�}�͞�y"j��#�m�U�-KQ1�
T0�y�� �w��,KD�M�w��H��F��yr" w�v�5j�j@��̌*�yB��d���c�w ���F�E[@B��0w"}���[�62V���,��"�B�I=\ZT�0�J�Y*fIsa�ߖ�B�I�Q��y���e`Z%ɰ#�(B�	%�.1���#-�T�����>u�C�"
,�1�B��w~V�a&�;d��C�<i���s$�,&�F١tH��KP�C�	o��3�-=3���1�E)U�`B�I�`6�L�h�2gJ��Z�(��8B�	Ez�SU�J�.�|D2AI6�&B䉸=|PR�B�Pzx�*�9IK�B�ɗ��Dy�AW�kf������O2�B�I;4���Rq7X$ڃś,a�nB�I�ˤ;��N!J.\��Ζ= �
B䉜4�:�Nהv�f��@��Z��C�Dh��:��'�0� �)��B�I�
������6I�� #okvB�I-Y�I#A�;=P�1Cq�^�%'LB�	@X`�y��ށ_e������C�	�b�~}���r1���@i��B� J���g)w*������}C�)� F�z�5��� %��/s��U"O|��q֟D�F�;�#�0J����"O��2��V%-�~= 4�
ڸQ�"O�8¨��U���&b�:]��"O`�Q�'��j�VK�5�T��v"O����Ո|V��k "w��"O }ۧ$[�#G��K�1LrN�S"O�hI�kY�al��Bw��4��P"O��E�3�T9�A�҃yX��"O�@�3��T�Dr7흭dXb%�"O*=��^S��}1&�U`K��5"O����' hA���V��<!`x"O,��@օL���H!hkʤ "O��yTƎ w@�i�:`�q�"O8)[NO	z�vQ@F
v]��"O��5�ÓU'���dQ�H��0d"O8I�g��
F%XR�CP&N���@"O�ȩr,Yj�
�c��fa��qG"O�A�BcžQ�f�(5�S%{ �"O�U��;l�B!��-ߒl�8��"O��3��^��(���T�Ek@H�v"O|yX�/�#bъ�Ӂ�-
v�Pq"O�t*v��4(�
�-A9a���c"OS��
�[\�`#��*j�ʀY�"O&5����1U�������E��@�"O��b6
�~��a�/D:-�4�I#"O��RTfآ~J�]���з.��y�b"O|p��!)��8��$����}��"ObQS`N�RO<��%^�f��M�"OP`s���z{4qӧ�������c"O:q�DAZ�`A�4��6l	��"O�p �:*�`3 �N�W�9�"O��NE�{qu�M<���r"O�����"H�PS�
.2���6"O̛砆e� �`�"-lɂ#"Or�;�-��S/:�KW�&��l1"O*PK jң=��9��V�Pm���$"O�5Sц@�5��1��u_�\	�"O����!��Pr��87�!+3"Ov�j�
 F�Z�!� &�C�"O@i�w�Qz��%��ݱ<�p�"O�(�B��t��/q���!)_?�y¯��h�y�d��s<�KѨ��yB�@�Y~$�rbeޖ5�2�iq�F�y2�I���@"cρ0\H�� 8�y��x��q�7��;q�,Y���)�yrő�>GZ��ٰ�ԅ�$ݝ�y�B���%��A�NHtd��yb˓<1e�2j�J�A1�Z�y��y�`��a�&| f�� n�/�y2�[=���l��o~�jp�0�yI4XXҴ�H�ؚ�����y�G��R�&ȡ�tb8�zWF�y�jR�Q���E�"��U(�+�y��ڶqR^4H$"7�$\����y��)>��-8���<x/�4XbcĘ�y�,�71��]��`�:�Z`�C��y�		�O�� �V��R�L�I�+K��y��S�(���,CC��YG�B��y򅞳c�t��� P*4�Z�o�>�yR�˙�Ԙ�LS5E����y���#[��`h��)��q�V��y���^��84 �?Pe�ak���y"o��h6����]�@�ƈ�0H���y
� X���gլ�x��@�9S�� 2�"O>i��"�	��{5JAP��(�"O�Ĉ�'Z�M����H��UC��S"O:�)�Gխxd����ܚi@m�C"O�}��c��j�iw�L�]6��q�"O|M[�M�b>�]�1�ZVŢ"O�����I�z�8QC�/ck{�"O�U�΅�^���!`��84Z@0(�"Oޝ@�O�n�8"��y=e��"O��
��P�K�� ktnP�=B�:�"O�� �-R����J)&(�9�"O��;�EލMƴ��g�~y�"ORȫ��Q�.I��&A��v��{�"Op�GC8E�r� �`II�8�"O��C��V5��J�� 9�(%�Q"O:)��Wu�J�@D�����"OTH�SO�|�B�ŃxBa�"O������P�bdqp�0Zf��"O&T"	U��"�)�(NixY�t"O
�Pb���'\8؇HX2��m6"O�]�C�&:�5HϾSz]A`"O(B�J׀TUh24'L,\���"O�\��ēLW<=�d�w�X��C"O�h��o��V|�Qb�CǱ;Q�}��"O:���O�8�	`rL=<��,��"Op��Rb۬Z0���w�,!����4"OF�A*V�0Z�Ԙ��J�J`�E�"O�� ���$C���s��#��W"O*lce96��#E >HT�D"OX���ƙ���D��N��	�P"OL��v�B�q9L��@ѽO~�j�"O�4B'h�訠�n�v:L�5"O�H��G98�F�Z�
I�)
��g"O�� @�p��j7�	3#BT�$"O
|��.%Jtp�AI��X0ʔ"O|	������C�K�8�y�U��yBĕ	~A��#nK�<nZP��yr��,8�V	��M�3�`����+�yr�^|^0	K�æ(�*���[��y"-Z�;�@4+F-Џ%�d�d��y�K��-�'�Y> m]U(W.�y�	UX��(6cEl�T{�!�y�E��2�QY�����yp��4�y���&3elp���&�203wdُ�y��G
B�p4r�A�X�@[����y�b�	X`5c�:M��%BO>�y"H����2�ʼz��^1�yء;��� �
7:�q2��y�`_c0qg��Y*�< �
���y��=&��᪤�Z5Y<>}� Cƃ�y�
۴2�~xQ�D��$<<y+�K��y"�.ml��ʰ!"���TF�5�yR��("�8``��)*>�5�scJ4�y6i���p�aĵ��U"sE/�y�ʖ	<><r�oF��(y#�b� �y�̘<-~�v��,D��#U.�yrσ�M�p ��Ս�����y��$����+��d�x���y�*��i�p���.WՌ�J4��y�g�'49X9`!-��T�D�� ۷�y��гX��)P�*dT�ȣ���y"�1ϮH�a��41�XЙ��@��y�F�	l��R�ޚ_�I�R*I��yB�N�
�{C�	@�؀rb%���y
� 0;�B�`dD4��I8?�D"OnM���x���;#厥X0�ęc"Od�ӤD�DK�y�RI׺H���"O�(��+m!��UhL	��`s"O�Iz�	ɡ-���)��Y� �Y�"OF�R`�p���+k��"a�/T!�N��9y�(�
N\��ROƿ~K!��JMj� c�:�����:>!�Ř1�4���P�W��iS�JϹl8!�DT�m=��EC��:������^�]�!�d�>�*9�Ş���a��'�!�D!n�
Y�s�޼
���p٠F��C�Id��ّe�T���#@�v�dC�I-?��C�+��g��u0E�T�R��C䉮C���lE�n��PY�GQ8LX|B�I�ڭҁ� vXX"��&_VB�I#F� ��V�5�4Xi`+Λ>�@B�	\���S�N{ `��z��B�5F���P�f�,��Y��e�1ҠB��t��)�L�M�ֵ��,��Y��B�ɜC�@��Äzh�Y`�`�,B�I27b�����ii��׎�@4B����2��U8�pqp�J�QxB�s��5��c��y2M��N?G��C�ɟ�\�r��2X�ɂ�S#�B䉻g�Z��n�:��Ā�j
�}[bC�	�G�h&��X�<��ʔ?E�B�4Q��9�n�M��`iB��� C�ɸ:�b)�b"o���g�B<'C�7B��i�gI�f>r�
�Hߥ(R�B䉿?��t��b�e��w��~��B�I"�m`���7R
����72ܼB�I�8���r��.oO&H�T.G.!V�B�ɩ/��5k�J�Jj�%�� Ŏw�nB�3_ʐ��>\��x֣C
U C�ɀ~��ʣ*Ά/|8�D�W�%�(C��5bŰuZ��_  ϸ<�G͖=%d`B�	�Q/����O8\���8��O5U��B�I52�<��M�<1� q����q��B��%�>�@�E�\�P��Bɽ{+�B��#	u ��� �'%�8�@��$��B�ɻ:`�YD�@&JD鶉سNjrB�'j�F���A�"cxa;�e�({�jB�ɪ4Wh1� (EF��]��%��B\B�I�>�rR��S�����̞�lC�	+�>9�W��}�z�a�)�VC䉪Gw.����@F�Wņ0#�4C�mo�A9W�H�)ȵd��H�C�ɊrF���N�i
#�*kC��l=R6�JU,�GiRdHC�IL�Z�#���wƔD���5D�NB�I�~oT-����)<a����Ο�/�.B䉷%��Lp@DH�!ްp��B A�4C�I#,�K�� ���(2&C�� U��Ee�O�����.���6B䉜"��@��!�x�C#"�!Q4B�	a��̲5L���x�/�5HmnC�I;I����B� B6�+2��5B�	"&�%%��-& uHf)ҭMC�C䉭_QB����T"MA���jРg��B�712�h	�iα?|�`�F�<Dg�B� q�$�h�E�cN%Ks�_DB��#]�>y�c畕L����S7T?PC�&A���F
׈|�ԃS]!�B�)� �Y1h݄U.*Q6��"3��Yӧ"O��S���O���B@Ʒ4���pC"O��ȑ�{�P1CVN�����q"O�P���!|.Bd���M��xb�"OJ1�"��8���kDHK�d�V9��"O�\J��HϪ�Y&U]��$"O��#��Ȱ�b��L�(�"Oz8A�,5^d�O�O�	�"O\��,��q|�y`N�� p�m
�"Oq8��\:
sTt�,C�(�(�"O:A@u�#X���@�n�m�LDa�"O���!J�9��������.�"R"O�%�Rj�5�rD�F΀_o�q�"Oz`F�5b\�bJ�Gw�U�"OZ�h���&'Ʉ�����+D5��"O�4:A�":E��*�gP���"O�`���X6\:D�����.>��`�a"O ,l�����N��{��C-D��S�̒:{zʆ�W�zF�i2w ,D���ѡ�t���F?x�*ۡn*D�<�F酤m���JaG	~��S(D�8Ç�Ě+����D�4w�=�G�0D��z�ʗ�c��������� 2D��a�	U�G.��2�#l�e��1D�����Ȩ?}��v��b�[�0D���sJ�?E����s(]E.�9�g-D���B/�4/��H�� �T��7�)D�����d�ӷ�߲	 9z�%$D�b�,�2��=b�c6!�V� �5D��D��(���Z!��7F�BD�6D�|Y˹ga��c�)}z8Ɂ�	5D��p�W���U𵇔%:Ш�V�-D��ɑ�!�<�
�Ѧl��[��0D�J�˃>�����O*]c�QѢ�-D�����>p�r5i�/ĺtx�*D��R ��5"xT��w���J� (D�Q�]�{NdL�@�!e\��$&D������\Y}95#�jx��F "D�i7'G%{wĕQ��LD*N�!�B*D�Ȃ���4��`�h��V4d`��$D�\����0ybWiY�f*@�"D��h�ꊋj�1����_C�v	?D��2��>��[re��K����=D�h!*�)p�C �sdM!0�>D�܂��ʵa��	Y��69Kpm�U�1D�dj�
܈Rf��ҥ֒Og`Y9Տ0D�l�"lVr9��2Т��"��B�!D� j��
�G�4ӷ�E�$�����>D�P`a��0L���W�3���;D���Sý
�\� ��&}��#�7D�@��hU6�г�є7b� �s�7D������C��9S�H�!���`� D�8�b��E�)��^;%ň�rr"9D�<P�MW!=�>�%_:K��!,D�p�G,`��h6ț�!MT� dH+D�{Qǡ*�{V�o��$*�4D��)aӏ%	αqM��T����+-D����hR�`i�*U%�tL6I,D�� PIt<��	HZ����'D����
oVP%�IF_�d���'D� ؗX�S�P�3w�>hu0P��o#D�xx��ӃX�ɑ �L�N��"e. D�x9�aA�W� C`�S��\oVT�<1d$�3M��,����c�t��j�h�<� 
�jTM�*N�0�vdC�K��X"O@���d�2!w�y!�c�0=d�b"Ob��C�E�G+��H�aϕ.G,@"O���@�U�^H	b0+�"2?�E��"O6�)Eǜ�YX����H�<A8>��f"Oi$�<6�P�K#��6�%"O�aCHǽ���
�,��j���"O�D�C,̀o�x4��	Z�	z�"O ����7{� "C膅\���Jc"Oڣ��!5	�p0���*Cw ���"O.�"p.T���3F���t��"O�ț� �=&'(U�� ��w���"O�ɖ�3�`,�w�P�\�n�3�"OV틢�E�U�.��WAM/=�4d��"OH�P� iPȄ!��Ĵ��E�"O�mX��[ 8xg�N3O�<l�u"OH���E��8�~\�Q�K���<x�"O�����ܭ6e�2B�R	U �a�q"On�!�e-"����R'�(ȈT"O
%H��	;ɜ8�rc�2~�p	�"OX�!��(�(�ae�� _Z�"Oٲ㋍$�^��Q�Y9\^H��ȓc��1�S�ٽd~$���J6x$��ȓ;Pm2&̉�W���;� �9e.���ȓv��`�A7��d�K�^�h�ȓD`P��OP�h$ɦ��;�� ��?U�H�E-�	�NUY�C�v3މ�ȓC� �A�Χ�$�HF�!���ȓ�h�K�V�@5F�9?\L	��z84}`�^$ng����P�I�PՇȓ4Q8�Y�h��a�E��
�47zhȇȓK���%�!����cL;r!<��r��Qi��'_���)ȫ1�ॄȓ^7>-�f�s� ��a��XYɆȓ$��Z�%��Z�	�Q%L��̆�u�^U��['D(�G'�s8ņ�"�xtqȋb#��e):/�݅ȓyȹ�Q �zP��%G��Ν�ȓ>k�C��Y'r��q��g������ȓ<u�����,�ڜ��� N�y�ȓG�:�#Dܚ
=��"�ⓓx�,��h�N��q�� ?g��(��UH����A2F)��	��!��0��'"�'�l�j�	N{n(��C����h�'�
��&�O,a9tᑇ}��x��'��A�OZd�!�$yV��x�'��5ؓ.ϡ
Ô�#p�ΛY��2�'�|��U��BAY�d�W`Pix
�'���#eD�|�tQW�Z��~-��'I��pK�+�Z	ҷ�܁��A�';�X�.�aE��ipÔ�T-Z�'I�x��ȤU��`�����'����e��:,�H�ר�|
."�'B�@��*�)$�0ҷO_�m�1��'C�x��o�W�X�&F������'ApqB%*�q�Q�Жhԉ�
�'ON �@�h�N�á`��F}�
�'����G^�^���B�O�:��e��C����eX�ޑ��酬n�z�ȓq~hdB#l��[l�Ǡ�>vv,t�ȓw~lmY��?V:t|!�

:EK�H��Z���z�-JdM$���:|fц�1/ҡ f�P�h�ܨ������1t�(	t��=g��0A�'c%���S�? �UjF��s\��ġZ*�
��"OR=��BG ?��0�7`ąx`�"O������jexJ[�*vʅ��"O�]�T�I<TZ|8Y!�Ԣ%�]��'�'��)�3}b�ֶ�Z���KP�5�v`���)�y�
ۚ>��r#�Z�^L��(�y���m���$�N\$�xE��y�R0�A��
Cft���S<�yr�^�e� ��@�M�ְ���y+�99� �h�㜾B��hX%� �y�nK�4Wy�ҀM�$�bp)U!�?9��䓆h���-p-T�.CjX�D�B�5!��c>茪�&>6�S-� U!�$Q�5���8sj��G�J:G��24A!��ؕPP��"	�z�ճ�Gˤ&!�D;T"��3-�9i�%�B!!�$��:|�,d@�
t5���˳0!�;����a���*dɣ���!�Qb��P����!S"��Q"OJaa"eԯX钸+P�V�p;����"O�$0���)����1'���'-���4
���0�2�U�R���3�-D�4��o��$��6.S@*q�R�1D���C(�)Qd��%Ƽ�$u�V�9D��s��O��0�D�'��)�',D�����F����3���/���P ,D��P��3D��3P�����G�*D�������hB�����K�)D��P��>N���@�=BEɦ$"D�tCu�)F-�tiâ]0Y1�08� D�໖ON�$�@N�X��L(�E#D�̪P˧~D@��d�1'2�b"��O��=E�ćC5d�B�a�%Q&�-+�C�~!�D�=�V��BEǄx��ƭ	�!�Y���'e��pq�A>u�џ�D��Y&|�|1��_-ax�3`���y�`R�4��@K� A]����f埙�y"�H�R���YT�� ��N��y��r�����)�"�
x u&���yB�KR1D�r���R����ئ�y���:��!6D��ȱ1�
�yR=x�1
�#�
���!�$��OL�$!�'Up8`�S�7e����z%��a�p�S�Y0"��V�-m�XB�IOVԴIc� �3��U:�G��)8B��*GJ��p�c��Q߮)��K� \�B�I�%CfApB�K��� �⋝��C�ɫ-2����Ĉ!2Tn-سhKUȢC�	L=�5H�-
f�ȕ,ĺ*���d(�\��A1-�#�Ψ��
X)<T�ȓG��8!7HEO���G��!�T�ȓE+>=����h\Y��t��ȓp�P@�I�[�b���!��NYx܇ȓ%Ft*� S,�LJf�B�-�θ��IO~��z�8�{M�=x�a.���y�$$c����]?0X�Wn���y��,޸�� 7TR��  �?�y�N�u��I ���|�E@���yb��(��\�D#x& �8g�5�y�)�7��8�Q$&��Â��d�<�������E2lj��Ԍ5?���)FV�On��D��FPj3���4)�HZ�:T!�dV|��jd#[>K��x3�*M�BF!�$O��(�
���	/R1!�� �i�U- �6O�0F���8y$"O��Z�e7Hbź��W��3�"O�X�!E���Qd.�(�.kD"O`�
F��9
L��̓�T��Qc"O�zt��'L*<�Z�M@+(&4�Ru�	�����"��#	35�śOd��Qa�F�?�)OB��Ҕ:)�]��ϙ�Y�>aH��[3K�!�d5?afUYH�0G����`
9o!�I�T�(D��N��5���U��	tn!�¡�HP��d��\�H�P!�-�ў �?��O0��gT&z�d�eoϘx��P"O�E�!�4��tX �Y �� ���'@1O0!��)*5a��R%���z"O.�w��&���	�o���U�1"O��²/�5G�9�N�|��TY�"O� R���M��pd��a�,�"O��ę@Y2|:cCD�)��zR�'aў"~2�뜋;�hrƅ�j��ņ[��yL����� �b��it˛���O����r>	�B]�oz�$�eC,}K�����OPC���QW8�P
�? ��%JS(�4i<C�ɴ	��X�D�s\�����͂�0C䉶m@ȼ��,��W�FQr$��;��C�	4+D@�
�S6B>�y[@ą�_��C�I�E��	�t	ï"���AB��C䉍:��0�u-���;G�@;�C�Ƀ1����k^�(�ms!�X�C�IB*�i"@��re$�K�K�`T�B�,Lt��i�V�(�BkA�G�7ΠB�I�LJ<��"��8Iza!�Ʋ#��B�	:5�m0�$J��Ny$��r��B�I:v!�@)��)%�p,�1��C�:C�!oz��X�!@�fH�x W�4%:�?	)O�������G<=;�g[:!�j��cD��?i���?)�cƊ`�3��e�,h34�C��؆�1����&�2�E�A�Y��i�ȓC���0��j�Q�#�}ݸ!���
�� .4����p���N�������<9�ǈ�<�z�rv�^�c�^p��'GP�<I�K�%�R�� ��R��"��H�<��b	k7 *o9X�x�(\Gx��Ex"�p�lY��LI�M��E*��y.Z�,� t��-�ư "�T�y򨙽���x҈�;c�i(��X��>��O�E���y�&@�U�Աy �1�'Pў"~��.A299�RbID�ZR`"��y�EJ8XTU��S�p���C��O.˓��$p>}�U@	9��3PS)8�`�c�O ˓��*�SZ��]0{g���ήXw�(��Br�<aflˋ$/*<��gi�p�@���B�	
)`��Pe�Mx��U�І*��C�	�/���a7.ǹ;��a+�i�E0��O��=ͧ��䙲O�T �hL �XjE�$y*!�$E�f0���e�%5f,�Ё#V&!C�yቭ@i��R�����t�OG�D�=!	�'`����#ő�U�\�i�L�J���~�tpڀ���N��.��7}���4�%"6�Q�{�|\@1���X�
�ȓX\��PE^9y���p�nJ����Q+�չ§W!�h٠q���z��ȓ!BnxxV�E=� I�b��#X�4E"U�|�'���4+���!�3$[�H�%�K�)5�'r�)��&H�Ā���4l�oN��y"�Ї Zz�ɱ�$�0L@�h��y
� �U)�oA:,�j��`cɟc7<�"O"I�ҭ[�Rv��BL���\v]���'/�O�c>�vɃ�aiD���)��D|z��sH$�IB����m�8j�"��$��A��łEG>D� )�B�,-h�w�]� ��[ ;D����̌��H��J[�|���X�o:D��Q��0y4$�B��u0tU�@&D�<�P,�=`f`�����s<!�7�'D�$*��Dj%nYy4�0m�����;D���I
�%kC+�h�[�q�!����QG�Y�}Ke�Џ �!�P�#_H��f��,�8<c��\6J!� �	���pd��+1�v�����e�!�$�!Gm)��X6+l4zӬ��0�!�d�0(�Q��Mq��c�Yp��}◟ЛP��B�Ԁb���7T�T�sc�4�Ir�����x=��"ӷ (� �EbՑp��� �N�h,Igo�	)Cv��s�],�l(�ȓ�@8i��G2�PP�K�$god)�ȓqR"@���\Hx��Q&}6걄ȓy
� ��{l�Q��tQ���ȓ%F�����39
5��& �J�h���Bj ۀ���
DU�#ML�t���?����~�Pc�#	���1"c	�T���C匌]x���'��I�1��YP'�$MUN=Zd�[�<{B�	&F�n����-��Yҷc����C� ;\<�ĩɳV�\Cx0B䉠�AzRɎ�wԙ�#�'|F�C�Ie�aC�ݍf&��ɥ P"-4�C�I� e�����_�OVD�Q�.I����D-�	����h��4��s�*(v�8 �$��,f�0c�'�p�āN5�ܑZ���?W��ك�'C,h2�e
(
�4��J�U\��'� q0D�'T����Fb���x��'ب1���L�=��a�!�
�'��Ÿ�'Y;	 ����Bp�&ĸ�yB�ʹ6�Th
!o��s�f�r4���y�f�;��Iӓ�˽8�	3h��yr��az��e�4~,��R�!U��y" ^�m7~�"5!2r��ѓK���y�cQ:|P�\�DlD|'����N��ybAӾ0F �3l��i��AЈ�y�,#o�� I���7b���$�#�y�芈+(2���C�0�Ɖ�F�\�yBl�<J�
 Eć�$^P�(Q�y���t)8���N�<Q
�H<�y���>�z�!�ы{�>�񂈘��'�ў�Os���o��dy������"��1
�'B�hOU��� 9C����< �	�'�0ԃǏp��4bR�<��'�L�p��Q��}j&bG��Ҙc�'%31ǎ�8��� s��d���K�'`�����۬|�"C�8���D$O��d��b�R<�6��8{ ��H�Il>92�BY�7�v�K��ǰ,P5�F+4D��z�*�!6^�bЈs��Y�B/D�|���Nu���#�D���AAcd.4�;G�|��u*���p+d0�/^_�<I�!�@|��B������æ�Y�<a����3�$�7ȉ6���8fN�r��?�
ÓWW`�q�
�S��Yc�nY
}��9�?ٍ��~��E\j.�%����"- Wbv�<q��/p�0�c���3#Bh���s�<�C��'%۔�`#ѭR°���]p�<� `"�?8,cA�Z1� ���"O.���M�0�f��"��:����"O�I�r+�������Ц�Z�"O�j�Hлc�|���!�`@A��}>��n��3&��y� ��"(D��8�_�g�mB�a���9��%D���a?���3TlE�<NN��&D��c�CI�N$�3�W(�Nl�t�&D� 鱏�2[G6:#��0T�2��.$D�X)�cH*A�)0J,*O���&D�`��P�v��p:B`L=&��ha.#D�p�'ܧ*2��j$�K����yc�6D�0��H�(QNi���.k_�H�p1D�<�&)B�| >��0��$ �d ��.D�,�3'G��x�`ʭ^#0 �9D�drBF��@I�����Ȳ1ܝ��$D�����:ky4=� �B2l�:�i"D�ت���4H�t�r	�7>!bP�?D�X�SF@�V�p����z�F��� D��`�⇏tN��R�;B���a�<D� y��
 �����D�%V
��Ć9D�T�d!��fî9�v(�5o(�D�2D���BG�c����1�T0@�*��.D���dY�F��@�I"6ĉS�-D����&H!P�2Ts���	�Ʃ�A*D�$qPbV�I���p�k �#dhX� "5D�X�g�U.U$ ���\� `�0�2D� 2��-��Tвg]3C��-�@�=D�\�@Ӧc2��@�[�rpݩ��<D��B];z���qm�U�(�0@8D� pS����Vi�@�U�.�;�c3D��"��� ׸Q �F�	�ȄXTj4D��X2�(��TI�Å#;��1��0D�T�F؄G:T#oo"2I�c�.D�$�aIH�zڵA�DǹS���s�,D����QѺ�S�I�Wp¡�F-D������3yW�9i�ڦc;X�cF-D�0V(�D!4�J�d1cڑؕ#+D��ؐa_tH���`��o��e:ǁ)D��*��"iK�h�������{�l(D�T	��T�=f�$s"!��-����%D���G�Y�~zԻ�(&��#G�"D��s7��	ob޸@�mR;�0��M?D����DR8�賌BjS�P�H D��*�o �v�]Х��3�ny�!�"D�|��e�ez:9���2R��'�!D�X�V��f�@ɗ� �k��iR+!D�<ⱥ�U�\p���5����g=D��Yv�Π��kUm��V���r�8D�B�ֽ	2���8f�"��uC#D��k&�� ���c���?D��YǉO�M�R��O.��1@i)D�0�W'�9K�bY �	ԩ�4��'D��B�c�>U�$}��h��~�[)1D� @���V�@�+[)*ءC�1D�$��"ĭ)�B�Z�Z0h[��c��-D�c�⟭>d(�Ԁ�$M�5���+D��(!�
�,���q����4�pc �*D�d�����C����(M�q�Г3 .D����ΖtOLYz5`�<|Q�xx�*D�$��L�a��	�`f�3@Zhh�a,)D���J�$@� ����%��0҆$D�d �O�����7 �ql]�c(D�|0�#�l^}���y��A��1D�� �}����,D����L��D��"O�� �KEr8��E�P�d�W"O��a�q)�)�`�:NE�v"O�{��W)?Кi��9N��	�"Ob��u�ݥn��HB"�@�a*ݪV"O�b�Eԑ�P��RM˹7#����"O��)#��^%J4aP�K,k��$qV"O^�� ΐ�G*2Ugl��:�"O�a#�@͞d�t%*0���I8u"OPX+��#Ȍ%�q��cD�:�"O� I,����oϪuG�z�"O]�V�W�,~�!UmX?!���#"O��#u��^��a�� E�"�j�"O��2�D҂qSf�*�
ɟ��a�"O�P�d3��AU���jW�t:1"O�s� R�̬�!�R�/ş�ydF�i$t���&�|��Ӂ�%�yB�".�(�5&L�v�v���+�yb��.������:v�B��b���yJa9��� �ky������y�� 4���q��2k�>���^�y� ��1��1�R/߆WrL�x�*�y���=w7t(:�熭K^v	�b �y@	)E1�а#DI0*d�e�1�y�A����ajY:$�IC�[!�y�,�op�t�Á)B��3�bԓ�y��If�貰.�s۰�����yBf�>2l���N&Q�LO�y���f�Zt��%N� �]S'e��y��B�D�y�H|�,��f)��y��!\D8%艶zUn	S�*]��yBlΔ.�H̰� �'sB2��TW�y�DΙA,�)�M�go��sћ�y�ʨ�T�2���c�Xa�Ə��ybS=Ky4 �Doƥ]yLD�R(���y2�@�3򁣦dA�B*�Ђ�X'�y�JНk=����˨:���w�4�yb��-f�T�t��0|~�x�L�y�NL E��8A�f	��&�Ό�y�N��+n>Q��b�C�<	�C���y���<;жt`�D%@+��z�c�*�y��0S4)���E���*ìA��y�`Х�2X"!�:rJ��Q Ǿ�y�E�3L^~)Y�DTSd�u2�D�yb��*O�6p�`K�Mp,�@@��y2���X,Ld�c�ȽE 6i�'ʓ��y�
�w$+�z�h塅��"Q��m��P္�Vȗ6Di� :�nS LZy��=�}q6���]p!i�%�}��m�R�Z��o���Y'bN
$Ʉȓr���'[�3=D�aD�Z)'�|���T�1C�;u���7�Q+i��M�ȓ �Lt���V��Jف;+��ȓ����G��v�i*�e��(Gv��ȓh��DY��׭\��� f#�%����ȓZ�T���|�$�f.h�q�ȓ~4��xǍ\� �{���\�ȓo2���&�n��d�(2�N�ȓY�b!��Ƀ]�p���c��m�!���\ș��A6l�Pe�F&�!��2Fs�P����2�n�� �ik!�Ę�6�\�����(��`/J;>^!�D�
�L@�n�'cl���n��S�!�ՋQ�R����Y�4=��	C�-�!�� ��N	:*��j��*�"O�e��j�!D��Q׏'�2��"Ot��ʄ�q�~0Y�-ܡ:LZe�v"O�q�$�E0Yn��FB�o/�e��"OҌ��+L4�PAq�Q#0���"OpiŵS��	á�w���"O�9K #��Co֕{AN=q �0"O4�iE�?��8��M�qf@x�"O,�zr��5��L�7
��'���"O2�*c�ýLȽ"��q*�]�$D�����K�I4DLx�+[��*�k?D�ܠf�,MU�9��N�$ ���t�;D���E��K�zm����R捓;D��6		0Iݱ��J�6[򡓰�8D�T��@P%KI��fǮg($��,D�0�A�3�����0A��5��(D��2i�:X;h�x���UC&D�l`2�	D�F��db�$X	�8D�T�c��7W�%RbV#�ҭҤ#7D����jĚU!ֹq�\��@4D�8��H;q8�pi�ԩ2[���Ub1D��3�^����OS��5�&�-D��"�a�#F����+ӢeY�M&D��9k��JEvI�BE3ڊ��T�&D�\yV!�'u��y��)���.}�B䉽ؔ�3b�'U�v�(rfQO}4B䉥
�l�$(J:rk�հ )�jCB�	�K.r���!�Ҵ(T��9�B䉴��s)�?4�p5����W��C�	��v�RV���ES���nC�	>a�%Q��\dE����^A�B�E���*�h�(1O�� f���6C��%a�
�Sp�ؙx�fMÇC�,��B�I�jm�I��/��).���į{f�B䉟@Dn��%]����!  �
;��B�I�j���B�E�n��;0��+�BB�ɰRj��ceZ5tT���F�%�PB�I�T�0l�E�p $n�.kB��2q���óH��#V,�B!۔ZC�>(��Y�D��� `)R�ŀ?�FB���zu�Q��B��u���_��C�ɍm�Thc񢚆&��y�*]�pC�I"j��L��Bp	�4+�OE��BC�I�y�L ���::�Jg��;oLB�I�DۦL���]#ִ:rE��&��B�	�,�I��$O�e��ʗ�b��B�,��y*�,k���c��T��B�@���k6�.3��1i��y�B䉗Y0 ����Jv�SA���C�3D����vɰ-���ٛQ]C�I����+�d?-XLe�4���b��B�I�v����Zi_�8y���)B䉍u%���-۱fH��pA�Z�X%C�	�"�����B/D��	 �9��B�ɌZS|�a��+$��X&�
�8�B�ɡI�ʕp2�<&�J9Z�ʣ�zB�I�l�N ��cȪ�$)�ăG� j B�&w���f��*1Ωk��� U��C䉚+�(�Q�(��^�{f���"�xB�ɁZ��e�1�24Au�v�C䉿J0�X�n�9s�����F��B䉶}�n,j�eϢ.XD���.@�B�ɏ�����'&�:� ��y�TB�	�R�:(B��S�V�(���	�LB�)� x���̏:3���1�h��"O�� �D�iw�� ��5t�����"O�}���E�Rv��YԎK	��l1"O��!���7|�<� U�����e"O���w��A�d3B@�h�t�z�"O��z�V�w�l����2Xh��W"O�iBA�Sux��G͔I��A8�"O�{nQ���JW�w���W"O�����	�����m��k��]�"O�c��v޸P
2�3z��T��"O2��S�͛{F�IYp���E�2
�"O���p���UOT�3���:���"O��ElS0T� \g����N�9�"O\�+�%����!&�A�0>��"O:]����u<Hj�dI/0����G"O�)KA,�
2Kvt9���� �X%Sd"O@��
�,4p�x��9i��|RT"O����V�+k�h
GO\9�����"O����@ćK�h+�\�!���z�"O:y@G�ʁqĔK�"�5^�(6"Od	��,ӎ-`�ǏQ5)ä�{4"O�����[$#��P�o	��T�1!"OvxB��	&b�-���I$iw�C5"Oj�"#�о� ؑ�R+����5"O��!/��r}3�lY��s"O�ẃ�R��j�+�[gPiQ�"Oh=�摠y�Ba���:5I�P:�"O�8���\�hg�hN�VRN`A"O��c+L2a<\ဠ��7P.t��
�':\U�@�>',qk�� `�^t��'��m(�[�K��B�%C�WM�d	�'tuq4@�:<	��#��M�zL�a8	�'}�d�
�4
�Y�
ӌ}/@h�'U>�!,L/#�l!SO�nԂ�k�'�Lt&J.R$� 􆘡w4�ݻ�'?T��疿A���C`
0q��P���x�/}���H"�50����-��Ǹ'�a{r� HE~�z�¥-�J�Fh���y⣄tn�3��^!n��)©�y�-��Yw�|�ȡhT��%���y���VX ��LT�J{<,��7�y�̺q%2���׉s�|�C�-�ybCLhQ��E&�<�Ì���y���
c~��j�	R�i*S�V��y���.��$�B T)(�����yE�g�&���H�8���`!i���y"��P��ӳIU.5����aj��y�%�#[<s�ʁVj"G	�y�G^� �ٳ�A1_�Lq	�B�!�y�kڙS���Z� �恛��y�I�w_>�0�n�he�T"�����yR.�`h��Q6lɦXd�biT���'b�	����q����Ŗ���j
�'2��X�I�8e�:�dEC�3�"
�']�ʕN%z���˂Z?
��M
�'��$	�-.Hu�F�J)_�d8�'7�Q��P�}�b�C�M�p�48y�'����NE�$@�����ݝj$�}z�'� %p7��$=�4n�([�i�
�'V�Ye�]���E��0N	�
�'p̑''B����K_�KC����'W�|)�A8J`:Q�
?8iX��	�'��eR�.K*3@�Y��<g| r�'h�<0���>'<�Hv�OH������� (���?%�P��kC'zn�i"O�Hb�ȅ<�:�C�jW?w_��8�"OP�(�cͰw_�)�j�,�l@�"Ob4Z�$"����#]$>��0�"O�-X��#>RSL�LUD�@�*O���r`
8OF���KI�nǶ�9�' �����h#�]y�eɆ<^��A�'�q;�^�I��9�b��&1tph�'(�j��7�h�c2^�� $x
�'&�(��mQ: 61�4d�
\d���'�"�1MA�*jR����ش���'W���%��Q���y�J��8!)	�'qJ�i�d-C��aa���*ȸ
�'F�] B��Bg�uyb����pb	�'(.�i��0sͤ=�P��4{�PA�	�'�DI�1�x�,rńȷn<=I�'=���Q���[��G�_�xa	�'~��r�$(RP|�	3�B<�ȓ*�(|�ҀN/?�6x�w�U��H�ȓz�lq�d�O�y��QQU�@&\N���¼����.]B m�pF�W!��ȓ,�(%����W�=�5���7�b��F�`P����%A�%��a�p�ć�tN4���rW�$�U�`cdm��Ky�u�c�#!��:���Eed���z�`�y��&^����W&���l�ȓ/�<ݱ� ���x�Xu���]G�	�'�ў"}ڣH)(|st�N�y�2��L�<�㘳!e]bd�r]��Bq�G�<a�B�&w�T�t��-��I��\[�<�O�Jj���91��	V�^U�<)ufF�9Ip�b�a9������h�<��oI�:��`�K3!'���T��f�<�&M�~�PBF����A��Pd�<	#dY�Wޔ��G����dA��D]�<YE'�?G&��"-�K���Qb�n�<Q�(]�6-2)��J�i�j�jG��e�<�4f�x���C��G���p�d�<A�Ǎ\K�Fd�4t
3F�D\�<m��6�qz$��~�� r�"D7�yr$@<uJ�1��;	K�y�"��yr��4φ0bq� |�
�Awm��y��ڐKJ5�bK[�s��h+Ƅ��y���p��pQg��h�փ�y��-{���]�^V��r�J�/�y�oڊK��k0A��`�v�����y�菾� �c�;e����Ȟ��yBU3��f�_����E�X4���?�S�O���KUBΌ8J��oߔP�>u3�'��NŊ\K�e@Oޔ�q�'���R�ٱ��U�t��,8Ƹ��'w�h��
��H׶��3��17c$�r
�';�d"E��e�b�A"�,Q�!I
�'�JT��o��{0��S�#����
�'3PiKf�Q�0y�Թ���=�<$�'��m�g�0�3���� ��)��'�t���j���Х�[�t��'#�ݹ�ȝ�R#�m���� hv�j�'�84��N�*xn�!�.�;c5N�'��1dfӧI��u���H'�	K�'ߴ��FA#v0p��=�\��'J�����4*������5'�y�ʓh*�Hٱ�R�};���m�X=z�ȓ7C��dΈ��5�îN�=�����S�? 4i���b�l1�0lK�`6��v"O�,�"FU*��H�D H��"O��+u�5��I2z)Ɲ�Z�<��
Z
DT0`�w�t0�\T�<���7�2pن��'_����ԉK\�<����?P����>U�����mAd�<�'�V'��\p�G�.�d�3`�v�<�7k�%.DH)�8h..\˄��w�<�E�Ҫ��,��1A� �TD�t�<�VN�+8\��5�1'�����H�x�<�gF	�p�a2A.�L�ap� w�<��N����Z��5rh.-@!H�g�<���	>X��fbA���qRĊ�e�<)@�4L�T�J�D��Q���f�<i��2,����^j|ݙ3�Z{�<�c�B:)	d1�E��Hy�XCnS�<�!eG�l@�Rg�

m�b�"�gNf�<i' ƺc��S cTȈҖ��a�<g�&&f�`P и~���P�a�\�<!�)՞�Vd�˸<��#��[�<QcٶS��	C�R�B���l�q�<��*C���hE���d�Z��]T�<閠�!3L��Vw�\Rt�N�<A���(~�[w�>/���9�L�<GG��}.ι�5�Ҕ����t�E�<Qq�v�}��N�tQ��1��CK�<�scTl�*e��g�
hx�a��D�<�F��>&�<*ԣՓ�Pa2��h�<�q+!7咹a��ŏV��)1��`�<iĮ4҆,�Ԫ�C��	#�A�<Q1cP2I�<�A�@6f�>�1�y�<���[���q�GH*%SV0��.Cq�<y��^/'�~D(c�F*1��h:FL^m�<Y��҅EpYrd�,y����l�<5���n�mc$�զK
�,�R�<�4
�<y��Ħ\�h)\��5	P�<)�Α�>@��ya��<��|��lUP�<A�b�6-����ňPdM�6�OL�<����L�U�6��8���Dp�<!v��$f{@s��ٜ���l�<! �ڟsךĹA�g���'�d�<�3�?Ne�����v���:b�e�<�ahD	Y4��s��
K�%Z��S�<�#�p���@Ę!S �ꑈ�J�'�4��%b���Sr)�6R�	�'g"�u��k�\[ǡ�t/�У
�'&֭r��I�Q��e	[�G5 ,�
�'
�H����)F?��@���#��Y1�'�X`;j}#fZ&�|y�	�'��<�T�g���'�)��H�
�'������PU�H�˓�I>���'Q�x������dHi�'?�\Q��'`5r剂k��U�#X�+�P8�'�֜�sH%��"�� �,�2T�
�'�h�ѪETZv�dfX��}c
�'���B�1QHH0dG�"��	�'�j3�[�a��3�]=���R�'R���p�Р�b-F3Xb���'?$X��!R�����oܝ��'�`8����1m��IIQ�H�1�DQ��&��M;�KūqIb�q)�)̘E���<�A5�8m�U�t���[5�,�YժX��ՂhoM�"O��D�3hPtB	�XH�pq"O�8�l`(軀�2'¦yj�"O� H��C���8!�FP��]S�"ON���g�K)LLʐ^�'�(�!�"O$�2f�1OP!P%Ҫ6�♐�"O���g�^�v�r 0A�X�>��E�P"O�q�H�gd8��`i��h5�q�"O�)ф`��خJE(� X�L�CU"O�c�ʰ�&��"�N���Pg"O�9ؠa�5�nH��l_�L�t\K�"O�d� ��_*���0Ny���"O�,���:م:V����́a�!�d	�P��eص�&Gz� h (P0%�!�$B�<��T�&.\	~|��Ȑ�H�8�!��[�sS���p� r�$��!��\97~9��dޱ6@Iׄ-"�!�$�.t�C�7[Vz}�7a6Bz!��6}����S�p�F�s��y�!�D��A%�ն�����$���F��a����щB�Ғd5�ոU��y2Aр.�Hi�2Q���qƮ\��y��)�e:�ݩR�,&z ����34J���ȓo�b��a�Ĩt�6�h`ǆh�X�'��}B*Z�)�`ԩ�L�7
L�8��*���0?iP�<�4(�<�F�8�J�Y,j���7D�Tx3
��/~���F�5\P
�Q3�
n�?Y�.�NC$:S�ҕn��Y��0lO(�T@���<ʉ1�P��P�K@�n����)�I_��/�?!N��U�]���ȓW�e��ӸP�,�J@�*N�O�]����QS�8J0TE�Ǖ5�B���p?��'T.6��V�՞p�D���d�J�<ib!���ȳ�F2]�"��b*CG�'v�~�C ��T*�8krdO�.�(r!bJF�<9f�����IĘ1.���e�{?9��)�'BUBY�� ѐ%�F񇩊�c�bЅ�g��kC�S5�0Y�]�@k�إO&��I�L��u�G��c��H���\,��DC?y&��qk,d���	_�^]�GOg�<Q5�J�����l�.M�d�0��\�'���~2a�Z�V����!F�\������^�<���F1%�X4�bE �YKƅ�op?��)�'r!�i�rHP>�(`�	'Ȩ��ȓe�8����Z�d�\؂
Y�l���Oȱ��+��9�j&&0]��Fÿ+�����J?��N\沭Q��:)fx�37H�e�<�W�N6��uѦ�J__�1id_U�'w�~�aL�w��H�rFɍ�N�ؒe�R�< ��Pxx�:���@(l(5MEV?���)�'>d�B��	nN��b�^<e����{�&�bCB�>�����0?����Ol��d�	W�SpF�,e=,4Jc��ur�~RR��(�iզo�Ȫ���m�$�h"�.D�dz'�(qk����BO�T��Iq>��9DaT����,@�!���q-d�����"=y� �"������8��O
<�a��=���邂F2�H�[��@���'��#}�'+&x��Eݵ�)b�M�0�,l"�B�~Y�AS1AQ#��� ������d͢[̜�-5Y6�)�f�	{3�Fk�rB�~�&ԸM�*����Ǟ]VX���`k@��d��]n���X[���gy"g֔�ēmӲ1:��E�䌲���C�I��ɜP�p�Q� �ܬqC�k^�M��@���Ⱥ�iU#0T�����3Q�I&U�Q������	.6ֱ���M��(��$Q&|_��D�?Bh��.=F[e�ϟ|x�$+>VJ~\!�Gr�� ����T8��p�̈�csl\�O�,�j�Je�]u͆�F'4<��|��/)T���$?a����U���*<��aE��\]��a'��H��B㉓a���� �
B����C�rw,*fkL�*+8�PD�z2�G��`������)� �aI�`����t�ƏHRD,;��'� ��4IF�KUJ{e��pL���D�6U�bq{#�V�=1ȡٓ%D�J�|s�hVwX�t�� M�K1:�ea;�P���4��B"w�8׫
����	�"4R�aъ!T|���%�p{�,��3R8��@G3
C��Jy0`���$��q���2q��t�B�,�d�A@O3��9w�Kx�O��!3'hoޙpI>Y<h��R;�i�	*$��Q��W-�K�A�VU�IO�}�F��«�b�YA�����\�Gkż.��p1�8ʓ;OX�'�M�y��M�M�; D��Ik�	��	�$r
8<�g��n�0љ��*��M�v�T�b��y�vNR�-��*YD8� �a�T
_B�)��ϛ0՚�"!g9�ӟ5d�-K�bO�7Ԥ"1ˉ0&O&�Asf2U'��S?���s��f{Ā[�TW�B䉖|��Щй��|�bA_(s�`t�Q��<������/�"�H�~�O����u+ �ooU�ʀ�YQ@dO�ځ�R���N�Z>>���,ѯp(;���P��0T���i`�B5ʓI?�0��/��5{V(q�Ƭe���ɨxo��hP��\�*Ы�)�`��]�S�l��3�B��Q�$a�!H�87>���l�}8��K���N��c�c�1	p!H
9��g�z*��r��)�x�fl�A�A/�D%�S�p[��Q�-�..�ʜ���)h9�L �{r�O���'��b�˜�@�:!��AH��r��,c���j�-1= \ل�ݰ*��j������ˤ�E��_�L�XT�O�M�8�f�G�&���q6O���DѕY`�A�&V[9b�)�mҚS �Li�VVmpE�5CGw�0�i� ]j�y��ğ�y�'	�I2���	6,2��������D��Y`�Q�-��
ѻ��ʀu�S�'{*�� "=&��1��9��i���џ0ڛ'��	e?�+O� ]�D�5"!S�L�hG�x+ĨC������ݖ *���ညf�J�
$
����	ʍ*�<-q_w<��E�ƹ?�E�g3O���~r���pD��-Y&`��D9}�9'$A�DE ���b��NJj}��G�O�4��7�t@�*\��������22
y��OR�֚_9��+��X0�����N �l����_>a܄�9ckY{�ᡍ��HOr��1�H2!갉�eW0o�^��1�'t������J1�=_5~T��`�o�N�0c�;Įy1���[���֪���>)q"U�?��]"Q��z	j6Ƀ^�_� 9������ORp�L$��k0:��%�	�c�݇lmi"Q��T�<�2)ƽ%��}�T"Y�}�bX�3�ʄ(�d�{�*�6I ��wLF%:�DD�t�O��&oGf�uT�1�vLi�"O��)��	�e�tb���9i�@�X�J	�Bz��K�L&ؔ��vn��D������i��<�0�p��*$�a|��6nrV-���4Z<8�0z�N	qG&¸ea.<@w�C 3�B��<�"��l�ȱ�eV�HO`�*�B
�V�d���9�S�Y��YQ*��"DҠ��e��C��-T}�$�!j�~��q'�+n$C䉞"S�D"�f�8(r6��r%%k�JC�	< �ju�d�V%GP��Uk��^C�ɒq�����w�A��(� C�5P��Y��"��	<�K�*ʳa$�B�	�P>4e��ٯ�0Q�c(U'W�B�	�w�2l��\%iӬ@�wF��x�Ɠ
U����n��R��	��\�F�h-�ȓAǺ��T͒��Na��O��Eb�5�ȓ~|�Ͱvd5ԞUq����y�v(��1�j)H���]&�01�H�Z`�ȓKp|���!T�4�`�CCe��{����'��~r�ز�Њ"�j���O���?a!3O��	�\�s7KS
|0���"O����V=@2�Jk������������9�Ԇӝ%D�|H'��x�R�@G"O�0B@�X���y�G�±2$H�"O��^�>�d؋SD�=8k�"O4i��&�{�0*C�O>xز�+�"Oƅ���H�v�C�d-y+F�1"O���'�(�|�yC��I* Q"O|�rlݥ"�VX���A� ��"O�}1��&1���H��#;��k�"O�y�4�]����FB�fAv b"O-Hg�Y�d��s2o�-/��y�"O� ؈0�M�*��Xj�h	�*�v�ȗ"O�|�tgjp���F�m��;q"O�y�$��I��]����0Q~�"O���ѤZ2P�9T#K�hJ��"ONx@6LG1|<�+��I�C���J�"On|�C㟹�����E�o���s"OA����hD8r� 	b�p�J�"Of(cr��&-jժ�X79p"O��Ѕ� �.��<
��R�$t,؈�"O�P���E/��1����3Bq2T"O�i���\��MI"@��1J�a�"O������,TNJ�aS _9R�M�E"O�d8@�J
I� /Рo��iR"O�I��!t�  ڇ�Jv,��S"O��(�fɀL�jšUØ�lt-�v"O&8j0�.K�m9'߷���1"Ox���'�=�č0�Ƙ6���E"Oi�6�N�eڔ��M��� "O��cQ��BѮ��*ĺ	��"Ot�q�<<�sG/�2�,#�"O6)�Q+��l���җȎ��4!"O��x�+@`L����ǘ�6�*s"O&QWb�l�QFEL�.ص��'�	�q�C�}�¢&J�(%z�)�'����CF@��y�w�Ǘ+�5c�'�V`�w�݉@����g�K~�Y��'�Ԥ�'���������<h�Q��'
hIH4�Jc|h���!9jh#�'BI��
T<P��aU�&6�p
�'-�L�")E$]h,���cC��h

�'� 0%$���z=�T'��~|�;
�'���q�&�:S侸��E�����'����'G>��9���ŨtB�t0�'�΄SW��'^�p��pll.�`�'�~�i��]c�I����
�'�V�<�A G$=����h!@� ��O�<�Hɛ`�f;�4�fY�¦�o�<��$|�:���oI	L;Ԥp�o�<�Q#�$o�汢q�
#%DXP�Th�<ٓEˏC�\�Q��ȼDPQ�g�	]�<����#uG
��jZ9o�q����L�<�*��a�ܣ��<�ܰ9�H�<���eJ�#JG�i�]9C(JD�<�ea�,O�%H�Ǝ)j��H�@�C�<�U�dG<-pw���z�DY��B�<�b�H��z�b�υ�-�W�	p�<QWG^�%��i�c�	�L]˃��m�<�rLV�E��M�@G�Q�ƴqGs�<��L������h�az�n�o�<I��\9�Nٺ$ ��4�B�b���o�<I���V�<#r.O�,��mji�<9Qn_3uqx�$���	�X�!W`�<ABM_,}�B���N��Z��]���RT�<ٴ�@0A����.�X�т�GW�<y EK�Fm�M �ŝ)�x �T�<����Jߊh� u|�Q!�OCH�<�S�-4����"T`�\�h�M�<� h n.tH o̜v�d�AO�<!'�1<1��#��͔
�>�(T��|�<i�.C%���٤mP��92��y�<I����l�
]c�%ɗe��#�d�q�<Q# �S�
�;
�i��� w�<QGϚ�i��A!aCxzv�b�Nn�<�w�P�9#�K�?-&� � h�h�<� ���$$�9Ql�CN�!�R���"O��ɓ�
+?0t��퍁;T�$٦"O�p����;`���B��F!)9�1)�"O"�@��  l� 	#��V
�\�C"Ot٘0��Um̼���	�y� �"O.Q��c�_�j�#���P�`�5"O�a`#���/Nh1�`�N%#�DQ�"O|{5 �0!�H�e�( � 1��"O�4�wI�1[~`���T��dہ"OxDhV�5�F����־D-S�"O�Q�L�=��r% -�Ԫ�"Ob�Y�bG,DjP�p0��(7l!;�"O*�xe��*�8ā�K�I#lyy�"O��'�¿;�jض�-\��u"Or��Fc�"$�f8ÖD�4H�"O>ap }۔$r�T�k�~y6"OXuj�D]2޵�e^�}�,1�&"O*Tb"h�"T�j��` ��Î�%"O6����>|�]�B�E��>�y���3�dh�)W-S�B3����y�mݙM[��tn^�Nv�X(�gɲ�y���6��ppJX;�>y����y�\�.e`�{�)*��8)��C=�yb/݀�&�`�B�'v��O;�y�ɗ�s]pIAm�%�6�1
���yB�H;m���5 � �dM��P��y"���-T��w�����K��y"�^�A�8q'k޺9ٲi��ϸ�y��;J���xUgн6��x� ۧ�y�N��X�!' R�!<�u2bc���y"N�D�h���Y�-
�>�y�Ř,��s�>r$X�����y�nG��`�����* E�X��ҋ�yb.P�@jXRP	U�I�� b�	�y� O*6��%sp@C�F),}ڤ%X��y�ꁫ/�FD��J�28�C�Y�y�ԎW�m���_�?l��i@��B�i��ˏ+(�e�a�f���U�+T�Ƞt��'Rv�� �Z����"OP9�MW�"G)*%C�/3�0��"O�L(�m��Y"A�ĉRr(�#�"O�,ADD�a�($�D��cݲ	�t"O@��u��7!�L*&���Ό��"O*�y���	Av���K&]L�ի�"O0�*�Jբ����P��'&N��S�"Of}�wHVY$�`� �
�p���"O�����v9�$A�/+p�*�cR"O��s�(�(������MR]�d"O0|�� �f�HjQ��;��Ē�"O��y����l�С�8$��u�5"O|LS5�Ƶ	�H�J# P�x>8�Q"O������-J�`�OU�~m2�
R"O45��E�=a%�<9BNͩ��9"O�e��ңhK�0Gm�c2xv"O������#.�UX�./~��@�G"O����j��8�6l�>zx�Z�"O�,���:����ʳn}�qBS"O��K7Da���3�g�7����c"OKU�AeLT�bm#5��:4�H�
�'	�Ѷ���#|��j�b��7p�=H
�'e���"����Q��g$(�s
�'�V,A#�ȠPɔ91K��=B��	�'\��p��*��k�ɛ�$f�i�'和�2j�n|��p����>���� ��`������"��D��]�"Oʬ��ށa٨Itfđ��-�D"O�L���
19�I�~^����2D��H6�-�"=á,�-|�[1�2D��`��I&צ�c�Ȃy6u��d0D���&�EY���#wl\;M0r*,D�x�2 �-��)��/E�����6D����#U8���mɛ<4�4D� )A���h�����Y�mSs�3D��q "��{�f Q��@*+=��@��1D��{T�C~�:�_q��j�k/D��#�m��+�*5���Đ�r�,D��`dKG7H���e�?-��xj�"9D��2t	�5e`l��d� *��{��5D���Fg�.�UH]���X!�6D�4!p,�s|F"��]��92U;D��a��˽N3��y�d � S�M�1K8D��#r"�U�¥p��7c�n-H��9D�4z3�Z<�[wkӖ{�`,Rb6D��+�B�HenE4��"�d��t�4D�@㖦�mD�t�M�2Aj �)!D�����N ��#�L�Lp�d@�<D�XA��	1�2q�W���d9O4D�`j��r����KF�5ā -1D��H5�Ļp� 1{�ʃ}i�ś�(D�����_��U�W�H-8�=Y�
8D�Tj�h_�{��,p#Û�1�4��S)4D��������h��w��
U�2D�xH4���WOzi��W�~oР���=D�<2���	�JX��JԄQ�,�8D��3�ꃱt6$�SӪAԄ`h��=D��`D8�n����,��s�=D�(R���K���EOM'�$��:D��(d�W�v��D��]����I8D�Յ ]f�X Lݽ
t�H��:D���k��B�<���	?�>Y���9D�܋��A�&����/��	a���h4D���0/�F��\���O*?����c4D�K�E�hЅv�LR��I8�g,D��r�S
�l	��̈�f6z<��n7D��d��� ͢�J'�K���|��7D��9Fh�AT�PW'�I!��>D��8�`K�{m6e�q�OS���To D�,��ņ�<��*M�0{:$ۢ�*D���D[)ih���͖d��S��%D���စ�f�q�q(I�#r��閍%D�����C�湓C!'%R&I��!5D����n_�{(�ȋ7�+�K k0D��&ƺ>MBU�R�d���G0D��rV&O)n}P=��'֟6��98p�/D���rس�0���L�'D����(D�H�Sk��<�d�㑅T�D��͛��)D���D�>wpfA�'BS,M��x�&D���A�SY!ҁ��[�@5ҷk8D�X��i�,�3�a_�Fu0$�,D�Rb"�0E�H+r,�M����-D���f�>/4����	!��r"+D�@1&��\fy����Nj���(D�Dk�]���q�A�� o\��S��#D�$�UBTr���B���LE3 �4D�¦%�B����`��]�"ՠũ'D����G�(H���j�7�B�`f7D���!�5(�X4Ǖ2\iD���4D��JCO�:#Dl�ř�EIl�	g3D�� ����B:i��l�jY3r7���S"O$K�hH[�e�Q�����"O�P E���s������\��2"O�U i�#p!�����Rx
�Hc�"O.���M��dIc ŹV��x�r"O�B�Dw�lX3iO�&�D�V"O�)��j��~q��馎K
x�pz "Oj9r�ǳ/<�l�q�[�Fż���"O�wF[?Sj�MC�kŮb��%�%"O~��6c�yДQ�*Z	�b0x"O�s#`� {��@�� �>�HX�"ODm�V"�o[��۠�Z�T�J���"O��i�O�x�T��NW�L6j``"O\�z���X��Y��MǕr��l�q"O����TE��@&Ձ璽��"O�@��	S��H�plV$�L@"O��+)�����$�ݿ��ؘ�"O̸���uh�]�B�:<�xLu"O����?e��E��ƁD���"O�EP�E�*��\s��ӜO|&0��"OH����v�K��(N`(�KR"O0��&N�Xnd��@�
a���r"OX(뵫�&b�%�t/U�x�:�Z�"O�L
!�2�p�*�N�|x�9��"O��{�	�`
-)`LU��P"�"O x�EL�0R��{0 N</� Ȓ"O&�h��"Gp�) Iύ�f�P"OH���)F.4!�3��~P.��`"O� W̕T��x�G��FO���S"O�p���e~��lM*�0#�"Oܭ�'�F74�f�p�җN6�"O�ۓ!BR�B�I�
�+�)�yr@̎��C�H��cO��k���y�F��B���;Q�G�^,�Q�'A���yB��`{�a��T6���'��y����(��t/I����&��y2d�
q�S��I����V���y����H��ؠ��Jf��1�fT��y2a�)7J<!+i�D���"��@��y⚳�a藁8?uj�¡���y �	Lh�t虒+���[a�Ұ�y&ؔQ�f|��%��"8�[Q�׽�yb(S�e<>}�b��f!30L���yB��Ӱ9k� J3Nlh,ǥ̆�ybBȽj�<LH�D>|����`���y2�ӌig͸ģ_�7�0:���"�y���:Z�Ó�
"^� )��K	��yB��;S�=��Ӿ�.8;���y���tÊZaJ�-t��J�[.�y�L��'��
��jGHh�y�)�)z(\�Q�T)u�X���L��yRg��T�*.@&lgҨ�W�Y���O� �d��z���-RI$���IP�F�|�ᓁ �Lu
Fǃ�I�TY�#�ί]�l��fǗn�S��3�.�!Š�7#5,5�P��/Zch�'Gh\bv��	�*:����n#Y��Y 2�D�(uB㟢}�bO��)v�ܺB>�:RB4/��M�!��S��}�to��@�|�� �6e�*qS��e>�C�$=TD��NS�;���Tb0�`t�@�?%?� ��gb�J��Q�v��`У }��#H��O�!��#l�}�����C*\UqC�O�h��;�)ڧUE�D�m�Ζ�E猛z	�y[E$
Z��O�?}Ȃ"U��$<�����6��lSF(�,)�O�B�'T�hD���ת.��+�P}��N�>�y��	D<?�dAf@8�	�?�fEv�󩅹?��h8�ƻ!���2��Q���w8@��U���g�1��I�W�� �T���b�P%#!� �k�E`1��K��"v,��I�0|Jwj0�F�R�߷Qg��#f�t�${aL� �~�`ĝ1*����7�~(�FG�`Â ����.��es��'?	 Iϛ:\8���Df�Z���� �4�v9H�&s�JOt�z�NK�L���)���exA�NO����nκ[d���B�tr�̈́�wr�S�O��A:3�1x@l�Q2ܱ!��e��32���F���S�O�e;���^)�ᡁi�����A6S���3��?�5f�:d��b��5`��E
0D�l��.�S��%"@유}�:��� ,D�l���UH�0�!�	�UԠ$D�p��"V%�h�lت��� �"D�x���@2e�B�p엪,V6t��G?D��2t��^�Z���� CP���7D� ��FӺo�>�I�:'(�H!7D��qL
�N9��%hڢ �L����*D��;#g�LZ��k��[$T�HL�c�+D�$�wnQ���C���4�R�5D��yV�� ����U�W!i�����2D�ر6$[�5���`b�[D�p��D/D�0�3�\�}�V�!$�R)lk��X�-D�X!R��<j��ܡ�d�C4�%D� ҤE(��K�3R%Hpa"D�@볨Ăy��1cd�'M�mȷd#D�أa	��0drUr1MT�&&��A�;D�l�G�R7]  Ks�5Tŀi�K:D�@�lI�{���6�J��
IJ�c6D�P�cS�W9��5�Ƈv4�Jq5D���cMܚn26�k��#4������'D��B�ŚA}�� �.��_�l�c�0D���a��j|a�$e��V����3D�<I�eN���f���d��B�E0D�0:���5 � ���.ҙb���q�/D��C�i۬"�l�#��P1l�`�L+D���-�VBN��E�#U�0�zn'D�8�s�:f�ԸY�.��c��K�l)D�Xؐ��?����J�E�Xͺ�E&D����(1�0�񎖬SJ�����%D�Pb���v�Z��0�U'>J�T�5D�PP`��"4"s*�d(HB�2D��5 ˙��v�W�29.pK"D��p��6*���+�/�7#�ʤ�1M=D�4��^؉ �]"zӄ����:D��a$ԒY�A�0&��7�eR�9D��@eJÖ ���� �<਽�PH;D�`$��z�t8@h�:pV�l�a;D��3�䄢7�R�$i��N}zD!�@9D�(XQ�λ,Z�z�Q, yjx�U�8D�����#�l��'`k
�c�#6D�0!�h�I�L4�E	-&Dެ3ъ2D��;C	�$t�.��M=`�*�e0D��;І�?2n0jD�ݑ�P7m��B�I�S/$e*Z0M�jQ)����M�C�ɤwN%3�GC�V'HQ���]�*� C�	�k�v����%�d�(�iIg��B��h`Bî~�����hR�B�w�l��㏼O4�͠���0MCvB�ɖne�9J�̢w������B_FB�Iie���M��Y� ����B䉂g
$C���P��y�e��B�I�I �iצ�:��1�c�5n�B�I�)����B�o��]�v��?�vB�	(�v�ڇc�W��0	�� B�ɨi\��ڤO�@n��&-��$�C�	�L��2oY�&�d���?+��C�)� \`��+����a%`D$<g�-�R"O�!���ЇJM��RN9\���v"O�u��#�� ����
+!�F���"O@�:��C�I�d�Pt���0��t8B"Olx���h˖��3��0ii�"O�f��:�`���P�h"OZ�����$�j)���@l�~L�3"O��x��OH$�q!-6 ��*u"O�lS�d˗7����L�n��R"O�`q��ɆDʱ�D�G�v%k�"OR�%�\��މ���V[��̛D"O��ô�W�H%A�-�{w�u g"O�i��@�+��� �&L9eI8��t"O��p��9|���� aD0��"O��Q$�z��0R��\���H� "O��s�!٫(+.��fH��&��#�"O�5��T*J
�\�%�	:��	�"O���C�u�Z�6dF=Yt䁡�"ODґ�N."�)P�E3^�`��"O��� F��v�V�`C�->]�0Yd"O�`Ӏ�N�4x��I�2T	
P"O�xQ0�!9E���<4F�=(�"O�!�@I;L��=�T�Z�e:�!��"O����*��d��`��e�;,�ኰ"O�%3L!�:\[�Dƈ4o�уC"O8}I1��=������=mX�Ec�"Ov1Q�)G!F�R0��xn�0"O�=hTb�*L���F ��R�"O�e ���w��fG%8��t��"OR��L޺!�`"#&�4���"O��Q�ᘢ f4]I��A8T]0���"OܘZ�W��T����,Z؀
�"ON� ��Ч4�z�h䬁+�΄p�"O`5�b@�U�p�cì�\����S"O`E$IQ:_Ѩa�+U�ny�M�R"O�p��a�1+I`ة�J�5h���0"O&쩶GB�)�y�wϛ~|.m�!"O��H1�P�[qAPIR��X'"O�9v+�9 &>��C��8�v�"O^����D�m�d��W�l��p"O�����E�(1'kޯ5�"O���B�5��1�"�ۢK��`A�"O�Q���. X4�`#U�5�0�"O��;pk,mf�!j��	z@���"O>�PG�\�ph�ǋQ�t6��["ON`;3o�LX�I�?(|h���"O
���R�IQ|,��U�xe����:|O�h��KU�a��� ���F����"O<����euzPD��67��Փ�"O:T�$���aI��q�)L/?��YPg"O�Q94��nژ���ty�V"O�XK%�F\� ����_�^��"O�u����j`pHp��[�J�<8ST"O4�J�-ǺS��X�#F�_�8��s"O�q�f�H�ֱcT<�tr"O�vKK:lAص@D�RW�Ld�"O��`�����R&ڱy:f`��"O T@�놰6[�1(�@ �I�"O�8�v@_��|I%+	���W"O,ܢ#nZ�f�A"k�#~,�@��"O��'`\>`l�	̨G"t-ZA"O��؆.U�i��AեҘx�x 8�"O�=�#	��>���r�wr�ma"Oq��FK�Q��9�gaZ���"O� ��A�E=A���'ߔ~G���u"O����b�d]�z�f�64��w"Ǒ� 	%
Iܬ�s�ˆ"����'w.�Hu�ș_p(� $k�m
�H��'&	��(8צYb��H�0ʘ	��'ﴙ2�H��)�� Ç	�VAȅ`�'@<��ɀ�k(�姁UV�D�'��ٓ�nBsZh�;TC��H��l
�'� �+A���ib�DoN8��z
�'�Ppd��[�b�bB48�,k
�'R&ͪA��6��m�Gn�=��']*Vk�";Ra���VtX�'�|At�U`���i�T��'C8|3v�W}ٰi�cH+
9VP��'�8<���"D%|�ܰ~��"O$�(q!C�0�$�Ax�d�C�"O���1�B�3�ܨɧ �:I�h�
�"O����g��*b8��7���%"O�x:��%V�Ÿ���X��"O���$�3�("�I�,"��X�e"O�1(2*��lX�kSH!m����"O�S	Щpl"��7F�:w�r�ZE"O�`"�!5e�F���ه2T����"O�9�Ш�`�d��(Zija��"O�]I�%Y7Y����Ej�f��ĺ�"ON�Bh�i�<ʱ'T����@"O|��FO�H[�M$L<���"O"��o݈=s詈��H:�`ysd"O^��W��&0�����#�?u�v�
 "O���6H.�*����f�D0ѧ"O*�S���;aD�&�դ��"O���� C�A��80���U���8"O�-��N�l�|iZ���Ns��Av"O�5��A�,Y�h��o��|��`y�"O�l��R��\{����B ����"O�ARP(��m���X�ü(
�t"Oh�ʃ�iA�E!k��5�N��"O��'�	��6��ۓX�M �"O�(W�ߖD�$*[��3U��;�'R0�3���@! �$kY����'�`�����3tr�y��B���|��'��Z)A�c��I9�b^" t�*�'��+� !�H�F��uxu�
�'����o��5m�9)�����	�'����	�7?^��!���:°�	�'�4,��˝�:^�QDs�΅x�'�J�����jYV��3�C�{��4��'���Q�X�kx�c���Aq�
�':����J�A��*�97/�-�
�'~� �k��:N�����5K���'�d� !!U-VQS6&�-�H��'�,���w�x�� Tc�:�'V�� ,�jY�9C��@'���'�R���;z>[�c�%�*�A�'�(A��,X%kթ��MC2�
�'Rp��/ȣ_v�$�1Hƶ>A�L�
�'���!��,_LԘ��X19�:��
�'i�� �
P�F# ��3{w,t��'�f�Xq�ß#�.�� *¸QB�'�T��ˉl�4u3
�"vDl��'F*�{�O�'0�*��NJ���'3p4���տH��$����;�*�a�'��Zf&P�c���17m�E�=��'�&hҠ�1Y
�����G�0��5z��� � 	�䇖gŋ6�ց�"OT\�B��[^hE�T�߼X���i"O؝)�@��Ԕ�s��|��hD"O�u���E�I��2m`��1�"O^ܻ���?�^09��ժE�|��"O��#A�ߛ7 ��C���K�2�A"O �jQ(�1i��:�
T>Јp�g"O
�I����e\��Uj�R�d�6"O��#��V�=�n�3��ӻ@3�ٹ�"O��i�\�'׆�1��rϐ�"O�(B�Q�d��m)pA@�"O���t��,�Z-��fA�~�9g"O�}�L�c�����g�3�M�4"OTPY��*3��h�Q�������"O�]	�*Pkr8A�g��R�JXY0"O-	�k�����fհ7�$��"OP���   ���^	)��I�%"}�}#�
��yBF�&!�z�����zW,�(�<y��Σf:��bJ�-1����1GQ�:��{��D� $�đ�aԂ.��`�#�I��!��2N֜�ps��j�����d�!򄛄����V��l!r�s"
I�t~!�d߮��� �.��𪂨�:5!�ć�k��؅�B%���Y����N�!��o�H �āG�J����0M!򤅿V{���ꏬ_�
��#{4Q����>���j�4�x�"�
�%r}BE0q��y�&�a�\X�BQj�L�"�
����0�	J��~r�V�C����B�l�*9Q#�,�y�/��Z8��nO�l�!Q�戱�yr%�(=�j<�#k�.\�� P��y⏋%`���J!�ӯ^h�V%C��y��	�p�XAc6{�suh��yB�Z��T���ʔx�i"VfT��y�'����͊E�Dj�p�喱�y�l�%�*�r�ۗC��<3ãL��'jў�4���t3*H�����j�$����I_8��4^�Kz��V�M�R6\35F&��l33u^���^2PvI�a�C)q�B�	�W��A�uʐ�R%���1n����C�	"��XԄƹ6���K1`�C��2	i҂?j<��e�G0|WC�+m����Q%S/V���j�.�V��B�I4�P+$�Xc���'��=�C�	�#�E����w �8c	ƮY9~D����(�+���0�̍q����F�u�fl��a�L�h�h��Т=�d BTE�HsD��V�T�R']ШpB�[-���ȓBy�%p&�/�L��
�+'wN��'{�dAm���'����CG�-������X�>ə)<kӑ>��S�? P1�*�P�8�k5!�2E����"Ob1`e����s/�9K���� "O*��m� �=��MD� <;�"O4���A�1*��U8�/�v��1��>�	�a��5�n��=8���&�,Yg�lF~��{4^D{�4kEХ��g�08 C�ɽ.{V-����P���Ղ�Z�~��'��S�OQ�г���L�V�C,�f�@���'��u�ω�e�|��H#��1�'�H0���s�4���S/@������Mc�OR�90 �j1�u�قgmʬBD�'���P�i��r*>��F}����� D�py�JF'sX����oՐ��r$>}�S�t�<�}�͟(�Jٓ$���"fF�#Q*0��'�ў��E�D�/�F��2�'o
����>����m맀ȥ�F�3%��)L �'��:<O�l���NM����$hm�X���Pq�<���X~h����"9v�8��j�'ў�'p4��PF�A�x�H �F�&B4��Lh��ac�)�BX�-%@[���'f1OƢ}��>�X�p�8Q1Jy�$똞R�j��ȓ3�]˕ꝯ����_�-Iz��<�	�wp�̳�!e��!$
����	�@��6M�<��X�b�9 ��ř��4 ��Zi�<9'K>KbY� �C���1�FXh�<ɤb !1ZB�UM���
$8dNg8�lGz��o��8�� Y��R��O��y��)�'l䵙5n�V���]]��܆�^�m��X�54�"��N����'@���b݇�]��_ 	��p���ty��P";E�<��/�"�z�*���y���XQ�P���+m$�P��\��yR�^1& ��NO<RR@�2�A5�O�"�D�G=��iq�A&��9�1��� E{����9[ ��)tE*��U9s�����:���5W�6�(�3� .A`��Y��<B2-ۚU��B%r+"0*�c�Or������t�:P�A��Q�Q$5ag�K�7D��;gn»?�h��2)� � �)j�0��	�1�
ɺϞ>
�|� ��p��B�I���u�c�s�#��K�lV�C�I�D"Pu�"LZ�`��Y�Vj,�l��<}"�%&�ȸ�T���u���QLW�yR�ͻk"Vt�g�l� ������٦���-q�<�S�E�� ����MV�!���	g�� �b�g$�H ��F&0u���;D�P���SHp��6,ȅ*F�T� .��ȟ�DP�A��~s ���d՛5\�90�"O
�
B)K�6��i��vg��s����=����JXPIRYr� ���0��'Wt�`��CFå(��&�3�'�L�v�P/s� t�̌c��Y�'r�-�#��cLyzO��bL�|��'}���fR�z�2����U0��x�'�j����
�N�H$F��E:$��'Ң���b�T�5 �Ap�(
�'�L([�O4b��T�Мs'J��	�'<t��@�^�[7��EM:V��	�'��;��G�S��tbU㚟FGe[	�'�� G�J�*�~%2H�L��UH�'2RA���:b�as���F}>|�'��P�7ς5 f�3��2Q�,h�
�'�z�(�Bʆ7��`�2�PG( A�'���OD�����p^�9/&�h��� ���F�M�@�6<�ba�
Gkt�h�"O:ȃƮ��J�B��0�ԅh�a�"O(� F8 �м ���O`�B�"OV�!��B� ��GiD���"O��D�@;��W�E1$$��"O�8��C�@3� �%g�*!~��A"O�xcjZ�S ,��RÎ0=�&���"OJ�qM��T��	D�ר~���I$"O��J�i�;��R��{���0�"O�[�"۶t�)�#F�q5���d"O��K���1b���*�ŗ52d��"O�������w�Q�#���2> �'"O8(�7j��
s6�7]ȸ)(5"O����ȅf�Y�A�t��M:'"O�h��Y�+��ݚ�%$�n��"O J����k�`a���Y"OnԊ���`�ԩ��؊\�B��R"O��бi�zw�ݰ���6���p"O�eqUH�+�hJ���@��'"OLp�"�_8;�dA���4�2S"O,�c��m:F�xfb��a��;"Oi��$�d�bP���W��%I&"O�=���ئ�"���ª5dĐ"OV$��̽x�t
�(��{]��[ "Op��킲1ud����">�Ca"O͂pHC 0��! K�#�ɒb"O��௎�-��p�Ϟ('�T*�"O� �0$�6tid,&,�,�8"Oȑ��V'3V.�AU,@:�.��7"O�DA���6�y���n���y3"O�PS��*J[l�/&�H"O����$f�Jj����e+�"O�y��l�q��)���Cd�§"O� +�JA�R"�'0޽���7D��lXFɦ�:����-�4�4D��B'D�VG`�*�ɞ8�ֽ��$D��� ϖ�����`O +^E�t�>D� �Gɦ��Y��<$��K�<D���f�XQ�4͉�G�Ȁ� �:D��b3�7��W턷:]�!�A9D� sS��2gW��j�Á�$�ZqD�8D��C�g������6d"dr��O5D�c��:���8��V�.�l�,8D�X�fl�Zi���LԽR����5D�P����T��#�%?�%�!O(D��3�	9%Tz�5-U�F,5��C3D�lx⪐�OLl�i�FQ 2�<�CB,D����&O{��[�5�R����)D�hB���@=x�#���T�.�1�&&D��aoBn��6M�?B��[� D���Ɉ�)I�@�q�̬�����2D��`@J(/"�bu�/��A��<D��z���w�%z瓳o}�ɛW;D��(���9A2��b�̃R�B�H��8D��ٲ��0��[��Ȧ= >-"��+D��q'oD"ǎ�i@
�h����?D��q HF�|��-H�');C��S& ;D��a���T��u��g��%N,<O(�}��D�m�j<��/ J�A�+����O#~� �4+�� ��%�k�(!��%�Z�����#�~Xæ��A�� ��K�3f����<��Q1�$H���`CM�o���'���#?Y����:m̰1A�G�%�L샃�����"�OF鱄\�%9��0Q�|iIPZ�DE{��� ��K����x�^�W�2���"O�ؓaZE��S���K��iV�$,lOH��5�9d2�h7F0ll]"�|b�)�ӆp����fK<|���b�-�?F���)��<E��W�N��j߼#TƜQDBZ��lE�E&1�bQ�
�$�1H���'p5ў"~Γ���@֮�=1r2��	���`���?	��-�0Uc���nq@��i�<I�t�^	y��މdx�r(S?���"�S�OΞ�G�	WE�up��&���1�'P�Q����}z�(`��&~����'����'��k>dT���#�Э#�'Vj���hV`�^0���6kΰP�'o�A��	կKN@幆	5�^�Q�'��-�#(�x�@҆�/	$Xq9�'ɛ�H�3a�ڄ�V��`�>]Z�)��?A�O���?��O����Aa̧;I m��Y?bfT2��$?�SⓩV��Q��4̈́�yR�C�(vB�v̩��D��JT�?��C䉚.���J��T�$x`�  �n�J➔���!&�@��*C��j*�PC�ɖ�V��E	�[����///[ C�	&b?���k��.�t�wA�I4ZO�7M1?Y��	����eHB�C �pص���(/!��7't���P�ф6���6��p"� ��'��5�УST�i��Q$F�R�'g*����^/3D�9��ި+�ݓ�}��'`xH��p�QXV�%W� �ˏ��x�P�~̧U��aе���t34	��F	&hvB���R�iBa(�.�
�h�#����'���Ey���Z-K��9)�-LU��U�g6.��{��x��u����Xƣ��h��'�a|���Q���c��T��]�q�B �yR���zw0�bE��#J�pUP�a�yrÓ�!9pö@��m��}�q���y2�O�,)\}�e�]�8S4M;`.��y�� �4�0RmC�0��"'`�"q��DA�M��CW�?v$���li{a|�|��g��uJ��</}h QC����~��)ڧh`��Iq��%4Z�,�)�Z�q��NT ��B�Wmw*th����א5�ȓE�Nt�SeT�-@��V.;��'}�'Jax��=K��bb�}��O��y��IX�ӃOٓ}r����d��M���>���AT�$��8�BA6���0�*;�OO5X�!�,���i ��<�xy��Oxd����S35����e(U�o��R�
���G{���>)�)<�� �յ=b���QH<a/�o0DA��¥pd��D	"?!��ea2�#^���7J:=�x҂	(��'	��t�§7�QR أBslr
�'�ԑH�o�@�j��"αD5����y �Ş ��5���ؑR�P�R���S�y�ȓ9"dM�4&�Gc��'�ˊo��M�<aߓc�1�g��
|<�`�_v�0��"O�����ԃ60(���~�B�2r"OZԇ��yS0�'M.r��LA�"O�uhs&Ke�P�"��Oﮰ�"On4r!�<3�t�B�N�C�t`AF"O���uj�>*<|xi�[���"O���o�C@(i��mF�,�\y�u"O*�p���:>���V�T��"Ձa��;lOX�ċKnź�K7�2�3�"O\���΂"b�v�!w̖�,��"E"O� 5� � |wT}J5�X;ۄi�f"O�A��b�B��P0��/-�29� �>Q���	̘M
��K���PކII��Ÿp�!�d^<8X�k0̆�+� �c�޳3囶�)��yAk�a:KSGX"i6�6�=D�h9ը�#J6 y`��7~K}9 ��OlB��:8ږ�:���2� �b�I-R]�B�	�fJ����D5�( ����(!��x��1V� LQ{���
1�P@�,%D�D����9�)p�_6�&����#D�h�ã��c}"�� NS�T�[�@!D�|�w��<UF�����5{�v�3$�*D�Pb�l�&]b�ˎ���G�p=)�y��<"/N)���#,�vP��i����>�O�  �Q�|�X<{�N��<�䅣<�:	��J�#L$ ��<#��P�j�Dy��>�H>A���)� �A9LA�1Ùy���"O�T���
E�a�����-:52�"OP���2���rI�2' A"O��i�*(�lP��E:C$PQ�'�!�$�%2*��K��_fąI��W T��}��'���ǶQ��а�"�wH\՚E��|�!� E��@��500|�CB�!���% ���K�=4���j��2�!���zL��`�͖t ����bka��O�HZ���6��0�Ъ]N}Ar"O0��BKU1T��ɳq@�IXP|#"O�y�J5:�����X����"O�����[��� +�;��9�$"OH�!���$@&d\BD)��s���B"OL�Q���%
��0�OX:�C�6O�b���I)�.�BE	;6��x��G'N��hO�>1�r� �y��(��� QR���!D��pBѴ�^!aAY1���W3D��"Ď�8�HUH��m>�}�52D�YW�5z4$��&��Q�.D�xPt�M#u�� H�>m�ri+#�-D����f6w"X{ ��h���r�,D�8:⡉�}<3'N
�&%�x��*D��Q�Ê�7��3�TA���
A/6D����љv����&�#����t��#<����i�X��5��O��ax�gF?4:�L��'�d�ːMѥ'N�豢Z\z�q)O>��~��IS&�1m�P�R`��� �ȓyzċ���8c� Y��2*ʤo�R(<��G���,}	�>,<h��s��r�<Ѳ�ƺ, �@�řNj�HxU��l�<yw��/s�s��P�FO��W�EѦ��U�x��'=�`S!�eU���(����	���'�B1���O�}�NHi �� �Zع	�'_dU	�	Q8��2��LlE9�{B�0�S�ӎ93n(��ȟ&�����KL.crB�	�jmp<ےƜ�Ptqa��b���<��8|!�!kR��E��#*X$�@�T�,��I&��P��b0Jw�*fȊ�\`7m؇��?���Zz8 ���=2t@8�@S^�<iTbÁ4�(����)�\���o U�<��-2K�$	�+߭@��8rUaWT�<��<xkՎ^5t�^���R�<	��_N RŶ1k@�dE�<1��j��(��/�,��h�1L�U�<I7�S�$���+!ȟ{�~��GS|�<y��"�n�*i��T���Yv� y�<ffS&k>�I�a
IVՑ�+�z�<� �qsP�Օ, ��rAWp���`"Ol���T70���e�[�6�D�t"O���dF��bv���T$y���G"O ���pc� a��E�fy�	i�"O$��%j�eOp�a�l�\c��1"Op�U��6;|����*H��T"O��K��<%|h�u�&B�P�7"OL$*'eX�U�����D
�b� �Ї"Or�Bҿ�x1��n!��y!�d�~����ٛ,)�{qIB�u!�$�na����,�Rt"#	��75!��)8~�E��Z��[�H�8!��:O'�yp��t����$͓�!�$#Iz؝R�#���za�G#̚�!�䉅I��zf�gH0mC����!��LF���������,T�F�!�D+�L@Cw��{���ЍǙA�!�J#?&p�T�:�yՁĭZ�!��DӀ��T��8~��t�Δ1y�!�X�1�XĒ�eC��x��lՏ0�!�$�y��T��!���p�!�^4�2��%G?zS�y�� +W�!�W�5e�����=4�ѤC�?�!�Ԁu�j�������G�0�!�[�����
�2#M�Wl���!�ŐB���B���&y^�"��A��!�$�
��:q
$9�0�@�E��!��6<܁��D�]��Ɉ�l�!�DX.i.&�J�l���ݱ�h�I�!��˯���#7�SU���&	��~r��(�d�@�Z�wx��
%���Y���y�<`σ8,�Ha��ȣG�^��CNY�<�D�F�Z���P#ڧ(��`I%�q�<ٳMA�M��y!B�$"�{�'�l�<��(�/ T��2(��c��S��a�<�v�����Ѩ%JO�6��C�BBf�<!�^�V�R����N����T�D�<�3f�(�|�"�N���P��k�<�bN1-��k�
p,2��`�<�oV�$U�l� ��u�0�c�<F�(-��% 竔�K rP���Xr�<�R���_����s�D-k� ��D�A�<�%
Ûy���`bF�":Y��B�$f�<Q�j-� �s3�ۤ\H�@�b�<��-W-
��m�'1��|�J�_�<��	�E��L�F�K�FpK�EN�<	C�R�`����DKG0c�V�Z��D�<)���$���3_�8���,XJ�<ipj[ph[��Ϯ~ՒRdCK�<y�Z852N������l�x��hCL�<	p%K�*�)��9T�=�3�N�<�a!�9	:�9���?C_&���v�<1k�C��# �4 ��ٙ��YE�<��k�C��a�e��(9�Y6�CE�<�`.�5H�\�����a[r� �c��<th�x8z��U��mH5�[b�<!q��C�jg�̕lsF�Xe��`�<�nVj	����ֱ��f�a�<���_
pZ����X���Y�<q2�|���`۬|�J��EZV�<	��'a$ 1S�'��D��I��X�<����0-P��R� A�x)�	A毉q�<���@�8 $�9p�%:]����n�<Y�#�2 ���>}�ܽ���r�<� $@:sak���?+18�!�"Oe��A��]���AgOY�'Z���"Ovt��e �t��A0>�XT�"O` ���)'`�B�nЏA�,�"O��S'�?�E �C�~���U"O�D�B�� j����W��Ĝ07"O��S�σKa$��3+x\�t"O�I[�J�-f�9@r��Lo����"OhP�e ��~���N;T�����"O���֫��%���'S�rh���'�pl�ъP? ;ά�d�M-"��%�b��Q�
�P ���O'!�dY�d�X� ��R���g��j>Q�L��#�)e�^�0ȅ�
PK1��L�4y�����'DW^I�R�ÕK!!�$҆h~��,�7b�$�G�+ e�����;�ZXcF�21����s����K3EP~'0����DS8�!��T"N��A��/<V,�0N+Q�H-���$8|r��3e����2e�O����J��J.����K6V��@��<lO<x����!MҀ��7Y�|2��X@re�Wŝ�_U��E��&Q�^���uR�E���ݨV1h\ٱ�*���=Q�5ʓe�PረO�h(�$u�1��L�\x�&"O���2	�H$b�hVd��Nb�����I�>0������|�1�K��DÞ�J�\yQBI�p�<�����
��	�ENP�A����*>r����>�I�H���ēf>HLٰ�!TduSQ�J��<ѐ��!֘'r��q�O���H�٧��<�#�OƍHeʎ~���f�1u�a9!)Έ6a�a��$�N7e����K�L扦;�D��<lC�|C$�E�FC��^�����U,B���(�D�㟀 ���NIEx�OX���S��s��k�$�Y�������?�3�@ ��r��m����(�t)P�Y��O��l��'�X��� S:t�E	�H�d��
�R2`��y���{+�DA��e`�t)��0��+�ļ��aEa�T'(}.Z�B\��pi�3���?���� �?9��ק����Op}���a����@�| ΍!�צ��'[�P��ħ+��ONti
"s4��$AØ������S2���D{Zw�@=���R�=��¦�!oc@5Q��O.��K��b���?U�"eZ,79� ��gO����:��.V��z���!P�n|��AC�.�@�œ�9;�B��:3>���l��{ �s�b3}*�C�?D�����W�Ѩ�zQ�*H�C��9C��$Ē�@
���''׮{��B�
6����f�_�a��i&��\��B�	�/F\���M��1F���䇣��C��=rI:���@8�XС�I(��C�I�|,{D�%�Ac
'�C�Ic�&}т�_-ud�x`���+2��C�I"���rtB ;��`#�X�f��C�ɕȔB���' �D��itC���ȓSs�5�!�Z0�Lh�CA� C�@�ȓE8 ���F1L��SbR?[�.��'�ў�|�Bȅ"QX\d�۲&�2���g}�<9�եNw�97)S�����w�Ii�D4-�_�ZjuO�#}���#8�O���|���7�R�T��<�5e�=�!�$�6M���y"�X>
z������<�!�Dے}3h��0k^� ���#4-�!�A�V�t@�s"�m��"�Cثb�!�dH^�dD�kX-iv����Z�g�!�UH�3sA��a�zb�͖�A���Y��H�q�QM�N�|d��-�b��A�"O�$�PÜ�!�1RWL� ��Љ�x��'I�lj���'�^�˄�<]9�$����~2�B� �`�	�o�O������y�EFD�F���@9��r`ё��O��~� :��O��g|
 ��f.F�9:"O:L����[��%�4��n�J�2�]��F{��)�cO4\@�K#4�0y�ۙ?�!�DL�!3`i�B��0����W
X�02!�S�n�C�Ŝ�-:�"��� .!��T U\� [6D�> y"�R!򄛞-��5��c�4~bE{&Z?llqO��3ퟶ�0|:�EW��=Z�BͲH��"h�Q�<!��$�D�4��3UY�i؁�BK�<	���\�)��)B��H�3�d�@�<х�L�F��\9�c˝8��, 卉Y�<P-��z Ȩ ��c*$�S��r�<Ʉ��':VL�6�r��[���g�<����+wّ� ^%C����u�<�B	�!n�Jl��R�}����As�<A��IN
��d�&W'd9��Nl�<�5�v`J�j��ݣ4}~�R��[l�<ya���>��$g۫.��X�"Mo�<y��3y9:=�b�� #B� gOWk�'�v�j�͋3x;>9�r�)0J��}���)-��	!�Ȉ�!�D�L���rf�΅vj �n����d\�f��Pp�F�1-���,�s�]Ybճ%�	N�%B,D�|cp	�@����%�I.	��KG�7F�H��ωX�����ٹer�|G"oZ)w�F�:�d� &8��PF	;�p=��ɎE�8�y�n�=k��e�cއL�����7ob�И�K'L2�u��z����%��G����6�̐h�N��<���j�D����.y^�QT�Ώi��O��HP��t36e͔�$�	�'��!�뚉s��x��J��L��^#<��� W��d��T�ϔ���O�"E2Op%��a4]XjI��K�!!���vO<xP2瑿V�,5�t%�(Xv�M��5&s�K���JP���'�2˺HCg�>�hOdU��5fzD�ș��E���<i�'2�����疩;�tu�u$&fN,hD�F�G� c��j	,yR���Gfh����Y�8؊�W�����*V���'���%�-7�%��X�_nԲ0"��8[Z�B���l��M$Ā����;\�B"O��`�I��HQ����D�Ia�.�r�@ٴ%�����䙔F���$?%�pDٕD��{���c!��%W�x�#TA��Rš�
=fi�p��0�t�e@;L����%i��Q#-�$P�S$۪-m�H��?ғ7�j<��E��mb�Ш��K .T戅�ɗ¾��3�_�+��`��f�;E0usQ�f�h�Es�P�b`E5��I��NX���r��+%4`IC��9���M)}���<~����ZT��u�'`���S��~��S-:|$E����.8��	_>N�.B䉎�}"¦���A�|� P�Ф$b��9!� �ea��įW���'ai��!�/w����<�>�j��H�1CFuH�2��A�똼q�`���� =Lж�b���Uw���hמh����, �ڤG=r�p�Ezbn�.Ӳ��K-��ԨĈ��p<�"�ߒ-b�8���� 
ޠ3r� K�8�!qK�*�0���)E�
Bh��DkC���R���)N1�O�]y�-W���q� S���#@�>�c�,��Y#����-��1B 
�3��"0J^�����,Q�6yV��!��o��tp���O>��Uww���<�}�тU$�\eU�
[�l5��IX�$Lm��OT5W����ի��+������D�V�(���̻o���
f�)V%h��,uRBԨF�)�D��vUV��~�'���:dU�p& ���Hj%
܁K� IՈ���D�H�S��=�dL�V��Dx�*х>��y� fT+u���{P�C�Vt�c�Z5d��\0*�;E���G�#k!.��䍅�K���T��)M��3FϘ4,HH�d��K�,�Fx2)^'T��-�W�>!3��l ���7>2qU�]F�$X.mtp2�J
�m���d�L������F�&!���'3�bՐ�X�#ifiU�
%_��U'��0r�ŗI�J�'�b?�K"_|n��F�	d�����
�g&�Ձw�׭m�lq(�=����}2D�LR��'7hX����U.~�PT`�%C��hJ>q$ F� H���ɓZ�h�%A&"d1PÜ�n��e�]8x��� 2y�-F0X�x�u�I_�X���`�z���G�Ġu���8��D�}� D|Bo�?{� �0�n^ ��x���J���2�!%���:���
,f�0��]�."��|9��{�B��Od����	_�"���k��"��$��j�
�
�G�O_��؅��C���N?Q��EΒkl�HɲM�wi,�pU�,��un"�Xu��)�� �Q�A��?O�8�a���!\�+�[�����Dӝ7*= ��C}b%ř]�0���pz��'AJ�.UV�@1��<� d$�������7$_]�Lp�dFK8	cQ
��}G����AFJd�?�@�59p=!c+ǫR������I���"u�Ph����p⇚
�"���E��(J'%��!�PRN<��D�'7T��';x����c��y�'�*���B'5P��7�闵.LN����2 ;�#� }�!�D�%o����&+��H�	B+;�!�D��p!�ꀇ�Q�hCFȖ*�!�dѱ!Ǵ���|�`�Uj۷�!�dK8(�pPCf�W��چ�q�!�d_�M��qT`\^�.X3� �.@�!���F�Y��N l��-���E�`�!��
c{�᪒��N|(�B��сs$!�H���4���):j�`�bS�u!�dV�Խ���ۨQ@،�F@�p!��ޠ~�%� ̄#�`<�&�?}!��X��h8�➗�.����=!��Z~�SF"�xy2ǥW.8!�dA���Mhe�,d�N �d�)rO!�D��3V�АDA�y,�RB㗼G$!��7<��u�$g?eQ}c��^�L!�D��Z�����1��p�ǦZ�H!�/%,� x�)R80��{eJ�`�!�d�f��K"�H�2{��M�J�!�,N�j}z��2Dh\`��N�8R'!�!W9J���'��)7��+D�!�$H�l@|����M���R��&t�!��>u:���lT3Us]��Z!�R����`օxe^LҶ�
>k�!�d�g�RP��5P@f0jE`Z�n;!�䐩B�(�$l�Σ��#�a��"O,HBuI�* BT�Ϗ�+(��g"O:��oğW�,mr���X���'"O:����A'-C��u��<֞��!"OH#3Ǒ�BRx{�"в>�xh��"O�I�$$��rP5�C�&:��՚g"O@��#�2#=�Ւ���M�L�&"O�%ۣj�(�1��
����"O��7�;xR$+'
!��h)�"Ox�wD��(��i�1iA��n��`*OF[�B�&v��Y$NʐYhi��'��Ds���<�]y�!��Pj����'�<��0MQ��Z�cR�W���'i�����	����tꄡyۤl��'"�ՈЈܬn�Ta��3m��+�'{�Q�"��N�����baʔI:	�'�� ��J�01���Zc P�Q�����'����G���ݱ����TJ �y�'W�"��;��́ �L��'�}�uI�L{��Њ�`NU+�'g䡚�E�:�P����}.�t:
�'x,{5$N�3�ؽ҂n۱r����	�'�ѣ��fȐ��R�&�u�	�'�����-R�T@��A )e�y�
�'2n�k���� "�������'qH�qE�:Y���,���(��'<��aƏ�(l�@PR-A�	G���'qd��fAZx� #J�{�@4�'��r���PY9�:~��
�'��b��X�mnBy�%��~_�ņ�5E�E�P���m!��6���f�����i4���!��;����b�"4��C	� �C7Nz�=�wh�5< }�ȓH��5�q�ÑlaB���O0V�z���s]� *A�͖�t�ʡH.Fn�C�)� ��Z�Ų_R ⓠ �F-�2"Olm㦋�~��� ���
q��=i�"O��q��	�'��26-�}���"O꽈�R6��0�ң�?g-:@"O4ya�@�c2��Y'!�BzZ�"O��!�M;/TlLyDA
92���@"O�\�D��8��3�I�4���Q�"O ���) �:`zрD�h�,�r"O"� r��V.��#Etm�$(s"O���fN)@W���!��9�t�"O�)`�
>>�"i{��=.]��s"O\��p	��&B@� �bɃ�"O�L�ӫ �U6@��M��p3��_u�<��MxZ�H�$�>Ey��t��q�<Q��S�^��B�oM>[J�]SQL\m�<����/:��,aCL�l���-�a�<Y#����H)B��7�
L(c�@�<Y��˨sFعx��^�#[|`d�B�<�`Lх+�*��1d�'yT�av.�C�<����,�^���-ơf�d���UF�<��W:i��Eа#�	�Dkp�TF�<�0�]4��a*��G�T������<��'�S�<T���w* p	�K�y�<y`���9���&A��Sr�� GNO\�<)"K�1�A���~Yja�f�w�<���V�j�&�s#/�?xD�&Vn�<�a�_?!+�q$i(fV���@�\�<a��Mˠ�@gH�$u��i�3��g�<	V�Nh ��P'Fu����J�<���7����Q�]�W-��E�<�2n]X�r��,�8`�/�Z�<��
�g�fm�х�>�#bM�U�<ѳ��J��3m�}B�3'��~�<��'�C+­mJ�zG����g�<���;�BQ�QiP=OU2ͩT�w�<�1��T�43Hٕk;��o�D�<� bȈpvZm��-��B9E*�L�<a�Ȅ�4����JJ�yvtY���B�<����}�>������(� �w�<�ԃ�#�q�m^�.S�)1`�V�<	qBYU���@A&���(��3��P�<qDD���ЊӢ�'�*�i� ^p�<!���v̖����@�y1�U&�o�<�PB�=j4���)�.@0��A�<�%�%#���+��Q*����"@|�<Y�!�ޜٰ�m� �`ų��~�<��`�o����re�+���k�'�V�<����_/ � ���$F�=�*�y�<9&L��dRn���@�*!~Y��	~�<uK+�Dd��`�%>Q��pǃ�~�<ᐪ��vj�E����@ �S!�M�<9P�H#~��x��[@R��`�O�<�&Q�) ������z��5��K�<Q$��#~tU�S� f����ςD�<9�^�����	�Lr�	���RM�<��,J?t�]h��[X$5@6.�N�<!a�$m�ݫQK�:8|\@�m�c�<�6���б!�w�T2@��_�<g(S�	z :�션����n�<ɔ��a񈥐w�L�pb�2�l�d�<��iȢ&~(<��#נq�,�*B��k�<���S�D��u07�F�2��ف�Kh�<A��S�4�85����ܕQ�Yo�<�%�b"h��N#Q�!36��n�<� ���#�$H�(�"�6ԃ�"O6u�0i�
v�@�w���P:D"O�Y��� z3�9h�ɐ	88��"O�ya��
�m1���2P�T"O }�`�.t���b��:7TP�"O<�Hv�bD�2��E���"O��� �+�]b�+M�|}��e"OD�B�ٞ�$M�V��;Oo�P��"O8���?��E�CNI3g�X��w"O�!w�]�� �"��"��q��"O:s���0"�5���ݪZ�:Q�"O�����	��	S�mΊ*�$�3�"OLIpEk Gf�a���} �"Oֱ��i@.����3��2D�"O�AvaتA��B�67����"O2$��Ͳ ��UJC˿jٲ�R6"OrQ��	�Uf�dA!M+�H�	�'��s����d� f&J
���'��9��W�D�R���gʄWX��a�'�d@�EK�c�6�8j�Bl���	�'\�`ŌݜloŃ�D"a �T��'�H�aF�Vt����aѦT1�'�$hw�P �X�"qi�w�4;	�'�8$X�G�J����.����x	�'8	�Fƚ;ȠH�gk��gU"��'��Q����M��u���ש_�P((�'��H���$(؝��)@E�P��'��=���%|m�]���8A�$��'U��;��P;79�I��M�9�J��'��}Q�$��q�Z���� fİ�'��M��hS$}tbT�#]=��[�'V�h�ת҅T<�A�L=q��H��'��T*���
DT���烑l�v4��'�$hS�A/b�ѠeҌl����'Z���iB�J�$\
��e�t��'�2���Mo���Y�v<K�'S>���a�8n��X���_F���'�4ZrŇ�uq�lˤ�4m�Y�'T!�T���c��S풧���y�'�Ƒ�&/1D�(R�e��3��']�Z���6��:Ci��0�����'�%���и+5\b`6(FD3�'�嘆��m,����+G&�`�
�'�����+�[���3$����
�'�*��O��g8�8�O�l�<�	�'r�����'� ����K�
 �	�'�*��NSk�Ƞ�
��	"�3	�'*h�q#A�/eH�4�rkѲwY"L��'p�TYg�C�s�l8��cVb�}�'����C!KH�IQ�1d쐵��S`Z��K<qń�e��: ED
i�h���&�^�<@�I�D�@8�7��9���b�[�I����2�&�)��.7Z�C�Ȕ�,lx�y$M�6�C�&��T��mT(y""�ؐ@�#IȾ�Y"�|��P�J¨b?Op�x�o�2������ȧ@:ai%O��;�N���<�#恷?�@D*��
��B�(�/�OterAŞ�q@ k���s��`�c�'�,HfB����"q�Ũ�o��MYFj̺D0��>���ڇH��j�!��<���&�؀㬖�=~¹'�b?� \X<0BnΞ�5hq�Q	�HC�I	M�m"���'cK��R�N&gS\M���|��`XJc?Obm���\���1#];Z����O@�"��S��pX;���Ӫ�p��� G�*Y���'�O�l��W{���0 A�Xtx9��'4���� )��S�? �8Q�gŝ0WbU�G ��l��)�"Odq�`�Q-��`s%�r�> �R�|RE[!q�0��y���:q�XPS@��U������/�yr��X)��h�ݤLp�qcL��b(��i�<q�`/}��y�ѧ>��(vN@�<��銤[�P3�,KE��1j	Y�<�K�VI�q�`�̕u�楩�	�V�<0�Qw�����W+N�`Y��V�<G�\�X��ñ������	Y�<y3�ͷR�་1�*E�}�f�T�<i���a��*��Y~br� mKY�<��"��O����	�?XF���O�<i \?m.�c�h�
���H ��H�<��k��S̜ɸ�ǎC��5��n�I�<Ib��tϴ�G�ɍL�(�2�-�M�<�6t%�Т�b�&B���Cb�<qk��V�$8@���.>���ըOG�<�@@L?�H�Hbb�`'[V�<i�M��09�P�2K��w�f٩�ʋ_�<� `�u 칒aS2KJ�0��W�<)#�>E��P6&
&�VP1�/AS�<�$CX�e.p�����Z���Y�ĉO�<��.�.0��b��;�\���R�<A���@��m2�+Qe.�"1��L�<1���B��ܙ�Ȣp:����L�<�E/�6\ 5�t�ƫI���JB��f�<�V�­	�@@A�� gr�y�3��f�<)���{}�u{�+F�-��4R�'�X�<Iሓ5M���%�\�`Ȅ��� _Y�<��9a��(Eǎ3`����EC�<١B�,-��AE)�Ѡ�
�y�<y��ԥigT��Fi�*x�(����S�<�����O"  RF�W�ys�h豬s�<!��I��E��Q?K�I��'n�<��iI4VZ�dDQ&جx��B^o�<9
�	��ҫ��l �D��q�<ѧ�C-6�5��>I���kSi�<q��8h�N��d�^THr�Wk��8�5
��4�`#$�`�n�2GV`�1D�@��?V�'Ub�d��<�'���\n�:L���a�-ovx���G+��n��͓��)�' n"�afd���T�"`�#�6ϓ�y"��9ړTuЍYw��^}a��K=t �%B���OkMǞNu�m�s�R����=�S��ㅙyô�(�ݙ,.*=�1��'/ўb>�Hs�T���kd��Y�< 1�m,?��ᓖ$�Ҕ�S��z���F�
[�|�	Y�����[@�(  �L�p"�?-�١Tęp�'Da��gy	%��jǁ9��Gl�9��'�IDyJ?B��=C��·jP%Q�v�`0�1�DP��(O��>ٕ����t�q��~���2��z?�T�������^�a�DD�7��e���\�԰���/"Dyk�&�~��e?E����'8���G͂,s��؀ѢN7H("<�6�w
R
b��*�-���P�6a�l��
�$�<��z�A�͓>Ly�7� ]���r�|"�\@���O5A��A_����e`�9JU��!�Ob�=E�4�A����t�T2#�r @�"B��yr�)�'W=���/	�9�4�x$m��}a��z��!��hO�)��j���k_9zM�U�(��W��`E{ʟ��*šΪ
}�Hqd�/~�	0��D&�S�'b����B'�!�fو D|�t8�'%ў�?�H����3�������-{���lF�<1�'���0|�c"^����;���1U�2%¡�H �y�>A�'}N��O��)�|�3G���$[���;�@�IŌ��M;�AB�d�VQ�b'U(�0=���Z!W�(�CDކI�^�q`�j�<� ��2/�.P��Ȣa�K(���"O*�(5+9sk�<�Fo����98�"O��CˣPbH%���#e�����"O��嫍<�,���"����`"O��G�"#����͈d�HA�r"O$��vf0l��?e�"qzF"Opa`�S�)ː���e
tP`�"O����$VHl�T�,G\V<s�"O�Q��޲^���0a�G�DN���"O�Ѐ�j����ЃH��_���"Od�����X�T])��C�-3m�b"O���C��,��;7/�=-�0qv"O(�H�@^�!������D�r+Bl"�"O̡�F�� rD�حq0�h0�"Ovt�#��7�(}�p�ރn��+S"O�U�&��q�1��X%!"O��9��S�B�E�#�ƥA�0a�B"O���h� o]Xb�J*�Pm�c"O��#!�$)� a���p��M��"OȠ�d�8)$�'�X:1Ϭ�1�"O��21�^�FUd�񣗮��t"OV�K��ێV�^��F�і����y�NP\������݄�̻ �G��yR��j�@�*h�?¢�W͙�y��Ձ1 x��2
��{1��q�L��y"�W	g`�5�%kٗs	x��B��yb-A�/��h�Gϖ�j�H`�6�>�y�c��D���z�ĕf����9�y�ߗs
$����T�H�����yb��/!'¼qV�#Hø��WE�yR���&@��jbC\38Ռ��A��y2���Sn��SNՐ�: G�)�y��� ?���� �[<ڶAې�yr�3��<q�Z.
r�#X��y���7!��<H�R,���ǫ���y"��e�U'O��0H�5o���y�.>1��9F��$��P䬊��yB�@&.���f����3Ռ��yr���^�q�t@��[zP8��Ź�y�`��XL���,�tG0�������'��(���~/:�+7�W��I�'[�,�2����t"�$W4M��
�'V��kvAY�|��g�s,�ՙ�'\��Dӥ{�Z��j��e���	�'ot-k�1"Qx�  �B)y�h��	�'f�HQd��#@���W�&k.@I��'U�� �n����G�u>��[�'�2-Q4C�1u�� ��h$�
�'j��
��1�@/���
�'uR���O�D� EԌ
��T��'Զ��%�^�E�8Y���[����K�'UxDa��V�w����y$|�����9TeM�m�D�[�]����N�H��,�d���;�PQ�ȓ�%A T
8��>7cb��k/D�l16,ߝl�0�Jb
 j �?D�+���G)挘��]�D6AK�>D���5"�d��q��,�6�����l<D��Ǡ]�R���)r��,����o%D��K2��K�B��Ua�K{��X��0D�ЁU�$6�
�rJ^�k��`��+D���2�K�Tp���4S)D�؈P^m��A{�K�PD���&D�@�#m��`�
���� T�0�2C1D�� Ll��]6Mꐡdm��,�8-a�"O ���u6���ȅ����"O�|�uD ,N�mx�Gb��m�"Ozl�j��.W� !�MB.{�	�'��A�,�b�H��^��T%��'�(Y��f$Eh��ӥB��T��'�"�hvlށ�Ri��'^F����m&����N\ |�A�]'N�nY�ȓ$��U�Ulɬz���Eh':�z���=�*�:�͔�VU�a��%Ζt�ȓ�T\�R荩5���ś�� ��XV�	P�V�x�l������ȓ�@r�$�=��8I��J�4����I�����4J���F��cr��:�t�`˟�:��0����Oxa�ȓ^7\�óZ	U<�hQ�*)���ȓ5�|�am`fl(��Mi!�K_[�<I�Gc��(��G�����k�<AQ�Z��*�P�N����!�
�O�<�b	�
h� a��g\�tn����t�<����%��"���
�����m�<a� շh_�d1�eX�#����&
�S�<1@�0��)#��W0%��`��N�<���y5�l��D�7%���Em�S�<Q��߁{b��8�%�>�V��*�R�<�B�v�:s�N0�%N]g�<!��^of%X���%!�~(	�O�e�<Q�	O�I_4\��A�7u��T�s�U`�<qS"��/�ת�4)�� ���[�<�4��<i���q����:�FXs�<��3 (|)h�
U�Y b+�$�q�<Y�M6x�05{`^* ��[���o�<�q��x"N%�T��iV�IM�C�I5i8�t�����J9AqX ��'+\�r�nU�>�C �K�6�8��
�'��C�� ���^T|�B�'h������OR^�i7!_�V��x��'�$�	'ǡB�p�j�'�F\���'����O��E��!�U)Ҡ@�۸	�'z�����
��|�L�7@� �B�'�(�:`ȜZ�a:�cX�<����qAS�R,5��wI�?�,�ȓ
�t%qtlD1M��X���Pg��ȓ`��y��MLe���'��ud Q�ȓh��cƧ�.}���AӠL�z�1�ȓ/�D�pO�� }��=0K"\��;x0Xڐǐ. 0��_�_����zr�Z�J�/zl���H��E��ȓ1F�(�$@��Nu U��SPl�ȓ^@*�TH�6�NĢ�j���$�ȓ)��x򀨎�
�Xd�5(]����mp|m�g&!s� s���`��̇ȓ#���f/B5}gt�;R��7��0�ȓeM �Rj�>B��qC4z|e��LX�A�f��YxH[2�,_߾��ȓ�����C��i���5 �%G�H��ȓwX�Pnޖ�`��s�M�{�Z���YZ%!�k�A�$�0��#�5�ȓ�0I���Lc��;� 	�vT��5��p�
SH�"7��!���ȓy^�y��S�R���uҿ%H	�ȓ@V�#�+V=ǆ�˕NѺ[敄ȓW.¡��J/E�Ik7Y�W�Pq���i��նha~�%)40�6���S�? �!p%c��cA:�@�3R!�x�"OP�stѪ)�FUѲ#c�l#�"O^a��w	�ei�I�O]���a"O�|�!��������o\ $�"ONt���]�?}ȴ�@G?RG:$c�"O�=���/	�L�ӀҪ|��Y�"O��J���k�n�� ���D�`�"O��b#]�B!��]�>��#"O,�qȆ7�T�'Fɲ4��Tz�"O>�2�l�/},ڑ�G��Q�Z=�p"O@�@�>?LU*56H�҇"OvX�q�K�U9���.����[�"O�904�� ��uX���x�M���|��'�
�@�*�*I��kv�L�O����'����պH�,�%KX5HWF��'�DWj�o�����$H'ze�
�'u�:e��<��"F������'F�)bפĘm�^���!�"�9�'|�@�ei߁XL�� 7$<2�:
�']�|���G%�LB�����
�'���xB
�H��P8�#��vD�ȓL,�����ަ���Z�K �q��P�L����<
�8\�V#҇h�R��ȓZ"��c�T#vU�=[���c9�t�ȓ|u8��sJ�K�&��ͺ'@ �ȓ#g�5r4k߄<�BԺ�K̬QD"��� 䬉*rK�����m+	'�m��Q��!��j#)��w��h��u��fֶ�QЬQl,�Zl&0���ȓf�X!Ъ�)䉁���j�t���G�����EMXP��'�Z*�|t��_U���&�7��Q��1���{�2(zA��4��x�	�3�"��ȓ?�Ux�	܄(&���̈wS4��x4h��Ğ�U�ze�"�ȋg<h��ȓ*R��e>�~�����mw(��ȓ\���g�oOf��.M �.���|T�{�9-'��Q���ox~��ȓc�������<M�D9� J�/Y�<�ȓ�9��!Z�{�R�� *�'�<Q��c�P����Ԉa����E�ȓE�� �Hͧg�dLȅ�B; *J��ȓ,�X#�I�S�viꦀ�m,�ȓS�*��L��pMZ��HUR��ȓ5�v���S�s؉�i˖n�ر����Zt���j��U���֕P���q��!����s��!�@	�P�Υ��?�ޥ`�I�.�x��E�/�=�ȓ��L*�
ـ|P�H"%��Ņ�~���c��&}�p�)�l�PBn��o�8$BpS޹���M#����j���K�2
�fP���I�W��ȓR���1�5aY������c�Z���b0Պ ��:F��u�VL+ �u�ȓJd��PE��(D9Z�3�>�b�� 6M@�%T)7��lu�T��ȓ?$A�����G�^��k�$O!�^5,J�s����}
#�D9&�!�$�>�u��ڛN�9 #cH�"�!��/`��Q�ͬs���C�0�!�d�)--�B���*&����Aغg�!�B�<ڴ�L=^[ZX�"!B�Y2!�d��)t����m������t!���6�h@����!UD�T�!�� ���� �Nѣfe�6v@^�+�"O\�Q��E�8����^9`CZPH�"O�̳WN;G�b%���^��Bh�`O��$�HP�u��#ph�H1-S�-�j��"!x(���	ß4��ݟ��]w���'�bf�6u�*F,�9G����a�+#k.��`&�2|�0	�'04�! �# ����䙱[���a��'2��,�0��.WӲE w�N�(����Ή>S�pst*b�4D��]3�"�O6LIv%>@AF ����!��Ec�K��d���'��O��$�ONc�
��	�B� #Vm�'[�pq���!�?1�O7��O1��Ov�K��HX axed	|��S�cW���
ݴ�?�q�i��7��|Jp�C���'����ʢWJ���H��5�4Qh�%A$K-����Ol���i�O2�d�OH�s�O�-�TaAգM�y_t(��C؅/�(ݻ5O��X���Ր>QZ�m8O�:�<��
^�0)#&���ddc �P�]|6`���,|�ͻu�ͿuF�HƅN8Z1����!o8 �'t�:��ܛv#��+�
Ň<I� ��V+�&uJ6�����I՟��?��'��G�PM#甧e�v����S?�q��F~^�"|j&k�%/���
%�J9x���H�h^\�t�i��ɵt^m�ش�?q���)ߵ=� 7B`=m�6#T�p���Z�r l���`�u� �{OI#E
�[=�I+�$TF�R?5�V��%`L����ת=�4�++�$Q4n[�i���*8�g�M�$�H1�|��φ��8�1��ݢi��(#��{��;E�B�ė��{ش�?!��d�	{<Q�ҩM�B�R�o��'BQ�0FzRo�6�X��f �hh��a&��p<���i�6-!��˃Qkj'��xF���2]�Fƪ5����O��_�0���O����O���Ũ="��r-��<����݊�?�T���*����"jC\܂�/B�6S �'��Z�t*K@ϟ� ��3e�Np��*-$G�D	#kU�5���E� 
{��Cf˗0��}!I��Q���'
2p��<�6=y`O�^/���A	��8*�� �i��h-O�������?����M��A��e@��S�&u��԰�L�X9�y�?�Ƀd�`��.�q�Z��>V���t�شn��|��O��U��qW& ���U	 �C�U"k�Kf����BT��?���?1������O��$�O.�p�8��N%#WR���Î�q=�t	С_�^��:P��<>hԃ7sQ���p�ҫsX�`�'3�~M�2�M�*6�RA�#k�K �ؤs ���F_�c�س�&=扷b�z=S��
��4��(8�4��O]�tO h�🜺Zw*�O�0�/A�!��t�� �|<�x�'�'�
$�Ř#[d��GB�����!�����ش��++�9o��mZ�b�Έ�B'Fl����m��.ަ4����?Q�D��?i���?�"�H��$�ʌ- �t��6�
5"�V@N��4��q�H|��t��_�Zl:,Fy�#��,�tL�r�ƒN����#�.GB(p�C=o�,���Ig�PkQ�H�s
�h��C��RO��4�'up7�i?��lT�~��2F�f_:�ppϓH?���?)�ʟ�����V�2i0-Jd��YtxDy��i>�	s(�:_ԕ�� P4do�A@�N,;m��x�4���?a�����^Xh �  ��SslܮH�FC��!j��u��C�h�j$�X*^C�ɝ\���`��L�_���`�?6RC��Q���s�e�^�9��F`�B�IE��3FI��!*^M���'�-�3%��z����g_D��x��'
�ӓS\ņD�4NʇG��'&h0C�I��/':,�����o�4Z�'_��������X�ٛ>���	�'"��Rm��(4�a��
�2-����'_��H` ���KD�%�&u��'���� �oѰd)wN@�Y�\��'�d��&i�m�Xa���X���'���k��Hm���e�
�x�����'�:���Ў�]�`No����'�@��-�.|F�@k\�
�'}�����Z�;�����]��|��'q�E�g2&^2L�4i�WR�2�'(���/��+��@�P	�}bH�
�'L�E�8Z�4h IzA��"�'=�ܐ����Y�̋�m�d���'�"$�0\��3@�hy��')`ų�bNE,}��][�$j
�'x��đ�tp�`��X,Z0R��	�'>���(ǵiMJA�1�X��4	�'Mn ��ݻvxh�a�� F���'�Ԩ8&�M+aS8Ճ��رA�qa�'��xh��8�0lɖ2P���'��cg�A\;��W�Ɲ#���'��4���F�g�4J���X(�',�a��<UUT ȶ�ƵM)���'���Ra*9��IcHJ�U���R�'h��CY�:e���"GB
J�޼��'���A�<R�J���/��RW�!j�'pL8�p�É!{nܐ@슦BN,p
�'�pX����!�b�hE	oF��*
�'$�;���U2�݇>�|�i��!D�P�@��%>� J%$V�z�1�=D�\��ֈO�#&<��iQ$�&-�xC�)� PiS�Пt�B�iЯ�"B˜qr�"O�|C#nI�<����M�(���@"O^���-N���aQ�0^��Se"O, r.B	���M+n~�!�"OLi���S�4�A�Mf���"O�9��"_�Jq 	9E�ԲN����"O�,C�!�`��&�+Dpx2�"O�d�2���oCڔ����5)���#"Oԭk�D�M*��$_�f���3"O:(��j�Hk�:1DͶp��@�"OD��
��T��1�A�}��"O�v��" �xb!J)lƝ�G"O�uZ���,odt����cK"O���m�{��Ȩ�Ƒ��O�*�y��M�8�0S��v3����y��C�P�x�S��#D����dS�y� ��R���[�>y,x۔�/�yB�R�p>��)&��7�ʩ�2aհ�y�R�G�n)����2�@1hL���y2��^���qlՍ
vf!#��ybǐ8R{����'	����y2iM1M����e�l*�1��6�y�_!!�:]�#.ǉ~z��5,���y����~�z��J�jY$�B�Ф�y�l��\�8#Z�dZ�1����y�
?U�XeS�+IM`�t���y��8�6�{t�KTZ�N���yr
�'):�Z	��nUb"JG��yr��<C��G�~�R�8��Ѳ�y" �X{��"�Οu��պ���ym��S�e�p�5�DzrJ��y��w�PY1����h��R�˲�yr�C�Ȝ��o��Ԭ;��\1�y�<㆕�AjSG��;qF���y���d�\4Q�eT�B�x0L�'�y��D#�bp��۲�S@ _��y�DѬJ"D����'=b�X�ӕ�yLA'ROB���`�`l�x�+��y�'�!E:�Lҡ����!fKE �y2�̅[������
�ʩk`$ϫ�yҢ�j���֋�\�zB-��y�ʌ[�����J��ج�y��G���H��Ɇ6�xdR��T;�yb٣A��#��_���%���;�y�Z>t!��3e�yp�eʡ�yBDߧ���(�	�� �F#�+�yb.�J�(QC��	�XtF�1�y"m�4���G�L~7�:ՏU �yB����S%���y�@`�$��y& ���e9JC�?l`��À¸�yb��)���k��#-ք���Z��yBK-	����C1R����l%�y�LH�]�P�҉�F��a������y�J�SejA�6�A@��<[��݂�y�ϑ�4$��E	؄�u! �y�^+,��K!I� �d�#��K�yr��"	�$!��(�q�İ���?�y"(ga�)�)pX&��#���Z���q�'~�c/�2v����ǓM*���'�BUS��\	�,)q2��G#ص��'%Hax&�fgΤ ҆F�X���'^ �sCj�	r�e��A_�`
�'�D�1��ے��03����8�v�1�' Y3��cu4�[k��5]�
��� ����V��c�΄�^�Q�"O��7JO	x��i�%B�V����"O|�TFҎj� ���I3Ov�q�&"O D��� �{�N�b��j�0Jc"O�q��ÙgQT��ÉJ�a���"O����U4��\� �K9֨���"OF��F@4	<��R�Z 
�v1R�"OI�@�ƜsU����'�'Ro.�2"O2P: ���3>�e`�!� gZ�2�"Od�rs*�
nB�9����> �ꈱ�"O���������*w�<A~���"O��r�V�O&�9�EEO}b h�e"O����Ô�M�`��T�ƥ�l��'"ON�3'3��)
F�#��� U"O�1`�CY�V�	�	�1�v� "O:)2B�W*|����=���A�"O�t0A'�86����֦D��B��V"O��"Ģ��u�HY �k��D�jh�'"O>5�ɜ�^i�y�
9F��)8t"O�(��I?ez##G{�Ve���/D�L�q����$p�f ��@�ܙ�V�-D��{���"z�zHy���$B��;�,D�$��[!N�Sw�L*�puR�<D��q�	�2iэN�c씁��"?D���BL].wnR��SjȰx���;��8D������	00UI��	b�Xi�)5D���ʓBH�=�n�;� J�o2D�d�a@۽(S@b��@ZC���� 2D���CK�<;q�]��Lə0MQȒ�.D���3!�1÷C�[-&��N+D��Y2Ϛ+�n���ǕA�Psgm+D��wk��[Sv��!�>��}��"'D�\��ϳk�� #
_�;���h�'&D���֙K �CU�ۏ:�<Xش�"D��� iԀ<P!�.Z� $�s�!D�x��A��N\ڠVƃv!�!��,$D� �/�Inҝ��-Cavt��c�%D�̒$Ȩ�Z,c䮂�=�@I)W�"D�x�(1_A�q�V���L�q�cO"D��!l�� �F���$��Q�VO.D��zP*�a�nl��S �I3�,D�P�@�͹��\6N� aA)d!��[qtMz��) 
*�����)�!��בy3v�#dL�d�BboT9c�!�DV	&8�M�P�	������!�dP�#C��:d*��+�Z=2GJ'\�!�ǔ@2�����"6�<�� }�!��,n�ְ��$X��J`Is��$x�!��I�;>LP6 �h�R�DT�!��0~EH0�t��1fp0�b�X�!��$^|")���O6.�>��5�ک �!�Y�_Z� �V*�%u�𥛷�Q�*b!�q����q�ܿa�Q���3BF!��ڛd�V���*�|���G��!d7!�䃻U��鹗gZ�4��))$!��39m���-�8Z٨�H'
�!��"{��!���+o��t��.W10�!��M�Bi�d�G�0؀<�p���9�!�� �j���R%M	u��4j_�6�!�DI� �@,�a҇^�zT:"'�n�!�3�Q�%iW;q�9�--�!�$Y
{8|��bj�N\���1��<�!���y�ҁA���@.<;�lW�b�!�D ���Q��@ '.>0�D,%|A!�� �t�Z�yw�huAI�|�F8�"O��!�h��9�G@׾�jң"Ov�8�� px�I����.�FhK$"OT=���
**X�r��	;��}� "O��y̢8���RR+�-��D��"Ove�W�K�
*��IζA�I`�"OB�p�j�H�X�"&������"O��a�ߗ������G�"�"O����/��%�2��8m۬�0�"O�$Q���n^%Q�`J�C�Mc"O� �KZ�HF 9`�H�"OR�� ��>0����̈́=I�)C"O2A�e�i�@	�Ĥv�-p"O��S�야`{�1ҡc��Jg@�(A"O~��4L�2w.�c*b]0��"O>����ӭW�b9�p̑}>$д"O���Xi�X�3��!'�f��S"O\$ � ��%�LT�1��(x�H�U"OD�׃ߕ�)�)�
��!�"O.h����-3
�!x&�J{�iD"O���4Փ�B�Up\]�w"O��+$�5} ijK�8b&�b�"ON�K$��.]Y���gP�'=:��"O�y�m�  �B����4s@"O�e�6I��Di��Vg�jZb�"OZ���ʡ,��D̆c��*U"O�a#!�3_�p�YQ��7}킹��"O,���Ã�	�d@Q�h��k��5br�'B!��D>~� bv�УU����Y�!�[<u���'�Їoqd�w�K:|�!�䚙6Ἄ��S�	kt��"ę#�!��bBp�w��|��}��b�'�!�D�
��a$�5֌��W�W�!�D��m�D
�!���9jR�$�!�D����c��j`��;�/9ao!�d�,�Z]���6lMa�U�xe!���:t}�qe��"g��V���YT!�"f><����>c��d�8!�D'pBR�B�!ѡy��d�d$��/!��W]耻'j@�}j�Xs�!�C�c�i��Eɺg�<<�dT�8�!�d25<�����϶@�����-_9z�!�dZG�.�s#�N)&�N���f�@w!�d�s%:����� -( b�d�!�M�h�<{�ڃE!XS�㟺F&!�D�	�d\	ө�'v��9a��n!���%l�܉B��:K�jA�CP3@W!��Dae+����)�ܔ�Ƌ�R!�I}��9���8 |�@.=:!�DUb�&�@�N��ba�ѹ�k!5�!�Ā ���F�g`���K��i!�D�'_d���k��� 3
MSL��d�3I
D2�������TJڦ�y��"Z6��I� �#{� ��^��y�Gۓu�t)�eE� V��y�Ղ�y��*XA2�"v�${�����@��yb����P����rdqpgH�y�nFlA����!h��"ñ�y�K�&/�%Q`	��ZA�8�e��y�˚�qu�0��+ټQ�f��">�y��N��8�N�2�� �ς�y�6�΍���	�=x4S�_��y�D��j�d��V��0���z��3�yB[!
X|�Ȕ� ;�nubf�I�y
� �ڵ��3����`���jf"O�����c����3x��"ORu�Ђ���l�㍋���B�"OpY�'�
��taȃbM�T=�U �"O&��1]�
�����X�*��9�"O$e�I�5�PE�e�?_��<  "ON�Q�!;+^��Q�>ao���a�x��D2ҧ(�̝��Z|W.1:��޼w`���ȓ
�(5���ߋd��K�$��~�u��X�F�w��3 ,�)K��̭g��لȓ%�0ݺ�n��S3�Q�� \�=@p��J���%C��L��P�F�hޤ��z����y�Ft��6V���Hab��M�vN��@5/�d+�܄�Y��yr"$�;ލ�iw">��ȓC5l�Yt"D zɒ��
�6��t�'Yў"|�D��-h�h�b(خ;���J�o�K�<��	*z~��a�
�)5�t��fMD�<�rLà.�iA�HЄ{���!�h�x�<Q�a�
�p��� ���c3��u�<�G�U	A�fyS���"�X�/w�<���0� C!�Ը#8�DH�Gq�<��o�(#��)��;j�!�`ąm�<����2$d�CgE9
��Qk0m�@�<�C�st���A�ش�N����H�<���]�����+~�bxℍ�M�<�E�e���jR�������L�<�B!�2<��-q�g�f|HYcFD�<!��^��z<h�iխUp��&��|�<a�+H�D[r|0�D�&W�fp8v(�|�<R��9�
�8E'�!Pq����w�<16Z�z�x0M}�\�!PJx�<Y��E�(��C��0��z�M_H�<�1���AE�@I��*�`�E�<���Q["q�'��"P�z�Y���k�<��I\�	��L#�H�=�ڭ�A�`�<I$+Y�N�԰X"���f|��i�__�<ɁA^��"�)�@M���@g`�U�<�!��3�9x〒+e��9��LL[�<���]O�Y�1�G(¡�׬�O�<����>�&a1���Q�P	��l�L�<A1XI1f� J �����1b�<Abn¾:m|�+DfV<LV�YTb	V�<A�A҅/��R��դl_B	8$��R�<�q�S�1Î�2HP����QN�<	e�ш&:�X3o� -�Ll���H�<)�Ր[,��1���3B�� #G`�<1b��oT��"6D�@5�E'FD�<��E"A�� ��.	��
��&�g�<�u��Yau�ƪ��7�0D���`�<)��;72��`v钲⪨�t�d�<ɑ�۱,�MpeB��>pk��O_�<� �� x_@�I�)� \T��CH[�<���'6P# C�
b�q�C|�<�eC�+Ix����H����x�eGy�<�5�K�Y�0`�#�@��S�*]w�<9@ۍ����nK3�R�KG]�<I��)�.%�HM+	�L�Ӆ�R�<�d
��|xWc�O$��U��Q�<�T�u�q���	=���k��x�<!V��8k$N�"�cA�j/u��@Is�<�!ǋU�6d�T�G29\|�`�r�<a%��/X�s�ĕ{n�u��H�U�<)����\$݂G��]�å�W�<� Nd�1�ްfG:���B`x2"O 8r�D���6�U�L�(V"OL��bEV��Ԝ��	_Z��!j�"O�����!Z���Y�I��Tv�mY"O���G�E�\��s�"��Ow�H@"O(�9%o�5>�9+��Y�Z�c$"O��I���H�&-8�/=lP��"OP)sR�G�ʽ��M�5J�@��'1�h#S�G�3�.��&12)� ��'Y�Ha�U�f�Ԅ�GC�/w
 ��'#�)�$A'9| ��� ���S�'�&aP�J�Mv � nV������'L���&㉊F}��������p;�'��!2Ѭ��@���SE@C�_��Z�'(P����&�6�JՅR�/0�0)	�'�A�S!]?ul�3���)�t��'�
0��Im�`=8$�Z�(�0Y�'1�T�g�C�=l��i���nf$ix�'����.U�#��u"r� lބ���'�fq�`κ	�h!��L؇w�}
�''��`⑄	PT1�%ŶW�t�X�'���$�U�w�^ȣG끠:�Z���'X��J5W�?��P�A�ͧ9� ��
�'����N�(��L�Ə� -�Zy�	�'Y/}��3`���wl�)hLD�<iЫY��US6�܊9d����EDA�<	��4�d�4,��"��EM�@�<�bL2��!CF˛���Y��f }�<It��@�V�c I��ŒQ��c�Q�<��"E�u(����X6P1X��Q�<���-����
=7�! ���r�<YQ��*U2��Q��:H].10d�<qBB�z�����L�D���&�b�<C����� ė�(�����[�<��L�/a1f=�!�I�|�H�r'DB�<�Bn�~��P��23.*�)�dh�<���U!
�������X��!�Ȗy�<yCB ^�������PAIV&y�<Ys��>L�&�3$'�q߆Q:�`�<�"�Y)t]F
[!N�d�W�<!@���tj()4�ʀ g��ihFL�<�GIo#��[�޵B��1�I�<��K�(:�SÁ�9E�A�<C�I a��E����#̀0-?߰C�� 3�T�@��!z�Yh��VB��C�I�7��	TN_�j����w��&�C�=j�ԸRi�/|F��r&V�e��B�U�X��E�� �9��C�I�#Դ� EE�|�l��C�'zC䉆B�B��f
>s��g V�>�dC䉥wO�y�@V"|ժ`��^2A'C�I*~l�
"/کH�|���)Q;��B�	[Њu�sKN;'J�RhΆ
�ZC�ɾW��*P�@�AZ�$ZA(� 9�8C�I&d2J1r� �f���ȡe�ZC�Irwh�cDAfT����)Z>�B� *��a�i�H���*5�'k�B�I&IE���5�6��x�5j<}ަC�IaS�P;"c=�����iU�FC��.~C4ؓ��E�utLCAɍ�,C�ɶ4�nqS�
^6��@᧙C�@C�	�����3H�LvI�4�b�ZB�5dV�0:�'^�iBn�
v휼+�B��2X1S`O�gr��8�گ)ӆB�)� hM��$��hs�8��闄��);�"O��XW�Y�B�. ���Yƞ��b"O~##�B�:�01�����*�v�`�"O��i���*x.�\��
ئMX���"O6��3Jߛ"D�U�˙m#��e"O�U��cȯW~��ڕ� 5�(��"O`�;*������+}����&"O��c4�,��袗	�^��=�"O�Y!%U�6�&�s�mw[.��"O����㉼!�0ၷ�I$GQ�y�A"OQ��*P��ų�M�{L�a��"O�i�O�.n�e��6=;.t÷"O��;�"�
k�tz�H�	7*|��"O0���ʚ)��q��+ʛA1~DX�"O���#��RA"l�rK� 9��c�"O"��&�L�Tא��S���~�K�"O
�2�팣n&�!� /��#}�A�C"O�%��#Pz���,L�G����"O��80�ޝD�Rr�,EQ%�D"O
����,U�8%����2,y�"O�$	�G���H\���U-(��)"Ox�XRa��7��AG4_���"O�2���}b\ ���C�z�S�"ObI*0�V�~A�u*�+�(J
#Q"OF�(��ڎ�P��l�7|*���T"O��A��}i~�I��C�2+ؘ�"OΡs�o�9
9��A�	�$k��(*O�I�@�/|���oلH����'2��QC��&v��p�3#X;@�&!2�'c��%d��k��R-��0$h8�'�v {e�3�ѻ�j� #�HE�'������̸]
��)�CUz��'>�z�K��D�܉2e��
�`�'���Ld��(�lW�\�s�'��%�KLi��<}��8��'K���&>j?���UnT�n�]�
�'�bT��/��.8�!EbCrx�
�'h^�%�	x������W��
�'��됩�+�>�[Ď�z�����'ɞ���k�=�,����n�^�[�'Ԝkj
Rl�����c�ʼ��'��X2iH
=-V��$�[�*S`I�'��Q�@O���Q�D�'_�dK�'��C슞[��s��W�s�,I��';9s��Q^=�3CRl�@��'7n�te�.c��+��n��DJ�'��4�!M�32�R�cc	�b��'���kr�����,Tǜ��&����&�H�B�d ֮qQu��aj��P�^28L,d`�%S�2�b���q�:��f	�̰��6'Y�E��l����<�炍&]mBM���3a8q��	�M*���xT҅�@��J����A���FF4�̐����I�u�ȓ�2��a��o�1��đW�r���\�8���N��e^���ؔ1EXԆȓIc���cb�D^!�P(�amJ���,.��	�I٭b��q�H؉5�dM��P�B|`Vh��y��=�
R��`�ȓ�iQ��W��15k ue� �ȓ�<I� Z ,���k7��
R�D�ȓt��)� � %{da�";Mj�ńȓ{�~�Ö�FsY0�@O�4���ȓ,��Y�.P!x��%"�3T�ND��S�? B���̌.F�HIDJڈ1�8��"O<���+TJh�5�0��"O���g�ǾV�Z)� f�w߲["OX�hG��m���E�S6;ն��`"O�H�
�$WR���I
��� c"O����ꆃ*V�}q@S#Ј��@"O(;�B&`�|C����rщ	�'�j���gO4r�Zy��b�<DBzY��'T��`�d���k���O�npx�'��$�J��p�@�ő�trj �	�'�����L<����Y�X���Y�'2���Rl�.f:b�Pb
D�;"�(�'��$�'�,FIY2�(ܿe���'��m���؆R2n�pP� c�"��'�`\B��-@�p�B��䢘8�'����W�3n�T�c'������'�T�S� I/s������C���P��'�);��˄,�������N4��'�Ӣ�l����J\���,x�']���c�K#mDR���@K��)�'�(x`,�	,�`�e���z��2
�'�`��2�N�:�F�8��Q�"6B��
�'��h�Eγ�`9���!�|�x
�'.��yw�χ.@���ň��	�'�\)�7���&�
�
�`�>e�	�'�H�xf�P�d��s�T;/�����'�X#ɇ?$� �R#I˔-oh��
�'�����G~	�'�˭W#De�
�'5��U�&͖���4P0��'�����䉀I��Q��JB��(�'��u�*�N�])�W���'%��1w�'Q�,�㠆�V�l���'XV��W�	��q�2�	�f`>��'���Y5$�8�%��L!W�����'7.�;w�Ɇ�*yʱh�� ����'�<�0E�������p욨#>A�
�'kh$*�G����%L�z��:	�'���ņ̀�p�GH�`����'3�|���F�@�YQ�RA8���'��K��N� �����5d� �'���3�dK����Z�CҮW#�1K�'�D�3���`?ڝJ���.Q��|��'	�H�(��(zlkp�;w�~�*�'N���BҚ!`�� 0���|=�'�Je��l�.�9�E��@��p�'
���뀞Tw�L w"͎*c��p�'Ѽe�����G�|=H�IKx	��'�&y:�/�)���g��x�؁�'��M�MA�̩� ��&T8��'<Ԑ�ҁ� ��!2
M�'q��'�TrE7�b-"ď����'z�M�E0v� �����7D��#�'sl�#��1�� B#-����'ǀ4�W���L��^,<��1"�'�ԅ3���$),��`R��>����	�'�� &�M�H���J�a>0���'����I�'JR)R6� ��:�y�DǋTi�)��T76�A��W��y�h �_�z�{���U�ސ�����y���s�0@�ON/0m*1IU?�y%Վf�j�t�D�Ӓx����yR"0�r��a3�V��AǴ�y�2A�*��dN�<} dp��K+�y�f�5-@�(cW�m�� a	��y
� Эr���:*
:#�C��`zU"O&�:r��R�6���H9@ H7"O��T��oӬ��.�u#|݋�"O�a�oR<� �R�>I��"O�U��aU9{[�a�R�G$���"O�Y�%	ƚ`���R%nÌHJl���"OR�%Ɛ�PasG�/P�}`"O�	�ݍ;��$��E֟=��u��"O�#�ɐ�j*e��˙$�Nl��"O�Հ��
|�HČ�_���z�"O�Yȇ�B�Oú�ц�4J��0iR"O���.e�$ث ��5�8�X"O�XJbfT��#�!�9~�0	�"O�$E�>v��SK�.y21˃"Of�J��Mk��rr��hz�A��"O:�zd�7�܁di�fa���"O2�2�!�#�FH��
<oL�9`�"O������o�(Ayd�K92D�9z�"OKϣ?F�3	Y��%q"��yr�D3o>y���\s��£�D��y�T�-��pi2A�$VQDMB�kF��yB�U)�pm2�J	�>(�����y�E K�x@)���9�<��]��y2�Ü�:�{�c��p�!��4�y�ZEC\��B�%���bQ)�y��ï{XE�B*�v��J����y�j.:�༺Pj ~�p[,T�y�j\�C&�Ã�]�P��A��y��r�\�D&~�*���eF�y���D�&��R$�^}p ӭ�y�l�e�� X�X�~���JЁߛ�y2��Z^e1deD�#� Hj'�T��y�NZ�C͞<�QEN�\F�1����yBdڝ��3T+���9#]��y�Ŭ'���`���u2���!��yB@Ȯ-�(:)�u��Hn2�y���m��Ir��]mEB`��C���yR@'��QALP8l��4!&�_��y���&�8��d��wV��e�
?�yN
�[�h]2�Df�0$�@�y2cN��tm-(�&U�6�J�ybm�N��HI�Ź7�Ľ�b�,�y2$Af�<�R���>p&�i����yro@M���'ئ� �0�A��y��Ė ���1��'a*=��<�\��0
�B����MH�OA��]0��q���/J(�BO�ȹ�ȓMhM�رM���b�
��ȓp>X�ʗ�)"8�	���
J�@��S%"�2L�E�蹣W�� W� �� ��dʃT��yD�ܽ�>d��U�fq{�ŀ0 �~���Á0ׂ���]b�T�*V(��c��o$��ȓ60�h́^Dȼ��0k�хȓk_�1��C�5V�Ո͑?H<�ȓpu
�� ��[�tLaW�P�dK���G� h�qD@�`ˆ`�i᪒��y����45��z�*�@�d�Iq���yrAD9��Yb�oI�4� ��bH��yF��h\���V�
	�U����y�B���Y��ɾ9�dQ��,�y��W�� p��:3Z��{3d̶�yreF8%>J�	�Ȁ70�$C�O�y�KR~��e�m҉,k�ًu@�y
� ~� � �x@00�T�V�`щ�"O�ͺ@�Fy� ��Y�<�He"OrEf�3m���%)Vn���"O����ڬhh�1��5W���R"O^A҇i�J�T̀1т/:��2�"O�8�Ï�(FK�[�T𛡎[�yRF��Lq0�%A۠p����-"�y�DS�x�L(�_��UXa#��T��^���`��ʬx��Ѣ2�U:|�^C�I�g:$�H%���;� ��qI\</|B�I�N�tBg&��\���g�4\�C�ɦ���B��~��h��A�F�ZC�Ih�������ywv��S,�pC�I�0�6�"�얰n�2�DBQ�LNJC�	�y�\A2��%9 d���7{>>C�	K'�rF$�P*�W7n�C�$whN81�06������?�C�w&d� B�����)%)�C�13F� Y�";���1�4;bC�I�(�D���hV'TqcV��3�NC�I���c�lİ:HIz�&ˍ�0C�ɍJ5L�a2DC2I�R��aH�cpC�ɤ ���y�Mĳ+�����+YHB�.I#�k�Ǉ�=p���Rl�6(�C�I6Y��u�D#��58��^�%�C�
�&}i��-C�py���&�B�ɹ�̝"����,B�N�+�^C䉚6�PEB�NE(M�Tq�`�[dlB�I0����f儋�X�%��B�����'��%S;�U�cY?
�|B�2|�y��M��e�`�&k:�B�	�iFd��	�T������
�bB�	g@M�v��74&!KU+��T�B�I<h�V�2�$�"F�
Cd��:s�B�	 ���	�m�n�4I��#D�B�ɧO�6��5cٔl��-�S��i�B�ɰ0�|	+S ��$�Z�	�i�83lB�	'�J�O�-[�&]�wC@0q� C�	�h�fY��. c��C���:�B�I�w�X��LU�H���o^$? DC�Iu���L��y�(#sl�mC�IMi4;P�>�
�r�/'!C�Id����N� P[��*���61� C�	�p-�a�D^�ͺPB�z��B䉔{�@! ץ|6V�x��[�H;�B�I�M��P��$9�@�%$i�tB䉴+�@�FA�:HX�e��z�B�I~.>�u��)#?2�+ө��@��B�	"%��ppNF�I�D�36�"|ovB��9���3�
��p��`ŏ��cWjB�I�,�J�8B�R.#�@���>�C�	 f�(Ð�DHz 1��҄Lu�C�7=\.�0%O�4E�j:G*N<3�C�	%h�ꌓe���bDB����m�D"O�B�')K���2���1D� ��c"On�2�JF*}�H�s`ڍ1{R�J�"O�Sb��/��]��O��-n�5��"O�D�r�α2�� ��6�1��"OPe�!Z</��4��Ѳm x��"O�d�Em^�\E�w� X`��"O���Ş=Li8�qǊ�3�0��"O�̩��F�(�4�tI�Q	R"O(,a�>.���Tn����"O كD$йO�h�q3-ɀY����@"O� ���G�U�́�"تK?�pp�"O�U�@A�<:��aX�B�,a�2"O&�DC��K�f�@�۾j�
|�6"OR��&��B��Ba]�4�H�`"Ox)��A���f����]� ��E"O�]�&o[�@K~D����0�
��"O���!��:� � פ��=w^��"Oz��Ќ_�"Y����_��|���"O���Kڰ$���V�c��rt"O2T��� &��iH��ѓN���#q"O�|R��H?/:0�qC Ӭ�B� �"O�P���SSLct�#�h�pq"O�HA%��8w�8$SO�3�謑�"O��
�8�.�2#L�&��r"Oh�│ȔU�	������Y�a"O�ԉb��?�iB��3?�X��w"O�}3sC�^P<
b��b�Hm"O�� �&��`,z�3ĥ� c�z�	""Oz\�D*M�g��1���c��I��"O>;��9?1���F�5a�	q�"Ox̪2K̲C�ћ5��k�P27"O
�"@s*�3��	-RB�PD"O:|���؊ZЪP�����Y<�!C�"O�sr��G�,��ԫ��n.F�s"Ob���jٳX�J��
Y./�^�Yt"O��&�E��}��N-����"Ob�[T�׉pH�@B'5\���"O�HX�B�)fu����>8I���"O��QIإtFJ�YEd	1nH2��S"O��bw�[#C�(��cC.n>�	��"O�����	2\`�2wB�2�!+�"O��*g�ı��B���1{Dh�1"Oh�yF@�(ZgT��V��4,d��b"OR�q`�N�WW��왷n���*�"OѪ�ċS���`�j��	 ��#"O.�`t��>e:��#�H�rK~Z�"O,ai�[�%ќ5c�(��OBP� P"O*��S#�(vQ�1`�F��H�Dd"O�#��.WX|@P'W� n�|�"O����L�N�$)b��רAL�8�W"O���1��8F<P�P��v8�"OPȒ��_5d��Q6�ȗR�j�1�"O���e�(|��E���v	x�"O��1A�֢_~ )s��>↔Z�"Oɪ��/95х!&P:f��q"O�aQ��0�f<�A0"0<��"OT�t�ݖT��M[D��#y@+e"O�H�k�� BJ0to�.^<�2"OP�,]'cM@-�W��><�4X�"O�����HEac�G����"O�p96 
���5�vOA2'ĸ)�4"OtHj�D]�Vts�$��Z��l[�"Oj�(6L�� �t\����	����`"O���Dl_jC^�Q�S ~��"OT��AB�:�2 Y4�
���{G"O�y8�5�lr�L@-*SL�@"O�i���)����g��(d����'"O����M��T
	@B�R	���Pp"O."�|?�T��J��)�H1�"OX���dP����
x��!�"O��X%�ӫe3����	�C�.D��"Oh钔&�(14b����b���5"Oh��_�S����
�S�b��T"O�AX�	:)�%�g� �A�w"O� ��S��שJҾujp�"�҈;�"OB��q�U�!g�yy���;1��8�"Oh�J_�@T�ˠ�D%H2Z��"O�ɀ.J�˂���1
1l��"Ox �E��-�pR� �G}u�`"O|̳�ߍm:<)��$��3�Mڇ"O�1I�`�0j�2H�㒍[T�V"O.���
����s�D�n0v�3"O\�,-����y�VɃ���.J�!�D`)�X��Ϟp�$�e�W%!�J�oϚ��e�@-Ђe� �ƫ/!��|��i���ɓM��P�e�C{&!򄔶k�x)��M�yVX��a]�=!�D��\m�c���"$��X����#!�_�X���Ƚ�,�2!	� !�z/Đ�� ��\�J�˧'I&V�!�$˔k� ��2��?���4G�+~�!�F�$�%C�&�R)���pOS!!�_���׉̅o�bI��G�8�!��Md��a��e�a�"瓭6o!���\�ntad��9lϺ�Dγ^P!�d��~E��l(��b���F7!��7����mH�by�@�J!��NrfF29rDDH��"I.!�D�Zg8��-p�J6��/9!򤀧7�=:������
L1".!�$ʕS#fy�2,�-�:��Ǌ�P!�.0V� &��*����H�1|R!�dª7�`� ��-����b��3!��N&o��m�����e������N�!!�DǴ��0���5VA�V0z!�䑌w8�ɛ�*�e=�xjf��3`!�T'"��m�M�&p5�
1|!�J)��$q�����S��'g!�d�Puƙ�$,I���Lc��]4Lm!�5���S(�?w����s��2@:!�D	�jQ�|��1���+�J�D,!��#u<���A�
I�,�����%!�d߳3�b�(C�Użiȃn��N!�D���R��Jҙ��E��-�X!�D��v!|$����f��H���3�!��J7���x��1#�L9�u�R�aE!�Xg�!��C�6%�H5�K�=!�dZ�nvTr�յ}���(e��"&!��g}B�)5�^���[��)g!�$X6y��y8��}�Q����<*!�M�/ּ��&W�� %��
	3p!��JM��r�I�38�AZ��Z�PyB$_J4H�(�2E�Cb��y��Cԁ��Ί!r�� %�?�y��[)V���)��)r�`(G�#�y�c��5�}��'T�	 ������y�K_�BA�C���T���ܠ�yb��!*�$�%�]G~�&ȓ�y"�Y*J���!�r2T���W�y�"�0X4tR�F=P��A5%��yR"D�gI|:��N+<X#"��y��C���h�b�DDp0i2B�/�yB"E�*,�AkvGQ 6GT��D�U��y"��V�V�2 o��%tNt��cU��y�j�3N�~x`1$J��|X�6�4�y$__�̭;g�P/&Y�e�V��y"�O�q��:�`_	M��je��yr�B�SH�g�B#{�	�1G��y
� ҄��B�QH�Is A�<
`)!"O�(#chM�j
��R0�]�4"O�uZ�Nǂ]���Ǒ�ĭ@!"O���!�G�=��f"5�l&�'D�$A�%M�|Z#A�0G���3�8D��օ�rvh��A8�=5
7D��b䭀���6�S�Q���!5D��*B�R2v�v�[p	ӸYRݫ�1D�<`⃚�#���G�ҞR�v�+#D���`���/����T'�Z]~����?D����7��0X���[@ ySd8D����<r��|�L0B�vf7D��q��:5�����ޘ%� Jqa1D����g��\�4PG�9S��$�Q�0D�ʦ1E�xp��`ٯd�D�A�:D�����%?�Bp���Տfk�˱�2D����������F=��J��=D�hk��Z:�%u���0��e+)D�d��FU=�������zU#I%D����ʓ0�F@H���|b�"D��*���.�(9�KȌ*���!D��&(�O�VQy�E0�����=D��@4
�
a�}jÍ�p,�5�(D�0;B�UD
�arF�d
<P�W�'D�<jD	@�R�n�S� �	�Tt�!�$D�2�,\�x���(�/ϩ	�n\��+$D�����E��1�$��<�6��#"D�01B�#3Aj$�^
T��qpC�=D��f�(=`�"�Ѹ6е���;D�heG�TNz9����<OΉ��'D��� �Wɒw��4G[(�y�N��^!��ZE�� !Q��ǵ&�!�$�0���ba^J�Vx� l�y�!�ڀ#�	���s���Ka+��_z!��_��~ȁ�J����Y��B�^�!�ۣS,�e!7�
�M�.]�aN��!�d��f�PnS#e�>��q���?w!�ҡ�^%���X0;�Z�au!�$q�L�˓
�]&�a[�Y�!�
���U�Cؚ��F�!��&k�,�"���\UP��S,�!�E;%����ǂ+6���� Q�-�!�d�6X�0�p7a>��W�!�R�G�eZG£q����b(޾c�!�θWWP�bU�( �,�0�\�!���<N���b�E,3���څ���!�d	����B](�c�я]:!�$�<��}�Pd�PgN�8��l�!�DH�V�uo�:[Hu��1�!���IR�j���N��'b�)�!�}t$�)��8�A�&L�!�ќ2�D�ҪѰz��Qk�&֌�!�D�3$b���#�Ĕ'�����+I�?!�Ši2<Xoͨg�5y�o �Vr!��b���qK����Za��4�!�$G+���c��"|w�h��K�%�!��T�Aj�L�#�Z���	Ԣ[�!��Ċ<�zHc#�ɒ8Y�pc��Z=:�!��>7�p�UP�MC>�;p��m�!�P	g0ؔM�8@�-�/ �.E�� �2Q0�"5Z��lh$k��qh����8�<��c�#^�^��q���Z�l��`�>�j�➐lc��Zcm^�sl�9�ȓ�����.H��� ��o�z��S�? ���j�X�4[��i�tay�"OpI�1�I�,]�%�B��5+ ꠐ�"Oʕ�C�?4�J�rs@_���0i�"OΡ	���x\@9���7�!:�"OX�Ӊޞ1'zx����Y�a:"O888+ٸJ��+Ў���"l�"Ot@����f��Nњ6��P"O�ܲp#�4#R^L+ƛP���"O"9����i.���cMd�h���"OZY07S�OuN\�&��	���aF"Odx9�ɩC�t�qR���\�X�3�"O�]������Ce	U�v�$q�"O�͓�)��/����S�`��KG"O 1����ma��b#'�9�"O��Z�m�2�8M��@�"�1`G"O�E�1��?t�$��,-=���"O�u�%�C�Х�̍X�%�c"Oƙ+�'g�x́I���˳"On�8�h@�~�ܭ
�a������"Ov=���<
������Y�20Ӑ"Of4𖯚�6ٮ���_���e�g"Od�@#�?��!�f�u����"Ox��o�o����fN�Y>̩��"O�a�6��&�.�a�儢�R���"O�Ye�ȵ`gz� �D	%VÀU��"OBTP���/S���FN%{J����"O�8��]�W��@�$�5L�(b"O��0��öV�X0��X�~u(�"Ov H&hP��Y��J6	��"Ol��š���캓.�*f@�Zf"O�hZWC��晣���&T��i�"OLt�/��|��-�k�,e6���f"O*���L	�/e���)��l�h!��"O�=�f�\�����P2JVRL�"O^��F��+4�B�'V�k��9��"ON�3��n���We�. w�pt"O~� ���aǐ���$A�}t�$r�"Ol�C"�478������0f"���"O&-�5�_�D5���KK��#"OH�{�P��Ɂ��v4ƵQ#"O,�p�ʁd�8�0�ޯ`��cc"O�|i$�8�l���U� �HR"O>���'o0�D2���7v�!�c"O 4k�
b�.���L�xqpeI�"O�P�%iŔ4�V�R*�F�@D�@"O���5�=�u)B�b}J��6"O�9���-e����*ʤ:`
	`�"OP�#�Q;$U|��c^,H����"O*Xh�m�:�;֌�0$ ��"O %��B�"�(�l��Vl5��"O�TZd@	�(d ��3JE�
Eh��"O>1i�o�=�$��HLHS��"O�0b�Ejq�|c��OL�=�"O�d�u,̤"ߦ@[t!D�<z���"O�8�B#�$��,P��Fզ5�@"O.!2�)��(t�� b�,��f"Oj|��E�\/T`ʑHW�m��u��"O���E ��z��ţ���#Y(Np@"O���`@�e���'�6S%V���"O��� 00:�"�%L*tAr(�"O&��ǰ�V� e�> ݰ�:4"O&1�����jw�<V�9�0h�"Oj�·D��B*��x VQ�(��`!�D� h�Ƚx��9\������G!�� =�Fǟ�d��!3퐶r]��	5"O䅱�^��@4"W��&~=����"O~�z��n[����hA>����A"O8+1oː|��!��g�7.�E�t"O4��D�z��p��G='��:�"O84�dÕ)%�4�k��4g��}�"O�<�ŀ��H�Q Y/t�J�3"O�x ���%�>}Y��
�uGB�V"OF�iI--E��@�,�<.����"O$�x�����ӕlR�OP��v"OLa��A-��p���  �~�{�"O8�U$�d��1�ꔖN�8`�f"O��r�)v\!;`����H�"O$����=�F|�Տ�5�9��"OL����ޢ �FY0!m��4��;"OD��$����:N�����"Oĕ�3�F�\OxA3�퓛k ��G"OD��1�(
�n X�̍�]��3�"O����>	� ��*�r46y�C"Oڹ�(�J��� �N=L,8��"O��3s� 0,���ES	3	��Z�"OD!qb��1DR]�W�̂��Y��"O��H����ƌC��W�بѤ"O<����'D��3�%
 6x2"O��PI'@���ã@�,(��"c"O0ˠ�"(�����_����"O�yy4��_�
@�2і�Av"O̽)H��e���@�V�"v"OXa&�%C��� ����d"�"Ou���[�>�*�ȶMD�Zlh`"S"O��HQE.z�Q�&m�zو�"O�P�� ���@��J�<��P��"O"�K�+#�����)��0�#V"O,���٣�ޘ����g��	X"Ox�Ad�;�zU@R�J�l̄��e"O��G�5OZ����/e��DXf"O,�BCD���b��H�,�(�"O(a��*��l$hBgRc�<��#"O\�'FC�cWĀ�0f1�T1S1"O"\ء�_B���0�_�<�c!"O69x�$H�i�� 1kȇLnr�"O ��M�0h�n�˒�խuj,�B�"O��U�O�(0a��'A\��u"O�,�Q�۵c)��B�? 1�"O�@�1�)wd�q�Az+pqK�"O���b�ƑP0f��p��3p�-A�"Or	��G�`������vUX��T"OX��#���f�h�I3L�9T Ԓ�"O������u�2�I'
��/@�s7"O>�����}^T�/� ����"O��顄�,=<3��E>J�xP�"O�X�AF̼+ bp��LRll�1z "O��³.��C4�M����\0�0˖"O�xc�d9���`A�_"�4��"OZ-Kcˇ��}��o��v�$�"�"O8 �v�U%�.�#�g��
���a�"Ojl����� �EsKܦ�R"Ot���
��:ָ����k��A1E"O$Y{���0�Ҵ��&��#�2��A"O�x	��	,�t!�! @&_��I3w"O�:ղ�q�T�^�NQ�(��!��p�`I�K*e�È�4!�D�`��=�I�$&�b��T�m�!�D�{��q!�(Y��!��@��!�� ��QT�Y�d�\A�Bj-iR��R�"O���%� ;:3���:Y"�9��"OaC�Y��
e� �^�{j�jR"O�Y�/�4��T���$Z5T�:�"O��$�$I�qh&.��f�U�T"O�
��Ŕ(��y�O�#,ty�"O<Y2I�C�`y+&�ݕ^?^!p&"O������|�p�I����^$�L��"O �!D��9O�Q�t�NAV�B�"O�D�M�#y�]D#H�"'d�"O�p�fm��1������8"`	��"O�yG�=w5���1F�,M6�!"O������@c2w��9*��%"O����Ï;A�j��ȼGbf��R"O�-�Iݧ3@ԕx�
^�;z�q�"O�������Nn,Zլ�;xGH���"O�<�pmJ1LXX`b��.*�]�2"O`i@���p��5Jp�X���"O�|'*Q_?p�ˁoA��[�"O��)JEP>�X����@��1"O�Z���)V��r°!9�s"O����¨�,Z��̗1�� "OvP�Ad� |�� �g����r"OJt�q/
0r-w�1y]�� 3"O]{$�M��Xtc'M�!YipeP�"O�<�ę�L��BK��),L� "O��Bm��t�����?X���ycT*r��5IR�ЇJ�d�0�	�yR)Pr�-�堑�5�x�sׂ�yrBL)׈��g�����mݩ�y�A<J���ŧ�!�`	X�ߍ�yr(N�s�i�q���5f@�dŒ:�y�`� �b�Iǭ 0\�seA�1�y��@=8�4y���l;�u�d���yh	�m��'�(:f��RÉ	��y!�y����+WX,Ks!��y�.2q�8T�킸x�����E��yb��!����S�`$t�Z#F��y���vs�h��j�
aBX�Z�g��yrǞ�M"\��c�Ľ_W�}k"+��yb�܍*r��ը +3�3����y�aQ�I�[��G�/���f��y2�!PHNjg�].�o˸�y��9*Vas �ͩN��usPD�y��J�N�#�	.T�J슧�ü�y"H�} �%����$GB�A�ņ���y�*�;�Ƒ:�C
5V$dI����y�/ �p�f&#�"i�t�ɥ�y�(˫Gn4�[C靧�4�+�/�y��X(FN����9?���Q%�y2�F�2���P $\�@Q0�����yrf˫N�X@�*�<~A��@��y�\�_x���X,F�8K�m�"�yR*J����@"(�@YC��_��yBe�j!ɇ	ÛK(*�q�G���y�'E�-hT���o�L4� R5�R��y2D�Fl�P�ު�`5A��E��y���
n��%��b����4���y2�T�G���ǉYl���S� �ybF�,��K�藖V%��S�Q�y��
_:�p�Ć ���9�& V�y�GȦz�Y�v��r|M;�kO��yª���Z��8`J�4&���y�悉i�F<����;5����e��y
� >d���Ȝj�HEG��q��c"OZ�IEfV*}�^�BF���u�P�"O� ��0j�.��e��u�"O���̘��j��5��/
�"O$��1��&k����ODS�H�R"O��[�ˎx``)<|�"O"���Rk6r	3 � �|�3%"OjT�`&L\�<����0��aG"O-���ܵ��]Ѷ�A�s�`T�"O�L�oެRl��s�R�Q�$��c"O�� �!^ ����'ОnTѺ�"O�d;� �S�h GΙ:_��y�"O.� f��t̬e贃���y1�"O|�w��,),\z!�J# ��$"O
�q׉�R�����J�BИ�"O�hæފm�8�qH�f���S"OR| Q=(v��Xc�	ڣ"OȔ1��C�@��͚�){��T�"O�ѐ�͞�\���6)_%[�̻#"O�$�%�D����-ݏa��=p�"O�=)g�O)i>,Њ�K^]ot�Q"O�	���R#:�<�����2J6�b"O���PÑ>�9��R�(<���"O������**��$;��?<1@a��"O��t� �K��@	�2*@��!"O�c�eS�$�~��?U,@�S�"OrzW��blt=af�Cm(@�96"O�ł�������<( uP�"Oބ
qS�|�	��O�}kV��q"OԨ+��.?&���BKV�X��"O�TEAܫ8��l1)�"\p���"O��xeB� ��
�2R���"O��9&�њx*�pgjZ
qpN��"O��#��?s耤kwI�"a���a�"OĄ�uAE��t�a�Ŋ�O���W"O�}�K��(4�%F(�"O���dca]���T�
�*�r�"Ol���$�2pze;���L,B��`"O ���]a��SU��2�(��'v�|CƏܑZ��Y�q�rJ��L�<AG�¥s�L+яN	���3�H�<q��Ű(��4��F�����z�τD�<�4d�%��<�a�	(�X"��J�<)�dQ
 f#�I�*D�"���LAE�<�-ͻW�敲S�W*@gr}*HA�<�R��<?jl�:�&��b��j�\|�<a"`� z�"��'�»q3�R��E|�<�3���������E�Nx��M�<�n�7`P5ඡi��}��ȗM�<A��5y*1z��L>K��C��\F�<Y�G�yq�cDM8�08��K�<i��p�X�q���*kyJ�x��Q�<���
����@�JqS�m`w+�P�<a2�O).6f�B4`�;D�(0p@�K�<���ٮ&��u��(�5B�H�<i�
;Y0�(��ǟ�V
v�hVLDl�<�b�� A����q'���s"Hh�<�!L��RC>|�-+֦ԢS��g�<a���(=��
�bG���	��e�L�<�!����јF_������)D��T�R�V�ne��%�0�.�i�J;D��*��ѩ-,��e��{T8����9D��"�!�ݻw�¬+�H5Pdl7D�8����z�!��TgLt���6D�� �$v�ިQrzP �i��'Bp�P1"O&8ۇI@�~9��b�_���"OFE�3D9 �����_� �=(g"O�������ܰ��\M�\��"O�0Q�&#Q>͘e�A�t���s"O��Pk�6�D��Y�y�&"O����gW��L��m.N�@��"O�$�Iu�D-�G�S�4����"O��׌ǐO���z�d�(z�Ȁ8U"O|�yw��0�jvBۣ;&F�"O�$���;c!���f�J�r"ؙ�"O,�;��	�B�����!*."��V"O�UA�%�!J7 ��b�ۚEa"O ��׍EW��I��	�;���D"O$%I�(�	�V0��T�~���w"O�8�e���$8(d�E�SD"�q�"ON�8��R̒��]�Zv�a�A�W��y2던9{�xPC�C|h1	
��y��	'L�B�b�DY�>s��s �Y��y���h}�d�Z�7���Ԡ��y���B}4L)4�=/��� ���	�y�I�� �0	��l��:��g���y�U��Q��*���ï\!�y��-~:�؅�FS�e �&͠�y�#bz4��bJ�GS|��a'�yB)!b!�T�^8J�}�G+A��y2/��V��tD�4>p0��bۅ�y�A�-	&@Q�#;4<b�VY�y���hfր�1$��Z�r�Ke	�3�y�jحZ�64:��NK��Xb$�$�y�A)sR�)��D (J�9�q%I-�y�o���a�g��jt��Yf"Ы�y�y���(�@������:�yeO�`Z�
�hֶ�25H�����y"��A��E�1�2-�%Q'
[��y"狪~�Ν'L߶0X�Pgث�y"�*�r)KOǒ#���[�)<�yRo�8^K�{E-Ϡ�����@��y���K5"�B��Y �QSL_��yr�Z�%��!I`I�8���BD���yB�P�TґB�O� :Rܲb��y"Z�g�\� �� �8��&�y���
 ���Y�Ȋ
A�x@`/̙�yB
���ś��ܧ�J �6�́�y��W�A�& /�=P�Q�����y�-��yn�5��a�<���Be@��y��Z
�����o+w�>��"��y�Ɋ�B�\�Kǂ�k�*�fo]��y���^*��t��,]��8�[��y"��#Z�����@�fè���]��yr'�<�f�Q��ܙ��G&1�y���&/��z��	(#��f
��y�"��G�0)wL��o��a�N��yBH�)lM�FB�x�"�Qa@���ybF����1�b܉td�����yr�Q9|DM���Z�r2��3Ce��yb�ّD6~��!SeX�=r��M��yR��q�,`T��2O�6��`_	�yr(���azEh uf�h�-��y2�L&g��!�g9i-����#�y"��f0��4 ۹[�&�/��yB�~�2�F�$�Ĩ�'����yr(�Q�`��Aj@�S�X�'K�2�y�֣'��K�k��9(�J�y
� *4w.5{L��&o���ɫ�"O�5��#ۭtv�����Q(հ��"OT���#M�Q,�T/]3�����"O�ˇo�)h2�#���J�J���"O�����2n��a�M�w:l�a�"O(����;�m��F�
&�1��"O�+)BH��BIנeg��b�"Ol���߇6�^0�2Cԫct��*�"O2A P��K�nQ���ޒPYpE�"O�E� KE�>N��ɣË!m�p�q"O:�QrF1}�4�� ĩJ�JHJu"Oyx�ǟz��id��$�y�F"Ol�a�� %Rܒ��E蒰6���8"O.�QtE1�٣��E�
t�`"O\#paB�yȼ����%��%�"O,�Z&�?��c�W���"O&�c�ņ��`@�LZ�f���"O���B�,u��8�� ��=��"O.��F�w�P� � �C�h�+�"O��@QHҧHr�AT 1��r�"O����
������O�{6���"O�EGB  wx�-\&|y�"OV� ǅŁW�v����{�TI��"O���g��-��5���]�"�`�"O$�"� �0���8�"oj}p"O��r���
@�5� �!0X�Dq�"O����)�D��+��Y�0�$"Oڐ��#�$��!�
" ݄+�"O�!�tI��J�ʡ�u@���z��"O"eٷ �aa��2�`ٓ�%b��y"�'�h J��݂���d�_��yr�1\|�U�ݡ{�x��K�yR"��Sߘa�v�z�b�(�>�xb�'��c�j]=O��x�"'�zP�'>���'P��zu�J��(��
�'j�����P�Y8�5��	ͬF]��
�'����˕]����7#v�&A�	�'#�q��-������F�R7q�h@�'�^{5��q���3�J>w�V9��'Z���F�2E�|���I�$uu �(�'Q���ԁV�E��YƌZ�Ü<@�'ORl�vAr���@� l����wn6D�p��+I���-Y�咳H���b�&D���	�$I� �s��&% ,�XPŅX�'����9O�4���,����*5Rk�<�'"O<�i����N���f�*q���t:O����ԝdx�K����d,#&���{r�$�)Yj�IsΒ:Q��Z��\#�
O^؛F�g*�QQ��+_�5���'�'pV��rP38>\��<�YC	!D��1aea�@�vW���G�$��C��)P�����ނdS�q���ޚh��C�	�L>fY+S�١A��Eh� �L��B䉀'���Ћ�7O� � TG1*G�B�I%/� <jW�2$=ƀ:Vo�6"�Z�	K��܉�o�,�F�X���5<l��W�"�O�O>!�o��a1Xd� �D�e�V���"O�ȣ��A79ȨE,�"]�&%���H��䓼?���Sm?�f_�QdL�C O@��ly�<�rGĒ��5t�\�?Ȑ�Ey�<��-W�=�B��Q���?�vu0�$�P�<bDJ�*eHP��D��̅��/v�<�bt�xe�"'RL\��k�<���6$�|��̝GH+w�d�<� �RG��v� EM�J�X��7"O��Pg(#'N�B�
fJ�L �"O����8~y�e%ɞ['L��0�� D{��)!{�����[�������r�xB�I)& ��g(�#TJMXT�[7f��C� ��[�)��r\ᡶ%Yg��B�I������O�0�т�n�v�Z�1Є(D�DB�i  O��K��`BX�!M(D�L�T)ݺNF�H +��=u$����2$��J'�&Gz���
zM@���y2��e@d1 Kx}z܋�����y���D�h( ���(�4]����y��N��"&��:^��h���'�ў����]�}��Ԡ��B�jR��"O�I3m�"Ev"d@�/$:^��X��d�<��4��1 �τ"sM���a�QPb}HG"Oz�	dgV*�䩗�_ 8c����>َ����*m����N�jg�aj���a�!�!,P��S��\�yb�]R���a�!��H�B=+�`����њB�a~�P���"nE� ��ɛ�,_�h��{�-#D�T�sgW5g�$��ҫj����d�LD{��	K�� ۥ	G.w���;���!�d-%0��GY
)��lC�d	���ɟ�HO�>y��L�5Z�>Q�/<JpȷJ><O�#<y\��P�k��A���ī^�-�PM'��#�l���+� �%0���O���q���h�INyR�B�KY� x� H�h0TD����w�<Q�#A�G� �sP�>8%"��*u�Iϟ��?��{�/B/7������7^7���L���y��Z���=�q��)f�R�s�Q��3�S�O��4R�m�,-�l$��^+&$�S� i�đ�X�2�"b�&<��aBCէ~�!�$L�O&F�3&T���bÐ	]�џF�.�8}�����MC�pC�Ў�>�yi��{Z �[�b��,�%�B�	�	|8�
WGWC~H1���B�	�fC�eh&�R A�jHQA惘-�B�I�yfj�����d��	H�-A�5�C�T@\;�M�(1������C�	w�"�q���w��eQ�ü#,FC��-�&,�r����;�Èr@C�Iv	(i�#��0ZA�A�o��N�C�I�0lZ '��*@�t�z�g�9O��C���(jd��E�@�y��1��C�	�?j�����F=�jE��M�}�B��.~iH\Ƌ��J����&�  DTC�(:N1�'.��5c�`u��)Z�8C��495����^ǀ� J�5$6C�ɾC��D��J�,�l9�s&ި'*�C�:)��Z�-�@q`�
5`>��B䉼|�:!�A�CR=S��٫U��B�	 5<(���a%�JA�R"F��B� >��j����J����!!)ߚB�9/R���#�k��Tɂ
6�hB�ɔg�y�#�	�O��٣$��fDB�(!6d����^�=x� ݿP�FC�I?|�!��d�!�X�g&�j��C�ɍ/|)SB��B���A2u�fB�Z��CN�%�� ��9��<�ȓS��(�A�i�)ϐ�y�D�ȓ �L�U@�$�8#��C�7����)��t�����A`T�@D��X���`S��;)F���4��*!����S�? p�x�i��|�:p(K�-��г�"O�j+��?~�a�! �3(�V�H"O�Ĩ�hѩi���,���8p"O�=YQnٚ*W��B�z�f��"OH}R郘[I�q�@�+F"^I�"O��Ah�-n^���aϞv�}p�"O΁:M�p����$OP�B��r�"O�I��	m�D$j�.�:D���"O��%�+�"���X�A b�"O�8cK��c�f������1in0z�"O�q�T�Ӄ,\f,۷�0\Y�uPT"O�TD!F������_�!��b'"O������u���lʘ>Hi�"O E��߰l�|1���{�:�8#"O��"kI:r���FKѥp�aR�"Oh Ç	"j�mp&K�O�䁴"Oh��P��v1�Siߺ~����"O�8�G9f4��AH�b0��"O�(��l
@\F��0c]�f(�x�w"O1��N73���8#��ʖ"O���'E��_�(�j6b�-xTZ�"Op}��	"�q�#+C�l{b"O���MA�hM\0X�H����s"Oq1��K)�M2�C��o��q�B)D���0$�'�Te�� M����c�;D�,��h\M��+�iO$Ş� Q�;D�ةr��z� 0���T�l� �&D���CÐ[�C�G��py��8��7D�d[&��;Y�V���<fz���O5D�,��υ&>�y��@_�]�h��3F2D�d�ecM�*�H��#C�C,�dCO.D���`[�D�I����TV���,D�,0�	|`�����1F�v��)D�TJ�θ��i+a�^�	j*�"PO&D�� �B%�(����?w�:�s� &D��2�νs�L�	�G�M^�ɉ�>D�@Bd�Gi���顯T�y�5��:D�P+F��E3�[�ҫ;���:� 8D�\���߻sx�s���6��x	��*D������2vG �ƘA,
����5D��*6��Ar4P"�����!��?D��r#T�3��W�lR�����>D��C��< x1�׮��u	� =D���`mĤQ��m�4�C��[�N?D�p��ܩFǎ���e�A�5���;D�;R��$ �Z��C��U���5D�Tc�N
]o�q37&�,v�^���K4D��C�x�F�(�m�>�L���3D�l�3�{�h�k�I��g\<�!�0D��v�� m"a�>j�,x��2D�����L�nH�����ti\� f1D�� ��c��(w�ĩtX8�`C0D� XA��C�:��G&�TL��G D��r��բD��`	�C�d�8t'+D���`��~n2$	c���9N՚#�(D��)�I�TB(�qc������*D� 	���Nce��j�����(D���#� cj�h��l�G�Qá�3D�z0�-\m:l��ח6*�h�r.&D���VLI������yY�%��#D�9Я��`�t������`!��*5D��RU� ��~]k'��)r�*9;G�3D�k��8B�w�0� ���TC䉱͈\�"�Wy��i�U)�* ^B�)� ��r䕩h���q)}��L��"O��t�Y��j�`�%�R���"O��KCb��f����րT�йj�"On��q�ܤg&9y@�^&��	�@"Oj�CW�M9n~�: R�=���H�"O��C"K�g"ECq�M`D��"O�C%'	@9 ��e0^L� �"O.�I!OG$K ���ɂ}�f�Ѧ"O6���gG8sid9xsCժ@: ��"Ot���mX���A�-a�Pj�"O���ꂡ.f��!�O�	O:@J"O���Gk��l|i��̉b?vuI"OjH �#�6w�dH��o"*�X�Qt"O�]��f���@Y"�C K�f�{�"O� ����y7^]
`��9�^P�"OP����(L4�1@��R�U��I%"O1"原�*w�mңm_�"��PB"O�(`6 ӽ&Td�S-ܣ!�,���"O�y)`��O�`��+ja�#ԛ�yr.��E��ӥQ�P��{��ٹ�y��WX�U;I�H��F�F�yb�;(��{�ҫ?�y6����y��X�m�X���@!h%�1�uN���y�ҡJ����3�4�ܭ�R�P��y����Z�pɪ�OX ̸�:BHͭ�y�Z��ӑ���pH*��p.�'�yr�N;y@b���:rh�0ӨӦ�y򬂽b��ph�䇂xv����醘�y����ZR'M jsH}�����y�@J=Dez��EZ:rUIs��yIU*3�pɒ�d̔\`v�#F�y���2[ľ �g�.T<*�֟�y�D\isM�,M��`���y���C&�j���4t�^������ya��B��q�n���!p��9�y����s Y�aSH�����y�j�dj���	iP��(���yR�H 21��$�	]G
I�����y$Z�5�Mʁ�$�,Mk�ƞS�<��_��>�)���t�8�QQ`�@�<�a%�T�d�1sL�b��Jf�}�<٠��^��2�	D�ڨ%CF)�]�<Q+�	�Bј���?<*�!�׀N[�<�6��Zr>E���4f��R`_Z�<�Ђ�'v�F�"��6>�T��Y�<���_�9�L�c��б�R��Y�D{ĺ�С�`E�2��PKŋ��yr\�]T�i�1ĝ 1"��5b֋�y�A[?c�\���Ȅ9����FJ�y"�ʷh7@	*aNU�������ן�yR,nvXPC�'s����ŕ�0>iO>�Ƿo�غ@/� BV��)$�B�<�
��W���`��Hbr�!��B>� �ȓS"�)�� g���R$U�6��ȓK�X�W��Y�
�TkǍTy�Ą�nͨv�$K���R�]����l-8s`<v�ԫ�D@+P����ȓ*���<����@��	����K��ix�FL�Oa�����(JS�ȓkʬ@@G�&Y���˝+�؇ȓ�M��ߑ_s��Y�HՑ=
���'��a�O�R���'�.�@	�'����"�wa�5�P���u:�� 	�'%�z$.��.�@DK�Mh$M��yr��� ��P	�Zh޹C��\*���B"OV%�tmN�#t��TE�=IyBU��"OJ�@��5����F�D�7Z���"O�iD!����pQkE%�|�kv"O�i�T��5sH�s�	�F�$��Q"O��r�Fbk�2�x�'�:S�P�
O�7���"�̱ȡ�K�,N��Mϧ K��hO��M�3B
�@r�yA焛�v-��"Oj�S�����AdA�zw
��"Ou�QgV�{dv��t��	D�̰�W"O�ib�c.hр*���d"OV=��(#���R��?-a���"O�=p`n�r�X2,�Yjy�'O0=�c�� �L��RE�E���8$%�J�	�Q�"|��'\"g�vE9wE��3|���`�{���<� (^�S/Z�i�큂7&8�h �y�<�t�--��d��JQބ�Q��u����d���E��¼\KP��b`�#X����Bݝt�!��hX\�����$�֨;#+�f����F{��� ��΀:P& *�/Y�8N��g"O.�����$���e��/L���B"OPH�� �q��Qr�+	�m�#"O�i���H�('EC+i���V"O��J��'��9���Ǐ�2�d"O"2�D)O���"@%� �b-Q�"O\�s��W�Ne#���(��	�"O$A���]�Y�d�%=m>�"O��v�@,#����)Y�f��4"O�M;�$�M}�i�bE* .R�x�"O��3��|�B�7��9m�!�"O�A5$�%j�Xc��t��d�V"Oz���P
 �e��߳}8`�3"O�1-_�)z��EF�4����F"O>�����>���@`�W>宵�""O$�E4I}�Э}�B�"O�H�K��M#���g�!G�0,;s"O������#�B�J�ƕ��`) "O��"cV�d�xZd���FNDD�"O>��Di�_X���U�*D:�"O&���G�4>���i�>T"O���EN		K09a�Ǟ?1�p!��"OZh��M
4i�>�;BH���F��"O�x�@F(DNa��m�D��B"OHd� �϶ �.i�g�Z`+D"O|�6�+)5@�3���]zn���"O����*�{�:4�W �] �R"O��)#B�Q�M��Ȓ�($�8A"O�:g�,R���ևCi�P9�"OV�+�k��2�q��.Ҡ��"O(af�Ƃi��Pa���Jr8�f"OT[���M��!j-�Ld�T1�"O^(��!��Iފ`�v-	-l���#"O���P�C=c��M�ąAiʆ���"O�@+�$��5j�%M0��5�>�y��єG��5CFA�?��U��F���y҇�8 ������4�qč
��y��6pT��	�(�{��E���yB,�[���YvG�4p��-P���y�B#P��L[�A�1k�vE�-��y���G��Q���0j��@8����y���P!0X��B�LcBT!fO<�yR��6@�M�h�1A�8I�u
��yb�ǰ]�4�#K��@��!�T爎�yB*�$Nrp	Ue�'�Ar$�M&�y
� ���L��to\e�v@��`Ԅk�"O�)��&��DnË3Z�}��"O���C�0G���#��\��"OI��*��u~��A	�li�L�S"Oҕ���@b�lc��\3Fj�*�"O�۵��#k�YB�-�k"-ؓ"O}���^�vZ����O�fV6��"O$y���V���d띊 7��#!"ONM���ʶ�ީ[S*�<J)�ј "O��b�IM�,��A��7/�<U*T"O pj��Z�98i�R���<�%��"O��(���1���C��@6��X"O������.MraɄ�J0u�"OnɁV 
!fe�*W�ڞ+9���"Of�ѐ�'(�Y�*�LQ����"OR���|er���ݧB�q2�"Of��r&K;\E�-z�*�G�hH(�"O����V�,�@[a�2o2|�"Op�s�D�&T�~�R��Zɔ}Z2"O�L���%����+��!�"O,�I5%Ngzm�B�5��t"O�L��Es��,3Մنl�-�d"O�\�ebP�vE�i�P��Y����"O�\aD,/-󠈊�c��;S����"O̹��/���Qg�ɧ6��I"O��XR��?^@ ƍI�E��xv"O�y��/G$� ��P�E8ST��6"O40�%#S�M0ܒSm80rj衢"Op1�%��_y�0�!���"��Q'"O�ĳq��iz�Ŗ��p��"O�L3e�g�X����K�S���0"Ob��B��Uv�iA��L�$�A�"O�4��L'��H7Б$���"O��@BbK�)������1"O�T5���t��%����2	��!�%"OV�Ss!6.�K G1P���"O�p�SH	/;��6 RJp	z�"O�� $�JC���i�oX�@��x#"O2��$ʞ97
 ���(H|�A"O�ykW�^�l��K `[6���y"O"��d�L���K�$2�����"O��S�X�lp���dV (�V"O*x#��	?R����EA�
"Od�7�,2�� �.�<*��"O4�!���T��K�|S�)Q�"O���Gl*������Sז���"O�!R��Pǖ�uK�31[<�Z"OT��Q�E�|��Ll�tQ#"O����C���m�P�5jQ���0"O�%��k�PI�'E��"�
]J�"O���Ĉ\(_�U�DÌ�fz��b"O�L�֯\ \�d$�փ�)>;�I�"O�9UMv����w�B�
&���"O��1��<b�V�ضHR<(
*�#�"O�����(9M�1 G-�0ܪ|�""OК�X4K�u��,�8W�^��%"O�%1#[l �� Cˏ#,�1"O��v�E!0�
�o%Z��&"Oȉ
fgȟϪ��4�S�be��"O��p7̎,\�|�`��y��)"O�y:�
�@���*��2upW"O���0bQ� ��W�X�6�i�a"O8���S�D'N�C��(�t�)�"O������0��{r!�;8�Hiy@"O� �a�Q�U�Ԇ "C�C�b®Pc�"O4�bN�3�z��t�� �6�Q�"O^y��B:H�Zu�k�2**��A"O��	���'�v�;B)ͨ}�)���'�b����9$�̰��O�5՘��E�a(���0�ܰ��X^M�!�ȓ;�(����Ҁtuθ[��QhZA�ȓ� �e�בB����4*E�ެ�ȓ�Ƭ�P!ӋY�T�[�y%Z���'*�Dʑ)��ADbA�S,~�8ez�'v\)�]��C��L�����{�<��@����Ӓ���p�<i��P����Fn?>��t�*HI�<��D�{쬄�0�G?D9�R^> B�	%�<�%�|}�]B��"�8C�)+�3t�4����WD�	_�C�($��h�(��^�Q���B�ɝpC��Ȑ5�Q5	�;3��C�ɰB��HA�̃w鲱�#�,{��C�, '8U��h566ni���_OxC䉕o���+(�:!њ���O��b��C�	�11�Ј5H��s��"��}�C�ɮ��I��^���Q�Ro*�C��38r�mY�Ch)����-6$�C�	�FF8��J	m8A	��ΈZZJB��`7� 1�&��zZT���k�+��B�I�9�񃃆,7^D�V��r�B�I8Yz�y�K>A.�uQ�d��xs�B�ɫg�F��i�)���b�	��B�ɽxU�@�$nا'��kW�D�O�>B�	 Gve@UL�#b �(T5��C�	�K>�lKB'
"�"�AV���O�B�	�
� ��a�U*	�� �@�<C�I�w�4Z�郌��X��I�RB�IRr��F-�7 ^�h׃�kp�B�7_�$��ʒr��8;�薈e�lB��$a@��'f>x��B! .6T"=��1 �bT�S���Ow����L�wz��@6x?�L[	�'0���6iC
:��2R��'j0�����l�0�����"Lu�󧈟��Q�:-��q�@݇Z%xQ�欌�5!�Ğ #�QP�Rz� �r�,���"��d�,e��O3-�]��ϨO�p��db~�YF�T>aΌ���'���L��!T�!�@���n�*#B�M�elD�1P��?��~�d!)��y��&�t��ܚӆ]!׸'Hj�q�.�*'�iy̒�5\��㴤�\��*�F�6�b'{�12saC��y�C�(ބ���Fݻv|��� 99��Z�M	�=g��+�a�Ĉ	���	�1@q�	l��i�Lw�2T�U ^"!���ď�+hn9X�*���6��&���>� ���&�7���b@
�+o��س��*kf)p���26�!�a
"��/�#bz�y�!�"��#f/E�gw�y����vr`���+*X\5c�N�4^�x�QG�F�H�����Ig@ �+!�	1p�pƦ؅*O���6t�@�It(�a���8������?����3OJ�����J�pMB&�:D�(�fD ,L�U"!ȩg`�P6�jN��r�'��:&��e�j%�v���A�	g�b��Z��M"A�������gB@C�	#a>�1�2��9H��R�٨I�Flʤc�*g�C��.�����I�$O=�%�B�P�'��ł�a�ٛQ�OE]�h�e�R!�WC�,��Rh�!�^A9�L��m�4���3۾mb���7�Z���Ǝ3�p>�V/x ���Í��\���M}b ��lڅh�☡avz@��"N�zѠqƜw(�B�ǆ6z ��`��ӎL�P36,��K1�,
U̓Oh<y�� -	��,g����U.491Rb¼=1֩:Z粉X#CQ!.
��Lڐf������ɼs�/WKܰAtEU�gi�l�'g�IX��/��t���&��I2j8A�O��ʶ��0
6l�(��c����å	��� ��J5zF�ΝŪ���Z�hr��K:L\+p*<e��ak>���eR�J�NH��=a�$���%P�����J�<'lD21�ʊJ������9���K��!�����,�*y,����䎴B�a�"K�1!�0�Um�
[��L3t�P�(��+�ϓ�Y�h��U���D�U��+�%�>���X��TT� XD;g�U�7	�L�Cm��g;�]�sA�q�Za��	=$���V�́
`2\��9mc̣�B�*l��8��FC�H��dA<#����LM�
b*p��8nf杨;�zL3�"�� �p��H
N����Ĕ�G\l�UU�m4���bD<d���G�R7���cB�8a.D�I�\<
�±MO�]�[A���EC�������\��U�v�\�Z&'�^�n��?��+���x5H�DȨ�$��լN$���Z1˗�LHl�"==���i�Z�^�1 �E$-T*���Z�U�`�� EXLڊ�D��<P�r�E-R�^=�
��\�`��B)K�O��(qe��/Z  p�K%z�.=J���6g�/
 s	?K*���Q�Т^�f$��FM85�p���Z����gO[�u�| ���̔`z�	��Ь�U8�, Y��dA'ړG
����ڇp�j���͖et�)Y@������W
(�����vg@-���:|O��A'�� 	a���SF�'7���HƋp;|�K7��y��D�Sl�lA'�F?r�x���M%2���`uK�s<r�sGoׯz���	5�D	̈́V��XeP�����2��nҹz��h=	����)<���)E��	y���*����H��|;�8I�jؑ\��ǈ�:}����MF��E|RޤU�.�I! �<h��ȫ�nP�A��Yj�����ۆɍ�9�8�^�V�"�aq��=j��ܛCNтD��}e�!f1�@Z�-�9d��]Bso��/�^1RF��$�0?�'�GG�UR7�8 �M�Cc��{!ZLHD�%t��{��<?�9���DCO�e"7h;�a�Ã��] �]z�R�kBgN�X)�4Q�����I&*H�(�eO ;�l̓u�܀J/th�í��;^,-�3�F<[-�)�↕9�X$l�Dq.͸�9 �V��B[�t��ɤm�j��q.�A�,����V�x"<���K���q�] "�0A$I �����퐍w��Y�҈U]�L� v"��J�Dp�ܥ/�^�E.�f/"���H�v�Σ>�4�R'&xf�צC
V�X�ӐdZ	M�(eBҧ�yj4�P��H�����''zb�ǆc��z���j#:��	��jٌh����<@z��b��C�N<m�֭�v؟t�����L��iBhJ%�aɣ���?�L�$���y�NX>�:x��¶N��i"���?��c�Q�5��%vݸ��:^����E(=�O5��P;�n�"���i�U��%q��#�Q  .K��R�AO��~b���qZ���Ԛ��4``��p���(&�@��5�� 2`�D|L��mܕ��_Ȧ��@h��#�	ƾ!�m)��c�\���4+��I��F��dN�hW�xr萮U<,��͘p�`�����DA�fiĀ�'�`Ԩj�'A�4 Th�*LB �X�����@��	�]~�=��'���pY$�,�j��N&>�4�2��^9H��aJ>!^9@���~�]�2c8�`&#�_�@9��N�ݜB�I�	.�IU�_���[�DO�p�x���P)h��i(���T��5��gܓu-R�Rt�ٌhnp S�B؇��-ivp A?O��A���}o |B�.D�z���*]��9@�9����&E�Š�-N�T�������@⑞
jb�~�(J��S�Н3�%f�]���M7{�t�`�'Q"DsGb�>=�e�w�@q�`�0����ҍp��S�IRxU夅�n9�%Jd��V6B�	&<�8H:�*�7ξ�Iv�����	$b�J}k�}��iS����[�m�����M8G8!��]�].�6�ۧk���D�_8!�dL"Cd9����#GH��͉!��խhЈ��rI)I��D�r��&h�!��	���6��@��LgK�P*!���tY8��0-�9RILy!�Ǎ`������q��l��iR�!�DX*�za��բ]���R.�<i!򤚢_g��ǈ�hw��V+�&B�!�ܨ0$p{���-r`��q�j�4f!��1���CHVg�a��U� �!�DO�# �-�:nF<ZwH�!yX!��=�lL��CKF&v��5���0!�$	!����菑1&�ٔ-��4 !��3<2������

�a5E��@-!�M9Z3�	�O�H�ID�G�!�Ą�;��9򲆘�[	T���CԏI�!�5.�,,+�M�"��p��ŏ'f�!��Zސ�##yӆ���DW%r!��;xͰ�s͔�jҨ �XKE!�	��tk��ɐm� ���ӂ@�!��[��Dd��#L"� ��M�!�D��7,N�3���gMt�`�)J�!��ÇH�`[�g@�\D8(ӤF�~����	�蘉�T"!�(h{W�0�y
� �pah7��0)4��4{�.�%"O�	"��x�

�(�^}ٗ"O��C4wq@�`��̾Q
�
t"O�����	� +��$��g�:I�6"O
�{e)b���a�R��V"Oı�7O�B�~E	aF�_�^�Ц"O%A�m	�7)�u�O�T���"O�q٧蒇9>t ��K09��E�$"OnI����o��q��g�<&�>�Q"O�C���1Q`ZY�df�5V�r�K�"O<DP�Q�o#�(j�E�&�y��"O� "'��%�~Y�TD�8b���W"O��q'"M�|�rdB#�22���F"OD�eBF�D��B��
$�4��1"O�!;Ć��Z�v�
be��)�"O��%���Tт',�"R\� �"O�j*��7�Hfx(�q�R�{!�"XD���CK�u���)� ۏ|%!�/*���@�Km��ӱ�E�!�D�(	@�+��כU&�=ё)ڑ}�!�$�Rc� A��'$*�eCi�)�!�� *��!B��	"�R)�hp!�䚖 7�:oX��2�8�N$Dv!�D ?>�\A* H���#�V�!�D
|Nr1�d鑢,o^3����!��OZ���(ٞ\M��T���!� ���)A����ɥ��rR!�ă�]���E�B�NJ�j��<3�!�\(F+��b�� �`��b'��L�!�dΛMX,y�@��c�������=#�!��Exy���W�I"6��q�i[�%�!��47ix�£D#?��q����+z!�d�9d��p�M�2�h!H�h9_}!�dH�K�p+S��X�j!�3�̫�!�ӭ<}�|bA��'=�`����:8�!�΂P$���1n�V�I�X�B�!򄟨e8�|�G)^'.���I�� �%�!�$W�C&���Μy�ڠ�E㕍x!��Y;.]~�;bJ�8+z�H��A�F!�$�z��Es�`�-g�
�CR�T�!�L�iǒ�J�a�4m���n�!�$���xb	�mn�K# �.g�!��$`yb7H�)_p0���U7]!��Ol��B���'R��p�� D'!�DY�'F����
2�����A(}!��-�}F툈e�^)X5��=�!�Dݰr\q�al���SJ� �!�D@�.��C�
8VH��w�M�!�$�	�nh#�&��tvȒ�IN��!���q�@������j54�4J�!�dK�d�\P���59^)�7]4�!��6+�y��͘q��+ ���!�ڙXe2w
	���LR�
�c�!�E����:��<x��Щ�K�r�!�$�uؾ����� �<�Ӆ�ٟ<!�D͒Yx�%0!.��!�A��3!�H5��u��X�g�9R!������B#�L�Vƌ) �!��Đ;��e�s�Րt���h�e�$p!�dY%)�e�l�?R̢ �aCZ�.i!�X���<XqB�*�r��ܫx�!�( ��P��_@�1� �!�d
?֤,z"+�X;"q�4ς*6!�� 2��Tn�		�yhRĒ4Q!�� �Q@ʛ|ZT����H=4"Oftx�G�2�t9�@N]�`@����"O�Y�׍�)���y��?C�v�8�"O@�����e���&͈!�lu��"OT��@N�.G��f/H/5��5�"O���̲s^&��h�2<�l��"O
��&GB><x��M )�tA#�"O:i�so�O��Y�@-��;&�Q�"Oz���BR()ؼ
�lؿ"t4��"O�B�T	O%���"�5�\HX"OH���WN4�7�5VĴ�C"O��`l)G+�	 v�U%)m�v"O�h�Ɓ6!��
3��v<J�c�"Om����4fw�D��-؆vZ�{E"O�YY�n�',���$I��Q�(�!"OF娤×F��x�'�!ĺE�W"O�\CO�S'<t�ܛ}�����"O.� 
�,?I���d��5p��R�"O��v�5)43c�X&yk�`��"Ot�h�@!lzT�����".�Z�"O�-��"�6p�X��c������"O6L�aE�,nT���"H &��āe"O�1�W�ǫ7������P?!����"O�mff�в�h?°�T�P��y�I�c_��A��{�mG���yB�H�Z�P#D6���x��S�yR�N"?���#7�̀?��a偎�yBlZ"� Ń`lS�E���8DHˁ�yr'8&.���!�� :�;��%�y��F|� �:�/ۡ7#��� �6�y�H		!����%�M�&��yCĝ%9��5�9ACfI����y��*@���-9ܺų��ҕ�yR	�4���Y )�>�~tY��Ҕ�yr���5	����nˎ3*J�����yR�ϡKN�My�拸8:��`�[��y�X�VE�;0"�>7�@1b͜��y���a� yC��Ո'�4�9�F��y��@7Z�I�&C�/�dX�NZ��y����:��\c d���P⠇�y"�у~Y2����&Eh#���y�aȇg�)��,�/>�F�kpAR��y"��YN�<Q��K�\p
G�*�yF�FJ��m�#zjQ��"O��y©�����5�D%y��д�_&�yr#M�q�m�Ќ�jΖ��� �y���R�<r Ǖ����!֜�y�	�n�*�h%L)����ؒ�y"JB�U��
Ç�p�&ً�.±�y�*�~l�3T�\<�!���y2+�s�����k�޴,�`�N�yR&Z�X���I���i(FTP�Z��y��Xav4uC4J��BCEf¹��'�41��fH`���K�{����
�'�N��� Fa�A/!^�
�'�x�2� @ĸ(��$*  �k�'���{E���vf�Hs�M
Z�&���'x��꒘n��ٛ������8�'���w傥K���,a�}C�'����E!�H�x�c��	����'qb�l��*)�$��"�����'Ҙ���B
*dH(�4c�7	��'�L�5%�3��Zw隅�|��'Ƃ�A`��HXRK����"��� bd`oD��
���Ч;JB�b"O` aFO.Ib�C����F;�M�A"O�-�ħM-|�8R(�jz(-�"O�/�-s~j�ئ-�"^����"OvI*ĭ�kIްZ�I#��ݠ7"O�P���39�>sBW����)"O���DMP�;F4��C��y6e�7"O��z�JG?i���Z@�dkzI�T"OHl����	P�f ���P0�KV"O���G_)M���XWh�!JO���p"O��BwOZ�h�=S�	E�w�$2"O�(�TH���,�eB'pe�+�"O�����;��+������"O��������*BG��%~L��"O$�2��R�V��|��& �3�걺"O�܉���8${b��*�y3�"O��@�OއM<HT�K�R�iS�"OL$�B�3}*d����B�� kP"Ox�
Ae1Y�r�N�"4`ʼ2W"O4 �T)C�r�����cX,Y^�)�"OP�pJ�>3X\1��*0RR�"O:�(Vn���M��L_�d*|8zu"O@�&{��\��kS�sh[2"O���
�aC�C�Gz ��"O:��Э��r\>3����Ga4M�T"Od� �5J��0����G]����"Od�X&�	�F���
���$B�*�"O� '��7�T �S�K�,� "O�8Q��F�JG�X�H0�|�7"O����,�I��*C5\H��"O|��BȑT����_
B$�� 4"O�!�"č=ut�zC�?M, x�"O�4:c儦(oX�9�dB|T�Q��"OƍR�o
8>&�e�2���LW�-�"O�@�醊	���1AJ�yGfM"5"O*m��E��bo�%�w�Nj��"O�M�2(U�E�8b5霅k��L·"O4�`��=:o"D�uh�Xk<���"O�����*弅�է״OW��:6"O�4J�=|ޅ"�(Ne1`Y��"O���¬��dOx�ևE�r5���"O��I��9A��<����r��"O&mBA֘���"�+�u�G"O@�{2��;;��bg!�02v��h�"O�qZ�'�1�`��T���p"O��I��vJ�Nb\���E"O4j0�G��9�!LJ�M��X!"O -�&Fԑ&�����,>A@�9s"O�p���F4$r,�Q7�['HF��x�"O�}Q������$;_2�����tB!�䌽u��Yʒ.ϷO7X��A�5;K!��V��ƭ���T�	�$�ܑQ!��SZJa�b��&y���2&�!���ՠg̝%O�޴Ҧˣv!���}'�Q����d㪅�K�<c!�dZ�%�@�꣪A>ѪTi���!�M>�уg�N�V���k}D!�$T,i�0k�䜰rvd�s��85!���
�d)�H�;GX��'�O� !�Dا �J��B�ɕu���ʞ�`�!�D*+�&�*ˤE���(���L�!�D��b�LW�X29�4MJ���!�$�j̬�I�%�X����N2r�!��
E�P����-]	
�&�L�r~!�� ~�Y�K�0/��V�T(.���%"O���dF76lQ����27Nj���"O�5�QDC������ Z7��Y�"O�eR�Ф�;@H
^�¹�a"O�bf��J=�i��Փq��T�0"O�ā�W�/��{eC�:6c�Qp"Ov�����X<�|S��qBlt�T"O �SO�Q��1��#ыF461pQ"OB�|?`���\8��Zt"O��#�Ǚ�=X�	��ˆw�D�"ON}�g �Z� G68�陱"O��I OW!���Ү�r/�@�!�G�.�t`������qQ�9[!��ڂt��B�&K �� �O��PG!�D�:�s�E��H�:�cM��!�E�.�j�hŧ
�(�<�xD�ڷ`�!�Ĉ�Cf�3�%�7d.t�@�)�!� d*D���9`�y��B?\�!���O�N`��$�++6�Ӭ
r�!�d:+u�e��K�-2d� ��=!��
a�r8�vhŁc-$5�j��4�!��Su)&0cE��&Q�F�b0b��H!��M>*�8��g�K+|��%JA89!��W�x����G����釼�!�DF�'�ށ[t,�7d��'G��&�!��(e"ZP�v��~s�r�A��#z!���8�yӧ�F.3R��җ��c!�DȎanZ������`�$��%r�!�Z�h��!�t�Ċ��Wctw!��\;3�jՑ'a{ǤZ+ӓG`!�d<q%�L�EÞvn\���*�Vd!�]G�,��V��=/#<�(�6�!��?T�0k@�ΫA.n��ꍊh�!��ZTɐ%���!: �
H(�!�N�^��4*m���uN��O!�ڌ>J��˵ ܦs2L��@�U'*!�G�4p`�L$�]�Q�ͣ]!�D_�m-zx�(� ppԏ		!�Q"�L��Kx�H �b�!���a��Nn���n�����"O�����g���p�k׉\�0@��"O�@i$+�6%�ݨQLV��ly:@"O,��g	�3.���A\�Q�za�"Of��oL�R���z�J� p����"O�,zw�_	(`5Y�	��`�u"O��b�n�b��O(���p�"O��S����D�^A����SqV=[�"O�B��҆w� ��%��O�D�1"O�q�s´B��`�c�ۅ#0�0I�"O\��!�U9RFp)�@�#o���Y�"O�ͪR���5������Ys�H�:�"O\��3CD1C�l+���+��&"O�	H�@ӗ��!P�����"O�ո$�M�>��Uх+�g4r���"O�<9B�"�V�zD�R�VL���"O⩱&Ü�(�I��J1t���"O�����G�Y9#��p�@�#"O
P{2��T&Ȃ�����w"Ox���\�*C*Ѩ�EU-:�ܕ��"O� ȑ(��OU�d���9O�v�Y�"Oΰ"�.kA�MJ-y?��"O~�Y4Kȏ(޽;&�M�f����P"O�������TF���g��'��#!"Oah�Ɉ3`� �B�ň�f?r�k`"O� .l�C�C Nz��%�I	x��q"O��e*قS?X� DW.��"O�Ѹ��9F/�91Aȴv�Y��"O�H�5�\�L����� +�l�b"O��[SL�*}Yn}@15�D�"OF�2�FԤW�PP�eɀZ�mpV"O�a�(��$�(�BKٴ��p��"O ���,\C�5��$A�&�:�A&"O�I�JH42L|�⤊�j�j��0"O��C�-@���D�w�9��!�"OEQ��ї1b8�i	N#vd�
�"O�]��@%t���@W鎫K�p����	&�h:W��s������8Ӗ�D
����Ó��2j�|�F�ڑ*,�	�<x��"~�� �M�^T�%`�zX4h��/� {
�$�L�l�������^4�>9���-X�p�y�&˻)��j�n�H��Ԋ��'i����-�!V�4��	Ø1����r �N��8��N�l�2��/Rh�d/�
����O���Z�m\po�ɗ�	^� �3�4WJ��#� ��](�kQ�x�a����#J���^/t���zF���{��9��I �O���JG��챏�~�w�G.M�$��4I�闸�2�`Ē4L3�H��1p����MG�4M� ���`m�S&|����;"� @�ˋFФ�1u�W�^�򄱋�Ě~Z#M�5��}�@�֥F26�2t�5�eP���lYb4CèCf>5���x��ݸ�Ā�^j� A����J����n�KI���O�D�:M�d�1�d��V˝�yl��4 �X��u�Vf�i�ލ��Hb�%��odQ>q�Or�|��L�.�~�@���Kt��3G��k���ڑ�G��Ma�β8ca�DJ�C��D�N���%cd�(_��41��Mà�9d�.�����?7��H��x "ŏ
*�[ƨR�X!�����;?���%����O��.D�p��!N��F���s	�'{$�S!�O0!T �Ыժ:4��q�'A����*��0��0�d�Hq��'��ɨ��"Z��A�P"�:a�<h��'|RR�K� M�0H�[�>L��'�412��#ZK@�kP��(�"�Y�'u���PϜ��pR�E5\>E�'���aF��;Q	��A��
 ����'���B�&sy2"r��FtA�'��Yq�=VxE�Q��#v�%��'��*2ńu��DJd�^�)s���'3���Bq�dz�+-+zL1�,D��BL�31_*u�	_! �XP���+D�@Kp���!qRLBB�,P��$D�X:tÅ?Rjh� ��f(� 3�#D�3���D�,�D���w�T2�!D���"E��r�@�F�
=GJ��C�>D�����;h�Ȁ��T�4Դ�&�>D�@J��,
�R�`�ԇ��}c��=D�����G�B����Q����#�:D� �Z6�����gL�e��c�9D�x��'�9��챠��.j���� 7D���&�@�.�.풴OũF@*�X�J4D��k����4���.'2�˔�0D�Hj�ͳkÆ���)`��0��.D��ಏơ@�%[�f� ���+D�8b��V�>�� �AW�0y�a�VK*D�4 é��cg@Y�Ġ �9�ҷ�)D�(�T�S!-<����b��$,���DG)D�d�0�¯F?�`�$ي�V���%D��P#GN6�$�D��w��J�"D�� `��`鈙��`Ɛx����?D�D��� �piD�n�6:6q�� �y�<����M@��k�'β��m���o�<�f%i��H���ǣ=�j�����<!%�$�z���`�Y���9�oU�<��]9ʜ���D��y+��Y�AM�<i2�n�d"k�0Q�~aAq��L�<� �22�P�n^ޭ�b�;'G�]�1"O�qq�/����ؒ�F�%E��"�"O�Q�r!я.�`I���	*R�� "O���D$:Z�4IvG� I �
�"O�	��cՈ['��+\����"ON		uh92�[BjЍNeB={c"OzXAd�Ă
�D�s��5$B�"O�"�#O�@�@A�&6Ȯ�9�"O�Ps�h�?F�TLC֭�6T�i�"O�8W���<f��Mɩ@T��"O�4QĨZ9a�F��$��� "O�l���1��u�&$A��)sd"O��b��m˔�
 ���J���"O�[
�~�d f�^�U�8:�"O���I�\��t��Y,=��aJ�"O��S�X �� sX���%��"O�B�*��G��9���=����u"O�����$:�H�/{ �`�"O����љsL�&k[�\#8�"O�Y:�@�6m~��t��q���4"O\Ie�Y�bO�xӧܿ�����pE{���_���Ye�}������M!�dE�,��L�(�,A�V9#�.�*}!���S�^��E�y���rm� ,!�d["�̍��C!Ʈ���Ɔ(!�7F���Y��V1H�ј?5�!�D%N �p$�(�ܡ�V���7!�d��[P����Ǉ�tU&��W)Px1!�D��^�Rq��c�bRb%�֧�!���<���qg�ެo���R�d�?�1OB��D�	L����a��)���!5ʕ{!�d�F�h����"�Ā&��,!��^c$�0�gW�x�t��&��;h�!�ğ�'����Sヮe��y�5�!�R�r�$Q�`A�	���:�k	�/\!�dT�bh�%��%p@�ԪA��3L!�d� Ru�a �N��(L�v��vD!�@��~��R
G?b`�󫄺	�!�ߚ#��D�'G0{�*,�hT�Ik!�$�)9t��b�	}��p�h�,p^!�$�1(o(�P��N1|s��eȄ5ez!����x�!�Bi��q�]/#t!�Ć9-INÒg�7+|���& H�2!����k҂θeV����U�!���H�����yT��ʄ	[��!���$ �����[W~��e���pI!�Q }����@%�`\�E�c!�,1�6���a�%ANEI�M�6�!�DQ�;$16�p%�@��/;���ȓza3S�ux���,�s)�}��1o�Q	�J>ww�xyB��|>���c����э�(O�x�@�lj���L�6�J��J�0���0,�����ȓB�V�xG�#�ً��_R�<� &ב�U�e	/���!��L�<�E�9\K�L��
�K%��9�K�<�g U,%hv�f�4�*H�2 �G�<!AM�-���r�Ϥ��8���E�<Ien]1�LT1��P�igBuA�nk�<q�	_/v`��d
E�j�y%bTp�<) !wE�����6V�Z؀a�i�<�fO(l��i��gݪh�r��w c�<	SoZ�c:.�0go�N�*T*NE�<YVI�9c�b���b	�*yL�RじY�<� ��b�/Ȕd��0������"O�upRDT�V�Di�V�ڣg���bs"Or�����=e� 4 �˙n�H��"Oz0����0D��ǦJ7��,�T"O�`�À��u�P��fD�L�2�	"O2h�
��a4��)�X$x��"O4I�V���=�T�ɲN��P&"O�iu(�[`���K[�K&"O�A��ዹu�j] ����eX�t�"O^�+v�	�y� �("j�k��E"Oh8��ٛQ�������)�L}c "O��ac0���,!����E���y��X� �d���ny��9�OZ7�y�1�Ș�`�׸7�����M��yb���6O��z��	�C���y"DR�n_8���#�B����ycV���t�A 	ȵ ��yb.oì�xUCP�'h �p�[
�yr�o��j%��>5�*�n܅�y2��0w�X�4�K�)`��Ɖ�=�y��� �x �3�Y
1U�\�㋋��y".ѣ@F|���J&鞵["̴�yrJ�=�J�D��2�zT9��y�:�J�Ô5y�������yb�^7'J��$[�(�DA�q�G�y�j[WD�����Rtx �0!��y�P)��B`�O�K�Ze
U؛�y̚�z�!�"9�2��I��y�%��j���a�N:+y�a'�y�a�o���2b6z:�uB�$�4�ya�0A,�BaF��x,����G��y��I2�<�V3wbڭ�6��y�o��\��50���9�f��FmE��y$6�@ ���/��8*����yB

&f�x�� 4& Tt���̇�y���e_��x�DY��<�"#�܎�y���k 5��W�B��R(��y�ܬ4:f�6@x���# �"�y�
gO�I8'#բ
s�p��6�y�O��Zh�C�����'����y�oF�=���q��<
��(X���y�3T"�4,&`���g�y&���}UMV� �0h�e�"�y�
�g���"���hu���h��y�$H%)��yQ�j�d,�9PV�y��3=���C�L�l%�����yrlݱxi���F��;H4������"�y¦�;ц\c��R�P̚�P�#�y�BJ����T��$sJ\��yCփrr��C`ǌ��T�C�y"���.V��@�HW2B��y��o��y�e�F"0LP6dJ�:~�H �����y�#܀����ێ/�	Y ���y�F#���%�]($$$Qxf�!�y$[9QfXر�+�j�Nq�B.D�yr�3v���n�O�cW���y�2F��P��!��`��C��yB���"�$���&'�����y�A�c_V�� p:4xuF,�y�!���A��8QT94mǬ�y��N1gLH�P����&��$��8�yB �3r6��x��}�<P�I��y"kǧ��l����g��m�����yB�V&V���2��]�5���NK��y
� 歱rGP�p6VՂ� j�:I��"O8�#�,�#O�H8�"@}��@P�"O8q�!G�(vJY /55|R<�`"Od�	w�ԑD�,CE.ϜD~
Y��"O,��c��g/r��m�1tF� ��"OFPÑb��:�f�
#)IC:��&"OI8�E�<��S(�RU,A0�"O����	,\�v�+�l��l\ř"O%���,�nš0��NB��"O�]x7bP�pd��dǏ(��cq"OZ!Q���`��@���y�x��"O\%���L>n_��q�M�� �q"O� RF�
$����V�H�n�����"O2�B�#��L0N��h�=�����"O¥�F�=��Qd.
8y+j�"OBx�V�ŐZb����� �f"O�}Ra��4&��]Бm�
�mH�"OXMraM�0$؄y����"O؜[EɏV�iC�̏����"O���v��V䘊ekT ��	ڂ"O���f��/D��Ո!��1�1"OڙH�w��%��bZ4F�~��&"O�[��߲u�x����M��p�"O0�A�t�Z�68p�=q�"O��$�r�Ұ#�F3��0�"O��)Z8��&�#Mo~m:7�	=X�!��Rι�T%I�&n�r�F�t�!�CiΊ�
"�.H�9A���=�!�#6��P3�\ A�=�SJRM�!�ά'�.t�5eϼV(���
G?!�O�P'@�{Q�?8�vt��N�%A!�䔈q\��
��5��e�CL�1!�K�!�y�a�0}���	F�_8F�!��9a$	H#uP���'v!���������v��`gf��!򤃂3�R1�� �5)�,�"'儓A !�r@�)J���2b5j���c�I�!�D�f���s�03�����\�!�$ǕK��eR&A�MH2ɑ�δX�!�$A�#6d��WK!(�H��Q�ƖH�!�$кX�	�� �/E�P�25axr�'���qc��Ħ������Y�Ι�Xmΐ�ƞ�~��2d _��?	�2 S��?��X!( ��<^"8g��9�^��5b3f|}�0GZ!W#�
��&jLZ0�U!\\�'W���V)oQ,�C���=]L�xҰDo+,�j�@؊Y-���DD˾<"�ĉU�r�'G. ���1*�6B`��6-�-0��B���I��������K��'l"��?Q�'��ʀ�N'��mҕC�3OQ�ٹ��D8��|�q*"@|��@[�$�qb��E�;���i��ɼ Y�U��ӟ$��A��@�>P��!QbB��� �O����I=P2��Ob!��Ȕ�7�FL��_X'�iA��x�j}��~��Ld�J�"�&�F�P���@�I'!����:)(�rjS�g����/{��
Z.x�abHE~���Q�?q�\L
n�$/@�I�~�H������)k�S!Mt�v�i�*�k���&%�������QGJ��&aqk_�GݰEh���~8�#ش��f�'3�6Mn�<%���ѵmd�Tѥ@ �Aqi��M����?9�3y*5G� �?����?����}{�]9.^
la�m�dv�0����?�E��%͞?�B8�ee�h�r+�Z�)�)|i���'
�s�Ep��S�L?B
��Cf�n�2 J�A��@3��9eq��H��ռ���ٿ�����O5H����̋���7-M@y�D\$�?�}��ԟ�lښ.�d+���ha���9R���i�R�'���0�K�$�(h�"�&R��aI�'[R/c�&Un�~��?A�So}�bڼ.��e6Ö���\�w*X�,�r�S�S>F���O��D�O�E�;�?����?�/X�V�*i�V"�a��s���3� ��*�CM�$y5^#'E�x��&D�b���Eyb��(%{|�� ��_� �[@hĀd2l���i8
Q*���yX�)1Sʊ�e'D)�#<�I�)H�e#ql["X].��sJ����؁��ONn��ē�?����'�(ڇ
3�X-�B,E�M���X��/,O�<3��E�EA
}0�Ú� ŀF�Is���M��i������ߴ�?��t�? h!!1�ѫ+�hr��ާ/<	�u��ٟ����w8�9������?G �S���;#C<�#6&�&�4S��\4d���bf��n!D� F�%�
�&ʓx��hKe��~U����)��0%�b�Ȏ$j�a�mj�0���<�g�|ШR�GY~2b϶�?aF�i�����3Hh�rIJ�T�0����1l���ܟ���b�S�';�fū��]f�B��P�Qd��EyB�*�
��!x!Q�*H�5��ថ�� 7	,%��Q��H���M����?a,�hiQ iӞL�C-Z�n4N�*dG�b�D���П���,d�m�8�|�qСW����*]�.vX���<��/�=�(*5m�wm�S�x��W8+�<��e��p�<� 1�q�d���c�M��	�zt��o�;s��p�!���� D'�����O�lڰ�M����O�~��`EֽL�@�مN��  ��ON˓�?Q��?�-O����O��2n���i���T�&���N���p<�7�ixV6��O��nZ¦90���[l��C��9���eA���?���䓈�O�A���  ��     �  �  %  �'  �1  8  [>  �D  �J  -Q  pW  �]  �c  6j  wp  �v  �|  >�  ��  ��  �  H�  ��  ��  J�  :�  ��  ��  �  S�  ��   �  C�  ��  f�   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6�F{��'O��V���&�;�+0:��x	�'%��"J�[�]�R�K2r��"
�'Oe#W烹�R}aC��z��
�'��;��7�������L	�'�:<*b&K"4����M����9	�'نx!c̓>�D �,ݻ2zX�R�'��@ �F�9<�m�7I�"+�a�'ր����>��Y�
�%&���'��0��3L�r5��M/� HJ�'U����J08fx����I$p:<���0��j&a��'�L-�I��w$��
��Ig�<A(K74~<X��.>IG�t2QI�~yR�)ʧi�n��EiY����3e��c&�D��f4���W��'^�4�KR"l&I��y���.��~#S�˩y��)\ ; \���EU"�D`A�w+ Q��\ ��/��i���bND��xၜ �.���+D������..r��nE"gp�`*�H)D���C���*����e��b���S$D�0�@%������ٰ �4D���HݦeF����� <����ķ<����,f�Z%F��T�:��4��4z�^C��*RA�C�呅[w  Rcífc����Y.< (��x5\;��*�ڢ>����*���?�Yw�6�MðQp4c�#��5>�K�'4�� M�G(�X��ա-�c
��� r��QIG��L�I����"OZ�����y�S�+�1tYL�p!"O��`qaʜg0�bj��X���"OTQ���[(�qJ2`ʉARb�H%"O"9 MP� ��#3!+L�"O�����@�Jl�2B�� �|J5"O���6f�M�0��jI6�b����'(1O� 
����8�bgJP2I�Ѫ�"O�)@!+��9tL��(� ��X/�y��'�=�����r���#�6�K�'�8L�W�>R\��I�6tP���?O҉#�CĵOH�p%��.^hpf"O�q#��p�4#5�۫ߢ��"O�<�bi�(�¤@�EL8#��R��[�����)�~�FJ%ᖰ'Ƥ��bC��y�m��Kk�Y��� �^�)��T��y"����<�W*:o�̩�l��0?I/O�H��kA�<P#�0C��p�"O���B��A�b�,B�@M����>�S�4g�9j<��UϞ>7�
t�T�_!򤑦nRȅI��Q+Lߴ$��삂z�a|��|� fT�!�n�a�Z3���8�yo�,1H���ǡh�8��D֔�y2�K=h�&�)[��$۵�	�
�챇�%�Ȳ���	�L�3e��K����?�����w�ɟUp��o�5w��Ԇ�In�'�*�y��(��Գ �U�vi
�'��m��C�`����	��Q��-�ד�qOH��c��,X$�� �ιVd>�pR"O>�!��<��;�!��7R�l8�U���'��#=%?u��k-@k�਷"B�n��>D�X0����bp��@6�0�􌼟p$���I'Nn�����T3������>���<�ґ��Puv�����.wBjq�CMY*�y���[�p�Q���!w��QRbQ���=!�{��5;z"�!GanU����ٸ�yb&�.Z����#�ֱ!A�*�(O�,��	!d�t�"Ai�9[�&�xB��FB�I6	:�+�Oʇ)�|P�N �2�D6-3��f,�7$�\#v��S��`&$D�X	dj�1~� ��5k���Ab4D��"���5r���5�#y���c�/D��"C�./����c����ts�1D��B�k��}��I�����P�^pPC ;D�y��_1Bvb\ägU3w�6��7�+D�|�Q��`"��G'u.8ʂ�?D�P��O�2(0�q�i��y�c<D��Qv�I�/( KEb	�rvx� 0D�����G�0�n|�� ��t��h@�0D�d;����#�4|Y��C�*����2�/T��{��.	�Frc��ukVt�7"Oʹi���G����̩ikX�f"O�\@�G���I.
�TRh�z�"O�@`�c4*��آ��\`pV"O|=� #D� �����:LMv��q"O-9&J&T_�ePL7 H��"Ot�b@�J34'��:K��-�A"O1�rJ�!.2$U��i�v�.�@"O�D��&��ݡ�gƥ|�ɰW"O�:�lW�nht`2`��gxN {D"O���W5 ��8�e �+��T"O���� )O7���@�jz|T�"OF,�L�5%�~��F`օ1wx ��"O��a7!��.ծ�fO\�g011"O� $���%%
���iᤋ$?yTв"OLRg�\�+�y �)G�=]*�ӱ"O���L�5I��9��(��<Ph0�"O8yk!���)�J�:Db�+�2x�"O*`��e�lJ<�q���!K�����"Oz�av,�� vN��o��r�"�w"O���W��\�Bq)���1��`�""O��`IZ�Mh�ڦ�ƴiW�|C�"O�%��$�>6Ac#��A%bP�"O�}��Ƚg$:�D�
:	x�@"O��k�kʱ2 A�u�Y:6�N���"O*��T/��p�  �2�K�����"O<pHpċ��u�0ퟆ9M��qQ"O�Q;���"]h
@:b-�mC�t�U"O&t�/ߨ�2��+1@�9�e"O~<�����*d�2�+'W�:�"O"���\�>��uc+,�lZs"O�<s��SD��CE����"O��Y���
A8�i�!� ���"�"O����[h^�Ғ��n�|(�b"O�@jsO��zUd��E�<����f"O��0�P7M�V�	F�(F��"O�&8�!)@$]�&�J��R"O���GΏ�+*�]�g�]�s{����"Or0P�&%�{$�"-4�I�"O�X7Q�4�l���?3 �RR"O� U�Z�kМ1j���j�AF"Of`���L��A�"��2w�����"O�X�A�)y���!�M�� "O&�F�x(qP7�U�R���"O���@��U�� ��0H��7"O�@��ߢ5���B�D�z���"O�yxqڎm��%��cH�� @��"O��� (UJCN�'|�pA�"OZ�eߵE�,$�ʫ
q�}�"OB�ؒ��a2����O�b�X�C"O*���M�)${�{pb�9,:�(F"Ov4{�*L��0�@^$n�s"OX	ch0,..��ϊ�!��)95"O���G���&u�p�6�U��y�Y�7����`ċ�f2)2q�B��y�"��XZ��	Pf�(�n r���y�f�%"�����)U�'��Q����yrh .o@<��!\!����`!��yr!�01�����K�����DѦ�yBH��%���Ť��,����'�3�y�)�
�5ӔR p�(b��"�y�f�Nh~�p�F�0a�ɠHI$�yb�V=+2��@ɚ�q:�$���y��0Y@�A���iـ� vf	)�y��ؿO� �ݺo����%`J��y�U������G*n���r%*O��y�̀/�`�3�U$k:�mb�L�yr�����Æ��z���Iԇ��y2���#���I\wj$�b'��yB��Q�D؊a�E6&7�M�R�Q�y���13�P�i �V	$@�I"�=�yB*vOb�Dk�/S�CB�L��y��0Tf~�h��͵O�����ާ�y��S0{���R�H�1նL�AMP�y��ٰJ�F3"��U�֬��R��yR�G#X"<�'̉�b�6m�%B�=�y�n���0���i<By�4����y�"\�&����gE�93�8�y
� �8��ß�Ti\�Q�΄�
uri�3"O&M�3��>��@���s��*4"O�4+Γc��$�U�	!
e��94"O��T
@�oN���H�=6�1��"O��8��*��S���/e*6x���'�'���'y��'���',��'#��
�*i���"��
M ��Jr�'���'���'e2�'���'(��'�r}Hq�?'�Da�A�#�����'���';R�'|��'��'��'�.e�˔a�Z�W͚��8���'db�'���'��'�2�'�2�'j&l��B�i�8����P9���:t�'��'��'���'���'���'���(P�<]Q���V�J�,�0q�'���'��'���'G2�'��'��� 2�Rx�hX� �ͤqcT�'�R�'7��'���'N��'���'�H�3�͍v�L��L�O�8���'���'���'�b�'���'Er�'͌}8F/C$R��ABX��hr��'��'���'\��'�"�'��'"�bW�0_�@qc�I<j["��'�"�'���'*��'I�'Qr�'�n��B�&U�A���o���w�'��'�R�'0�'c��'��'*�hI�0d`2��h7m�L�"�'���'���'���'vr�'���'�D�@�!�j�|F
Y��Q��'gr�'���'�"�'��!yӰ���OJU�����-���Tֽ1g|�+��EyR�'��)�3?�q�i
n�i�*D�x24�P z������d���N�i>����SѶ]�0��ҥi�H```���Ms����<޴����.c[���Wl�5��6�^;b�,T�c E�Ͳb���	syb�ӠI�B�N ;�xli���68~��ݴ[���<�'��'z��w.��J��{�|���B>Q>�J��Of6�b�P���'��%8�4�yBG�X�>�y�IT)U#���"X��yr�C/D�H��w�: ў�Sݟ��W��GQr���AA�sX���$�l�t�'��'>^7m��91O
p��◭\A�(h� �9�-z6��O|�O�p�'���i��ĳ>a�υ�*���(Q�{(�=��D{~�nQO'\Ѡs����OrP�1��4���7������\� u2�ݖ!�>��'U�֟"~�7�h] B�Կ}�}:�Ҵ+����1t�����������r�i>}�㉸��q)�4?��m����@��ͦ�I���m|~�͏q���H��ȃ'�z1#�o0�(A�k�;O��:GjY.�z�'�$�㳣�g�g�-�i�e�T-r�t�F��z�B�I^�4�r� ��	۔��#`�|��@����)p�\
�,�6�I!��Q�t,b�Ψ�P��b�h���p�E�y���
�+.1�l���0I!��y�G�	��E˓t�xsԣ[�Mi,�q`�=i�̩v�:]	��UD�~�*�p�+́1v�,�b`�k�uY���J�*��`K�)� 6M�O��$�O����D~���:s��$X!��>�H�2 M�����O�H�0!6�I�?�	Ɵ�3���5Q&H����Ͱ8�@(�+���M� !�
���'��'��$,#�4��Z�H\�$[ꉠr(_�E4�I��Eۦ��e	}����'���'��Ò�\>r=`t�J�.��;���:���O��ư4��'���՟�	'r�1�lY�P�\�@�̂_[��{�4�?����?��ފx���ן���ҟp��su��b�W?WMz郳�D�&@��ܴ�?I��,s�'���'ɧ5v�֍?�R���쀖,��AQq���M��
:�����?���?q�����OF5(&gS�hB�S�ji���w�Rl&���������S����i�N����d�JP�B��$ˮb����՟��	Oyb�J1M���%im����a��5��]�@BO��$�D�O��Ĕ�@��	�B���7l�C^�M�f��+~^��?���?Q(O�9���zⓁx�R��q+�?r�HB��=f2,�ܴ�?q�����?q5�M[��9)t�*peka偾�L��2ks�6���O��$�)�f��d�'��d��z�Ʈ#
����(Ȋ=
O���O	�#��O����O�OrQS��1R)�ѳ����	��	۴�?1��D� p�ih���?	�'[��7d� �Bg�s3ȍ9���kH�ꓺ?a@�����'2�L<)�gē]x�+d�׸RՀ���%�զ���,�M+���?)�����x�O ���pOʬdI@��a�q�p�P�dv�D����Oz�$�O������ʧ��)��*�@Q���>"�|��a��04�l���	[��fyʟL�'�Xq�7��b�"D��V���JI<��<?�����'�����|�Kwl�%�a �+�K��F�'5�$�4P�4z���⟰ � �%�6*�F�|,xl��M���'�@9*N>���?I���$�7�` �VD�l�8k�lϣ/��,R��B��ߟ����L�'~"�'���`êL�I��QzC��5"�P슁.�<5��Z���I����	ky2d� �Ӫv�|�H6�WS�\�)�$�%�&듋?I��?�,O,��O�Y3A��O������,�ZA0v%�F��+�Nd�柴��Fy�`�,A��Ri�#�&���a�a�)fM Lӱ�Lަ��ߟ�'g�'0pSQ�'=�Em���e`G6�J��Pi�-��m���\�	iyb�17��R�D�k���C��՚u{]��L^�\�z�CH<�.O��!���O�����3� |��@,ԉ/�0gɠa~�%s��x��Z�� ���)��� ���=�����ە_�0B��(m� ic1�R8�J��a��-4>����Q5���`)V	0�yxb/}�D�C`	���e�2c��1N@rG�րHr�$R�i��������
�"�)g�C?3��lp��X.���@ѫ��d*`D�l�	���`�� �R���	n "���M�0?���
S�V<@��)�'�S�� @E�rI�Iן��Iğ�[w^�'P��1�ަO�x��%ġ&2D����OL����=0��*�O������Z�,I�a�;eK�hs�jCeP����t
~	�2����d>Y@�z��/'��@��0�d������D��%��A9��z��OVUu�'���|R�'��]��1ҥ"*�T�#�=�H���<D�,9���0h�����C�db�"�& -�HO��By� =W�7�B�E-^�s��\<�1� ݧ8�:���O ���O8x�/�Ot�~>�H�&��7��<YU��S>��D��3 8�Ks�E��ЅYv�ĘO �F2�@%$�"�;t`�H��4�ToE�	���޹�r���|�VD�#�	�z�����O4Cd�_���cun{���I��(���O���+�)�����"�����e�); ��+�b�<�c(ڷ,�>9�NI�d�H��0N��<1%�i�_�� �ɘ�����OJ�'=�d��b�0Oc�M)��'� ��r�O;�?q���?�"��4$}~������~Ԝ�FI�>7r,P�A+C��<�Gf�L�sŋV<G�\as��f��S2O$r��f��~Ř5��� >�ģ<�I����c�4hس!\0D!l� �u�B=O����O�fX�1�ǂO�t�9�#b�a|R,2��N}*iɳ#�' ��ͩ�����B�0)�x�'�rR>�s�����	ߟ|�U�M�B�� �3R^�g�ϳ{���е�X�+�V�1�H�H:0<�Oe1�B�Z��$�Ӊ�(_���y�Ç8�*�@�Ȅ	���V�ΎCW�x�Xw+�S�N/8ʶ�
q`�|�]�?~hxX��M/�=]�p�kL%<}h �	��M{fT������<A㈚�~s�ق����6IȰ�_S�<�ԀK/K��ӄN۬H
myw��N�'0#=y�i�҃ G��s�*~�@��S�o2�B�I*Y�Y�I�f��%�Ǉ�=~��B�	)),ijb��}��9"��fB�ɭ���3`A*C���t�O�}�nB�	!20*�k�O���5�SG-Q�B�� FjŠ�G�[���S��ۖ2АB�I�Fi�E�r�<=|N@j�iF�K�,B�Is�&e��c^+d+,��6�I��B��T`� HR�����qa�T��C�ɰD��Ḳ*��N�����z�C�I���<���M�(��YF�
Q�DC�I�&�R3��u�h�P�d�&ks,C�ɉ5�>E��W�,�v3�+ˬ[�4B�		9��4���� � h�,�NC䉅
L �T�`>�y����:�~C�I	m6���!ԡȠճ����eqHC�)X�j���/�K�ʔ���
3AQ�B䉨[8�*��J9�t��IrH�B�ɀ\�+������*^?C��/�lC�k&KG��`��]��C��3m����'�Z�c�d�P��>ְB��3Zw����.A6�jD��a�jTrB��W�Ѩ�#R�k�0QdAK�7�:B�	[ؐP�ω[Z����4f0B�4�����2"Af��DĊni�C��8^���;���W���a+C��C��	o�$ I� :�b��ǈ)�C�>V�����jJ�4��H�@D�b�C�I��,��8�� �E� ,~�RC�	�<"}�HA�����&Y.d�*C�	���x23��:�NE{d��0��B�	 _` ���G�?UN9�s�T�I�"C��/Uu�1���B,|�0�g��~�C�I�_ls%UZ�HiȳT�9~�C�I0ZE (#���0�<�y����4�C��*�s�J3 } �3�	:&��>!Ԣ��H�{��Z��� .�^�#����y
� x�Iģ�,5���굡Y 1�f�=Oz�P�!��������Pu���@x��� �"�`��T"O�u��oU����H%Ό�*���8�E��L��z�E�
��%ɲ���Fi��녯���0?�S��8�
T𢤕3!�j�C�v��u�`�<�5�\.�rM0v���l�@����D��'{Yڀ�1��)I7���#�C�IF�S�4APcb����,h�<dpF���y�j�#�н)Ph[�3,Z|��=.��9�ͻb��:O>��X�� �
x����i��#QHZ.^èL�g
+h�!���)����4$[:�V��g��+>D��Z� Y�K�QZr��%
/�0˒�>ʓ1q�U��hґi���	��� ?T��H���e�"DبX+*���vs����@��)��IG)9!LNXb3Oغ:��|N@��6�7p�Ƥ��ߑ��dP'.`��Ks�c�@���C�����Ċ�i\�]1!#�`D�쩑�Ɗ�y�T�����FA�I�6\�3	 /�H� "�/���=�O6]�7:�y7Ô�]���tc�9s,�)b�uEC��,�v�r�KՉ~Y^mZ)F_p 1��$?ٲJ�l~`b0jE)Nz�8�';ʓn*P�Pb΁�lCf��`͎$w�L@��23�le6C�&+�$� aJu�L�H`Q�z0as6�ٶ+yꈨS�Ϊ�䛥'��|�	[�1B���$�c����e���DY<G�����et4`�7jZ��������=j��"s��X�̡i��G��y��/om,�7��^���e�1z����	���=�O��m��ywk�m=��iS�^�Y�HU���D�xrc�-7��s��&P)0��rAIh*r<��O�aqE隢L�T�z���9��È�DFkbS�t:��1�+rAax"Ȉ�m Xɢ��i�ܐ$/�1\z,�f+�<A����AR�a�`h�ƭע.6�� `8�4�w7�(�b��J��Y�@ -?A�hǵn�	��i�l\�ȕȺ�O�'��xc��[1��C#�Qt�C�ɀ3:a�L�;Q�L��E8	X�	�Q���D�.�T ���Šs��g}���5����R���a�T�/%���!�'��4��
�:�Ɓ��V���ɨ5�ނ9��p��`�n����|~*��c�P�U�B6���C+4ZDJ�%%�������7��7�F0k�{}��w& в�ȨO\t�
s�%דu6p�E�)V�z�ѢH�0����'�L���ßv�S�� V�*�����U)Y��i�m�5��y5���"C�I8�M2ro�Y,���>P"ZO�Y4e�+=�D�
㧇�	��O���	x���P��(��AagL���)D���1T�^�y��rr���B~��#�F������j��)�/�B��ԟZ8�d����:-���028�}�Sc�-5 ���ku��8u@�D_�-6�⡳i���C��]�T�C��ӳ~M��	�C˟0�CD�8<��	#��A�H� �� XE=>�����@�
jh���	,c=�@�u�:���0k��/D�!#��O}|� �g"O�($�M�
0���ҰA������2 2�E���S?��'J��O7>\2�Μ_��]�E�PI�s)۴8�)��H'����DF�N��`w	
+`���h��m��* ��d?�'�d
���3��\��� kd=؉{�K�k���iF�n��0�`)F��Ox\)�L�5�Zt���&�bA�!�i2�=q���'�����،�1�#k�7��{6f�1ji�̆�	Htb)r��ͮA�$��c(ư�t�v4/�=\{A1��z1����~�Ob!�����n�~�YAL	h䁄�*D�T� U"P�J�� �V�H��U���T%2P$ ��D8�~r�O<�韠�Ǖ
|��̻�aBTo.�.9����:2x��ɞH��`�`b�F}H��VU�LT��͏�?d<OnTR!�T_�7��&�u��S���'v&|Qfa��+��41dL�h��KSD\����O�ErDc@'{��))L���t�sq`^�v�3�lL�b@��DGW����Z��y
�a�(Ww&�q�o��i���'.�Mb� �1�ҁaE�F�:M�{���(LK2��dw�T��Oԛ�j���m��1�F��&?��ՃڸL�X��b�3a�j�kq�S�ģ�1��0�w=0��5
�mFx]�Q�ĳR��	�'�0����A!v���rHE=l%�d��L���:XJ�$ቢc09*���Z��t���e% �5ȖZƬ�yѩ��0<�U ��6��0b-ޫ����Vk�+a��X�Z�t�4�����#AP�nެ5���JE)��=��T
L|5�s�'r������Pt~"�DdpE�(1��H�a������@�Ώ���}�D��E��!�>�h���iR ie�,ؔs��F.&�RF|H�L;7��1~Sh�g}r֟� F�BN QtQ����N5�`�$
O��S�NƘe�a�2G�<b��r!k'tld�YR�m��1$nM~��O�a�k	vL��	�(>���1�'\�Ț��/��<hF��3W�� x�j̝�Ɂ�'ø��e�V;7����ú
L!�����vh"}*BK3�����kX	v^&1@��[�<3��,(A�����:sV�S�F^�<1a̍.C��"��C�m��l۔$�X�<����4k��4���A���0�z�<�����M\��ʱnӕg�)#o�q�<�+��ް�:�Ĕ/0�=a��	m�<!E�1{�y���\�U������D^�<�K_�M`���C�Iܮ�+���V�<�',�?R<�����9ό]k���S�<q�/�^%aS��O�b����Vw�<�g�K�0�#�R��%�@L�t�<��Ȗ�FR���4bR�:��a"��x�<iUk�5�h\+�7X:��لiQt�<���	 H��!1��/s����J�z�<����zVii�I�������z�<���b�\� 	�\D��u��o�<y��
�V��dс���Z�)����i�<)��5D��2WO�0MP�i����b�<��j�����Ái����E�'œ]�<yP�!Q� �C�� �$ѓl
W�<)T$�8,���`�hk�!�V�<y���D��S��R�ow>�x�@U�<�����w�]B��B7{0
 B*�x�<q6�+c��X���'lMÐA�n�<�ƪǧUʲ�q�l������n�<�E&%L����U�z�F��m�<V�Ź�2@���E�Da@q�<)���(ۖ�{� ǚ�5i'@�i�<�k�#-E��	t&͘M��-�P�Z�<���NB�@݋��[�L�I"a,�U�<�4�P�j!(�s��(fڜ��GQ�<�d��2>��黃�#�Z���!�P�<9�À,Y�60s.��3��S��CU�<I��C�)�ڵ�vi��Eru���X�<��l&���'Z�s����	n�<A��0*AHi�Ǒ��^�"WA�j�<Q�dYx�tc��z�̽�&�Bg�<�A�d.(Z/ʉ!kF���Z�<�w��N|�����ńM�P���EX�<���� �S��;<�JD����h�<��)T@�p+	�)��q#�e�<�cN�m�0* oC6W�*0���Hd�<�NU�[� ��F�Da��BnX�<Q�g�fMpSÞ%E��2��^�<�&�+ k��@�c�d�du2��Q�<�f�}N���a�P
 ���z���Q�<	�Eڼo�����	B�(����O�<�&��i (�:� 6���c*M�<��eیl�n�p�-N=&�(��p�<���I.V����5&+� ���c�<1A#�g��x�a�B�Ha� e�<����=X�����b��d�`�<���9�>�v�4v�-(UL8�ȓ�DqҤ�rlz���G����m��0�
���o�	x�t�*��$a|��@(Na��(�Q�2�Ȣ�̛{`�D�ȓ��"����|5�l��.[�E�ņȓ;�88�ဒNCЁc�ӧ*|8��ȓf�D;���$Ĩ��Ԟh4�9��S�? Fĺ"�W�:�� ЀQ�NOd���"O
Ij&��=G$�Ii�f�[T|XF"O*x1�]�|g��aҮȄMc(�"OV���H:>@�a��P?���A"O�e�e�=kB�Ѣ+P^'��+�*O<�"0�ݗ�൪��߲�
��'�<�qׄ�91�T��J�0>ꖙ��'1��K���7[N�ICtM��=i�@�'*�pXQo��D�Za@u���X�'�Z��G��U�%�I��T^x�x�'>�����=�p���@�)x&��	�';� U��]36xA�� o>���'�,ܑ� �	(tq�c��i�D(�'E�� � Jm��X�BE�Z�8��'��u�悈2c>��jg�.�z���'�֤[U)��}h` �Jڕ1=h��
�' ��3h� BJ���L2:�� 
�'̖(6�Z�]F���F	�.�D�	�'x����&$��[FhЯ*ܺ�S�'�n ���	�|F~qN�?*h��'�ne�De�W����*m6���'K� �U�ןY ��R߼v&�r�'�>��UM<uW�X�"T0q���Y�'WX�$�/�� Aacŏ3�z��
�'m6  ��	 $9�ʂ�'�T�	�'�B��O��)G�u�M@r����	�'��]���ݎ|�f��VjG�j�� Z	�'�I m���:�#��ُi���'`RDx&���#<�h�G
h�����'8T
�ŝ6�p���J�b�  �'>����H�#,�\@�+��r5��'r�
��M�.`p���F��D��'�����R#ެ16����
�'���q0 �/E�*B��EW�1�'�vTs�����"E�� xk�E�
�'���X���n�.��d�L�h����'m�}��'e۲X8A_ D�8�'�"�lT3{��3�G�(ZZ��G"O��`wJ��f��%��/Q<޽�"Od��2�69u��۵�CBIQ�"O��w��]����煷~� ��"O������"��� Ƈs���ۃ"OPDړE�1�:Y;��A"p���"Ojd ���	
t�q��.P`c�a"O��W��{��y� �M x���"Ob"B��	{Pz���9:���CG"O ���MG'
��a�Q�<�4�P"O�X�A%P���-Ş\��SU"O����$��y\�����]6{��=�"OH�y2�
(Net�XC�� ��A��"O������e�4��5cHIXh�+S"O ��"���|"�G$R��`�"O�Qz���Y�I��O��1)!"O��ె%`r@G�q �� "O��uSk�FUA��V�G��D�R"Ov-RG*P�uvx�����n����V"O� 2&�	it,�ӋS��q��"OJX�����fߐ���ᄂ<v䘈a"OإP����H ����	m��c"O�K�g@�r�`)����4X�=��"O�ʀGG�<Y�ZP�E�mJ4ݒw"O�u�&/ǀ6!���ت|�ر�"O�hBUn/+�t�2��1�8\�"Ox!i�5�0��,I�X�is"O�  ��q/ή{�\���I�d��EC�"O�b�-�F�z�3>�8�H�"O�3b�ҶN�D���Gˊ>�R��"O���C�4NQ�UR�����dɓ"O���!�L�B��)>p$�b3"Od�A�
�{x�̙�2�
첅"O���M��������"O���"��YKVq�D�;S�Q9r"OԈ+֗@[�\�s��<���"Ob�!�HB@V�M;S��3�����'8^Tʴ����y��['o%v8�	�'� �(�
n�>q!�]�7
��'6�e�f�8}N�E�#�D,�":�'p�h9�JXj2�ask�Bq	�'����a��͢D��fY(}��ܻ�'��d�L�ۀLr�BM�{3��1�'Ul�Q�]�2��8I2K����'����lX0����h���`�^�<Q􂂺ox>��b���K&�\y��N]��hO�O��U�b.R���ې��+Gv���'hp)	�hG���������P��'�r	�Beԇز�!��P���
�'(��ۆf�*&��y �aK�\�4�'8��r��R��� �!At��	�'�
��7�H5yw���ꑚ�8�'xD4�K�i�"���mV�Z���'NR%ɱDO�K4t��ܨ9�X�'�Ĭ��� =�$�y�`	�M�
�'�Х*fGZ:3�۳!��14�����'���yN3X(i�6��w6F-k�'��$��䀨�
b�M�/�ȡ�'̌��V�B���"�jB K�'��ͺ#�ϊ#,�!�DU�+b$�'�n=�� �&���A"S�'
�|��'����B����:4mA�j�us�'��!6��)��8Ӥ׵0a���
�'�$Ȃ�Ir��@�ȬS�n}1
�'�B�Aá��.]j��R�ԚM�~ �']�!24�_� 7�=`W�HZ��	�'�d(C�Ƀ�B�����A;�(�`	�'Z(u�K�~K�.>���'���Z��Կ>F��i�Z� ���j�'!�Y�JW�FXd�!V�Nl�P��'��xoJ	W[2�+�M�` ���'���BK�6V��e�?^L�
�'�@�x��-�q�wi�0gX� �
�'���K¼0�F���i��Xj�-
�'����r(� "�N�k�mM0b5x���'�v�c%bì$٬`���C�SI���	�'L6����J���B�X3Wn^l8	�'����&��:|�)�eG%WB���'I���Өة�`�Wޮ�Q�'g��U���`���H�O�����'��	�'��6d*�q�Ȝ0ܖ��	�'��@�u��B��xe�	A	�'v�#1�!k΁r�#��Y�>HR�'r�(&��;�P���-� xVE�
�'	l̓Ԫ����\"�E ��%�	�'���P�#W(~$I������m!	�'�`�[�eO	���B���3)��'(�� /-�Ј�0�r�'UN1��I��m�1�,�LU�'���K�])��Sp%���p)rf����'��{�,�J�(�E��m��#3b)�y
� z�0Ac�tf�X`L�����f"O�@��T�+�B���վg؆�0�"O�P �.N�4 �6D*h���zA"O�@r ϵXN}�IE�>�`u�S"O�\!�,�y�����;N��}S0"O��I �N*a,�m��DM��I��"O�I���h�`�!�j�5��<p@�'Y�$D�0� �V	�W��D�rK�2!���#��2�h�
��3%],x0!��L�'�@) ����{e�����/�!�[>�(@�3�ӵ[]0���+��.�!���Xۘ 8v��!o�<��+ ,Dh!��ƻ=?h�8�#�MaF�pbh�Z�!����r�EfU�옖g�$;�!�<��=����_&�$�v̉{b!�$�7
Jh1õJC�3 �T�`���.5!�� �l�{1&�{,����1�!��;F�č�w�<x�Q�ME�{I!��J4	�f%ꇥ��<X�-�;1!��Ѭ<JL
��P�s��%�
3 !��2�D�R������lY
Oh!�$N�u,92ׂ_S�050�.�O!򄟼c���1�O�ɬ�C#H�D!�H%,��P��1͒�C_��!�DR3 Ȇm'�l�����/_'�Pyr�#-8"�\�R�8��̐�y��E���(2/@a���f"���y"�����d#� �>Gg��f�H(�y�%:Һ�J�ӽ�ǣ)u�1��'�N�����Yaب$*Ϝ �ti2�'��(jƉE�!q2�mϮ�{�B�PK��!���B.��)��� hz�B�M��D��I�1,��bV��$6�|B�I���Xc�̈{҈�9�,B�	�T��(�5LՒKXlc��܄&�B�	O%J��$��58�`��V?~�C䉈��Sb⃛���y�/�/@b�B�I�V�@U q&�#�5�4��_-�C�I5}:B!��/?�X���+#(pC�I.2���� �p5d�� ,C.Z8C�	)6u���s�!'�P�j����C��%s�(Zg�Dwq0�q �3~�C�	���i�{�&����x�C�I�
��4 U���84 AH��8T�C�!Hl1� �\�p��d��I�.��C䉦B 嘰�N6��"�J$(@C�I%z ��E�I��h����k��B�I�[3���2�Sz���Z�dH~z�C�	2.�!v�7D�<rg�J�L��C�	0	��5�%�9�p$���	�-+�C�IMZ4[Ѵ\��I3u�G�U��C��T��jBB_�dŊER�=fC^C����)���t�PY�c�VC�I=���5�.kh�C��K�p7�C�I�n�� ��i\�ق���-)!�$ l��pR�k%�\H���1}]!��

R�(P���>D�`����!�Ĉ%%H`�TQ���p!���1�!���UiL	��
>g+�d���+Bz!���A"�c a�!=6��U&K7\!���=?��dyׁ�v��QT��HE!�D�%I�v�2� <5��`��e�+rR!�DOZ/���I��$�L��B?o9!��,��do�%fOt����=A�!�� Tܩ�	�)�R(����\x�t�"Otm�Tj�$bN�趌�
]z���"O��������
��!V�@�i"O�(W""P< �rE���ѐG"Ob�	#țP�4p@0��"lxp2�"Op���L�����Y����`�"OdSr��8c,ػ��߮I����"Ox[�ψ�8�<�C���+���S"O��Ff�[�(��"Ǜ#�0]�%"O��R�j��4����!Q�4�+�"O�����K�/�!x����Tve� "OR�{�i�^�0�(2GZ�h��1"O��y�.A�+�0����s����"O��@�Q�n��eϛ�8X
�h�"O�WJ��;��`��R�p��{�"ON�`�mN�8��$��,�9���E"O�T��X.e�6������y ��"O��p�čK�<02P�5l�X�"OF��+R�h�FA��O�
dM*�"O�M�d�6#�r�ф��,R� �р"O��h1e\7J8l��� �$�"O|���D��X�1C$Ӧ*�Z=�"OD����
�F���CQl�mw"OJ �g�	(&��q�h #s��p�"O޼A�,�X��lH

5��T
�"O"U۰�B�T2���(�	{�r�c"OP0 ��>U	0����M6�Q9"O@e#"�N:��s!��E�R<1c"O*�3G��mr���↷#3�lH�"OJp�p��P�
�l)��>u���"On8���ѐ(D:�,b�!y5"O"Xq�
C�Ě���*
 ^��%"O��gE_����4)��y&"Ol��L
	�H%�P�:#����"OhA��؞v��`���x2��"OP�*� �_C*�"`�%��"O�1#�� m���kૐ�����"O�-�Ʈ3|"��i�ZlP�"On�Ѥm�#��C�q�����"O�I� ά2	(|J���H���"OP��V+�2U¢@���;�����"Oȍ[���2D`����?��m{�"O�Xi$�N>���6��;<j�"ON�0'���fq�キq �$X�"O�ؠ7Ig�4��UqҞ]˦"Oh��$�Ѵ5��M���&�)y�"OĤ��n\8,�<!7��j�zQD"O���F��Xv\:4��9!V��"O,��P�U0�04G�28��F"Oh���3�Z��Ƃ��,��"O
��4�ڪ0y�$
4��o�ʤ@�"O�a��C��t6H�V�7��� �"O�M�r�M�>�`)3��5�@}��"O@�PtG�`��M0��N� �"\j�"OZ���N�Bgn�:��Mu�8�"O��"��]$�JE���N?r�ԫT"ObC��
4��a�%B ~�T�"O�𛤣̚S֐U��e�2.l�"O�B�L�a�<e��%�b&��"O.股9n�����.�%t�="�"O�)S�)�T��Ǝ�=*LxRu"O�Ah�å^q���mW�

V@ۦ"O�$ɴ#Tk�d�1V��3�.�г"O�h�2�M�\a�5�e+�Q��<8�"O� ���,8Kg`T8gj�;R�R���"O MRԮ
(�ĳDɔ�J���A�"OLqr��Ir��p/M�n��Ph�"O��2PN4V!p%(��O�i�Y�"O�iR�O;A����Ä%�F"O��#�鍡	�Y�G"�J�T�#�"O��YC��i:����"�B����#"O>��b�Q�-B�-[���!~�|�:�"O:|���������L� �+D"O�XG��=p0Ը�a`)<�Dc7"O�˅�Κ5���7i^�ob� "O�ػ�(�;��4#��)p�8h��"O ر�+@%<z���A�;|��
 "Oi���g��-��*[�\_� "O�(
�n
3k�6A���E1�P��"OR�z�K�*O��d��bF�?M�l)�"O�@������:��W���_[�`�"O�(�^�n�2�s���;�l���"OjTb�%��Ѣ�AN�`���"ON�9�ы,��)��lθi+�"Oޔ��gː�숙��N�.�" "O���-��Ie���)uL�2"OH������$i6fO�oH��t"Or��o���qRB�%b'(�	1"O�y)�`�=C�:q���wi��a�"OL�jD�V�@��	(0����2"O�3Ƃ�5�����c��?�U��"Ox��Ȑw�F(�B	�(�9"O"Th5
š%@z�ې��=�@T�P"OR��UT=U���̞/���"OLL��l�;"��9��EA�L��F"OҝpOE78��K<u���d"O4��W�ǀ�:�Y
�"O��#ԃ5���q E�/�VD�"O�0y�^�{��A�A���"�n`�'��*.�搬�J�+B���'�4��,	�K�D�C��!d�<���'ޞ�$DI�r���r�Ѝ`��\:�'Kީ@�I]�j��	��!^ذh�'��xS� G��$s��/ZF*��'�n���愱:�% \'�mS�'��8�#�ע�;T�\>M��'�nũtm�79���� �(\��Q��'��ҵ%۞b�mЃ̛��=��'���#�L��D�#��6�rH�'Y��3�a�~��g q����'���ǃ�<�3�ߣp�zA��'72�BE��x��H
�gK�m-n(��'! ����J�2,�s�_�h4$���'��I��ꍋ([�c醽ao�H�
�':�J��R�?���BT#U*�J�'�1A��,ǔMiF��x�'� ��J�d��g�+(J��
�'ZHp�.L�Z#0�����%�h�X
�'��I��I��wN�AO�6R�š�'�ƌ��@g�����V�R�z���'�Z5SE��& Y�W"V�R�8���']�|Z��2�
 WH�wXt��'d"\/�b�:�O�>"�t�h
�'�*2�O�	�P�R0�=ζ��'� �w�͵VS��bb���|x�'A��U��>~�0)R�7��0i�'lj���Q���1��r���
�'ո$Ӥ�#6��Q�� sZ�@��� lSIġiT��8&Ç�R*�kg"O`q��_b-
(i��E�U����"O����(�?@68��ѴM2԰%"OLu*v������A�oI7DrIb"O����F�=?���Q�ҽ&?����"O�Ͱ��=k^�]iB' �ي�"O ���%�0H���t�J�z$�E�""O�)�B�֦P�Q��K��@0T"O4��c儱OA6\y
�d�$���*O ���$�1�6��j̰-��m��'v<��Q�S>� �M� �6��'�e�VcP���ɒ"��7R���'�H�Ф�V913dpQ2郸
~Z
�'Q
��ݭ.נ��M�	p�ȨZ	�'���2b���AY$��)n-��@	�'+\Uh�FU<w�l�V�=_e��A�'�z��r��'
��cu-@�N��A��'	쐓�^�H��@�㟝?|���
�'�� i�D�f��q�kB
1�HU�
�'�^9�M�O`����8��;�'�@�y��U2#'j�K����byDk�'PX�6�\�1��}�5���V�����'��4�E	M	7�>�Y�!���"�'� e���@x&U��Ĕ-�����'+�'��&	(�����(`���'3`�	�bA�G�Bi:#VS��'������3Hf����C����']0�fm�C�h}#���?�h�k�'w����L0�i��)9۠]��'��a(�M�	k��H���25�tr�' �=���W�^Td�"�oL�J)��'/l�B�B�:V-���y�y��'��I ��ӈ1�<�i��~Z�8��'�ẗ	��) �z�I��d�j�'�N<s��%h}0�!�E��B	p�'d�4�v��hL�c1b�l���'�J\[���/����ؘ$GB�Y�'3�����D�ӓ.��r�`�'+�ER�
	�@/�!�c�J�-~i��'^��z�'E6Y��\)V�V�y��J�'�"�b��1��]ڐ�*h~���'�L�c�?o�&�[0/�8��!"	�']���aU2w�rI{�Jߚ�1"�'�bT�3ㅞ.LDyK'(�P�  ��'�d��$5���g�L6Bn�3�'�����01�([��͋5wF�Z�'Q��B��	fxI�AJ-ni�'r�)z�X2f�ļRĄ�$X�3�'�00aII;cRl�K�.�-�J���'���@"�}Nr��b��u���'�\��&䑒V��"�^���LH
�'a�@IU���h7�Vb�R	�'F��q�� �a���*�ñQ��	0�'m���i��9� Y{v���B��
�'�"�K�+�Sf�d�
�&A����'y� 1��tӪ1��ߥi$(���'[�+�.\�>C��w ��c��Y�'N����/�>�4<��C�*M^���'�ʽ�g���6��` t��*"X��'���PU�
�J�0ٹvBϤ*��%��'�x-ɇK�%�V\06�X&/�`0�'4.@ɓ���%�>����" ��'v����6AT���L��FEY�'��`���V�v춤e�f�,l:��� <EPu��=
�5a��T'�%��"Oj=����F���r�[1
�L�U"O8�7�LG���ՠ� k�&��"O�TZW*?J�h+�H��<-p�"O��T��m����f��f|xr""O(�a��xpT���ϟ� ���%"O�0�6Ξ#@�c��Gg�I�"OzL�p�=g�V�{W`��bK�Ѡ"O�e����'x�*A8�iI�I���0F"O\BT�1�%0�!��J�{"O(Y�MK-�~RP΍%=��D2"O�9�2��7@B���@D�)w]�yJ@"O�$��XY`�ac��KM^���"O���́�t�nu�t!�&5\�p��"OP����-|$D!��D�Vu��"Ov,��R7B�*p@�ǝ	���B"Of !�Qh�@!�i9Z��Y�"O"i��&הAe�p(P�j�%"OF���l��'J�8�!�%L �h "O� ��dI�+�^��b��96 ���"O�	H�T:���0���w!�*O(L��C83�h��amY�E��h)�'5��;@�A>"�Fab�ƕ�N{\i�'�R���X1,��U�@��Fyj��'�
�3�ED	P� y�%МS�]:
�'kl`��e�W�����T�QP����'/v��%��7,0�QH���H��II�''nͫ�᚜Gh�W��P�D9#�'Dq�K=���h�@�/~1H)h�'�����鋀	Fmce�
/J�
|:�'3�q�̖H��i:�nFĲ� �'>�PY��K274�T���!A[`���'J���%���d档RG֢c\�r�'=Fq��/��S���Rd��yֽ��'!��C�@#	W���cE��=�2B�	�'M&�A6ŏ;��{�Gʋ��B�H\	٧A��.�8p �	5K��B��V�N�:��Q#.C�0�%%F�of�B�	�3dP拣h1$Ԃ�N�u �C�I�;RLE�e�9M-�i�1�Z�7p�C�3��`Y @H�i���X=�C�ɘn�T|q�FPQX� 1��Q�RB�I.���Ы�$1���R��ɖI}�C�	.K�x#� ���0/�	%��C�ɦ}�Fy��ƬX0�{@i�x��B�	U3H`y���hX��� �O�jC�I(ȡ����/4LT�q�4iRC�ɯgU��+�j̹z�h���C�C��u\�h�lJ5D��/ibC�I2=��*҇�.gD�3���B�-, �\@�-U��ԥ1��"V��B�ɔe,^��
�-'ض�q�ܸd�B�I�`�E�ElV�J�r�z�Z;H��C�	�W���"�'�-h���?�C�	 Sx�XŅ����s��3ec�C�	/Ѥ@��F�b��q��Kҋ vB�ɵS�.����5�Q
d$��,C䉱,P�eW�4y��c4㐧a��B䉑Q
,}aPN;\!�9Ч�P�0*B��I��Q���ڙP=`eA�D�t\�C�	W��e����|���V�I2c�C�	h���s"�Qz��Щ�aǕ�dC�	 LAZ�OՆ<ʼ�3��Z�^C�I�Ms��z�����1p��ukJC�)� ��K��M�1��'Ң�p�"O��Sb
�$��� ��4li�H�'"O�*�c� M{���Ն%e�EIr"O�1i��
��v�"�χE}�(p�"Ov)��
şYŜݰ礜���"O�1:�I�[�Z����ݲD�H"�"O�e9.0*`���!
'�A¦"O~(�$�ӄ@EN,BD���Ƶ)�"O��[5�[�E��9�0��9U��0*O���A�W2�:i��F�����'h��k�ŉ�U ^	���8���'��qSBϒ�D�z���.F
Da�'��	;�e �]#<�j.6+Fvy�	�'���� �����#��9�,H��'eVA����AFH��Q�O�AH�
�'�<�-��'��q@�!7L4-R�'��1����/#���ŋ�/�!�'���Q�Y�=ΐ1����,�Ή9�'2aA�c׉Ps�ph�m�z�z���'�n��`���yb· �U��'A2��L?"Q.���e��f|	�
�'? D裀ݿ0K�s!�P��9
�'�,5�`�Z�n���"��Zn�-k�'M�쐱lX�,`��Dŀ2K�&��
�'��q�3�l��H��D#H��U�	�'���ڄ5iآa$nՎ?����'�A�a��[1��ӏ��<t>�*�'��@ C�d
�,8S�)��1D��0���!l�� "V��h�!-D���Q�~�<!�ʏ0��4�f8D�8��
o���˥,3�Ʊ)��"D���0F��PY�`�Ǥo�z@�!�?D��kPC�ut�1�R�p�B�
U.!D����g�?~9: Y5j]�?� ���"D�̻���4��Q��+[U��+E%#D�XӲ� ����s�%ٳ�!D����@�rnJ�@$!q
���g#%D�h cTઁ�hC�����i$D�$##IS��4H�f
B2No� ��H$D�Њ��P&��K�(<�tH��=D�x�*C$���6��y��9*)D�PI���8t�ݢa���1F�<�+3D��[�F9[�L�c�۔òxH��$D�d�P����0����% �T��%D�L��#_�O-�,���Jdr�#C,%D�������D�T�'�	4�80�5�8D��@��;#��}�'�H9}�,0�o8D��ՃC$@|�\K"��Q�
���9D�؃�C=?[�.�2�΁Ss�6D� !F��5�������x��� D�X�2\<W-�� �� eJ�)�$+D�İbd[=z�đ�"jmi�9c��6D���L/P1�� ��p��6D�Tr���= �N�0�H:ْ�$3D�X����k�DR�k�Z�`1D����'I�����Jӡ(�$����:D�����$͘��aʍ%x��a K6D��r�`[6c�p#WD̬�vu+�?D� ���I϶l!3�H�uYx؈��;D��*	�) >�(��;7�dlR��7D��� �"8A��gyzP	��'D�ԃs̤��x�����a |, Ɓ D��Y�o,-z�����e|&��9D���!mO��8l���(#
a�� 8D�� ޔ�C-�	eA���H��S�q�!"OHP�B�?#���ђ��-��9p"O���M3� Ȁ%҉&��!�q"O��!���4N�8���U�(p�P"O4\���"�������̌b`"O 0�/�A��)�B*K��ڤ"O��L&l�i�aB�[+�L0�"OFY �Ē1Rb�q� [�%0-�W"O��it�ȠS�L�BB_4Q��p�"O�L �@(;��-� �I�*S���"O
�a�	M�p|.���Ǎ8yCԵ��"O��iV�^��[�U�-�b�"*O��U.�$rJ �R�*:E��
�'�R�!j[��R0�Ƃ�4ԑ�
�'�����(!`v��{�/у/5���	�'m"9�3iP75>�I���5,�H��	�' b��l(o���d ��*���'	\�s%F���4�4<�"�'O�(��N.7��hQg�	���I�"O0e��ܥz0|�P6�1V�r"OB�BtK��p�ՠ���V��"O\�g�2 ����f�ȴ`��-�c"O�ty6�#Zp�QǋF�6%�!"O��"�Gt�r0��X<��H�"O@)���QRoJ|Q6(J�StD��0"OE�D�:_�2���'��%{�ň�"O���7�Ǚ[��m�'�,0�*�{�"O������x����_?�,-+"O2����~��ݙ���7L�8e"O4��A��|I��1v߲w����"O�i�BI�F�
5K4�?*~\�"O�e��y
����x��p�"O��C`�ǋy�r���J6R�*9Y�"Oh�ABJE)s}x�+2��7}x�`�"O6y�4)Ƅ�>\����F��3�"OP�g: Mbh�/�/Vc���U"O��{'Y0Kp�q��Ȓgb� {�"O}��¼dl�@j�,�Yw��t"OС�/
SlR�
㊗@c
{s"O�e�!M�?�9�	�+vG��Q�"OZ�j���3��}귇΋v!R���"Oܬ��lJ�b��UYG,��$$�E"O��k�F�+t	���]g���A"O�3��@�XS�����i��
�"O��C� �rt���H6Jb��ɡ"O$D���8P� �A�6WX2q�"O(��3'N�QQ��D�d:!�E"O��憜4CTʹꧣ��Hf�d��"O2�1�H�dY��f�ŇqR1��"O�!�B�����
Ƙ7k6P"Oj��g$|7>��V
I�=,�*"OL�hR��.�XI��+]�_ɎM
r"OT���+Կ�h��l��"Ol�sqA)�Y��j�&)�2�("OP|i�'O��LiW)W
^{4�!"O��[!��.]���R��wx��t"O��QB��H�IY�J��K���"O�a���ڌ>�
\����*b9�R"On0*� � ���9b!Q�f��!"O��إ�ǵ	n���"z����"O.h�r¾J�����ܪR��@�!*O�`p��@�`�fU��Q7|�4|�'�fhґ���&:�H�Rf�%i�j	�'* �
f�,*�`����d�|9B��� "E{�� s��y3d�D�s�~�3�"O�i��]�v!kGI�'��S�"O��`�$շ<z%h��ҹ?�0Lp"O��@�LS�<��'���8�ʹ
�"ODha���bعE�Pd"O�ɢ��ݺz@
pp��T���;2"Od�����C�^!�d��='܎���"O:`�U!C�*I��ǯ6��h�"OB��D��2�� �D�$E���"Oh|#���<<a6�:�F4�"O�5�"I�i�\8���$���0c"OZ�¥�V�b�R���*A�.n����"O�i��&KZ�15�S�"k40�3"O��Q%��+[�\(�b�<\^��)�"O��ʐ��?B�� ���[uNM�T"O�҆�:6�z5��U�C�,CS"O�@��N1�q�H�'�	�!"O�T!�GUu0��׌� qB�I�"O�����&�&���(�bL�2"O�U���~��G-M�ͮ��"O�heŜ�L�X��NĠ�@�"O�x�k]uĂ�ۗ U-
�:|��"Op)�5��<7M,1����cF"9��"O�tIU�P�QT�p��ᛲ����"O�ĩr"6�	�`�L�J]�"O����~,Hj�o�?�@�Ȣ"O�88�O�|�l=�x�X\2�"Of@s-U/
R`@�JP���"O�`w�Q�����kӪ^��t
�"O��)�f��J*�C��`�e"OZ0KQ�Z`=,�b,4�2`"O��"�O��Xʨ|�P̂�]�2���"O>�䣓?vp�]��
)�M@�"O�P٣��:��U��ʞ�G�Z��"O,h�� ����GOU�]�<�u"OH�3+�-w��[��9��Eh�"O�@:D�Y�Ѓ�P�7��a��"D��р��g݂i�c�·2��!�$D��)��<-�����3l�<)r"�>D�x��i�D�,9���;x`=@I8D����?9��0�l�1qS���7D�T�p'W$|#�-H��[�rH�yt�1D�(:�e72�ݡ�荾b"��뗋0D���I�]#�\�P�)z��}٦)D�����>+�\��� ?;�	ª%D��a6%�R����#|�p��%D��X§G�{�y��k0[Av�36O!D����X�~�V�!��ؽaf=PB*D���Ɔ�s".ف5Ҷ,�J��N-D� ��bՉ�H��(M*~h{D6D��+tf�!y�4X���C JX��f`1D�`
��1Ð�GDE)�&\	�K.D���O�Ac�3�	��V�b A.D�j�$_!3�|��F��c|��x@D-D�Բ�o��X��Ո ��a����*D��A�.ݙ�Y%-�2v|��4O#D��Q@�'�R��7�
4U���4D��u��K�4,a�!ߴ>)R��`>D�
�&ɑ/dD�S@�
�o�@q��G=D��`��1������ڬ@a5D�T�7J	�[�	��7o-��a�@/D��2`(E�^�j�pd��9P��hi��.D���c �q��x
ql��3�N ��:D�L�`�=r���jـ";H�c�4D�� �!A��_���t���=X����"O8H����0:1�$�$J��`���"O$܃RSX0�c2��'=0*�"Ox�SfJE%�+����(U��Q5"O�%(�!� �򑲆�O<9:��8"Oq���5Hc|�a&o�CBD��*O�pw�U#tt��G/����'���ȳ�	1m���cP�[&U��'�̑��RKi:q�E�1p[���'3<X&M#U�j���c��UB�'�8XanS�V�N4I�i��i�d��'��2v�4Y��L"�(��_�^ �
�'~��Q��\���E%i! �@�'��}�1��X��v�ԪO��`Q	�'�x4C�D��7K���� ۞LC"��'*1��c �0����K��q�'�0��p���.=H z%��8�R���'l�+���Lc�!u&]�w@���'y�سQ$�,� �X�dZ?ĭ9�'�&CCcXL}V�X�k(p��
�'�:�HC�6@x`��|2��	�'mD�)�H��5�$����{��(	�'�����9V&P+�._>z$Z�'�����L	���Lb��A
�'�4�r���pF�ܙ���|M(���'�Lu���׵!��c�7 �z|��'װ8�CٵT���A6N�g�\e�'�x̋��o��� �$h�-{�'��(��	<�8��F[�HЪ
�'�`�U��"
Zq�Q�N�e��J�'�5��c��
1�I#�EAu��]
�'�f%�g�E�Y�*�x�>q�bA
�'�*9	%��{x�O@�*$
�'#Ԁ��+�
{����O�1T����'�v�۰�U�|q���f91��MK�'
:�7K��
ަ$��޹�'2��eiJ;^'By�fۚY����'�$�"Ț1�z�ρG1$�q�'�I���[���@��@N����'o�8Jb��h��GA�/4��P*]n�<QW��j; ̸����$�r�yS�P�<aׄ�=v��(�I֬�L4ID#H�<	C� ���k�伜���G�<a���"	p�"c�r��+d�N�<a gV,L��)�bL����Ã��U�<�*nm���L�,���S�[N�<	���z�ei��[�5�h�7F�P�<�5 =;����V+}`�Ͱ� �K�<��JLMÎ���@�%<?�d`6�YH�<ᰯ�6u�Z�K�<�Q�w�SE�<@�бs�0�� g��(�N�C�<a�Ô�XĩvCO'$	��ƌT�<�t��$� �"�ϟ�3���D�O�<��E9gݛ���pq �h7@^S�<�#G�R7�%��(�-�|�r�O�<���υ�Q��	��0���Z0�A�<�k�h�`	Ca]�_�tڦn�s�<�R�2`���s�ُR��M���Io�<�k�WdL�"��!A>��/IF�<!s�g�+�ꋚu|�A �j[B�<�I�XhZ�R��sn��cs�<)�KT�:p��S�k�I�~!�"��f�<0�=��7�PL�椹�BZc�<as�W-d&(�'�Ӌ��%ig�U�<� ����՚+д�btA�6S&q۔"O�A����F@�	6�C�"O��3��$K����aЕC�x1�"O�)� Ͱߔ�HǁV�Dz�"O�!A#GEL��
�!K-����"OH�Ʋ~=��Q�`H 	Z�"O���&�ǚc�^y�FiO�j*Ba��"O2�ȳ�ߴl�h]rr��(f�D�7"ON�q@��)-^���%�:�t�a"O���7g����{p�Ե~��{�"OT��”�8��t��2�N���"O.%2�GC>vH4i�aR�l�`Ԁ$"O`q�H��c��m�/�sj"�c"O�,8%���><�*1n���1B"O��B*y�j�S� %F���+�'��z��5b��R��T�	�'M�� �E�8i �a��@TP)��'@�q�)L6�T�! �*a:�'e�I �gM>}��%��]���]��'8�t�S�L:�\��&��h\n�q�'��t���K1�2�@�T�g����'Ili)��BI�nd2/׺X�r�[�'@̹[�`�%���Z��Z�[���'�Z����,x�Q�+�V�p�S�'ߊh��m�e���P/��C'0���'���w��PW�J�#΀i2�A�'=b8i�h\�:������+N9 �'2�uU�7�!)�
-,�� ��'2�adD�i"^A3 (�t*�'0$�ӆƳn4iz���ت�P�'zZ�PȝF�
�����At���'�T͈��
'A����J��	�\	�'E�!���s�fy�a��<{$��	�'��e[s�;"�Nerp�Ng~����'PT5�����j}����,�_lb,��'L,���I�y�Hy�W��(]��{�'���c��E��{7+��,��u��'<V����Q��}�5G"#X�	��'�j	�v���q�8�D��m!���'�n`��dxhڤ��Y�Z(��'����\�k�D�-`��)b�'B�]������TPe�Ŝo�4A�'u||�$�P�g�|1�A��p�����'�P-��͒CYr�r����o�^� �'A@��gF�D��n�`��@Z�'�H�ծB�i�j�HY^��a	�'��$��mΞc"d���[@���q�'�f�Ԯ1�*)Я �On����'[ s��^�).�MS&�$F*h-��'I$]�5�/	�:�A�D B[�'hP�h'��)}6ݣ��	�2ۼ1��'�$���R/Mm`��!)�)��E�'$�	2Ɣ�>�0T Z<\z��'�`=��kn�f��F��h�����'T�9j^�c^dB֯B�_}ة@�'�n�j�''"��y�f��3$�Y�'i�
�E�-�8�l�4L��"O\�acɘ[��;��ݧ���V"O^� �o�/<pG	I�9�6�y�"O�,��H�w���G&Aq�X�a "O��3S�G!�|�i��Ѩ���"OH�9�	W�F�DD����º�"O^i��KC�qh����Օb�P�"OD\�᧌ d0h-:R�I�=�zY�"O� ���c�Ҭ<�Ҩ��h �EG�p�"O6��g�c���Z$&�3T4~��"O��3p&.M�>tɦ�T%B	�3"O4�@O |�C�
.E�@pV"ON1��d������ҧ��"Oz��,H�P�زI__�@5x1"O􍫡֞(ɴ,R1�ȟrv���"O���'�Ձn�=c#���Zr� "O8I�U�SEE�Mĕl8p`�"O�h%��su��*�Z!iW�IQ"OЙCa��<��r�[Q69��"O �YIv�rW8!��0!�͛�y���
���5�\v��$zpȓ5�yB���h�)���G�sE�4�עF:�y"�>#yn�B0�ϧdr�rwFT5�y��N�B���"ֱ],m`-͚�y�*E�y��vN��_�sF(��yBD�9u}`C�Y@�t��y��+--"�
�N�]�.�[K~C�IX9�c
̳c�
8��	�`�B�	p���B4�K��3Pm3et�B��&�����'Z4혧o�o�|B�	?��Y҃��8@���{�pB�	�X�<y#�_�br8�U��2WŮB�IT��qR���Ah��J[PB�	q� bTG�8h$B�x��:EaB�	 <O�����ZB� 	S�d�B�	5���7G�I��hʐ�Q??r�C䉩8���aG- E�jQ;L��C䉽
7����?�V5V�hC�	66��P�h�>!�F���q�bC�	�nV�%��+F�V�z����>@B�I�X����Am�gʰ�Q��78cJC��(u���JP�>�tl1�%�;a>zB�I�-ބQӐ�P�]�(��e ��o4C�	�`6��xg��=��i��-M�C�I9.��y`]�n0�|9W�R�C�	�Q�x�s�Θ7|���pG�E,o7�B��<�2<@Dɒ�6�5�i��[h�C�ɏB+�eQ��t��i��?A�C�I7Xf����nߺ=�2%g�v��C�^u�$�6d� >�$��j�X/dC��,�&� T���*���`T�_�XC�ɘ8����F	s��TeZ���B��M��0�䪛�u$�t2mD2fV�C�	�#(����,�#.�eP6��0�C�	Xh�����HJǤ���IǢv�\B�I�?8��@�W6)�2�;e��	��C�	��:�K +o!Nyb&��-�JC�I%K����T�[;<)!�ۇCbC�I�f
�y�C*�� �dj(/|#RC�	�>�`���)I�!QO��CGHC䉞��%QG�|٬�8�o��U�FC�Ɋ<vZQX��5ol
�%ǰ&��C䉣.�ؙ+���	3%^�{D-ȵ*�`B�I�F����NH<&��dB�/*xB�ɛ!�d�)Pv
�[�	���pB�	!Q�\�
g��8��׊�$-~�C䉺9W�U��C�i�Ҁ#iU���C�I�"��%h��|1z����"qzC��<54���D��dT#S�S lAPC�I3]%j��ƉE�2��S�ÐZ�>C�	�4�v5��@�"`��1#ĭgg�B䉊i��0�cߢ&����*{OTC�)� �Y�''
���N�*�T�"O�8��ѣ'�4���ω�?��E3"O����nF��X)� �;� �r`"O �B�mB�{��ʚ2��س�*OF8X!D̤t#�%(��K�]���i�'
���	I�(b�`v�.X��Ͱ�'�1�Fݺ:,�j"R5L�h="�'�LL�tE>h�2� EEL'o��@�' $9��E�2h%���d�x�X�'ޔ�[d��7�j�:�*��=(
�'�l���͍�z5�ڐhE���'�X|j&�Mx�\mۧ��/�2l+�'�̩0 HSh�D��p�`�'n2�:"�@�k�LJ֋��,#	�'Id�됏�����P'ç��
	�'*>�iÃ·��)�Q*��\���'�0l�D ����bql@����c�'5�u�Qi&0f� ��"
��'��D���áXAX���)���rę
�',�8Ҏ�?=D�.�#7����	�'L�%�w�պPZ��	��¬����	�'���I@ۚm�.��'�;K�M��'(P󠩆��BI� G�N�<�b�'A� �C�]!|�eq�	E�y3�'R�\�CE%�&,h��&6�6��'v��5C�<�t�{��.��ȓ,_y�3C��?t���@��*C��a��l�<��?*�!�%��$6%��ȓzv�}���>m���f<d4�ȓ&ж$�b�B=(^�A�w�ηcC
8�ȓ0z ���+��vA(��W2x���ȓs�b�#��D<irV�s!�T.��ȓ8� y��k�X(KF�Tb��ȓM�� ��Ȕ7re�B  ����q$e�Diۿ���#���,A���,t*0Nޜn�)5�uΨ�ȓf��pIH9P���W�=����P��uA \Vgxm1�8���ȓ��54
�7��]�t�F�8̇ȓ�-QGL�gd���SB���Y�X ��C�*Ā���d��p�ȓkРX�bĢ���Jκ3Aj��ȓ]��a�d����8��cC8Gb`����4�U�V1X!GH�^�20�ȓ,Q�)cA�_�;q�TP� @y��͇�1,.�+��<�hАR�1@��`��m�~U��HH�R+2Ma�-V,w#ʝ��L��i	*Ċd���f�A�'d�ȓ)"�!*aʁW,@�&O#*�̅ȓI�A1Չ@M��8��@"#7:��=<J�8��V�`��hpq�M�D����>�p{�.�m&�JA���(��O�l�yT�S�>����@�Pąȓk���r-��p���! ���U�B����Pъ�D�y��\�P+J����Y��#
�2_���s�*ȓ��`��h~,�3�.?�t[�jA+?�@I�ȓ	W��0���<5JVS2��'�Pt�ȓo�2����
`�����T%=T���J�Պ��XWh��-�9O�,��M��%�baT�h.�B�!�#�<��ȓ[%jtgX��� �/��H�C�	�x���ɡ
,tB�� ~dPB�I�f���A���#�J(#��pXXB�)� PyXg�S�m���BX;j��	0�"O*]Х�LѮ4����,�T�s"O���H�j`D!�䅯P��yA4"O�I�����"<���	�0��"OMS!�܈Ix`C�!ˆ���"O��TM^���J%��t�5�"O����c�%Ғ*�?k��A��"OV���E�#�4����t\&)zE"O����aӬt2��� DW�Z�"OF��N��=�ΥE�[%d^�y"O�+.�v^d��#K�Q���;�"O6h卖"8��@)�F`��C"O��Rq�½%�F�D�wxxS"ONHx�X!Ou�4zt�J�i�q�F"O64Pa&�|�`(d'
�_��M0R"O��X�#��D�@��4�=׎5�P"O<]��`�7����W�̚`���pa"O�1�_b <3�R2v��q��"O�� �JJ�Q�ڐ�w�
����{U"Oԭ�`I�4M�����:*ird��"O��ӔoBX(J���#?��p��"O�����n�r�K��V9\��"O��X�X�w��i��Ȗ�&訴"OD`� � �����,�R��t"O�Ie#��
��-"k�!���R�"O T��n�
m>�
P��F1�"O<��O�O)�s�)D>b��e�"O��y��GX]AS���-�$8�v"O�Ի#苺_~�����W�z�J,c�"OL�c� ȮR�ĐPc�Z�U�n��"O4Ix��φ�<��fY,_���`�"Ot��`�l�x��A�F�&c�5��"O}��S%����}Q���v"O��#$�J4A�L�R[Uq��"Oj��խZ�Un���`��SV�	�"OJ��Y0m�Vl @��v?x@	w"O��ۤ(��_ht)E�NF�i��"O��ӒBڬp��c�O,q�L��f"O��v*M�:���rWgՉ:��|�%"O*A	��8V{��&КLpz�"O���c��N+ȵcD卽,F~<�"O(�� ��}.܀�vnѲ+�Uّ"O2P�Uo��,J�9�1.0G��`�"O.1�u��D�Dpr�M�� ޠ�"O{d�ӿ%\���Ɖ���p��"O��Q�F6O����A�O�_��q� "Ob�bQǚ�ylT�&J4.尿2�'���K@�O	x��`��I5oT�'��YZ@��[��1�h��^L���
�'_x�ip�W#Hnd0�P�����'� �� �x(���#9�"�"�',H5+ф�F�pZΐ�DXR���'��l+"ω�?�
i�Հ/8��@s�'u2�{p�7P
���n�� �p�<颫����M�C��G($|�'�Qb�<ɠD˾e4�P�dA�g`N 9fHGa�<��虳? ^�K�S�c�$P�x�<Ib��M�t�[�.]�P���c�AI�<Yf�Q&b��XҒn�?+��h��ÞE�<�c
�_�燆!��%+��	V�<��JA.^�h�2oЖ|� ���S�<��"2n `ˆ���Z�j�ÜK�<Y�	�:+F���� 5"�P�jV_�<�` U=m��0Z��
@������X�<� h�ӂ�ķA����� �m"(#�"O☉F��^|p8@ŝbbxrV"O���dB��eLˢ+o��)��"O:��U ��(ږ�Cpe��Y��� "O�bQ"��]I�ꎚ0�8���"O�T��i^�r~8�2���:*b�"OFi�֢̹I�|�5�-A�1"O�����1j��X96 ��/�� �p"O���eY�jQ����o��
�TY�a"O�v&K�|;s̏h�tQ"OغE/F�&��Ȃ�	��	��8C�"O� Q���;:������*�c�"Od�A�Z��]����"0��h�"O�y�qmY�z5`0���=��3V"O��#�@�!�>�� $~��q��"O��BF&8�I@�^923.�3�"O|T{��2�Cg�,"�v5��"O�u�V�Ј�"؂#hW:7t1@"O��yfL?X}6A�Hך~b��"O��p��Ӯ+��	"�#��h�"O��R��� 1q� F�j5n���"O��K"��@!�6�W-q���"Ox���nċ26�i��G/nﲜ8S"Oyh�N�h� !a��/�f�+�"O�+��@ǌ���J+k��I �"O @BTn�H�N�0�̔�V��� e"O1b�O��d��Ɗ�&l��!�q"OV�"hĨ0М���
��@qұr"O<e�#��
W�P���]�lh��p@"O�q�g��wkB��Q�LRL��""OL�zҏT�n�0sCEQ�`J3"O��{�.��f���ᢤ'SmJ�3�"O� ��ַ2��D8S�D8s�h��"O(��\+}�v��&��B�����"O�(Db^�~���@1�lM�v"Ó���ӃOYTU�р�2ky�1+�"Oz�� ̰?,�� �wi�<�W"O�d( 	�W��"#MW�<�Jl��"O��0���"k̞!C�pU0!
""O"t�@e�Z#�`�p��%G!��"O��p`�Q1_&�$o{:�4+ "O�	�U��+T�*C#�6@)v}S"O̬��"��uެL�d��-�I�"O���d�PO�Vi{�e]L���B"O �1$ؒH��J��D�L��"O�V�2�Y��U�x�$��}�!�Ĝ"���o߮X�\�[�C!��6@����EO8$���h�!�;�XM;��7c�h�sԡ�	�!�ě�(��I��6 ��)	� �6�!�$
T��;Ac��s�إKg��~�!���N�P(�'�=�8�e���!�$C�b�x�"�%9�|Q�EADY�!�$�+$�!�3B&Q�����Ԇw�!��
�Yڔ�1 �FB�Y��N�.B�!��1�X�I��}ٖxi�N�z�!�T?;�P���
J�8������!� a{��XC�	C�,�iT&'W!�D�=bT��x�^��;��-o!��W�����hS!R�5rW��8<!�D�B/&\�6�O�"SZ����S��!�$T�\�fM�eL�v@��2a��)�!�d�{�Bj�5~=��jw���!��S?wf�K���, Jx�1$߈�!�� ��k�ES k����0��h��"O���ĕ�t*�z�`ȩ.���"O����
 f���_�_	TP3"O�Qp0oX�c��p��ɐ	Xl�C�"O�1���02�����I�5oWV�Q�"OT�*%O�6{r���B��/����"OڈZ�I0q�eA�bG�'���""O�m0��C�x��݁s�L�$��4X�"On�b�+�#�`UȵL�1�HXs�"Olp�ˊ*zp
$Pq�/_�,�"O��!�O2}�A���ӂQI5"O"� �e��Uv�<H��w�i��"O~�W�L�N����B�ڪ��S"O��kՌč<�^%��#چ5aB���"OU�V��@��_�fU�A"O�\K@i���:��*�.?��e"O�a�槉�(]4I2�JI5+��a"O���1oy�}�5,��W#��r2"O  @BC�O�i��K�
�e�F"O"�rT%�B�����H�0��*�"OB��R(F��D�&aY�A�����"OHJCiW2d�"�9��^}Z�"ONq;�G�-�n����$y��	��"O�0�&�C/� !��ͼm�`�t"O@��E�g�`�����n�� 9�"O���r I�<m���5��b�XV"O�xp�j�AZ��Bad�f��@A"O�|*���G��³��%2�b�"O&0������d����a�"Ob���� z1dp1��B�|H(��P"O�Q�@#�C�Va	�*Ʊ03�pA"O08��ŗn�P�Ï�T.ڠ@a"O�"2(}`��e��v>l��"O�)cVlA�*R�J��3AY�M�F�|��'�l;���2��Q҅J��7&�
�'�Nء�h�.�8��C�:��0	�'���R`�N1���u".o��uq�'�,p` �!�l�c�o��#�'&h{2o�J��nV�~pD�X�"�'j�>�	�P����ߣEh��a_�Q��B�	(p���B,DR�H�nȟ@(�B�ɀ-d�yU˕����J���|I~B�I�_"��1��v7H�JE\�\B�I7h�𰰥[�o�.�d��!�B�I�,�(H�S�D*b��0S� �t��C�:��)I�OC*T��Ă5\��C�	SJ�@�W+��x�A�k�fB�ɡ7�~��bc�&nБp�!�&b�`B� S��AB���g� u@3&�P�C�Ɉ#�6��5�_�5��{�!t��B�	0i�^���@CK\�S�O�2&��?�����3l(�TA��Ul����c!!��
0��|�bK�3#�|Y��βR'!�d��H\,i(��v|B�c�P3h!��ƫ\0�i���}_����1]!�^�<�b���I�}N`�%���!��<����$����Ny�G��(A!�"tGȅ��@<�H}���F�	o���O�� 	�֥�c?������-!��U��1;H�aw�]c�ة��&!�H���Bg$�X��
6u>��"Z���IN�f�Y�Y�UCgF�X�f���{b~es�۪-I!ctc��9AɄ�l��{ ��ʘ�t.�/\!����S�? "}:���P0q�K,��8�S��A��)擓H�f#ײ[O�Yu�^����!�?�y�̏;I�h��'Qw�y$���HO6��Dـ}����䅹k�\��RgJ N�!�D��"mѹ�dԩx�����t�ɩO��kL�D~r.Rp��6BF;.=\<��j���y��!K�:l1B�[Z6+�f�6�~R�'�v)z�@���Z�f��J����'�ޤ3�ǝ�k���z� I�F�0�'��,�@���S��A��*����'��L5��!��DQ�ƞ6\"Y��'{L�PP�nc��AǪ�T5R�'|FꆗgEl�b7ϔ�	'�T��'g(!ᜮ.���-S���'�-��MI�X=^����s��i:�'��9�P��?~+�)5!͢ �l��'u�0�ǼP�Č���H���'��|���l����d� �z��s�'ɦԫ���&^�j4����z�m �'Q�����M��'�{��%��'N�����P�*����!1nvֵx�'��A��7R�����+��K8���'XD���'�? �d/�a�ES�'���sf�M;%VX�CC��X�
�'�FIyR�Qz� 9A��\� b�\�	�'Ǟ����ք>�ֱ���Y | ə	�'v�3֪��X��(�]��))	�'�,E�S$>����Yi�D��'�LQ�c���0,bAhB��S��\��'�D[�MF=Im�!�"�R&@�
�'U*l�sc����U�y$�a"O����f�J`P��ԦNtF@�`"O�$7�و���JP�_Jo��is"O,14�	6U*zu;�� mVv�2""O��� �wY�x��#@ZC���@"Ofъ'�J,�f(��OկG���6"OL�+D�J>'�@��ĕ04\\� "OXa1U� �*���?ʎ)�0"O���	��P�8v�E5/er�P"O���1DT�n�D5���Ų(�Lp��"O�9�gԷ{���2�P�<�p,�"Oz��	��yzhL��O�4"�"OL �$#�>Nn|��=���q�"OZ�1f���0ӈ(�)Wa����"O~2��=4�(u��]��H""O�h�Z�3�G�>ƽk��[9U!�ē5G�8�P��=�����R�	D!�$�v��m���
I ��x�I	2I�!����l���)�mZ1j�7�!�Đ�DR��#%�Ʉ���f"��A!!�$��6ܪ=a�c�%4�s�`�	!�T� X�X�kF%\m���  �]T!�d�-���A�\��Y2q�S�^!��U��0��F� �n�3W�|@!�DȾW�e0 �̠F�\ēE٠E,!�ɰC�`!��A=@���*@�_!��ʡ;��u���XQ�\D(�+��D�!�d)io���g���P�JY�I�!�d�`�*�%fįŅ�8��+ "Ot�V�[l�"7ĝ�",���"O@�C����z�*5DɅ!�ah�"O�5v�G�;��)��:?�t	2"O���fJ7Ŋ�������"O�s�O��w~�]aF��R�@,��"O� B���Ԛ)��ɕd�if��"OpIu�]�wN�`�I�P�ི�"O��AU K�@�"U��뙐��}g"O0�%�N|Ƅۅ+�9 ���А"OA��՞iUص;�_mhb$k�"O^��u�ƙ<:MR�č�;��j"O�K#g�cʝ��F�7�Mc"O������{5�QA �T'5�`"ON��mѠMw$�h�,i>D�"O��)cL�n欲���0l�ܫ�"OP�� >X���b	�]�lD��"O��8��I�h��a�@��H�"O�ɠ Ǘ6�y��""��4�"O���&��	��h�2F�b����"O�y�w-5����eW�2]��"O^��Ed[bJ�5�g�\�"}���"O��y���!N�T�H`G���1�""O$��R�
xk*�"E	���e"O�$KaBǙV Dȹ���&I.�R�"O|mQv�^�L}(PP�h�
~�*�
�"O&��u��5*q�r��V��F�2f"O�8��LZ�v�:���sȈ�(g"O"ܚq�ó��y:C�֐;��)	�"O���aÂ'RAԴh��\�ru�E��"O��ZU�ރ	�Y;a��GB�"O5�V�٠8�|=a�ω�~d]H�"OJy@񪖩F��ر�/ǰ��9�t"O���
�Es����m�.+^R@"OL�Q����}X��*�gҝb(��"Ol��fBݰ6B�y!�DsY*p90"O���+�l��借�&@$ T"O��Q3�I�K��!�OU(Q^��"O$)�fA�8�`��� ��M^���t"O�@���g����!B\+��`�4"OD�S��� �xM�堎�`�Q�1"O�������D(�0ǹws��"O�݃BFB�i��P�@�ʀPp*��Q"O�� �C�$�\|`$dڨW����!"O�H ��Wh&h0�Y�N��9zd"O�8q�Y{�c�l�8F� �"ON�3m\ &�hV��U��A+�"Ob�BwdW�(��ܰ���b(��"O�a,V�A�쵫�f�'@�d��"OA`�L�xV	��g:�F=�"O�!Z�&�>�P �%F�;R�^ݒ"O䌘�/�7Je<@��e�|y��"O�@��|����MMUDl��"O� 
��|��壶�L;6�l�"O"L�%�-(��YrէT�8��͡�"O�5�dK�!e��p�F��E�ȸJ�"O��0A!�/Z$F�.!�$H�1"OZ� �R��*�rEN˥�f��#"Obi`.�%l�	�pL�5MxxȚ�"OФ��e��(�sE
�< 9�7"O΅��
�)ֆ�1��vT�-��"O�5���C ��"��C&]�<h���_d&(x��'�2ãnP�p��
եHiV�*	�'r.�A�+��9&Zk䨎"o�~0�	�'��!�G��>a���⋇o_pS	�'cJh�W#T5a?+EO��9��'5 ׭����D\�r����'���˴.ҒA��j��՟m�d$��'�|�9C���h`K�+0�e��'��:�ǜ67�MK�%�S������  �y��f�$|�����-D^�"Op��K��j��ɐ�5b�"O8p��D�C��T�A��'H�TP�!"O�	A��>7�M�C�IQu���"O�(PbK�z{؁˴�֞S��P�"O=�oF!m�!�5"��a��MkV"ON�R�O�ȩB�O[r¶��`"OjlѠ"Q0J�����.��v���p�"O"}��G�,2�r`��Z�,jN�2"O�I���>%��X�" �i�r-d"Oh��U"L?nf�� Q�7Ѻ�c�"OL)��/թ<�>X��V���2$"O�h	FݬN^����%�!t"OF��ċ�X���J�&=겤��"O~���,�!609:��M.c�|h�"O�l� �Q�����%:(hj�"Ov%k��'6�0�RVL�4��C�"O��WG�	q�Z}h���4�|�k�"O����Ռ<c̈y ##��M��"O�����ǨkF�h����X��`"O�-�j����]b�!$V:`EhC"O�UA�
%����� #�DYW"O�pyŊH�&�h��7���"O��"R�}(���+o+z�yq�O��`�� 7-ZqS��/,O���E'��1�����!�Rl
p�'k�O&d���e�-��T��K!r ��)&��/)E^�z�O�\�A	\�-��	�ň֫>�h��@��/.�3�$r���@����E���C�,EzR\���Γ+y8E��N�lu���Le�pP��6\����OV����x�$	2qp��^�O]��/3��4Xm�)�0�ʳl3]s�B䉩ʂ]�$샏X`�4k���0
�
�LؔN�4�e�o� Rg���F G}"ER�V��q�1i�2.�|1	��<�)V2,�h#Q�ȊU(Y�ھI�5����!��`�Mݥ|��������0?)���+[� �b��O�H�8��t�	�����!b]�jB��A�� T !��ɟ)&��?N�V1#f�W�(2�A�K�2e��C�I(�ub Ԯ%����&���|��� \%2	R�r/�n5����+hܧ�p`�;�,*�g٪�$�S�k�!T�
�*�
O�sB�9�`��CBȮf��`�v�O"!��3��֩=-��"�jN$nO�LB��8�n#=�4CL8Ql>� ��+_.hi���O8�����	q.�\�0嘴46�@�nr��%�R��J��0���r�bS*^Y�T5��kX����"��	���Ƣ�x�<U���!}�ͅ�'��e��t�Hȋ���F�VhkR]�k��ӎ>���X�6ĆY𡋠�B�	�?�0����#�~�I���8c�1�C@ΑN���Qb��A@|�3F�ޱ��EHr�~ޭ�pk�'|�����!�ɀl=�O0$S�"��R4B ��+�y��G
���!R�(��Y���r�4Kr��� O�v�^,z��_�.�M��ym��-GX�P*;;�P�c\��hO�M��W�6�:�.>4+��pw&�7gF�4ѧ� d^� ���
)��#���!u��f�8,��­����<����J�z�14�U�#U���� (�\x��)�A7R52E�D�!�B)ĄM�b�a��� S����!*�V|�� �+�rݚS>n�`u�G,4^����_�j�C�#M��<�M@�j
����G?^	��(K�g�<J��0]�`�8t�T"M�� !�� "lϻm���Q�"^�i�������	�n��� ���K[t�P�F��y lO8Hm�T�����fִ$�����TƉ�o2a�0�:B����;Na�|�'[P5˂���99(hE$}�Л���Oxv��*t><B ��M6����
)cS�(� 댦3:fL�u݀	��P��� ��|��Z�-�/� W��D~�,�FJ�'N��JYI�Ћ_�z�P�$�z��yѡnw���ULV�CAԴ��N��@My�'�V��<aK@E��MQ�/����H�ז���'ئ��cD<��`�!�&��R�m��:OZ��� Gd�/��Eд��;��=$�"��b\c���x`� 5j�f�+��دH�@x)��3lO��E��+�D�1����<TP�cw�-,H���g����<l("�u�!�c^�x�T���
�&8f08�A��+3ꁨm��\��M	q�R �e�)�%�%�6��Mr�Ս�1+�M!��/��t����_�� H���qx��*�&2 �mc��K8be9�g
�&g�k��е�p��CV�' -Kn:�Ya�D�W`J]`Eb�`��Г�|^�RUfT'1sf�̓9 �y!G��Sj\i��1aG>Up�'+K����5A^ ��䒄}d����#n�氛4"�� L��O7>)ʖ͎;H#Lݨ�o�x�Lk�#�k���ۄB���d�ׁ�59�7�� �ͰE�̫2�*���>#D�P��'���Io�����˛�1���B��AU1�y��%��=R�lrS��/C����_�Y��sɧ5���b�lV7�a���ɰ?V��R ���i���x<�Pà�&�O�8p�	��Ot,"��P Jc�)���d�@��� !k(|�u�R�v�hbrIݖbd�XJ��B7Y� ���'H�#��Ii6F�$h.�>3ČPfaY����Dg��0gJ��E��@�ɨ�K@8Kv�0s�č TnmA4A�����G�4iR��T �#l<�i���6OET���fłN,���'(r���/�;�LPSFGܤ�|�"�bW(��|�J�7`~�i�a
G)q.|��WO
�:�H`�g�&�v�:�;~�VU�Hzh)����P b�x#l���ѢW���F�K Qfzͳda�/
���w�1mS�0FW�I���`��������G�B\���_����'y��	0,�;2�����c6sq|�
gg�L��9" ظ��':B��cΨIf�$,0�YC��C��?�Co�Kc�0�S��4v�8<���< bC���|��͖�_N���#�� 4�Ԑ
�J'x�lA�d�N�'x�jE٥�>#���2K�"(�L=HS��P�����͈�,�!�$�V�؁��
�t���L��9xE�I:���P+י)޼e�l]�U�ԙ���_�x�=�A��J.�]� �V2+P�&�6�O�ͣ�G~�8��V'R�*%�E
����L���y��nu$M�҂�$��ov,]��ḑo�:Hص�? T��Y�9o���g��!3Ƿ�����7e
�Âi�]k� ��>� `ߗO,v���ɭ����;>:<��5g�#<YƦM�^ړO���:X��ƛW.6$H��7"����j��!�D-���	�sg0��3J��E��̀��H��m�b�@���
��b�L�zQŸ6�]
�y��S�W� �@B�%$̬��ə?�M���S&F x�<���Lt�>ѷ��ʈ�(��A|�����v�<I��E����PuKſS�䙹��z}��F+X-���ۓWD2$(�통�����2�>���I�3�6�k����P�F,p4d�Ĕ�E�����f�H�� ��:�4�%J�;'����$�XId�D ��s3d��>h�ȓ3,{�$�*\���Lg�.a�ȓr���IY�=�|���M�A@�E��P]JTs��Z�����\� [���ȓhaN���.D-8q`!3�9d�p��m
|�X��.+�9�$�EL+��ȓdK
�Xl����@�F)��	��vfHX`p@?xG����i%MX���ȓ!�I��a�6�t�Cfk�#fĈ�ȓm�
UeB�fLP�ۧ��k�(�ȓ�`ѐ���S��+�e��]�`	���0s��L�6[N=sׇ֬P�dY��C��P�!�$d�܂1D�<.6訇ȓ�I;Q�ɬbK>(ac+T8���':BM	v�X�0!v��4"�/����ȓ��$S��P%=4��g�E�J�z$�ȓc�~�� �4ydĠB��rm�����I�5AQ>�z4�.Հa�Y��F R�.�F�$-�&
R�C䉯O�\� G�Ts�+�]��C�(�J�R��c�a��� rTB�ɗnn���ˆ�V��C&�M�B�O:�YKs�τ��1a�($��54v�H�?E�$�]!f ʴ�#K۴9�e;��P��y���@��l�v�X7��Pf�yr�K!<� �(
� ��*P��0�yrkX:^\m�åӟ���hE�U�yBJ@�PDr�� �M�|�����9�y�h�3)Ԩ�d��9]��)��&�y�Û6J�,��OU.*:z�pC�M��y�	D�K�ڼ�����)tf���%_8�y�FA�����&*G%(��M�����y�̙�.�08��ݾ�c�j�(�y��H�5ɨ) B�7�%�6�؛�y�c��~��H�dJ�~EĘ�� �>�yb��/e2V���m^H8R�D��y
� �p��7W~t:��i�
���"O�l�$[0=���Q�˖.�R�"Ol�r�
�(A�tyv�
�XF���"OF�S�yH��[7#��uN�ys7"OpT�g��5	YZ�r2��SV�!("O�a�D�Q��;o �u�0"O.$���_r�B���LO�o�5�W"O*�i��"] ��!M#.�1�U"O��p� �2"�x��D=R,��3"O�����E2L?��������1��"O�س�CAUP|�3�|s�	�D"OJ5K�֝3n���'5j�H�"O   Q�R�b����ab��}͛$"O|%x��m`(ru!��X���"O�YV!�TZ0yt*#I1�]�"OdU[�<�zxCi��Ѩy��"Ollsr�.@�nL£nAV�4�p`"O����HZȪU/�;&ô��"O���q��7./� �1���<�b�p"O��!��ߣ?b���k6ҭk&"Or���'Z�~��-V:���1�"O<�2'�\�|(��ߏR6���"O��:}� ��
�%D����"O�57#$qf�@T�]�DL:(�"O\�k��1,��Ppp I!$ƌT"O�t3��N�h6��1�D�	���:�"OQ��80�|J7DN�:���"O�:��n�����R�x��Q"O���q�G�Z+&�Q)t��i"Oj�{d�����B�C�20��0�"OR��􎋶�*$�g)M$8e��"O|8u�ĉv����S+E,��i�"Oh�l�5@���"Mޡ�l��s"O���o 6�B]rmS/)#����"O,��J 1b��½�0�E�T�<�E%�����E��5�*0{�C�R�<�vc�2h�c��Ѷ�*���Q�<�%��ۈ�2�N�T�	"&dHy�<��(�;�i�$i�fNH�<񠢟�1r���O* �"�H��I�<��	I�L7*�p��)A�tu��UJ�<�Ɯ�kʪ]���� d���y�<�O;P�C���'-G��+D�Wm�<�3��4� �[Dҡ����b�d�<�g-�Ph�kp�ן$�R��j^f�<�U�Q�n�*�:7jR�j�P!A��X~�<i�(�V��F��̀ӉQf�<Y���4���:�#?p�|��2̏]�<A�*�C�h���lQ�SE�����G�<	P�A���)rl�
n���RW�<��$#5��
cY[\D�t�f�<���E/\�]�č���e��u�<a�jTOBĵ�p왐rv���
�J�<A6&����p1
�+ �.�jD�<�o��XH��B4AC��D�<�v��/.����`��\b�}��ŗE�<��ʰ\�쌒wd��P�(�����_�<�di��K˸(��J�4���q�/�V�<ɦB�2�]+���8�
�BD�_�<�"�0���#�L<J4��A�Z�<��(C�fo���� h����RcP�<	�g�/߀���X=\�h��w�Xt�<�"؄^醩k�����U� u�<a�/����İ�%7v&��$!�l�<� @�hS$*M���뀌Te�r�"Od�H7�?x&ڰ�%H�;d�$���"OR�3�l�-�%BӨS<u��l�"O�X�Fe	�/���gɴe�j��"O��ZG�,,��=J��Ej���Bd"O$���'2��$�b抯6d|���"O��)�Z8B��`+���7����"O��w�KH��P�E�r0��9�"Ox�k�����9 �"Rt�Yv"O�����~d��jݗWf�B"O�]Bw#**,��$�سa*��KR"O�<�c��.�j�R�_r2�U"O(��˒�,0E۷n�!�BĢ"O�U�%��	p85����h��<;r"O<YBF3K���s����VP@"Od���˯\r�h ��6R	��"�"O�5ȣƂ:g�h0��E�xl���4"O�hQ��/|9�	p�B6j��*�"O$�@�$T들��dx���a"Ob�!�n
W���P`L���=Xs"Of����~-R�:a���ً""OVu�bI<%!�$k� F��:�"O��R��B����J���L��T"O�QJB�Z�dĨd�P�0^0� ��"O�P ط	q�l�GÉ"2ft�2"O���+�',�ʴ��i�@��"O�T�&/�3��=r�W�&P晒3"OVY2Sk�pߒ@2B�+,@Be90"O�12���}W.�@E�**ry1�"Oإ�q������b�	U�e;�"O��:�%�!�����!P�	���"O�u ��J7Ix4( �}�LS"Oڽ���B5�P4F<wK�H�f"O&xAMzƈ�Qt�Ğo
 �Y�"OL���6��B�mшhԻ�"O��ZՈ��/4��F�c,9!p"O"�2co�8�@*����{a0�"O�8�"$м(&�,�Ӄ�[��$�0"Oڈ$��!6 �[FA�E���"O@�aEHT=T���룦��KM��K"O���a�ODk�Q��FC�
���"O�����@�s�T�FD�&W,`{�"O ���.x���EJ�`I�0"O�dZEo��iˤ4	���p����"O|Yٕ��'/|��΁0K��)6"O��0A�%s�f���Q Q}�,A�"OB����c�PD����QQ,�"O��i�K�1)�T����B\T�"a"O\������. ŧ؟mG��)�"O�Y!R"�f�Fi5��=4��"O0(���$H�pH��_����"O�]�#�:<��t��,O�h`�"O��`��T�n��Sb�L�B��"O6٤�� S��AE���'=f=0"O&����PX��Z�j�#q��<b�"O���=�i� �S�2j��"OԡOŔK'^@�!f	!B���"Ob}���T>3�� ��Ɋ,�h�c"O����	M/&<�f:t�>T"O�=����ERz��CEM�6��U�"O܀0F���X`�QI<����"O�0#Y98�������#"O$pᇪX�DZ�MI�&�g�bQX�"O�t�J\�o���ㄜ7o����"O�  Ц��3=?�t+��q��j�"O&�b�iǍp��T�1t��ɑ"O���eC�� QB(�dx�"O���!͠~�y0�	A�8�vE��"O��+B�+�LDòN�'���q�"O&�K�	ϩ`���#�/�8�"O.�(b��"|� ���6@��W"O�A���V2��(1蝖C;��Q�"O���C	L�"M3�J�d*�P�"O@��ץ*̸��U��|��	7"ODS����=HzPrRc�d���6"O&��+�~����XX��"O��֦�d㮡
�߲L%*m�!"O��R-W�o	�u�$c�u�~�Q"O����QRA�uZ���遂"O�d��̵qO^$�֤(E����a"O6��PI4'������;M�"�K�"O$�K3NL+~�Ȉ+�,��h�"O���풹]�@�a0A�>N:�3�"O0)�R�F�R�	�j�D",Xj�"O�^ʐ	�(��g�1X�AD��!��8���A�\�Y^Ƅ0q�g�!�d2	k��X�ND�~�`%���!)�!��r����H�/!���U�ķ?�!�d�C�Ze"cK�3|v@��d�̈́8�!�d)9K|YI��R5{䌂#l��!�$G�SVH�C��ivkXBt!���%�q�UT2iG�I1cXO!�d��*�E��M͑9��3�#TA!��\����P�@F?�xS�R	D7!�dM�
vtR2 �	g'0$y��1�!�ҋ>�h0@A�1��%�
! �!�$
.-�m؀h�?CTH�-y!�%n���b���JPT�i��Ӫ]!�DY�^{&�: �J����K�!�X�)|*�`6�T�Y�Ƽ�EԷ.�!�E.[Df�`��r�<����)t`!�$&`̄ZS@�6[u���jчS�!��ă9p�@5`%5��1H��!�L.3��Q�0q��%؄ag!�d�u�Xܩ6`��Ien%cW#�Bm!�DԀQ�����%|~hr�c��f#!�䃪X�(�g�ξ�t���,!򄓆���#�ʝ�@��%z%`�6	!�d )�L�%��7i�	�R�ø=�!�K�5�e�
��)�S�'!����*���2��|���S6u���ȓ3����Cm�\�(�9�DY0b��-�ȓ�f�AB�)H}V1IP��2e/���FIޕ�t��'ay����	3�8��'K�����TW|ɠR K4	$^��ȓ"�V�5gӕO ��F
aa���$� #�26p0`3���xj�(��v��is�f��>�X��;���ȓa�,Tӣ#B,i�A�	�
3�|���NL*HY1`H+%��"���Ն�/B���/Ȱ*¸P!�Ș�)�ꥆ� �h��gbC���e$1!��ȓX�d`�FE�q2�,
E�T Rղ���8tF�26F=�l��3��,��<i�Ub�%֖,�A��ܟ9Р��ȓJ6�cL؟Kc4�D��1�⌆ȓ��4�۶1��)9E�(tFl �ȓq���@�F�E����C�|��S�? �]�c�ˣE�0ق�\�,���"O��*U��M
V�g@�k�e�"O� �s��lP�{� #yi>���"O�s����&\��O�T:��"O¬zT A/\!A�臁TCn���"O�L�D�0�����AN�{7��"O�����LqLm9����Y8Ĭq�"OĴ0���y�-6() F졓�"O��)��$nJk�Y%x2ސɃ"O:�A�ѝR���H10 �xg"OT�m
�F$� ��<4�<�"O�Jp�`d�;1+�6|:�	5"O���F�D�W��y�$ˍ��k�"O�qQD��t����@&|>��"O�X�b�P�N�z�ʑ,��p۱"O]Q"��	ވ8ځg�,M���t"O� �K�LX�Iyg�*s��"O< K�}�`�xS!��b��Ia�"O��y�*J�F�J�A�*�)KA"O�=���7Na��y��p>	�Q"O����Q�%���(� � �y2&K) f��H�a@=mF����ۻ�yr	׽Ka�� �Վb��A2؜�y��7h�LA嬖;Z/,�r��y�,�6��h�䆋V��l�A�O��y�U�KN����ŉ}9���)�y2L%	���y�2�����=�y"�[�ut�ݺb��!q��a�A%N;�y��V�M��5�W�Q-h5$��pO�yC<g�|LQ�-�,;��u	0(N��yҭ߮\T4�H����:u��w
K�y�f�,�p�g�Ĉ�����Py��S�x�̨�6!;ID�+��GV�<qpa�~78� �K7��C'�Q�<����p����� ���s�(R�<I�(�]�N�z1 �}<x=��I�d�<	��?pFR�ZB,�'�=9��NO�<1��@��h!0�RR��x�H�<�0�J�BD�DXl6�`�n�H�<駬K!�@�
�h�?[�:m���]N�<����"wi�L���?*l�[4�m�<���]?�,�ॎ�>R��#�R�<�P�\S����rj�'�<�Is*H`�<����_�Q� �8D�ysLX�<�0J��?�Y�^$c"Ly�s�<!W��`Z`�� ��&�܀��Q�<����HN�]�Gl
K�^�y�d�I�<�R��>
���sp?$C��N�<�d���P�P�+��Zs��Y�Wo�I�<1D�ŤԪ):�A-��l�UE�<��E�1B
�ڐcP"��k��Z�<��B�;sg<��פ�;���@W�<��
�O`Ld�w��>�8��j�<)P�����Uk>m��Z"ȖC�<1U�Y;K �L;�A��A�����W�<�i�6J����p(9��#EX�<!���>����2	�A�lQ�ӥ�T�<���#
ZF�:��������2�^Q�<���M.R�m҃Ꭾr@��r桍Q�<Y��2j��D_ryҊ�N�<15L�I���4���|m^��`�E�<	��\�v�����JK����{0Ɉ|�<�'���Faԝb�$��o�Nhӡ@|�<!u���t�b�N��V���ظUH�����cx������<�  aDmؽg��ܳ�e[�����|�E���Oq�t�yW-�s�Z�31ԍ%��H��FGw���0��ջ2B�P�M�����Q�U�� �t� ֢,��JX�ĸuY��I�IF��q�'����ᓖ���T�^�H���FO�V�m�����N����l��%cE@:���
v��0 �p��^�b������+`����	�WZ�a!��\��a�tA�erZ�3�b�t�jl)��tF7muGP�)��-��i����,G��Q?`h�e@��Fp�p!�C��^���iI<���iF�����~��O�r��q��`I�r���Xǒբ�'�[��<Yr�.6�,�e�jxP)��'`q�5�%o[1Ԍr���	N���[��x c��G�*��$\N>q��Cư����t�2`��/HN\�� DL;z�EAWC�|����i��vv�a��(��.���a
�FIy¾i�l5B��˅75tA���a��o�)p�L���	uh���"H�E�g�$9o��H@�֍)��Q�':���c�Mك"C>Ac� c:8�soȺ6ޖ9l��h���n�OQ>�u'��K"��g��9	��E���dbM?�xr�N��]�%�A�A�v�x���y� � I��=��K�;�H�2��-�yҩ�o���*a�M�g`���p��&�y"cK�W��˗*�6\2�"�� �y�
"3b8*�#_�YR�I�IA��y�g]
�4I����P�N4���
)�y�k�(֑��2Y��ԫg!� �y���1a��ې A�R޺���
�yrFD�ǞQ��.�MX��X�� �yi��;idH[�� KH��6�_)�y�`�24,��+���9;�.�k1E���yr�P�sXy"�
M�9Z(���bK��y"���R8�Ce2ئ�@ *C'�yR#��[�l��0�L�.V����+�y2�'!���P揌4\�|�&cޱ�y"�(��⦇N<,��9fή�yr/ɐmhh�O��*!L<�_��y�'ݑII�P��$�rXJBa��y���(FHzv�"d�S%���y��^Pl�Qp4X�[a`2`1�y� �SVa��J!S�^q����I�<�W�
�*�x��"W�
���N�<�w��nZX�t�E1�p����A�<�C$[@ǒ�9f�&�����^I�<�k��V�xm  �$pT��(HH�<�LŹP�<q3G��L�T�5@DA�<��ȅ8z7�� AQ��0��D�<�v�>��£@�3��$��@�<�A
�:JtF1��I~�$,�A�<���T�4�p{��r��� �^T�<�g*����� ST:=!GI'D�`��#Q��2$֯R"�0��8D�LY���`h4$�3'Q-L���#$b;D�0˕�]&'t:t*����dD�9��,D�\k"O�Q��ak��
#m,�� b.D��0�T2�Lm��^I�l�" 1D��YS�U=*r�y�R$̋.��Z��-D�tQ��­`�2D埦��xK`�1D�̉�C&r�H "f�m�xpC��#D��yR.��3�y�4K� q^
�8�7D�|�D_�etȹ��\t0�]3�$*D��1JA�qJn0@bQX|a�f3D����+ə+g.����:�n�p�k.D�4�S�Nnt�D"T�Z"4a8���!+D� �c�u2�c&D̏�&�
� -D��z�?�4��-Q���C�)D����jUE��x!*^)�ڸa�d'D�XH�B�7q�]c�-"GK�l�'�&D�$���Q8?��T�R0�i�ed'D��$���&��d��O������"D�� ���O��Z!�L���I�t��"O� I�蛶r8ndj��?)���"O@��#�ȊC�m��b	���"Onp)��LE�����A�̰�"O�� "a�,���è��xt�T"O�%�D�
�\����!�R��2"O#�H/{VXz4��]�%��"O؄!S����0A�K~xt��"O�@Ӄ��9��Y��D[�'J4�1�"OTcClX���1�T��)X�"O��Ptb�u��,�7��-w��sq"O�h��NC�,8��蘝-�i"Opաsh��!���cgN�&���!"O�� L�dl�|a�*Fм]c�"O�%I�Ȕ� ~�@�5��j�a�"Ob�Ig��Sk�q�dE�.�	ic"O�]��H�m�uI�A�	��x�V"Or�H$k�cQz9�%���u�B�AR"O�5�TiR�Xq蝻�Iϼm��Ф"O��i�郓*����ӄk	RqK�"O@IH�IS�P#JL�ą�/��"O����H�;j�q �dN�e����"O���#aP����EF! İZC"O�"g 2%�A���@�"O\�
�C�[>��� �І�2e(�"O�Yef�#n�Ѷh��wT���"O�e��S�aufq�M��eR���"O�j� <Lp�)���<'M�xx�"OȔʐ":-,XU�W%YB�$ �"O2�X��\2c��yc�5J8�,9&"O.c��U������Ĵ��P"O�L[��.dk�X"v��0�P�"OD�kX]�n����RX�"Oܔ��ፏ���`ťS*.hڕ��"O�lqf$A�q���%��}�<""OЉ�MC?g�v��GJ�k;��d"O"`i`g��$��z��+} (�I"OV�CcP�a��C�����lx�"O��!n�i�9"��V�v�Ь9�"O�I(s!�z�F�f`W�+�z��"O>1�"�E�_٩��7�� �"OR��a�=X�qx���,2�� b"O�HC#�S�an�H�Q���e����"O0l��n؆+��PQ׫/�9��"O�l�S�V�5Q�r��R2��d��"O@�0v(K�{�j��3AO�;�8�s"O:��%�ZP��{vʈ.@��"O4�R񤅢Z���0�)����Xs"O�0�ҩ^;uRJ���m���""O��׌B��>H�f�]":���� "ONa��7�(� ��#N6A�"Obez"@��l���h��8HH<��u"O�lAQcX�#��tт
׆=tua�"O<l*h�<'`�[�jA!d��Y"O����e�b9 ����A�k�"OL�RL2m�,y���\�
�I�"O��B#]%U���&ҦV�~QR�"O���@`EU0�cpn����"O��p�O�|.͒ @��?�8I0"OFv��L���o 7Qnn��"O�x;�(�s��q��H�9kX��"O� Q�\���!�h��h�@�"O�Ԃb��6K�������`_��"OZ0E�W�aK�ebF� TL��P"O� @��ҬW$�����4�m�"O���k�>#�����-A&�ဦ"O�Ѳ�_�)bB��`J� �.9�f"O�-;2
ݻ(�BP��Q�0�ҨP�"Oʵ�4[�2� ]��NРs��pz�"O��2o�j_���P�����`"O�%ӕ(�
A]d:�gSB�|���"Ot]+�t���$\?uzv��"OST
Ց:#D-ء�V�Htv�u"O����Ѵ2^�"�#DpL4��"O����/3��УE#[?�J�F"OҘ�F��+J0�/� -(
���!�M/ ��1��H�GD�ᇈ��q�!��8b~���8
�����h�!����mD���?XM0mց���!���Z�"DZUo^ g�ޱ1�BVc=!��/Na��U�-�(e����9 !!��Z&~�y �\�0�bRC�X�!!�DԨO��y1��>q[�*�w�!�$�7I���V��28��(c�C�(�!��)4��q�0g�L���� !�$?c���1�܄5=��#c�.v:!��˖T:��DR�R7|���ᘽ �!�� �.MI`�1f���8�!��V��V�Q�	j`Ȅ��n!��S(PTp	��$؍H`HR#���c�!�N9%Jʉ��ꈷ�֩	tV�N!��T3D�,��.ݰlS��͏)L!�]92kliD��/�%r��׋;!�D�!Z�u��8*�� 
�� qơ�dM!�z��5���'ʙ�rNB�y"��$Ȳ����t�Dh"c���y�f�?�A�u/�]c�L�1D��y�dϖ@���'H�&r��M��y����O2�\��/ێ!�r]�oP=�y�)N>p���i����l�����y"��x�X���� ����ʌ�y�ƞ�^�\[u��)��!�p�V��y҄�<Lt�Ac��J�t7� ��؜�yrV����1��d ��j��y"
�h��Di�d�D�z��W�_��y2O�'=3xL�u�J�@K�4r���y򄐀.���{牾$��\H�����y��E5,�v!(򀋐k0N�Y'�L0�yrDHӒ�	�G �H��3c�r ��B��{�kG��ȳ"�p�ȓ5��5�5��k�����ށ��fhz����[=[��3/��*o<��ȓ/l�i���D("a �߲����ȓ5;��m^���Y���YAn��
�'h ��B�L�a����I�x
�'Z�Ԛ���.{z�I��F�G6��
�'�D�Y F���1���V!M�>��
�'Vx����.'���ˡ�ۅ����'����X=%��쪱ٟ� ���'oX%؃�P��Z�W���
�'~���J�h�J@��R+<U
�'�zH�@�X(&�u�� :�̕�	�'¨3@	��p������2A��z	�'�:pBDD[�sN��4��%5}����'�2�ӏܶ8�.[*�ڨI�'��i��c9!�%oK�|���
�'6�()7�[@���5�ز	B^��	�'NF��SA��) ��O�Rk�Ѡ	��� �푶�a���C�
/+�4�"O�1*dmD�j�f�KC�V�4�v�I"O0]�5��/���	��ŃV�ƙ�"O����c�L��Bԋk��Y'"O� ��Ŏ@lܭ0�*Z�8�Pyya"OP�;��J���1a��v�����"O�����)|�ްQ�i�d����"O��!���z�������b���"OT �E��1@XL�u�]�X��XS�"OZ�a�C� 5�p#�iZ p��@�"O�U�[�h@8c�I�?�N}��"O����F6Y��a�H�%�(u�1"O�A��I����s��?P�蕒�"O���'��*F��J� j`�"Oܨz���U'��k������E"Oh�����ڍ�jس�H�XS),D�ܡ�*�<r�x��Ivt�7C<D��9��-vR��4��-p�B''D��ZW�Y��у��w�Z��� D��2Sْ�@p���	� ժ"�)D�4�üb*��
՜M��4�I)D�p�eƁ�Ah֘9�HԡGg�$ʷ�&D�xs`H&�^U�ŏK n���H&D�̻���(�\�q���4uh��Q�%D�8sbď-QT��b.W:R��?D�
����x,��g�qDVjw�:D�8e�j�L1��ўL�2��5�9D��* &�vd�'J�6t�GF7D�L�&M S����
����6D�4��g   ��     	  �  '   �+  17  <B  eJ  �V  �a  �g  Sn  �t  �z  !�  c�  ��  �  *�  m�  ��  ��  7�  w�  ��  ��  ��  V�  ��  W�  ��  '�  R  z$ |+ �1 8 �9  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>b�ږ�;K'DT`�^��@�IE<��T	�����	Z��(9ŦL�'�b��
Y�<ڥ��-QANZP�[�VB�I"��9��(��0�Qj�)!�B��<�@�'6�HiP ��N"�B�	� )*�X>2B��!�@�,FD�Ǒ��!����B��ID�x�fφ
�nB䉺V6|i6�]�zq���3nL� �B�?nR�R����|�� J��^�>�f�'���t�)X2��r0f͇ڬ�x"$��y�@M5?�<aU�W����`��y�b�����Au<�l��i���yr[�(��Q��;���H�ѝ��	ٟ����',�H	b ۷_|���-F3du����'H2bD��(`�̪�9�� P"�y��l��!�t�W�����p�����O�#~�!��H�Ī���3"i�Pn�B���HO�➠Z���;ܲ{�*W�1B���LF{��� ���GEȓcX���I�c����"O����Y)u!�5�������D7�	P�'�^Ʌ� ����r&*�%F,���'@r��d��4 � ���/K�`��n�<)7�)�'b0�Ȉ��[�\X��b�/��<C�Ʌȓj�
AP@�/"��A�_�su¸�<��)��#H��D�Ph�?G��ҤL
�  !�D�O�!��-��p�NL�`�w�Bx���I����,��v|�G�7O��`��	�L�9`�gO�J�}����i�C䉳U��X�⯗i4]�ej؁uR"C�	%u$�`��x�F�����@����$?�	�N� ��t�Ⱥ'\b ���H�$�C�,i`>@"b-��1���	�~�c�(G{��D�� rCRX{!BQ9��J����M�'{`s�
F,�X�W��{#B08����^ܓu�����H%���in\N>6��ȓB�0X����!}�	����o�>��>1�����L�V��ik����sQ�DzVǅ��0>��6}g�x�(���G)���%��y�����K=tXX��Ђ�_��ɺ�'������=R��l�)R�H(R�'�|�k@蒳d���駡�R'��	�'��8T��D�b��?0
I
�'�~4�� �@�"i�-���"�'�tY���<]�i �$/&��[�'��8
�ʠP@Z��#�C�#���S
�'�и���5"Ĩ`���$"��Q
�'����lN������)G&��	�'�$5z �88�(�j5g��LMv�8	�'�m��
�5����dO0D���'�Ԋ%O�b*�����3B
12(O���I0?/*��C� Nb|�Ȗ�[�9=�����<Q
+Kt2X&+�'|���X>�IT�)�?AF��0E����IK�X�X�z� @؟��~C;�39�H�W)-{�����? ��0�����ʆR꾙Q�R��hO P����X2�.E�X�����v�ޙRw"O����Q7!�ib���u�j�Ӧ�'��d>���'!T��.F{��#��Z�މ����?�4��TY�f���&�������y�	MA��Lj�k1T�L�&�J (F<0�'-�	0�?���)����qzq$��<X�*V@G9!�$�7$*D�{�g�<p���U�	1���j����F
+���CaL�2(`Xp/D�����K~Hc��<@<-�� "D��	�e� - T�y��̸k*
Mhw� D�(�@�&�(�t-�~���  {h<��F���4$k�+O�#��0�,\x8��Ez�M�'m� ��H��V��)'�;�y��W�*�8�c�M��aQ��H<�y��E�cw4P� �T~D�;�O���y���1C\�@	"ޣ`V��1��=��'��{�
	����ˑ.	~�1y���OV��G'BW�	��M*�z�b�J�z�� *�ўl'�<��Ģ�se�X;� 5��F{�4D{���k�|a5.I g�����.%�E�2��#<�	�	�d��L�!օ�E ��� �ON˓��d �T?����%�=H�n�)��XrOW��0?��O �q��D�]���p��A]�L���i*��E��'? A8r`��.��ň[=%����D�\�O�r�&�R�l�u�@�zm�<��O����Il�婲冲~�X1k��H��x��v�����p�@���E�"K@���Y:!�� !�/ԥ: ,�%M��,6�Rc"O�e:�h�X�d��)�"O����I�8 �$�"+A�X	���B"Oz9K��ӱiǠ ք�W��2�"O.�%hE>DR�P�\
?�4���"O��4dL咍x0c�0}�8 � "Ox�bf��|��dZ��N ՜��"O��!���b�&��סM�Z.ʄJ"OJ��#1�%�A�<t+	t"O5����. ���ρ�DT`�"OH�k��"6�@�q�-��W4@�%"Oj��AD�#q���0$�Q�#�<��"O���v��x�b��ޒP�����iw�#=E�ܴR���ț-3�hTp!�B)E����iL� �ڻ}0J�3&#�(wa���=�ش��<yF�"Ap��2�ܵ~� 5�¯�C(<9�bՕ2&�� ī�n�����O�aA�]1	�'�x�;�	C
+L:$i�Dޠ+`��	Ó�M���$";��=rw*޳��TQ�Y/!�DLS��\���M6G.:XfP;Y ����ا��ҩ�BD}���G�6f�` b��y2�$*�,��5��!p����Ь���<y���<��-e�x � �t,�A��W�EC�I=dqn��c��@�py*��Yj>b�\���)���CB�Ã��K��j%�J�!�ā"]z��Ѣy�PՒ�ټ,�أ=E��'��L���b���P�l�q�Î}��)�IDr��b���3n�y�tfRR�qO���Ĕ�n�Le�P����$1���sn!��r�`M�0�X�DwJ}#1�\�J�!�P(�pT!� �3�Ș��OH%h�!��}��[%!�����@d!���Q�����|�p�3	�!�O.l_"����X�6���"�4�!���4k-� 2���(9q��$%!�d�9Ey�k�(ґNp�0cʓ�!�$K"m�fH����Mbv�B'B
�n}!�D�[� }��a�:��Q�b��@!���"l;����C�b���	�N^)P�!�N�6Ҹ��^������.�5U!�$CV.̨��iډ#wh�G��qO!�DK#%b8�#҅*Wp���-�@!��͵t��ɋ� LD��sG]$2!�dХl8�v� �~�)�f\�f!�d_�C,�<c$�<l��ϑ0!�H�~m� "%���*�r�0�J$J�!�$6B $��d�
�R,9B�	�`�!��`q406�
1ͲP'�a�!��	$$V5�� �Eˆ�B�DY��!򄔳'�r��u�S\�"\i����G�!򄖚{��ltmP��e)��± >!�B&����U&��w�`X{6M#S#!򄖴^�8���h��vB*�X3d��yl!��	f�
P(O�.'��xV┫k�!�CF;�0	2Ïzњ���."`P!�dS�g��i{@jž	,�ա�	�MJ!��̄�^U"d�U�.F
p 1��!y;!�D�5��%�U��>A&�	���S;!�DC0t��L��`9!֬�L0-!򤎫R� +��1	j]p��b%!�ĉ���=���!k�Q8��S !�đ���Ha��D���<��%�^!�$� $��[��?$��!Z�e�!�D�5 l���'K�*�}("$��!�� DԛS��W�����Oq��E:�"O<|��$M��p�lB��0�Q%"O�EA_ zJ��@k�+��yW"O����J�(�D
F�H�@ۈh�"Oc M7ސa���	R�z!:��'��'�2�'���'���'�b�'�z�8bH�!ΰ9�'���?�����'��'���'���'���'�B�'�Ҭ��苆6��T���	FYz�*s�'�B�'WR�'�"�'���'x�'������J_}!��9i�eI��'�R�'$��'���'gB�'M�'��L)Î�$ӤUaGϛ Ŧ�:��'���'���'�b�'��'�2�'���DO1~K�]+0�\w�4���'���'P��'���'d"�'�R�'���"����)N��"^��?����?9��?Y���?i���?���?�G�*�����N�3����,�?���?����?���?Y��?!���?�� Y�$�j��ʌ�1�(��X��?���?����?����?i���?����?������,5���H�N�¨�4�R��?����?1��?!���?���?����?�`��`��� ���3���Z��?����?���?a��?����?I���?���c]�X�րI�#\�0K&
���?���?���?���?Y���?���?�&a�=]Ͳ ��ڧ.��{���?)���?1��?)��?Q�q���'#r`�
v�><ط!(^��dS4 S�����?Q*O1��Ɂ�M��ғ.�r�jp�F�c�&�#��	-'��-�'B7�<�i>�#�MSo�0/��`��188�����[=U��'̄ݨD�i2�I�V�JP�����''[()�gaE�`������\���<�����?ڧoT���*�_���Ʉ:�ly[�i�T��y��I���݈mIn����3P�:���+:-��޴b_�&5O��Şgވ�Q۴�y�E��~��%P���G)�Q�̈́,�y�)Z�2����"ZA�ў�֟Ċ$��L�d��!�]��\�!{�<�'P�'�X7-o�1O4�kMZ�j=�4���Jn�4(i k#�I1��D���b޴�yBW�౵'M�Lٕ�ڍd���3�+.?I�+˶^Q�I�h�ḩb[©�Yw�����H:���D���_�y�J�Hj�˓��d�O?�ɯ%�����#��*@		�~����,�Msu�PB~�g�d��9f�P"ᄤ��#��]<�扱�M�³i��gۏ;#�6�� #I�Y6l�S�+ /@/ P(�(ݺ8�(1kP��9�,���̙;�2�`	ߩ1B�c���7qN�,�b����m*Ѡ�39��s&��o״ �5+�:O¼�ȃ��7=6 ���`����JƋ6|��bďJ�$<�g�	*n�<8RKyyR�ީh��u���@E��@�3\���V��W!Zё��S1VLLC�D�x����T!G&D��B�9d�Q*��?�\��5*O��Av%F=2�@�PPJ۳k�*��A��oKZ�����	���/D���Y�'C7.�0,�����&t��z�Ԥ���9m��+��/T�]ӑ�8�M���?����0��\�tmѼ	�0i��*	 �gӬ���O�`*���O��$�OV�����O
��J�ʙ�q��2��?3,Р��4�Nm��i���'���O~�O�S�o�Ia��պlr�Y$-)��4l�k@���0�9O�����7>t�Y��G�B��iQqL��Q�Լm�ǟ��I���[�*� ���|:��?�@FP\8����?T�4��1l�	Ο��I�u6Pc�T�I�p�I.�65�c���084)���m�T�z�4�?��IC�RF���$�'�ɧugm�=���SR�1&G.���ۢu�1O"��O����<�d��5(��˲@�0(^�%j	!x�E�xB�'K��'X�I�(�	x�Hi�VH�+|��xk��ʊH�|��@3�I�����˟��'�ڨ�pgn>�[`,Y��``F]�SZ�X��K�>����?������O����S��u�D݉��η{f�!3�ϓ x���?����?�+O|$�&�Qs�1Q7hp0��K?���k�=,XҔ�ݴ�?������O��$��jt������L�m�m�#�ќ"*�t���i��'}��2�*eCJ|
�����Nִ�
��]q�9+Ê�
"`n�vy��'���\��O�"��Mc'AD�8�T;ҀRtM&�H���ަ��'R�ò�d�>��Of��OCJ�BɎ�bB�F>�����]b:�m�џ���>�L�����'	�D���Q[�E��5{Dt����7�t���4�?����?��'!0����GZ�W����D��6Q@��k�3"7�7Mφ\���?�����<���%皡)֥ľY+f�E��6d�
PKԽi�"�'�����`a�O��O��DR�F��Ο0��	B��i�'���'��C�yB�'	��O>�`�
r�V�U3=�4 8]�@��iJty��'-�'�qO���T��N|�����>E[�U�8���Ŋ/v��?�����D�O@�CᎳ�9�f���8j�̓�1�ʓ�?���?����'m�tH�(�b�B��#L�g��h#�A¥~p܌��O��D�O�ʓ�?��X�����N�(u+qK{�H0�/K,�M����?����'r��NJ]K�40t��6k��	��[�Lޤ��'%��'*�	��|r��Yb���'�H�8����RR�1�V�Ailӂ��>�	П������:O�!����{6�I ��wx�J�i?�^���8ֺٕO���'��tU��3�YC¼}�R�L�9,c���2m��ݑ��3�~� ���(U�=ks��Zg|��2_�@��� ���	ҟ���՟���yyZw\���J�)G�\
RI٫O��d�^��g�����?3�T� 	�',[�M�!*b�V� (��'
"�'1��S��S՟@�Q�ێ?#h,�t��,~,�/ҏ�M��i:n���<E��'/�,�2,M
{lU�O�&��Y�CO~�����O��Ď�%m���|����?��'ν�V+��~QȌ@��^��xb�#0ӉO��'I��ƒ_Ti��>�bt`�icm�v�'�����V�<�����	_�<�j�1���|܊��G��nW(�%�� R`+?����?I(O*�$�rv�E�_�u�jC� ^�mF���qF�<����?���'��DG�oM <�өK~�R��b��FN�B�;��D�Ot�Ģ<���d6��i�O!^dC	+~����wŁ�p����4�?!��?�r]�Tz�z�v<���4܎�3��.I%��R��	ʟ��'�R��Zb������-׉�Q���5��J�O
��M3����'G�	�J|�O8�g Ts�		�$MK��`�@�i��W�\�I� ��ݗOh�'Y�d�@. X={W�r�@!y���Ai��>����iQ7D�S���� ]W&���h�K4( �ʖ�����Oɳ���O(�d�O���\�Ӻ�0׹fU� �$@	ʄg\i}R�'%���������O#
��7/�=����l�'_鎰ڴ:ܱ����?�,O����<ͧ�?q�oΑ<�v�@�˅�e���W�P1}&���܉��DK�y���Oj��NQ	M�L�P�A���!# ��̦!��˟���Ε�����'R�O�uX��	 f琰#`��>r>�)��N�x̓(�"mi&����' ��O"` ĊA��\���Z���Q�V���ʗTy2�'�"�'BqOt�ʠϜ�Dc�P��� n�Z��r_�2c�C�R���?y������O���杅O�BAр.)I�V��v# �wx���?A��?q��'	��JpʌC��-��K��@J��BۼX2��O����O"ʓ�?af�]����%��H��K�F#0�"�a�	�M����?i����'����A�*�r�4?f�B7���Xpy�LM�Xd�u�'h�' �̟L� ]K�$�O����$��� `�N?����i���d�O��b_�D�'�np��O��SsD����-.��&�'��	���iIDg���'	�O��x$$9�U0W��,fq�C�.�	Ɵ�\/�c��'W<.՚�"��L*���䓱�ک�'�2�O*��'���'�T\�֝?*��rM�.[����!@�H���?����~�8u�<�~b�G�[Z���1iS6%(#�Pئ"��Iן,��ß�	�?1���T�'�!rM��.���K��%M���C�t�ܵ�fE��v1O>m��:)��b��U9e��Q�*�)/\5�ٴ�?a���?!4I�.��4�����O��*O�$����l-���R�V'�����'�"IZ�o/�i�O:�$��Ģa
35:�Y��˛A02 �mj�&���1^Z��?���?�{Z�,�2�N�� q6,�{+���'�p��%�V���O��D�<��A9t}Z�h��
f���s
�h���"��d�O����O���	s�x�֤�x0nL1eB��}+><��eB��d��?�����D�O�)b���?i��ɯRrI(������q�,�d�O6��8���A�c��;%F7�ڦvP�%���^����"���1N��	ן���Wy��'���C�S>U��;({Vf������>zP�i۴�?!�B�'v�yǈ8�ēEB¦�2�.�e�P�JԾ�mZ��0��ş���t�$�4�?���?1��X H���j��u���yiֻi!�R�$�	{>���˟�����4i�}*@Z�X̼�c��ҸqI�n���L�ɼ1o�� �4�?����?9�'�:���x1��WU�{�l!Ǌ��W���I� 8]�	~�i>]��6ܻ�#M�UB"J�48�ub�izj���|����O���៌�I�O���O��BQ�ݏur�/�nɺ��4EԦ�� Ο�&��N��؟��F�{b�*WDϒK����"���M����?�i�B�2��iQ��'J2�'�Zw�B�p��C�d��BQ)N"X�x�O�˓u�,����'�b�'7\L�fT/}[z8�!��x M��p�����V��ilZßh��۟8�	>�����p��D[�rn�Ң,~"�BD­>�����<1��?����?����?9��.SVl�RK��h�B�b��i�����#Q曦�'���'B"˼~
(O���G�UWn����l�PIĞi$�|�C2O<���O6���O���lȃCǦ�h!�ܚs��
c������CJ�M����?i��?�����O*e9�7����!�ض)[���0�o���G���������䨬����a��Ŧ��I̟0۶�ئ�⵹B�E���g���M����?�����d�O����3�����8���
Jn���)®K���	5�q���D�O<���O�(!!�٦-�������?�"�-X}����.�&�'Ȯ�M�����D�O$I��=��ʓ��i6�e�q�܄:�,���Ƈ�E���4�?���nM̬d�il2�'�Oz���'�`d��+ج�4�)���ajbx�WD�>���R�Z��?�-O�i-�$a̕1h\aPEm_>�zL��>�Mӣn�.^����'�'�D�O���'��f̨sʜ�2���Q��9�c�r"L6�� �B��Of��|
I~���C�� *a(Ĭ���d8�D�7<ĕRD�i�2�'���V0Xr.6m�O����O��D�O�.�(B!:�RU�W�|)rmȧ���	jy�(��4����O>��P�e hps+�<\��I C��4.�oϟس鞅�M���?���?1Q?y�y�b���ː7*�����ݻB[(�oZڟh��~���Iş ��⟸��y�TB�8r�pA�-ŷ2\��Ad��=��A)�HlӺ�D�O���O4��OU�I��Ct)џ:�ĭ�HN�y�ؕs#٧W%~�����Iџ4��՟������YG���M�S�,Ux�p���LP�e���z����'b�'�B�'���џx�t�{>�� 2*Vl�A�'� �B`hE�Y��MK��?I��?�V?����M���?F�2:lĵ#4,$h�����m1�V�'��'=�	ş$U�w>�OqSÇֳjEd`w�@j��z��i;��'�R�'b�J&�oӨ���O�����VM�*F�9����-|u2�)�(�0b�F�'d�	ɟȁ�K`>�%��s� ���f͞4�@�Aե��j�@+��i���'�����rӜ�$�O��$��*���ON��
�8G��$kc�>e�`t���N}R�'��,���'��i>Ť� U��
�)4�f��`�&	Є�ƼiX�鐅Kz�r�d�O���⟀D'�X�IVmDS��'0u�ׄF
w.�Pߴ<B�Fx����O�)s��30�p���5���9�HW�9��ߟ��	��6	�M<����?��'}(0�b�ڴ}<-rA��]r Cݴ����\	������Oj�d�Ok,4+Վp C��5j�!T��>G��v�',*��b#�Iӟ�$�֘�ab������xv�[�~�
�r�>�������O��D�O��'��e�/FR@s�o��((��?,]�'Sr�'H�'Rb�'5r��B��/�X�G�ޒ?�����#E�'���'s\����	���􉃹Nx� ��j��M�(�0�ē�?H>��?Qc���<�I�0�B��-y�x����.T�I˟<�	ʟt�'z��=�	ǟL���!R�F!�P�B��#���l���&�(����+�,�ޟ��O`0c�Ĝk
��Bj@�Cw¡�ӷirr�'_�	*�rJ|2���ӄR���T�g�[A(Q��K����'�"�'�
yQ�'��'>�	C,8�|�j���-?b�!����x�W��q���MˀW?9���?�z�Ob�&�!18����I��9����i�2�'��4��'ɧ�O���P/�~���:5䛽z'���4H���9��i�r�'�B�O_�c����K�h�@[$�P��|�v���MS��9�?�K>����'5��qŁ��F#x��%P=`t:���`�D�O������'��Iԟ ��@��`��4V�L��$:vuo�I�ɀZ����N|J��?�����[1R=4���ň�>��]��i*�B��Zc�4��Ry2��5�%�W9f}��#��Wάx�F4����
U���<���?����DN�6j��6dG>~
D�R�Z)�u�1��^�	��X�Iw�I��\�ɣ{I���a�ђ��<P��?x���Z`m[���0��џ(�'ئt�Ba>��4$̢
�y�$`��� _�8�'2�'9�'"�'ch Q��O@�k�E�9,e���@�Π`�S�|�I۟X�I{y����D��m��dٝ?��H�ɉ�d��"��̦��Is�Iß��	� wZ=��R���*p�8C�!�d��PaG$v�F�' 2T��ㅨF��ħ�?9��"p0I�0i����Y�l�/k���x��'��EY� �O���N�� j%������6-�<�)�=i����~
��ҁ����(M5�l�a犁
��ъ!�>�I5������?Y,O��)ҧ	ոF\TȂք
?�`�qP�ix� ���k���$�O���Lq%��S3M���y����4���M�PH��4(k�Xh��?)(O>����G�R�aKϰ]$�ܣ�����4�?��?�t��y����>٦̗yPTi��	2{���ڢR�q�'O2�[��
���D�Ov�$̗��c��9z���Uc+T���'��1xS_�4�'�R�|��?F�( ��8#�����(Ur���\���" @j~��'���'���'}𴩑(3f��c@.UӅ�W�ES7��ON�$�O��d�c��y�3~�h8�
���ʱ�ӬsD��ş|��'hR�'���'�F�b�'�h5ҀΟ3q=jYE-�r:����r����Oj�� �$�Oh�A�ʥ�S���)q�>4�ǎ�b��!b3������O(�$�O����O�)×��|"��R�Az�A�8| `+��ii���i���|r�'�Ba��6���kO<� .ݡj���.��.��cY������ �'� ո�0��O(�)�!^�����8?b�� ���dnZX�=�L	F�ܴ"��LP�A��~Tʶ@�
1\	nޟ8���U�<�������	ßx��KyZc���@�^�?�4�+�H�:��H8�4�?��42=·hj�S�)��롍O�>� (���\,v]m�$�)��4�?1��?��'9��'��	_+N����F$Q��)�S[�7M83�"|��7Try��נ2�x$��,X����¼i}B�'�B�ʴx��O ���Ob�I� �$�������Q ��+(S�c�t@5�&��ӟ��I����$�[`ي�A��O�O��a�+���M3��]�L�)ęxB�'�R�|Zc����$�AdQL�s%�$>V��r�O�ȗ��O*��O&�
_� RP r��Zan�c�	F ^T�'��'��'��'?L�H���qӠ|��$M�g�.���g(��'�"�'"]�0�rj�%���B��y�<8{t��i
�� �����O�D4���O ���'B����`l��saj�q$�4�����6����?����?!,O$��d�YW�ӛ( ǩ�m�b���Q)u�8�޴�?�N>y��?��JLg�;7PaJ�-N�RF���W��7�o⟔��Uy��@6��D�pa����r��s�Ҳd��bFo	V���	�*`"<�O�h+�fB�M8@��E��> ���4��d��N�*�m;����O.��_~£	�� Ū:L�T��+�0�MK���?q�O�s���OqF����f҆xk��]4'�&Xݴ�PJa��W|���V��p<���**tz�0E�q�M��aU{�<9fÅM���  Ɖ6hV�{�LF(jLtq�k]	t�8#&����TǀY��E@�Ŏ8t6&<�NC"~d$���+W�9ك���T�2��
<�P�����3�С����"u\�c@��!C�B�yj00�$\����
� Lj3�� sv����wkVQ��K�!�DQg�:�?����?��r�S����'+*|��c�0H0�-6<IQ��F�X~�xPF�5�p��e�׬d�=�Mc�*�TY���y�T�tʴt
p�D(D�:��&j@�La��:2��T�l>�p���Ï�xk��DI�%l�����t�ߴc��F�'�����?1�K�<��3�a�*����G�[J�<!w�=���&�''Ҩ�:SÝH̓L-�f�'��ɰ3x�j����$�	1L��4C�:Mf3���o�����O������O��q>��w�ԲMK�23/P�Y��oZ�>8z�Bwm�~~��7J�P���#>&A RE� y)��
vA):骐n�'L80 �� Zw��!��'$:a���?)*O�����,�Ċ�����*|O|�E��r�h��J�$ɼɉO��n�-����j�N�ȅ����7c�\	�IXy�c!tٌ6=���$�|���ب�?15"أ;�"��$ 6Z�~�+ a)�?��ܰ��(��5v���&���<�"T�)�ʧ;�d8e䍠N�̑	V��!1�4�O2%��J`,��)&!��3�B��锤��`F�q&�] aٞ);B�L�4	��k���m��'n\Q��?���I�Oj��ȕ�$Ȋ���^(9���"O��*C���V~E*A䛶��q�4�/��|R�鉖T�N�+�㏳`<� b��4;I�YAݴ�?����?)���%W�ީ����?A���?ͻd�B@��H^+�ȺG��#?�r)��)=�+BFӟ Z�NA4nx�c>�O][T��%DN�5B�������G��|�ԑCt�!�N�G��}q�^iZg[��TK�5{�|S_3�J�sA�i7M�Zybb���?�}������I��ZT��Z�1D�"S,�Ear�34�T��/I�T�����
�"���'?��)�(O~��*M�P��g ]���'�@�X�H�_����O ���O����?����d�ۺn�:�y@
B��QZ1���UB!�լW�;�� ��R�"��y�	�L�ȹrd�pi��0*<к਷��"�e��ּ0���$[�7�]��$�2D�(��e��8��L��'�"�'_B_�X��r�[���BS��&/�e{��S�F�Q�ȓ�T�3w�Ji���F;(~�E�<IsR�0�'cJ4�Ƥ>i��G#nt����=�^I�3`NILl-����?��ۗ�?�������Y��f��Pf
"��#���E�~$�h�m�M��
�` ;�ɠjb~
��.�谋��V>+�
����	�]�����Ģ6�"�%�p�'pj�J���>aD5�P8XB�]�В���P̓�?�ϓ �&9R�Xi~���b�ʔMgrń�_-�vCI8�����5K�@	2G���y�W�вA�ʟ�M���?q+�-S�D�O8�c7������A��B�/1���Q%�O����T��a`��/U�4���J�V0]G`|�ϟ�I�R�_ u�}��䙥g���I����ųbt�2�c�+y�h�Pc���~��ז?��@�� ^59TO�>p��spL$}B螘�?����'��S˪h�@LA��8aLK3��p�<!���<�k�#a���fL�B�(�j�Hi������M�Ey�))5��%w�9J,.��P�'���'�(A�%c�>:���'j���y�-����(�G��D�BB�D�,0�ތx5DO����'�9=#�}��I>�@5����$l��æF3ԜP҅�(w�H���o*�P����n���&a���	V@O�i�v�!Y�*��)?�������S���?�gl7U��cR�DC`Lb��z�<ybH	�{���┈�M��Q7��J~2�.�N���byRe���A��\� �x�B��D*
�����a��'
��'̀�]۟����|��ME	;��yse;~E�%jHA4�h@��2���c'n�n���B2t�<�A��d�(����~���'�Xq�,���W,�����D׈Ai���]���a�+��~�0�'�@A#u�M*b�7e������ȍ��?1�i��O@�d�O�X�wJŘ5�hV��4-)ԬK�g<�OؓO� �� T!K�G��$��k^�E~T������Ihy§��~�7�O���_�9�:�@@���y�T�ȵ[�|���O���2H�O���{>�Ic�@�;�6����l�9	��ӛM�BP�d���%q���R(æ9��D�))g��hpi˸�*��&]�z]��PeD*uנi�q�D"�D��������[�����4�?��aɔX�"%����q^ �-]�����Op�"|JV��?p'2�	�&�?�.aQ��[<���i���P�ͧ?b�,y��^� ,�s�'��	� �Ht��|����)��}��ҽK��s�ϗ�;�.� ���:R4�D�O\墠O(b52!@�%ra�mr3�!���]>Q�4a�	@l1�f(-\@�C��4}�ܪm�� ��J�=��Hr���r���>Y!��	r�.U�%�X�	�p]�"m>}�+X1�?����h�����/?`L�-�y�ta�e%�PϊC㉜^
p	�@V-�r�j����a���d�w�'��ɀ���c�� ��iЎ"��؊�x���Op�D˼}
��k�Ob���O��$��B�܆��E�#NJ�O��1��ڸ݉R�W?�@ �g� �q������D�xb(�H`�i�w僄Lj\8�C��0f�=�G@Y�L#>��W A���������x�EO�v
,��a�R�P�0�J߅�6KBy���?�}��ʟ��I<y���%!��B3( ��!P��ph<i�B�,Y҄��n[\�j�+A�AD~� "������6X�D�!#-�"U]D|pQD�&BV!�dV qf�zƃǣZ\t�*���7%!��ݜA����G'k@�#
$~!��=F���q��/4��t!�:t!�2��m�a;"�~A�K��!�DR�cO�h�h��x�˦EI�!�Ă�"݆I;�F�*|�R� Z�!�$3Q�(8!�ȊD�X�cq+2s!���nI���E��1`��)(SJP*%g!��ʙ\���H�aH�z�Y{�tR!�ڹo��<	wb�9e�0[���@@!��;we��{�n�^������!�$��X�D��֢�6)�&́�&@�F�!�$�PA��i������%���!���>&�a�r
��m)�e�8_!���k�dѢ�K�X0ɑ� |@!�Ć���%������&���
L+\!�d�gl�ЃX�?����ȗ"N�!��]�d�By�#�4E?dĢvH/J�!��G3�M��bZ�aO�:�v�!�d�7h-�3�֛]Kf�J�� )!�d�<	 t�2�|�� 1UGƖc!�ȻbP��q�O+G�<��&ԔS�!�DA/9���Z��#�@9�� ]�!�D���T�Ad���4�e"�?t!�7u*�5��/q�����a�S!�~���)��P���:�A�j�!��}�dQ��lz�,�1�ח]�!�ߢ{Ĝ�j�#[�PwZ�S��<p�!�d�?"�hфJ��[@�3�L��I�!�$��0��M2�l�1(I^�k4���#�!�d�y��E:�	�P4Э�tm�:�!��,�D�`�	�) ��sm@;o�!��©Q:�%���C��" �V��!�
{��@��N� 1��	�p�!�DŌR����u�� Q�:�yQ��#�T�*�`�7��þW�a9��O
Y�*%s� ��ɷHY�I��"Od�b�K�40�D��Fj�H��%k7JV8dM�BD8)$v�@�N�6#�I&�~�8|���ɭS�r�9CaF�5�@���9J�J����?�>�ᡇ�U��D�&aJU��t��Z�z�YQ"Xdx�X)NK�^�t��pc����b�>�x�LбV��X=T�z��pFd��/�h�8��؛M.�I &[*8J��@�"O��ٴɕ'=ތ����QC�Ԓ���LX�g�ܚT�-1X9]��}�;j���d�
�3�| �0
��0�ȓ?�N�DヿO�&ږD�wY)��儎I�>��pf��)QP�x�M��|����/QJ��B���dR�}Ȇ�-H�a|��S�x`��
� �C2��28,�rUٴE�a����d�<,���)�O$��Ä2{wr0������0{��	>&��i�U)�+!~��bBG�;r�D��Od̓T��{������G����'l:Ex%�A1�t4Pe��r����îC��
ES�FV!��(���~��>�ݗ'�%3��A�<�cG��;բ���AL,	���J��٫�'yp���$��&Te
�D;=	�$S�Ǚ*K2)hVID��䑑�^���\��CN.�G�����"M�"р��cmR�A�D��ϓbQ���eC�uT�1���m����V�W$cs4z��ٲDܝ�yB*�vG�@����H'�����/n��Į?n~2�გ�O2}R֥o���сMv���`&�|"��L��΄�':T�{�kr������]:;�y��IU�g?��G��T�|[`�ʄx��C�]NXRSNϗE�mj�A�x�ʄ���ue�#~�;v6%��	 -T�<UIQ�[h�pU�coC � ��B�P�D�G��O�t�5 �y�a��G:q����u��O�s��y�l�Q����zP�d�N�?z�l}0�)� O�)Q��C
<|��]������2��<��M�B���t��m6�� �Yb3�U�@j����nӼ�MKGd֘J�h A'Hݔ^6�L�S}J~�À}�� "�m����E� H�'8H���#mr:�@ JZ�O���F��	���c�C�pO�	E��,l��uc�<y�.$���\�؄y.O���p͌%l�\H����%Tn�Tǜ?IW�y�Rǔ��ZF��O�>��Ox��)��<�$���$�G�G�X�SU��#K�yC��^2:�џ�a��6�2��j^��^h��H��0b�"C�?'�D��ԡ&Ȍם:���ߩ}�F�;�O���hV��9�#-�9m�1�g.�&Z
f�%�'��0�c&��y�F]	J�� �H")/�����7M��1ӑ�T�O%��
^8 8|��O%�)��\�v����؞X3���@��<um�P���]�m*UKG�S�}1f�%?�R�ôJ���T�CO�YSP��e:M��)
���DQ-�ħ8&�x�Ū<yQ��r�NX"�n�M��q�&�WuH�)��"hV,� c�.r.�ק�����-�(��$ʶYi�}�@cJ��L��I�Ϣm���ȷM��CU�=��}tZ�K�JI�/��T�d��0�vq�C��]yRM�n�����g���_=$��7�S!��#����&���Av?<O�!�Ȓ�f󎀴;x"t��	݁^b���E��c�I��/R'��D�>UG�>��I?m9�eX� 5F��T�oL��a:!�0M�v�ېl�j�p#��N�ޙ�'�(�"��,a�dC#�T�[:�ѡ��2j���DFtJ���=J�>a�'�Q��<M]r�"�F��X�i 
�1����-�tЪ%�E����9�FP8��:�`�k�	P(����g�S갨�ƚ& ��d�<y�F�?Q���/��mP�	M���×	N��'�4��gO6L��� !>��p	^�6%2q��N�Y��D�%%��I�t��(8�E�!-l�mb��ɜN�*djPh�,����P%�&����p�R�F6��Iբ�?�T?yJ(V�w����P�ű+����$c6�Rd��"@�o��!s�H�#�X�'�X� �M� 8���R �>}N�p"��U.`9��jŒ����'�����4�!�y�LБn���V.ټa0�LƐdO낃�-e��YNNHdK*Oq��n^�}\<��9�8l��	�x���ͳ!^A���i����aN�?�\=��$ҰX�$�ȡ6W�0*�_#~"��X�\�Ơ�:<���ϧ;o�$?�$3S�Z�hV�_� !��ʟ��0��&�P� (�8/�x�cb� s�ڐ ��"?�֥��L�q.H��'? 0\,�GgMJ4�z�4)��E��M[�
�"��"����4/ �a��("�^0{pzxR� R��OA��`N pC��S@"�� v���Z�P��P|�c%�C:��ZSg�A�	���@�8��G�q�8V�5��2�y���h�yӧ^�U*"�(�$Ùl���h�.@�w��X�*���2�˒S��>�."z` h��E͜Kp\p�� � ����ͻ �E G������考�I>�5��A�c�/#�Xq���[��9o��l]�aL�b��S��<_�٠1ŉ�����Q�>Q���#�����y�-˯f�D�����_�j��:�<j���H�҆/٭!�)[��ރ��a��(͓�����:I���x����G.H��c��	�`۠�+�O�òI��?p��J�m ��|�;AL]j��� ��_�"ZP�S�� i�%�0��!	�"�	�u�J�JJD��m;�鎅PJ47K���� ����Y
��T�13��R�	Nm�O����+c6���jOBPP��D.�� �0b�/q�8���,u���A���k�6��򤄤:0��+fUb��&���grJI��|"�~�T�&{|d�Ŕ�8?���Bی>��mѶ�_�/�������j���ꇅ�6-;�|#��[�)^  ���$Ҝ4�VA-OJM��=��$���*꾐���\w�!S� ΦRH�xId!#4z�`�Nߙtn@�D�%�A��2?a�j��2�±��_�7$B'̍F-�X)W$�.��eIsGI2T\Ib�n�<�)�-E	�ʧ+-j���ER�$h�i�/E�U�$�֪�.�$)D�V�&R�YABo�8�a�˽J|�i!2��T��P+��|6:ݩ�_���K�����m$|�'��6���!�D�I8���Bʗz�'j�H(A��}删Un�f~k���;�B�8V\Iǔ?B�:d�CŞ�sq�%��hյ��O��!P�S�}�k�L� AV��τ�)*L�RK0����'�DLS�h��*�z���$G�`+�L�c���O� 8P#�9l R�P&�2�J���I)b�>q�B�$2X �5�\q�b�T�b��SŇ3e�Vt��*�%(�
HA%&�p�� C?{
�@�-I\N�Y`��0�A�� .$X������E��O��'@�C�y���v�2���P�<I��ه0r@*r��2}N<Cc�Y�D��|&�<Ag�I�|
�(�bH-1��4}2@6%��5��x!aJրp����2���X�A°([Fj��?��J0�!Y��p�*Y؞�3@*�_nP!��Ģa�P��@Ķ2)h���ǑX��\ڎ��̼[(����-�R㟔���F3+A�Y2�ވ=B$ój)�I�$�V,+���&ւ��l�Q��'V:�W��);�b�J�φ�K�8=�f���1e:��w#��$y�زq!�'X��3��ٱ@�MV�0�"KC�1��5K�]� ��`��i24e�Ǔ��p�� t�R�$$C��Ey2L�X>�F|���k�x�͈8'����Q98�݆��{�ƽrP��`��9
��5�gX$nC���h�I�����(� �;r̃}X7��#[���a�	�yj�bG��OR��e��6&�#�� ���x�����$�f�
�"%� Z�d��Q+qr����Y$:M �uM:}�E��u�*�=��!B��U���<�ׅ���Qa�P�t�<A��E� TH�S�tz�P�W�~R�+Š^DHөG.nz����	>R�d�'���+L����8r�Z���Ә'=�U)�b�< GӚEd��>˓"n��5CڞcWn��DK�$n�(�6\O|<�V/��?��Ϗ?Y�Ő!�Tm���
4O�B����HO,YrH$�"d���p<��;0'�$�B(��������/���Ex�-��~�NEK�@y�񟈽!3�C4K\TcaE�K��RuY�X�&�
+k���YD��Dޑ�����EAU��*��yJ1��Y�$I3�O4��)�fb��T�^���B"��<�ӧT
Y�� 䂗�?���BUJ��J����Y, .x���#%�)&>c�X���;q�T	# EFY�4É�I����@�"����Ul��	����[�S��`� W�Ej�F
f�u�Q8�v	u�J�f�`�b�퉇3�B�A�tޥ�Q��(	����b��fv �wEP�Z%*���XN��|��$־S[���o
��)D�I)jp;qH '�ڄ�C���k�<q�k]�pR��r� �p����S�T�_� �ȭ�r�W�v=��P���d�;-��0㐚(*��t'F��h���C�Q*`צHȔ�=a�ى5�� �@�e����Q"f��3Σ}�;o
��!���d�2���I{��u��	\���ˀD��k���0�Lc�'3�	+�@��cƼj��-��(�bq^��ďP�f���� ]�Yb��d>��O���,�麳��N�8tyc�*��B�>T�C�F/q%���K�r "j �3ړ���UCM�#.�>]ӒH���׀q����`�&i���1%yӰ�4��]�Lq��,]��uD&h5�90E$WT 1�ӞJ� AzԆ@�{��MJ @E:(�#<I�y|`�p��,>���H����)����(�Pl�	]V,��k®~����ǟ2JE��Pe� �6��`'��Ou��Ӥn���1iG$�y�FY�g��I�p�a�p�	���w�d{2Ǌ�L� S��T�p�{���O�LB�Q=C��H;�vT;���a�4�z���10�����gW�A�	XDR�C�<A���Y��Ҹ a�H�JH� �g)�/٘Ĩ�"�+R���� �9�ؠ���''u:Al��x�hD��^!H�x��'=��y����-T5�������]�wi�S��=q�l�'�`,ce�T[�8qr�Κ�x���d�F�>B��Wm�#�;&n��)�n���M>Y�)p�+D�L)f���L�؜��A1/ȴ���H��"<���2[��;�'�"�(�k��
��)�7Ӻ=���zR��aF4>��s7�ˣk�jl� 'D
vd��-�2s[���%}�BI�4+
?�y��� fBs�Z?rL�|�ĩ� �f.D7���!ì٧�����O��)ҍ���ԋ�'��M�fD�C�2��qᎍH�P{&��t�V�{�!­Z��������:<D4�!��D`��R�"3}���KD�Zr�XC N]E��0������u_ �4 ��=h�u�
��(�sM�b�(U����O�]C�J�_�( 	�J�h��	)��iHG(\���� �١����玦4��y�������:$�a���)�Zq�C�_�l�
v��P�@e��ÕG�<�$�W?Pih�"�
>�D�b'G~}bH4I�pћ�j�6��`�@�H�O`h�l	Q�4�� �W��Q��'ܢ����#A%z,�G� 	n�Aq�%I�81���$��4��g�|�d���$�;,�:��%̀���U�̘r�`$��	E]�,��@"O�iQ��\v��{��XZu���"O~|�A qL$�i��FPD��"OZ��/��z������
.j � "OV<3�40J,���Γo*@��"Ohi��A�nʔT��>{L�"O&����.Z�l�*���O��F"OX0�r+_=2�*Q+�[���!�"O2���Џ|
q3�j$Q�X��P"Oа�%��P^\r���0$*2��"O� �4sR�7'd>9h%��'���A"O�+tۜgf�m�f'ϣa�(H*"O]k���n��(Ph�X����"Ozy#�l
s��C�g�=F~�	�"O^d*
$ܪd�L�h@L�rq"O���s*Ǣ��-i��,n!����"O���l�5�T�b�K��|�a"e"O���pD�{6��ڝ^G��rD"OJ��R��p�(�ɰEI�s��D`3"O��x.��u�L���L���E��"O�Y�W�;��-��舲5���b�"OـE�L��N%V6H�G"OBu	�EN"u`�Z��;4+�x�"O�]Y3M�@�2�0C^�@Ǽ��6"O��:@�0���֨R�h�X��"OF���˗ '�Xv�Q�*��)�"OB �*��Ah� ��@�6�<E؃"OyCnT)L.�!�)�;�~���"O,��.6@��=ȱ闟��j�"O@�x�@(z��=���Hy��"O�U���� r�q�tI�0��ȫ "O`kg�Y� �V	��gæ ��'��X�C�s��� ��]�:���'6,���@F,
�(�+\�<�b�'�J�+�lY�C Iؘ\�Tѱ�'���3K�G#VMچbPP���
�'z�����V)q�L�:Ʀ�v�	 �'fv���S�z�Pa����dS��P�'n��S����d���b�.��
�'�"Be��9����E�^$���'��`����;o|�iԱ%��	��':�Q��0#�rE��"�Ѝ�'���q�T:,�9�B�H�'ݮ Y�'�$��GN�"T���Ҏ�P�Z��'<����%�1a=�-�n�E
D���'���)�DL	����D�P��e&4D��QsN���.�@�A�)#A	�G1D�TQf˻B�Tb��ؚ8�����,D�� 7�Z�gR�a�%oQ�]�쒴F)D��:�W�d��Qo��+�b��U�(D�4� ���^#vMI�aȢf!��0�.�!b��94P� ��V!�D��&! , FĎA���QiL�!�Q:ɫ���k0��Sf
�nE!�6P
Ёďȍc�]���C*!򄚥oR u���J�SN��b@#gw!�_���Q �F�5�f���"� N!��Go�(���l��9d쁻t@!�$F,e{��Qj��W^�!�ŋ�'GR!�dZ;�D0��)Z:<!��R!�Dk�34���=S8���$T$!���Ql��㇎8 Ml(z��^f!�$߃n���Zp�f8�1�)�>d!�䉱�j(�#h	�5��ըT�T!��FOl%�ʉ}pd0���0(=!�DS2a~�}�K¶0a�����s�!�Ӧ��*�m�`W�\��I�o�!�[:"�>H���Q�IB���ț)z�!��4Ԇ8{��:���a��Z�,�!���r�n �"O+s�Z�	'��1�!�$��N�4����hQ���C�!�d#5�LD�����*�S���do!�ZJ80��T|6�Z�F�	<�!�
)61NH��)FO q�vB!�� P�a�"��x�
�(B�$sw"O�h�HڑgpX��	Q��j�8�"Oµ
#(�Q|�A��ҙ5���!"O�lJ��&1.��ȧ:�f�ʕ"O0Laj�/' ��d�U���xC2"O��qb�*/L�	�$�_�RySp"O���C!F�H���4"țg�Й�"O0Q�(��	�L�2�KԬ��AI�"O� r���$��sUT"܀(��"O�`*1�FlZ���o�!y^�+�"O �6�G� /�4�ԭA-M?l8e"O� 3��9\t	�G��HfP���I�"��d*۰K�4A$%�C� -��a�%)Kx� �  w8�C䉹	��8�����șb�����듁hO�>M���	�q���s!� w��a`�9D�\�q��,y2����h^33X5a�C#D�ZP������8(b�1"�#D��	��B������-w�FIK� &D���%�@�3���Q	F�uvC>D���%LL,t���-�6	@����1D�v�Xh��I�Y�
Թ�H�8j�B�	䟀"��&���H�4w��Dc�,D��	E�zĠ�!�0I�r`[V�+D�4�`N�:NA�����)��٤�?D��8F$[	aU�g���>f@����>D��3A8%�h쁠%�x�`؉�%?D�4x
��X@����"eB�RS*;D��R�З0�~Q�P�\P��(a�
9D����όig8�ZÁV=p&h=��!D��!'k��bO���mӂ�4R�?�L���I\����\R�*!�V�B~!�C�	�r���ao�>^P<�{qI�@ېB�	�v�V�B�@ŋx%�4���hۄB�	Z���&+߳2�
��K�!Z��B�ɷi�p��&�:a(�"�@�o�B䉐��p�B�+��1j�n�0����?�����	�\�A�Y":���3c�<D�4�%M�jN��r5n�wU XHq�:D�)!�'|$�(��� �1���)7D��ZPjٴ��r��G���y�
_���IC�1sk���'�y���k5�0�C荅�q	�`�2�yr	L�<����_��`'  �y�g�'b-<ݻ�nՆJע�{vA@�ў"~ΓT�ne9��šr��sX�14܇�D���M7,j�`K3�,y����_v�K���"�"�BU<^�Ȅ�B� skȢy}��B��9(b���q������|XB�� *� r1���ȓL�HY�(�mndD��L�5��ȓ`��2�$4�"�B휯���a��ɒO�'04�R�d�rQ��A(��,�*Y�,K�-�Z~�U��g��s�4R5t}�c�������������e�7쓬9^"�v"Ombe��6�"A��[�^����O��$�5W� �c�AΛl�f�:�:F.!��6���r�£y��%��d�#3!��WV�%K�X��S_�a}R�>Q1���q�� 4)�Ma �FF�<�A��,�j27-�85��\ ���K�<�4�C�W��0�Q�_�P͉��Q�<�(i�*�R�j�6���H�v���ק� �b�Q W\~}��O:~֞DI�"O�E�3Nڣ"� d��E3v�:X0�"O��"S���J�a�ȡ@8N�R��
g�<y��L�5ˎ��� 6n@�6��_�<	���w�� F!� �*���[�<Y��� Mфp6�Or�͙ %F}�<��k��-q]�5����)�^������S�����Y��H�N�̄���x�՚<*(ŨʞB+��ȓG�]���$8����1�Tg{l��J�F�+��-L[����ED5X��V���J��x�`��6� 9��kG\��W�H��y�1�
^4l��ȓ&��A+�JĔm�f-���,u�Ҕ��\�x��4S[r�F�<�0s%"ON�`�L�
f���f�\<\A "O��Cv�v�����΅���
D"Oرꂍ��RaB�2d�F�XS�"O���bY�;|�Q:1l��1�"O��uoΧ-��!�"� b�"�"O@�86�2{2�02צMG�Tف"O��Z2��K���D��I
<+R"O�ٷ���R���PG���e��aK�"O�5!��4	!�
0��9Gܞ�I�"O�s fZ�>e4i�2�äS����"Od-���֢m�H��EU����"O��S��^R�e)%C�4b�pA��"O�<��D5�M��,� ɂ"O��c�����t2Q���r�@�"O�7��6D����Ɓ�(��Yڄ"Oȝ��eڴi� 1qAE%`tY;�"O0d,�q/jј!�:�,�v"O�`�_�U@<`��U���a""OƘ�a�	�Ac�쐋� QPu"O`�M~F� {c�Жz�^P�4"O�����-+�pb �����%"OR�����V`�i���09(A5_����ɰ)�tmg��>�`�d�W�C䉙m�"�9�݊&��ɇ�O5�B�"�jh�T��'��p*�P�kvB�$.8����,f�t;U#B��C��$!�*�&��nô�C1�$GԢC�/r�!�-|8}3�5OJ|C�	�~aV���	��+�*v��'1���-p��H�cY�5�5`��y��E#"� s�\0_����J��y�a�%)Xl{��9��Ļ��	�yr)�H$$�b�^�\M�x�,�y"�Z�P�H4�EW��ثA
̕�y+Y&23�\C��W��z(;����y�����X���A	/�4�%S��y��*�Թ�����#��!FCR��y⒑U��X����3�>И����yb���e�¨�a�9 ����_�yHVy�V�;�	�Pn���y͘�JȨ #�މb�83��C�y�I�T�R�i#��V�U�6�[��y"��42
0���BI�k&��y��1e�耂bQ�$ B�H6n��y��Fo�<��"kɳ��yB���!�L��i���V��3�ة�yB�ۛo������� �U��y2`
�f �)�BS�^'��S�'��`�&i�*� �+g��V-����� LC �� )�a��5z�E	"O(�
��Rn�,u���c�Q"O*��r͘]~Z�V�y}Z�0�"O��d˃�p b�!X
hUΥ�&"O����*�$�(%B杀(�B�"O���,D6yR�����7���%"OVpʦ#[�2��ń�����`�"O���I[uΤ��cL;h���X�"O�q�ThY�{����4'زsV,"a"O���,2o"n��H�dU�C"O�����T�p�����
.)� C"O8TǤ©a��;������a"O���F-I�?r�(k�K����Zq"O1J��7P8@�{D
��hu�"OX����+j�ՙ IZ����zT"O��KA�sz� �h0]�)�"Of-II�(}f�ꇧWa,����"O�5���2e��]Je֏�¸J�"O�Uc�?��Q`��#v��,b�"O�h�&[�5�)X#$	,R�@�P�"O�%���W.��HUm�.9��i@"O�+` ��H������ak�֔C"OVy1GF�b�&��&a+$ސ�cV"O2x�G�7u�������<�I�f"Oԑ���^�.���Q�䚫(��P�f"O�lڇK�Pl�@��ɒiP!�e"O4�0��Õ�e��
_5
K!��F�<�����2�.
�Q3}�!�$Q�0����[:S�&	+�I�
X�!�����9&M��]C�)P�!�d�i����䇩���a�!�T"I
2M
!�I	42�����!�$֓t���αe����Bx!�D�s�V zqR4W�h��e�;�!�6��M��Z[�ڤh��.�!��Y(U���3��1"���Tc�,m!���`�Ph�7N�"Ŵ[Ub:Y�!�S�\y2%�L1�b�ܬt�!�J�aQ��b�VUj�߆/�vC�?o���1F��B=��J�LaNC�	(5�4sq(ф:<Ra����4��B�ɺw�!��]8o*����f�PC�ɾ�hQ9�阈&J�E(ѵ�s�3D�\��IR���^�IQH�e4D�� ҍcX��bV&s����e0D�h[V�5i�Z�D��l���!D���Ǐ�7Q��y��Z84����>D��P��0$4�⋌��lmAQ*>D��B�M�Fr���.x:��ѵ�6D�`�v*F�h
r�i��ʇz���4D�l�����$�9Я��d!+�B-D�`2�ƚV�2�J�f�]��ZA� D�o�C<6��=�e�X�aӴu��;D����/H$D��e�J�:��9D�0Rrg�3C���b�(�X����U,5D����I�=`>�0�IحA�4(�ׯ8D�Y(�-�l��t���Y�I�(8D��P��
o�! �W�i_�4�g7D��!��k_��;wDJ`�(�1H3D�� q�W6e4^��&J��İq�$D��6����P��;��L0�%$D���f̬aU�uXDB�&�Z�%D�*��kH�I��d�#!�m;��>D�d�B��g�� �AÍlv��s�9D�� ���ǋ�2��I� S"(@�"O�I@�ݘ=����0�A*5��+�"O|��3�ƵP�X��@�=%(�-S�"O`80��J+g������8~���"Ox��U*M8����nǖ-c2�(0"O���oO��#\#Y*9C5"O 8s`�)wwFu��$B�!Lb�� "O�1!2홗(0����җ#@���"O�y	��\�h�����!$x�3"O,�i�e��y�<x���"�U��"O�Xx V�'���c@E�̨4"O:@E�"s[޴� �9/��i�"O��C�7�`aR�K�q�,!"ON	��m��Xc�}P��˹2:4zw"ON���?/��@�$��)�Y)�"O���ݖuI�-����J7�衃"O�RJS�+����tb�D/�a�2"O�pQ�e��1�L�3��M$ �"O�	�QВ`=1 �E�^�f"O<�*P�R&s��9��F��Ą� "O6!��B%W4ڽ���G�#�2d�"O���FJ��j��"c$����CC"O��ѧ��kn"��%h�u�R"O�@6���W�B�H3%]�V�D=S"O�(���Z~��(���j����U"O��T�%*�A�	G�䠉�"O�\#�(��>��0aY?S�L�S�"O��q��A�rs2H��Q�O{T`�@"O�t�uJ\�2" �ɰ�
:v��"OH|p��#<�3Fl�'< �ų�"O������.�`���LǛw�8��0"O����ʀ7�a���=����"O�lx���%��qu�ub�B��yҡA�du�c"�b2)���6�y"D�#)�� ��m�"H#���yBm�;[�e��ّgu(xKTNL��y2h�Z	���g΀v���Nݼ�y��,\����"gĝmkR�+!ށ�yb嘄���ס�R�!t���y����$w��W*�Sj�u4i�y��:wF\<�R�ϩEhʐ�L�yb-ҭ�>�sl�!R<횰�O��y�MM�������Ys�7�y�E�S����CA�#Fd:�(��y��\"z�<��5^Ŝ�
�B��y��F�XՐhk`��OT&(J��	:�yr�E�kB��T��X�J����͗�yb菲ŀ����;hy��(ϻ�y�e)'���J��0�֌1*W�yR�_�Y�T�8�N`��9�c��9�yI!׀��h(W��c�қ�yb�ݨĶH��Oq���O�?�yR�#p��$� �B�(<S�IW�y2Hͪ��H0�	c�F}h$�ݮ�y��Uf�ؘ�D���f�J�;�ybd]1-�I� �^,4�7̇�y"�S?�Z̃���Xnx"M��y,���t�uoĴn��,��˗�y��_�m�@+�1jҔ�:P�ڎ�y���,|��"���(\$�������yB��-o:��XF� ~��y�!B �y"�M�q�4y��fW���a��&�y�DއdG��ud\ i!(���y�c0!f@���>Y�
Q '���y
� �eHѥ�&2� �u��0�e��"O�Q;�@}�h����S'�
��V"O|i�d�pR�1D��0�4��"O� �
 ���1%�Μq�HH�"O~�4-߇ �P����_�lz��"O� �!b�n� ��o�SG@(��"O(9���
���H)�(įZ�"OV�{��X��5�g��H���H1"O,z��DB��pE���"O6�HC̎2?�F�!NU�*4�$�"O�9�Є��'�����jB�L��
V"O����{� �*Uѣ;��|q�"O^$�� ߹> �t9ub��C|��aD"OȬZS/��/��U'�mw���$"O��(�"H�}�>�0�9Nܩu"OH9��×(Y�Ɉd�L?��a�"O���-ȲC�2�Y��%k|4��"O� ۡoE�ATn���F��`s��� "O�����K��Kd�#,X~��""Or�#���H�:X�VJ
�D�x�t"O�T�4Ǘ�R� $	�Xm^�Js"OL8���Ie<Z�?J��\��"O�4��� 4�D|R��uc@	��"O���,��97��Pp�ށ���"Ol��O���Y�h�%>�^�U"O~���e٘��!Q�aK�Q+��2�"OxQ��b�/�����.��]��"Oȩ��&]�	(}@5�U����"Od���������##�٭iӶ��"Ohͺ"'�Kиp��g�y*݇�{
li��$yÂX#��װ���� H9�/� ~��ό�"Eb]��zB���G�*q"ժ�@[�1��I�ȓX�+�ES.a>(r��H�xL
@�ȓ(>�eFMX$`�B�@@�1�Z���|;\��w���,�4����is��ȓSJ���~<��7	��T���(�zEB��J36�ATe�S4����q�r�����:d q¥Y�/��X��aĴH�'�+s�b|W�ƻk��Ն�2��R�$?���jcg��r�X����&��T�xTt*R�Pj���������#J��� o~���-�L��t�M�Z��]a���&����d�D���MsZ�s��)}|4�ȓe�!9�b�+�8����ҧJ_�$�ȓ.D��P&���Y��攢�ȓ�L�:�o: �<�;GE[�]�H��ȓ{+:D[$>�Ȓ���d�q��5�4 �R�O9����Z!.Q�ȓ|~n�+�G�?B�q��L�-,0��U��i1D1M�V�z%���,�R�ȓs/�!Bա/+]����?݄�'?���+ȃE��#1)�3V.D�ʓ]�VEbSM\�,T2l�%��*�jB�Iq�z�d�\�[m (!��i�C�%	��A�"ڴ����Q�
<�B䉝U�����
cn��b�=c�ZC�	&c����"��U��4c,'J:C�I'�1"%�g�|�Gi@(yxB�	�u����`��m�ٰ�Ӻ|�C��6_�ʤ@w�ѹw5PJ�ܲ&��B�Ɏy���B .N	>R�p��X:ki�C�84����E߲W��c��|F�B�)� `�7I�;Հ�)����2�����"O��Ce�;�ȷO��q�Hi�a"O�X�� :RJ��f	�u}D���"OҍX�DؒO�z$��$Y�����"O��9�8&G����4a��K�"O~�s�i� on���� p���b"Od48�G�R��-�*��=]�iAU"OP-�+����`�$M�"D�2"O�	:��Ѵ�4���F�Y&L��"O�2¤Зmm%��8|���4"O���g�I�H�59C�5��*�"Ox�� DƧ���a���; A �P�"O��1U�!C�l`F�aF(�q"O��3���T� ұ�A�G-���"OMZ���k��C��B'�h��"O���a,�~��x`w��!.���"O�kK,hh �!AZ�P�n��"O�i��(з<YbQ����*�v1�"O�Kp�I�p*�m�(�*��A"O~Q��(�3sb��@l�dY��B�"O�0�c�D*`E���Q%�	J�Y�"O$]�cM�M���oӸDS6t"s"O��pJ��r�niJb��Y0�-!���JRi����(-�6���1sn!�ۦ0�p(&�*m�(9k3�áE!�;��9�6� �w�\|93�Ԋ�!�$i��D��"D���[�.�!�7K��	��Ȍ*,0������!��L�)��+b���q��74�!��V5�Ĥs!�5x�D�0G�]�!�d��4����@�XceU(m~!�D[�m��c�����`��$�!��΅.{f��Ǝ�F�|�"��	F�!�$]��~$���Yܠ���3�!��_S#��!���:l�P�@�i}!��&V��a�7��.@��U#���1m!�D=-fa(ra�E�(�i�
�8�!�4츸�*�Ǝ��!	�!G�!�=YOd)b���*{�r��!T�6�!�$�:m@f�G�z�D�����*�!��/�����P's𖐩ң�%W!�D6,}*�t^4~�H�ʴh�5]!��V�d� �[B��$����H@4$!�DH�@���.F/;� ��f¥'+!�� 8-X����� C�)��գ^x!�˃!pj�SF�ϽB� @��ǫ�!򄉕.抑0��ŭ뀥�g$�%�!�dߢ1�jd#U#E�Y�d�j"�E�'�!�D7g��4) M����Pҩ�4F�!�D�c�0%�A�%U���9R�w�!�dӕ~f
��ː0ӎ����C|!�$ݬeA䁄(t��#M��Jg!�d��Z��)�DF�H6)�&�ىyc!��jV�cDΑH�bod!���	��E�㧏�60x�-��<�!�ě.|���dl�T�"��*֦$v!� � U\�n[�{����+�/L�!��~K��4��D����e�!�D^�;u���Gk��!36	2u���!�d�7H�����ת|�6�WտT7!�d��FN���iYq�����g�1#!�Q�V�6y�+�)����I�=!!�d[�f�|\Y�kĄ'G�����
	!�G;,[Z�j�%&O�i��F;'+!�� R\�AD8;ɾ9�$?m8@�p "O����V�����y!N�b"O@X@���v��e�%�ܟ/ ��C"O�4Pы[H�!���|���RG"O��@���O�r���ɺ� l��"O@P��g��3 �URB��ഌP�"O��V�	�0����L��2��`"O������>zξm[�F��	�t��"O��0� �TFڹ�Q(7m��,��"O����`Ѧ|jv=��畭 =֭��"OФ eÜ�HX�(�emOeh�"O��n_ɞ-�c+ԧ[L
ԑ"O�*�##T�����i_)x���Z"OmS'��-�(���*ȁP|����"O�x�6���cz�eh��=x�}s�"O���L�$[6��ֆX�x~x3�"Ox)���B|T��0�<M��ɰ�"O�T�5��}b�(�b*	��x�?D�̩3�H*]Pd-ҢF�b�}��.+D�<�2LC#A��13ᑌ9��I&D�<�$�ȯؔ�b��ھg������8D�(���Q��dn��j���G,D�`����6�hic���<�șĉ+D�p��7<�0}0��֊|�<��")D��ӳm�%��X��Ǒ�Y�Ԃ�'+D�T����#����c&�6S��18��*D����$LT|�����B����'D�xH���5KT����3VT��{i$D��C.�f\��A ��;Rۋu&$D� �׏N3(�L��E懆-��k&�=D��@Ԃ	;�$B�ƿ>�X�E�&D�쁒m�^ܠ�j�E�s� I��$#D�p�#���w
X@��+C�����"D�C�N��/��ubԤ�	=�s�"D���V��v.P���+��zï=D�����3���d�� R��(u� D� �U�W]�\��H~� �%*=D��*1瘭<�̴;'�D�h��0fC;D��CLJ�7H��1BBA�?�Ai�=D��#�F*���S' !t���"4#.D�t %�,C< "�a�FI0�Q�&+D���7O� +y��J"��G�4�)c�'D���f��h�Ȁ5�BBZ$��'D������J%j@���.w�꽋�&D��!��v�h�$"_�_X�@`&(D��#�N�W�d97`\7
��":D�����4[ӊqP&�[zj��a	4D������F}�$���L)O4A�.2D���l� v�4 ����
c{��)1D�h��ϱm��f
�Ot�ҩ.D�����^'�Y ���7h
T�w�!D�X�c,�:g�p�
�H[�m"l�N%D��!�AN�"���ȔkX0����4�(D�tKƩ�8`*�P;���\�a�w`(D���A���C�j)�
ΐ�V���(D��@6�}d0�g�
�|�L��&D�$��\K�a5H�e���)2�$D��� AϓU���U��3Oif��G�$D���	��6�X�,tdQ2E�"D������q7t4p�Ή�Etmʅd&D�T�nΒR���[f�8O���Ǯ?D�|
�� �x�e�W�C+5����9D��J@k/P~B��b�aXj�j�6D�H���!^�(�S�L��	�>T(3 D�� �0�HP%7��E��O˷l��`�"O�	s�#@6L2��i���s`����"O��2͖w'
H����26Jl�i6"O���U��/-�`I1p�XI��%"O�`��̆:dI��0�N5ֽ+"O�����ڍQ\ӳ �Ј��"O�8�k�5
b��Ӑ�U/P8�.�yb���+2J@։E
}fpH�'��X�2��p����n-A�j��'�a`�M�]�fQ��Ϝ�O]F�"�'P�x�#�P�2L�q��G�� �'�j\`qg�{^T���I <rn.���'l|�)%-$�<�j���|��'�xyiB C%"$���E���9
�'�pp���E��TA%�_	��0�	�'|��$+Șek,H�'�XVl�a�'���2'�A�l���U$!�����'����)�6;�0�"%�X�V(�'�*�jS(Y2����)͐J/�\�'������(r`p��$�=��m�'��%�v-��^�jH���S7���'�tC��WaLy�� ��0K�'
  s���	�l�Z5ƝlxAb�'R��,d~JLB� o�d��'J`�Ku��=F�f(IÌD����'*���'ͿM����Cg��U�`�'��)	�Q��
��
�Z���'��<R2H�=\�Ԍ�o>�K�'��d%@",�a3FP����	�'�b����@�(�ؑ����p`�'\.U�p
O�>m��A1���
L@�'E8��ՔGXɰ�H%�\!��'G��t�����`p�����'��ݲ�":�]�jR�&��'∽:��A.���K�! [gp�C�'D�m(u�řh�d���nH!ڦ�K�'K�0�%�r��=�C�BwҌ}�'L�|z3�X�`UP��aeć<�zlj�'�ڕ���X��Pi�O�.��D	�'|<]��a��lʢ��?)
�ܺ�'�BM�D[� ���R���@��'񊁻�d�=���L0�c�'���m����2���ez�'�>x
�/E�9J(e���2p�4Y�'B>d!���ʐ0�b�ƃX���	�'7����NJ�9�&��nah	�'&)!�
@�BM�a�֗Ca�)��'{ऐ�`$�x���E0����
�'#����� N:�=�5��Q�{	�'����@ߛ�,���4$�p	�'��("�D�wd( �T(Z�W���Y	�'�\f
�0d�P��cG���}��'�u����2pKL��6�s3\ ��'b�2�(<��u�` H�jy����'L���R�М3���1@�)9�֔��'��\j�"à#nb�0�'j8X�'7J9C��e������^%&F�3	�''<t �ʷDj��������'�� �rNT(y�̀ȃ����'�0,��,q��	Q�`O W��o�<q�(�|)bA�#+]}H6�hqN�I�<Qw�א����#J��1�츸d(�G�<����� ����1�2xĄ��׎	x�<�B�N�]����aJ2;��B"w�<� >�����_!Lܪ+��ْB"O<tK3J�9s��rRZ>f\��"O�-�ǣ-)��dM�~|��"O�Ȋp	�Z*��0S�N+F����q"Ot�Hѯ[;/��S�� �麸Cb"O���)�C;\��$F)���1"O���#�?�]��,V�H��!�"Oޕ��_�\B1a'f9A�!�"Od�s�a[$#ܤ�#6'ұM�D���"O6��$JI��8D��|��"O6��Vb8�x�D��U� "O؀�����kf���tѴ��	�`"O2	k��8#�-�G�N�Ό:$"OEk'f6:�$���ݼ�LXk�"OB�c�����j�Ǜ�1�R(B5"O���K> �a�L�$cl�8�"O@�s���6p�YQW��4On�9�"Ov��g	QBؼ"ʐ�~A|]�"O�����1x���f��q�(�X�'�<A��!F@^d�1ɬ&jd�!�'�HD��ץ5,la[�h��r�0�' Z��S�.C*�P`�i�)���'{4��R�0i��oߐ
捊�'��93�/b��f�X�|Ӱ|��'gLy㲫O�N� Ȗ*�@�4m��'D��1�fPkH0���E	=�L��'��;��ف*ZZ�(hG]��0�'CZ0�N%�$l�E�!����'�DP��I�8=���u�T�x	�'4t-�w���,�g-S>�rś�'5��"�h����@�� +�� ��'�`H�d K��A��+Y=x�bL��'�tu���+O9 
��Ps��M��'�X-�V+��t��4��!pV���'��{�ØB�B3���i����'oHXSE�0m���B@���]�Da(	�'NZ�9��:5�ƉPU\��	�'�l:��O*6]�x��玆D�8�c
�'���J��E%`�`��`A��AS�T�	�'��tX�ʨv��! a�+���	�'�l�ĊV������ ��K
�'���0f �:}�
��t#L�
+�
�' �\XfU	WH���#t����' u��9I�� 
��G����'������F��^��C!�9<�S�'w�x��ӟ9S:��铩/J
��' ��#%Ξ(����%,��c�lP�'�n���j��kQ`�X��؂"C�=
�'W�ZF�MU��і霄P��d�'C8A�!�ؿ#`���%Ii⩛�'�I�6�{{�$A��ǉr����'�2�*�M��6q�er��ƴZD"���'d��$ċ�i��S�R�"���'�$�+�&��&�r ;gϖF�pUJ�'�N��6�̙���6� ;����'&~�I
�ilB �bL�a��q�'ƶ�Ɇ��&�c��>#n����'~ěcO�'*�xXRN��U(�'�����ߐ����a� �R��'Ҩ�6ₗL�tQ1�_8y����'�dU��kH6�j�1�M�?�V%��'�p(��k�c>ة�p��.)&��'��@X&�úq�r�R�ז6Jh�9�'
��!ŧ�Z�|R2e� 3,�ٲ��� T�8�o^�\j�}JU�R�era0g"O���CN��9�0:S#�,C�;�"OTAPw�P�oW ��UJ /6�92"O0T�����6��A*�k�~0\���"Od�Q̛B�z�G��*$�(�1"O�i�c�~��@E�Y�P��"Oཛ�D�#>Q����e�
Y��6"O��t�h���0F%m�*s"O0Ћ��D�v�*��s�b�i�"OYӰÒa�������J|��K�"O��%D�D����D��2b̥;�"O<JtG-&�F�7A�>R�p�"O���P�
<�r4� ``"O>%�V�K����E�e.5a"O���6�e���Ʒ*
���"Oj��VQn��JE����i��"Ot�sCZ�HR�ȋw�*�4��"O�l��i��9�Ăp��C���"OT�BkF�(�kQ�պs"O�Y  mW�P�H�!UF�$R-Hu"O�-`t�K{�(=��ـ+@��7"O������������6-�k'"O�ٙ��|| ���a̓�T<�0"O��j��2A,�k��Й�0�"c"O�x��j��G�4K�*�QM���c"O�I�� W�f��@*J�
���q"O*�3q�DA�I��r��"O�h��/�z�<������i%��� "O��x2��O�����D|�W"O�e &�W�:ՠ����X�@�"OR(YA%�5�\I��G��Y@"O4DQ"z��`5��*g�rc"O�x��!�fH 8ċw4��!"Oju��,Ы>�L�R
#ǐ0a@"OL�����F�]��C(�~��"OT��6�ĭYyz4���0�е3�"O��#�a��x���ʄM��= %"OΕ�#,��|Q걑0�͸O#4t#�"Oq��L+��}*&$�T���Za"OT�Qő"%z�ъ�)��Jj �u"O𴪀�֟p�h��#B�#e�E��"O� �0&���$�8�KI�hF��w"Oĕ�DOB�mӒ뇜Y,��"O��t��%NC2�)bJ�<���"O��s�_�<�̍XQ�U&���S"O�����`�Ie�|��"O�P���Ӂ�m�e�Z�le�LҤ"O��@��gn�u�3$��wE�M�q"Op���Hn�������T#����"O,�a�H�:�N�*��C�Y("O�Q�-[�0%�����-5"В"O�Ȳ������UH�V���1"O&�9'�t�f�0�Z3^ D�F"O^U ���.<�>���	��\�A��"O$)˦�Ǟ������ܴ/�t��c"O^�"��a\�X�%ɰw���S"O�|8�O�e�yQ��Kp*��W"O.%�����#�vA
1��"U�X5�'"O�p#����*t��O�]�r1ۧ"O�A!	Y�وx��N.|�`[U"O~���
@o�8�HH�	x�"O���/��M|���BK�q쭫�"O����"|e`� egX{ܙ°"O��󳎃Cz��`%�]3 ypU "O� ���2�	l��X�& 7����"O:�(B	>��W�T�t��9`7"O<��c�Z�Nd�%�߁@�<�"O�Q���G�i�a"2�͋8wt��"O`��JЧd�
- ��y��@�"OV�un��v�x�g�ХZ�tcs"O�iab��1Ҋ�"R��  XJ��"O"-�W��i@�r�ǌ&_9v@h"O|��F�q��!��_16,�t�G"O�i�(ϻt2�ě�&	,��c "O4<"V J�|m�L�&e�'��qB"Oh`Z"��)(��a�O�\ P�[�"O9*���'yGfe�qe)_g|p�5"O�J1(�0mX�����/"���"O�����ԓ�N�r"�)�B�"O����o�L{�P�$+�1kΔI"Oଉ�"]���"�dJ��ĸ��"O"�2�k��|�¢��|�4�"O�}!��Ԇ\́�0"ՔPČ�"O.M���@�*��1Š�Ci����"O��>
�nx�B+.&�{#"O:�0I��x�2ӕ͗�aw(�aW"O���%�6e?4IH���Ve�!�"O���R��,G�B4I�*�HR �g"Oޔ�C��ϰ5Q 	��[0v��@"O���T��!t"�mA�&V* �K2"O�` �KR�G�^�b1��/g���8b"OL #%&��!��
TM\�5J��P"O�	��W����RSû4�$,:"O�%h��ȉ�JEP��lh���"O<=)�MJ{5q&��fi�T��"OJ��C%�<��i��0S�"O�AS�_/ ��(�Y�R���)�"O,I��� t��P�
��Di��"O6Mȳ��~��x��l�#
���"O�G��q�dtr�+ߠ}^��G"O��# C_}'v���k�?����"O�Be�ŀ��,/��Q�"O��Z��*J����H$E:6"O(˔�ë7f�M���,Aʉ�V"Ol��G�ʎ������zH|�B"O]u�Q��:Ф�)=��E@Q"OEb�b�B!J�gR8�9DK!�d@�k��(�f�Š2:�
�-� S!�DT�u�����F&Bx��͑�5"!�D͡wG��yЃ̑uR!	Њ�%I!�$�=>��4
 ��R�TT�ũ��<^!���g��
��ӽ&�*���O�:P!�D�X�
�2��� 
^]PU-�[G!�$9X��8�aF;tZ���6D!��N�ޝ��ȋ^vTb�**5!���F���4˞
�89���t!�$Ϙq�.<��H�6�&��c� c�!�$Aj@�8�EbI�(VN���e�!�9ARl�shEKS���rAƯQ�!�DH����4�8O���ͫ20!�S(*L�����:H2���41!�� D���c�F,t�nL�D��!��╰�&��R�@���-YJ!�D��r�a��A �5�!����cc!�$_�H��v.�b�0x�ȆT�!���:U���c ]�Q�g�j�!��J"U��T��"�l���&K�-�!�d�^�a�%ʳL)��'�9B1!�� t��cA6@�¼���ƙe� �7"OP���ِgM�L�SAT�`hB	H�"O��ԇ�K8b���mϢzb�a�G"O�� D�əLx¢�:e���1�"O��a�D�v����V}�W"ON,���1[�"4 ���5}��"O��!2�_�$�r	P����/B�0�"O����i�U�5��*�ʙ�"Ol�6�E�ER��*�t�4Mb�"O"x��#<pP�P�OU�j�q"O���2-�%U�F�bF(�f�*��"Ob��M��
��Y�t��9q��V"O�0��&sDd: �H�6d �	A"O,��l�&�zز�
+4F��R�"Oڼ��g�1*�Hds�ѕ&9����"OB�"��9�@Y���<8n��U"O���"�}�ak���"Ox|�Q��uH}��J�:~�`�"Ox��S��T�D)
�~�(I#"O~�A!�4*�T�K���f���j�"O��bM�&��(���7�`0Q"O�ũ��#s�r)K5-:mB����"O� ���H�#� d�q		�U2v("Oލ���)h0[��Y�p���K�"O֜UJ�(���ąO
��刷"OL��kF	n�����fŀ4��˗"O`<��A��̭+Q�A�A�9��"O4u�Sg�+I���7U���12�"O�HC˄(oM�H@��!�ڤe"O�0 w��C���r��O= \�"O���c�ŧu:����I�&`*�"O�$yU�ޗV��Q�ш(C��jp"Oj}&�h�C㞹/��`� �2p5!���i�b �!�����"�!!�$�I��%CU$֟�|d��a\9W!���^���i1}�����F�!�D�j�^u���6LC-���?!�!�A�5��d��*݆�j��Z�!����H��#.����/
�*�!�X��Z�{cj�1)U�h���
V�!�$�PE����U�;4(Ĺ!�!��I��5�ؖ&�<PPf�);~!��]�'!��� Z�}�t�Ң�|�!�$0lh��v.+�́���ۀ}T!�d�C^���w�[6"y�����
�!�$�h�ظ���~1lbG�M�v!�O�L����!�8��^�!�$�/\�8��D،q���Z�!�5�d�2��M�z�v�OU�Q�!�$ߣi�h�J׬�C�rIq"��v!�䅬n�*�4�A(5���l
X�!�P�Ҍ�5 �Dh� ��!�d�
RY�hs����D'	.��)h�'���ӎ�?�Hts���4ty��']bQ�iS"M ��Y�x��Th�'@�� o�!$:��V�]�X��DR�'̦�w�Y�]��'٭W����'j`I��9��ݒ �AA/
<h�'�vqÓ�ɟ,^�afO13����'����B�J�4|��A�-{���'��d`���i��$�pK�p���'�>�uª ��	���
�c�N�p�'�V��&g7R�^�W�	a�:��
�'zy��ޮ<Q�Pr&�٥Y��8
��� .Q�"��6lNД��A�4uh`*Ob(F �"jzd�e�E�
i��'/�4�%i�l�<�f��dEH�'U�,R �\!B�B��-F���'��UZc�O�Y&<���32TU�
�'^�@��L�*�"gɶ�M"Oj�1@�ȯr��XG�'IB`a�"O<Bǋ�@L2Iy$�%F�l!�"O�ͣ�_&�d�4B�,�i��"O�Y"��A�,=�������pl��"O�8�ҥ$���R��(�m@"O68 ��*�2��U�E+'=��hU"Od�+�
@6t�jW)��;>9��"O���,.f�$V=:���G!�y���~W6�#�o�1��d(p�(�yI�^h�	�5G؉��Dp&A�y�	�6i��y�`C�rPh���yRl�7
�D(���?�:��1E�y���1� �4#"���0��y����m���P"ؼ1Z�/�%�ybŘ�H���g, ��槞�y���?1��=��.A8QL�=����y�ȏ	 ����g�K�X �6���y��B�,����MZD��.@bP�ȓ;�:�I��Ù*�$�aFq�݇ȓ*'�`��_�J��*
7D�&u�ȓ,J�����)C�)�Ŏ�5s["=��<�p�A�MK�(��TZ��_�{AՆ�y�(Q���9M�:T����p�,������@'"�,[]��@p�Ū`)*��ȓSm�a��	�F��� �I(2� h�ȓ,=Z �sMUT��3��_
Ob��X��SiܾL�xL҃��.� ��ȓwd�(��qԦ5r����{����4��H� DA�V(�a�H���T|�ȓH�@�`�
W[�MA�S7[������lq�Qnǁ	P\�X0�5Ya����^����#CP���N�]_�m�ȓ]�Q�J�f´S��Ư'��م�prY��~u�d���;����ȓ*S��$�
{�
��K� E�Ju��(�MQ���<���h��u�@	���� TK9ۺ+TK� �T��fG�� K޷b���E���m�ȓB���X0ʡb�����M͠c6^M��Mn]�h�-�m��fڶ┱��$���B�n�&>
p�$���	�J�ȓvk�鱷K�	�k��Ķe��ȓ@k�ϲz�u��L/�*��ȓb<�M�I�c�(,A�LP�V� �ȓ3cJz���^UVŰ��7&��|�ȓ^��]�#�\��
�b�Μ��Ω�ȓ,%H�+t�(}u�tz��	���-�ȓ�r�����"z�Eb%���w��ȓɮ�2(��@���)$A
Nzz	������/�Wr*�)q�#p�d���nD�ч%9m��Ń$ɏ3A��%�ȓc�ttj���e��D��C	-kv�=��6�^D�0���p��@�*�e�>q�����Aj�K���D�5\W��ȓ��<����Y���{�bZ�P�l$��r�䄚e�U10�	��(�N݄�Y�t���� 1i�̨$$�-�V�ȓw��a� �j�q���-�L���S�? �;���:ctT �c_�3���2"OhE���Ű,��9�֢7 ,3�"O��d�ɲk�*�q��8v�H�`�"O���!i� ��lcuhS��uS�"O�5��!/x�a�%w��Hz�"O@p��.͈=�����˕n���`�"OT���h8Qp�i�6�yf"O�hP��9&8�H!���o�H�"Oȑ`��?�^�x�,�:\�D���"Oz|``�O�b-�͚W�0%}��"Oɹ��ǹ%d��ɟm8l�b"O�9�U���8XD��,w[�0i�'�T�	6h�Ex�*��		z-��'#���L�*y�HzG*�t�
�'��љ�n�x�.L2��	�R��	�'��1s���&� S��W�`��!�	�'���J4�ϲ|�Y�o�\x��z	�' Z��h�6T,dՂkH�θ�	�'�,��X�q��h��h��x�t��	�'��Eb���&b	d܂ք!w1�	�'0	R�˃XYf@�7m��tWp�K	�'��(�U �
 ����Z5B]
�'?��;u���I�ꏅP��R	�'L$�k�g,Fs6IB��@�L��'����L�ٚ(��	'$r>�[�'c�$ɴ�)b&L@W����`��'~<T����*B
�rƒt,��'��Ԓ��G�H������k^���'?"�Kw��J���Oɑ^����'����&ؗSq`;Gn��B"
9�y�A�=L�a	��D7�H=C`�Z��yr�^�`�0|�R�L4-�^)	@�V��yra	��a���c*��!���y"b�B���R�U(z���6+��y�٘ȼ�r��D��5�dM;�y�j^����T�!��h�se��y�D�#�6�*�
��vMP)�3LT�y�,K#�P�!M�2v�l�RT��y­eȈ�u���w��$�.���y���(
��%� ���D�bd�À�%�y���g7b��c U�<��0��͔��y�	(XZV����2���℁�yR$�/zz�h����v��	5o��y���z�T$V�s2d�D�B��y�HI�S�XI
�C�-�R(����y���=(�H����_'~ϊ)Á���yb�W<P}�I���yp��T	�yr�65�~�1U"N�T��a���yBDĹnu���b��`�6���K��y�-9EXv�V��Uو!jX��yrÞ7m/Fl�2�6HU|� ���y"/�����G-X�8+d9���.�yBʄn�P���I�'��q3#����y���#p�yy@�wڲ�%,��y⯄�I��'M��.�������y�l =^`Dh֏��B�� &@ħ�y�&��i�LL봩�&
��q9D�I0�yb��`6�i�J�J������0�y��!�|a��؍Qe"�� �$�y����R�l����%E��(�H��y2��텞)`�|�  ��x�'*
@��Ve.��a�,Π)X�')��6l�)Gᎄ0��ܥ�H���'�$4Z�kG�s��;�,Ȝ�c��� ܙ�W���=�RT�����q���1�"O�Ms�M�-�5�e�!g��Ae"O�[��
$S�%�%R��B@"O�0���g�	�ף(+���@�"Oh䑥nԾ%9 ���  _cb�1`"O�!A�]"���3"ܕV���+"O"��j��Q�D�S�U:@�nX�"OT�Z�I�<atf����
͠��"Ol���,_�S}�xK2�B�m�x���"O8�m�vU�,rюF-2u�3b"O��'��+q�؛An�)MU�\Ӗ"O�q0SH�-��0��!I�d��"Oa �bQ����1�fPT\��s�"OJ�c#%�"��4C�R6���"O�	�'��N5Z���	� �̊�"O,@y��C$c&���{E�X �N�<��C���j�@�(��KG�<A	��*��+D��V��aXQ=!��
'o�0u��3�YZ��9&!�D��7�\��d�X�3����-�!��`dX�� _�xv*�8�//W�!����mb�c�(`w��F.�7z
!�d��Qł��N� Gnp���G�!�D3O�zu{-G<U �	B0�Wr�!򄛝c���� ���($e�)h!�DH^�0�%�Hn0l���
-6!�3#�TE�xD�L��Z�L!��D/OA�� �ƈ�<l5#��oB!�V�3���X�N 9
}�gg '!�D�'Y6��3���>�B=(�+A*;!�d�����Sj�&dV��k�'O�!�A3`�^iJf��8�Qa�I�;h!���1��-y��D�p~BL����qe!�D͵a� �9C�?j�>���HG�}4!��1Fܩ�h�$x�@Hۡ_%!�D@$����P
1�*�9d��=l!�dF:Y����kȽ.�F<�ύ�N�!��A��Pi��H]�l	b����0�!�$ئ�%��b����
�
@��!�$�Y��%�F�0~��9��Ω3�!��<-�,,�SM?Dw`M�@�%u!��0Xip�B�#9L����go!�Ā:�z�T�@/w��ѐ��V!�$ޯd���e�v[�Ԛ����GN!��)/D^XsEI6<I�ɢ��ҥo�!������)ބ?O�uҎݱ�!�Ę�}�U)tBX-O?��s���!�O:w���6�{�H}i�#<!�D]8Y}���qa7n\R|�6���!�D�*��a�&�/��q���UO!�$�3�bA�rj��w;�	P,X!q9!��PIY:6@	"p ���H_%r!�dP-SUf���¼7�"P���wc!��R�b|���苽`�ڌ�p�N;c!��<L�����<o�|K�F�10�!�d0tl����F�W��L��T�o�!�/Z.�8�ь:� 0bmرY8!�$K����J�"��`��+�Y!�䎵Ҍ`Ξ@��P[�Q,x�!�$T��Ls,ǫM������O��!�D�2:ئY�dC@��@�Zp�\�!�D�=_���d�<S� �2$a�u�!�䈵)�*�j��Ԕe�P9[�o�f�!��)o�a�҈�#�<u�EN�9m�!�� ^��a��6�\L�@H�%p��AV"Op�{OՆ����l�t��0�"O4ͻ��@
5<HŌ�E����"O��@�8\�� ��圤Lr	�4"Op8�AҜ\n��"4��b��Q"O�a��C�Y�|�(���}�&��"O�xA�%Q
SHl�4D��/��d;"O�x"��ޕ:��l飈�<���	�"O��Y!R�Al�J� ��� `t"O�� �K8P=,�+�j˹�<"O���U%Y=Z���;-��qC�"O$8X�H�`ONQA�˵Y@�� "O��Q0A����TJ3���"Om�Ф�%)�:aC���*���Xt���G{��i��-/6i�D��5V��Eyg�&�!��$���/��U���{�f��C�!��9�y��@D�@|ȑ 7�]�3!��^�vT�	��!�l�4���O�%�!�$ �=�Ș�SJ�:H��I2䎝3�!�dބ���J�	O0Ԫ�p(V!�DJ�
�(9��͡,� � �悯IL�=E��'TP��D��!' �T�ɴ2_�U�	�'�J�	`�UYn�1�U��|�^m�H���C�'�����ho����fݐv��)�㓌�r�lڷ��U',�y�c�>�d,��'$��x�"�3�h���+�6Z=9�'�*�	�gɚY�F���������'<��v��
Mpn({A���}�6�2�'���ˡ�Q�5RA��M��<3�O��Ě�	&�m��'�'���6/F]D!�d�=�h�AɄQ�J���MB!�dʪ	�����C"V��� Z#��!}��)�)�(��h�̍�{�V���`D�!��%̀�z�&lUܬ���r}!�$�.1 ��fm؟,���H�]_!�ܽ~d�����;4|��ܘJE�9�O,�p	5*`�P�&A���"OxТ�ɟ�"�^��w#�� -ZY"O`��A�]�d�I7�J�=��"�"O��[�BV� @��34���"Ox\��f0�^y�#'� *z;E"O��u&Vni�	e�бU�9�`�'p����r� �����B�!�U�Y��B��d���I�M4��oQ�*�&��$a���'����ǅ"_$9���-N9�)�ؘ'��`!�%L9>�N���m��a��|�ȓ���`U)�m;� B��X7�>p��K\�SPk�R�6��@%D�'|=�=�������J6m�&%Wl��x���#��OV�D��Bp�򄚤*�e�t�b@����O2��2_�M�7G<Oob�Z�)�=7�b(����V��!6�j�C%#�3
��t�eȝ�+��B�ɶkx�$�@�a����2D��>�O
�Ig?ia��O�S�Dd�c�"8#Ƒ6����C3�0=ъ����l�P�B*hn�a����#�S�Oi�Hy��ĦG*�ْ�ݾf縘����(�'2H��S� do�9��5W�ņȓ8�A"�&X6p�#΃2._4�ȓnr
|�s'ľ�P�ǖ�:�����\�z���L2�m($��4TJe��l<�R�Ȁ	� �D�9h��` aL^�<�@�!��-z���&H��kEv�<9v̊�[+.p�C��4��`j�g[t�<a��<��i�V�U����oXF�<� �E9��G4>;���'�[)Ϊ�#W�� lO��SJ�.0~�������S�\<�3"O����λ}�]���_�!�h�S!���XE{��"��M�Z�f�U��X���k��I�OUFU�v���m^�Q̞'l�,9�'�&�y��,S�����X�e-雉�$2��)┈@�؈}"$x�F�^@�$�ȓT�j���-f����E��؆�k
X�6��+n���3(ٺ$$����-x�"" 'y\���diQ�,*�l�u��~�K8���M�<���y�!1P�� �KG�<ٱ`
'��i��H�;���+���j�<�#%�:���K�62��Q��h(<��4����ц�$a� ��0f�;q����r^`�a��4��"��N8j�d݅����J��7�~�:�+�/	I�ą�b�(Cf�
:��P�� W�e��3��q��.׸G�D+7�\�8�V\�ȓh����^�pΔk�M�P�Nd�'X�}«¹J���e(Ɠj�F����X�ў�j➘��h�EF�Eb�he�0e*&D��c�΅U�Evߙu�����6D�i���:t}�aʉ4[�}�I4D�ܑ�,��SrL��"�
UT�HT�1D�B��>0 �u�\([��!@0D��З�� Y`��QF �E��AѰ�)D��[A��]Ÿ����U��D
d�����䟠:�\�3�^��H]z�$ #3!�� �TZ|�+�*/��k��P7/�OX���p�JY�����qDJ��!��[���M����>�L,$��#�n�O�,!��T�>L�D��,�c��J&DW�,YJl�4D�(m��),*e�����<@ʡ�%D�dK)U�n��9�M�(I��(��"D��4��"S��B4�ӵ-��M�sm"ʓ��<��Q��!��Ѭk�	s2,�@�<y�:� z�K)~~Q�$��@�<I�fV�G��)�عIru��~�'n"8��CO�UĎx�h�=O^���'[��A�J�?����	=D�<`���9$�(��"Ǭ0� x:g�>.78�-���D{���c� �5�ۮ7������28�p	2D���veI;)��;�g,G�]#�M.O�=1�b�On(�򗈘�kFVX+ VO�<�0���F#�)��B:�Z�z���P���.Mg��pY���� L�F���/�؄�iR�x���.�z��sB�*�%��guWGݢ},>� F�]��"E�ȓ;�.�)0́(˒!��C(�Ұ&�����+Lep�Xu���F�l��7�P;7xC�ɪ�d�%�ֵN�|(���9v"B�I�M.`X�ٍ<X��T�":-VB�I���ɳB
]�Y����׋`t6B䉞oݬ�э�.a��L���z�,B�I�,�P��i\�# � t�Ц~�N�D{��9O�@B�\�je#'��
R�9(�"Ot�I�j
�P��D��Վu�Z����x��f���J���	&��]�!�4M�ք���!$�D�1e�~2�� ��	3j��2 �(}&U���'"Q?� P%��l$�8�`	�,o5����n$򓼨�� �@O�-L2	WC���@Z�"O�9�*\kf~��d�&������P�˄3M0qO�O��$L(cM�,)v�I?*��s�F1;�!�$�UG~}�F��u��iflB<s!�� ������:c�����e^�.�� ��OB�%�KH��{qB�Z�U�@w�|���R?6
�DNH�m��Ͱ��M�<1!��):(�af݁tmʬ��IH�vz��.�HO>}¤B��l0�B/I�oh�m�����>��s���%�Q!+��tj��Z�8��%�<��' qO�"<�Q��2%�!o�%Q^�1I�O(<9ܴh�̰�eG��1w�<��u2lAYtLū	��%��� 9kQ0��ȓ*����#j^�,��	� �˸L�bԇȓ4�&Q*���6fw�"��gS�IFxB�)�ɂ�;�� b�́�(�@�k�c�<�vC�q�v�3Sʄ($S��%�_�<1�#@&,��BBH#mdR	�q�F�<�C$�>W��9 Ǡ9L�!��E�<��O�{��12�Hذq��\��@[C�<���=M��H31�G!G� b'Uh�<17�KX�X0� V+P�jG��z�<ɥ�U�v�R�k4KO:y��XR��v�<��e��VD`�4,A3����{�<A��S�V$ʃ�Z�M0e���L�<i��h�0+ĭ3Ò���L��<A��Zjʣ��'~b�gLE�<A��ܽ5��P��&�����D�<�"�Ī({�	��`#��}ꡉ[H�<a��ɐW��c��5\��@�N�C�<��o]������I/ ��Dh�<!w�P>�<�O¥"
q{R$�o�<IF3>�yHK�"D�b��d l�<�n�=IRQ�%��`d��"e�<14�	�J��ǯ^Q�R5R��b�<��[8c��eI�X���CcG[�<��(\�|����Ȃ1b����SO�<y�꒢KN4E��-jt�i��M�<��ϯzoRQ8�!� lM� '�T~�<�#�)���`�	�'S�����^�<�6,\n���&���(��icE�W�<I��ٜ3f<���%�-!� K��U�<�&���[��Q� uR�d �M�<UKZ�b���c�fՊ{� ȓ�Yp�<Q��r��h��C!�T�QG�<QV&�$JU��ƊN�:d"A/��<�&��R���I�2@���h�r�<!���'0���@l5�GfYs�<�a��G�H �5C��e5�XnGg�<Y�bO*t��G=. (�0A�I�<)��G usv	��&"gĒ��P�K�<���,�ΰr�a	�c�Xq	f%WE�<2�Ɓ�4\ c�=��9�p�P]�<��B�tF�P��j9����_�<�4�J�Q�ژ8�n�u�]h�n�V�<I�n�8\�4��g M$6�@��U�_�<y�̕�S*ԃ��̦@:��k��X�<IeBʑzcD(y %͝K�j�0.�T�<�V˒/��ͱӄ�='��5�d�N�<�g�8BBc
;"�`=�%PH�<����%�؉S� �'M�����E�<��lN�+��ـ�8t���C�[B�<��Fq�,�RI�$:)��MB�<'�>"�jxG΅��Jq�W�|�<	���S�������5����Y`�<U��C�LY��<8��I�CB�w�<���Ԧf�����
4l����FW�<��K�J����:L!^9�`\d�<� ����L�8��i��-�|�<,Yt"O���Q�;ml�8�O�Z���ç"O`���
�w����̖�F�,L
"O� ���"Wz��� �� .�,���O����T�и�h��8�+���b�{�+��,��)b"O�<�D\�gq��k�k]�l�F A�Y��	F΍.tʴ���'�س�jUz���픋-���Y�Yj�9���y225�a��+#Ru�f��*b����BӃ�PxB�X1�RIY�NP�S%@@x��Ĕ�(OLD!h؛2�\Qq�.�ӘO��h�#�� $����D���#�b�Y�'AJl��)� � t�������2�6{��(�CB�ͩ��_��(��	�x��ur�!^c��vd�[��B㉶c��\���w�Z�rsj��F!k�*\�U@���)2��� ����O�d��'�����O�F0���HX�L1e�T�tX�,V�X�V��<�X��\R��} %T�c_j����e��D�蕽d�|i E�ǟ}���db0}R�@�=�j!	�	���G�-	��裟���?	������<�p��QCЈ�y��0�ZI��?���Q�4�9#�'I�:��X ��\ ��$���YH,�	Q�6y �[�Y��Z��`�I�X�V����'5@��T*G9d����EL��(\���%��	�d�X�p�Wb�(W�Q� *;��dމ!�P)v�(�Mc$�S}
Yу�1g:t}�"J�� ��8��	��ʽsF JF�Ϥ(5T�'�W�r�D=DF/�*l�ң��|�z�d��B`��a	�'.8@��7§f��`�ø��j 2t��'.-BU ۼi(ĪsL܀
PHw�ӡS
��QV>����	�V��r7-�4|\�+퇚K������K�v� Q@��9C�x�>�O�q��	72���+�暈u�!��a�@Ch�Gd�� '.�{�䓟��p�.�0y��i��Z13�������[�@1FH�Q����o�n�����aax"m��\	P�2�݋c�ۀ�ž*�zܑ���)T�h���=
�L���|D�R�Ldś0�E>)�tԁg�ԩT�(͈��ھ6��P 2��d��I*j�p$�䢂��`RR�)O?�H����f���'��y���J]',��`R�/�>x�V��G�z��E���$�u��	A9P���j�x$���DՂ��I24�F�q���)�	��c�w[J3��Ŝa����O4�������<9���_?/�|)q���.MĔ��A*�	��鳲�b5�z�ON���<��Р�"֘1Cƈ��k��N���iLo"x�a�dL�L�'���5)��1C��Z�����>I@������;�H��%� )X��[A��=LN�5����, �0���A��u�,�b��t7��{u
S{���)�T�i�?R�8�g��:u�4�"�u0��kU�ҏ{zM�L�kG�!%,��-�I���7O,P�+e�L�pΊ�v���V	
�o����'�j=�|���܎8��<ඈ=,}����
�9����i��h���W?����NX`�*G�E̒Q�n�8Z���@B)�Y��]p��Ճ�dҁ16D�P�(ٳ ���0kZ<��	�)V�I6F�3��p�1�a�x�r`n�X!�ȶ�8����IպS�Gٙ7Q*��|"ڢ !���Jծ6-z�J�Ǫ9* �K�`�\�"��ӣN�D�1LZ� �����Fp��HA.h(�672�����.`!���=R���)�C�;]Ph�A��@�����$۔���B�ya���j؀r�T*��I�\� 0�g�a�R@nH�I+�d���T�� �$`� �h�h$퓛. n�Ү��#l(b�'l��%lK�~.�8��=.A�Wザ.b���rn1�f	W3~1<H����9�������n�~-�'c·/b��S^�	vh9�f)��|7,l3��˜m��9W��
q$YB�A~b�^,)�l�$�@�l��R?Y-o�&9J�f ���1��A5T�45�D�� ������1OTs�)RO�&tQ���+/��� ����V�$��$Z�Y'���`Iƣfl���R�ЖV-�����۸�f���:+aY	"[�]/��� )F�go���F�T+���b��Xq��Ꙑfj��C��Z�l���)�(��a��'4���tnT<t�x�-.��� ����X�kaͷQ����r�ގ�x�A��=t�ts%��,.��V���x�J_�-����R��+F������I����Ic�PR�DǝZQLh
�P֟pH5̆�!�萁s`�2mH6l�6BO�W�xp��9<�&�×o"�֝�����f�����Ż>	���������ݜ+��b�dD)���I;;F �`�W�=S@#�?�A��-E\�z�N�{��0�P�a"�(��|��Ӯ~��pʍ�/��bqo}�>��ɃU�2`cih���A_�Y9� e��# 3�U���h���c� S�(b��Y�kl���a_Y;�`�@-bپ4��	�5�T��C	:�6�2��[ĺiY��Q=d <9�6Cԅh��(�ć$��KvBӂl<\I�V��c}DdPBK>b/&�v�T��d��Y��=E!)�8(��΃'Nvz�0E�$O�����B8�(�ёB�1�yBB�'�B�:����<ӓˏ% �H�IĮug��@!�1>���Xw;�x:�˝srT$��h�L�m$<Yu��$��`�C?}���>sL�ూ�?N�M�Of�7-�&`�Q��5!��J�F��>��ch��I,�A3il�� ���B�wu�Z	ӓQ���z%��'�V8S���;��)3E*X.V1>�kr:O�d�U���:UC;&��$E�n���]c�r�eV+=��x��K�6Z�����'/r�qÌ�X�f�E�8W��%�E/ǟ4�2���	�1N^F�{�'�v�i�쓛Z�l��%Tx≷E���g�ϓ_>��0����Cy�AĜ�|���>�Ń܌1n�� 4!��F΍Y�	��^0����ZK��HÆ�����5��+i褑�D��˦���i�|I��
ںhg"�]�M�{�? ��)�G�;m̆ͨ��Z
!�`�Ď��A�OO;<��es�'un=0�hC�xp���!��D��pX$�A�DQ��>��B�'C8����g�����)E��|@�S�?SKZ���"̑y�bm�,B�PxJǤ��9&�8��ַ��K��vJ^���l���-F1
$B�r�ɝ�� ��
o�̑�`�d�©+�*�Ap����
#F�hvL�;0���ӷ]���:��۫<]��S�+@;��- d��/B����se��������C!��
�h[��~���o�nZ.A���d��G��"�$A�"!��g�/K�P�:4�@)`L"<95,	�vOT�����Z���Jĉѧ�U�e��Gf۫o�Q"t)�b�z��3�Pu��8O���ΰC�s��U7Z�'A�Ir����<�1��+ߘ'�%����Y��ʤP-m�q�BE�`͔+Y)�x���F�;z��	]&�H����i�:��'N�}�$��$��R�F�@�Bs�<�'L��2E�]`|�1���W"M��jǢ�:l�yh��1M�p1z��'.촓���Mʖ+P�#xj�#��0�( ;1�T�oRT�z����F���N^�%,2�:,��I�u����,nWX�2����;rP�r�U�F	xȰb�R�G;���'ă)kN;D�Ǐ/L0�㌒;D4��0C~����s�l�A�=B�)�lԊE��a�ׇ�ss��C�O �t�V�pd�8��*�F���'������	�\�@��,g2.������+��x!h����j�'i� �`��B%����.b94��"�΢+���"#�� P��ɀ�&A!M�a��㞌���P� 9�ǁ#]L�����XIv�T%;E$�W*������dQ���[�a���V�TZ2LK*L}�h�5ϐ�|*�a	$$�J4��A�f�V#P#J�Bg:(`Ģl�Avű�~�i�A�Dę������Q�J �3��ۺhb�-���^KT����K'��۶�ܳ*���T�ԬjB�h�����!��@�v��ʅ�R��蠑㑋+�L�vK��a�T����>���A&l��3f
�����#�
(�6�׀u��-$l */b���7���bL�E���R�Z?۱O���`o��VC��R��kڴ]uZ��#.X.	�hp3!
��o�6��է�<�����F���9�&*/�y���/�dlQ�_l�>��;R,##��9}
nI#����,�^$�OԊ���t^��`��
�h�����'&�8 �4��+l°1s�Z���tjڴ$�$Esխ�7 `BDo�6�����ҥj���V��j2&k3��c��4cҫW�k��b^3��, �%ئ*Μ��C�m EV?1s�+i��j6��)3�@VP#2��Y�%�[�"4s�X�^-s�^�O]�5�e�2eS�y���0��c�D8ĸ�衢bj�tU��d<P�f��s�_(/�R�	'�O��;�V�8�����JUrT�����Q�l��kߩ-�0��)0�V]����M3�kӠ]<��
��7Pg���i���V��O�XB���I�z�꣉s��K���'@�T���W,=��	hg�ٸS��D�N&M�r���	_�s��<��5�w��fȸ�a���h���7��x�"���BK�/�=%����O�h��
�!{��=�'�V
0>����}��ۓi�,WEp�p�1:㢅��MP�=���:�V�44�0�n��
��I.ROb��V4=�����;3�0Qc��D(�va s��L�D�5�X��7,�69��ڠ�U96�,q�D�{�bM C��%hB�!�'#R�kN0��˒b�6i¦�Y�}42!�FaŁ<��i�'nI��x���I�C'��k`\:.�<:���/-�|�B�b��cؕÂJA���ɲ��V/E)��;&`�:+� jAݭ(�`�t�I�DR�j����<���=+�J�� �)�����}b*�#)8, �2�W�`���2e�'g��Y��"6�,5�J�Q��������:�,S38���AՎH�o��!L�#7�$9�s�P�4�q��q0qz��QOV*���%¾I�`��O�\%Ky���R��N'L���<ɄJ��{n����0^XZ7'\xB�G��� � E 'wr���'!�#vt�Q�H�[D�G�~T1n�(\��a��'��D���3{UH��2!�)e��	4o�8	�w�Ԝ-N��1f����t�h��{[V�2ᔓ!O��!˞DI�XBF�ѯ��8BI�W��	4�����Ȃa�mS�41��$I'��\�t�U2aRM8R����,��J�j�)���#�Ąѣ��.¨d����S AI�M̛:W����,˶IC�81�H� W��y3��ۜ8j�+�k�;$�ЪW��J�JٶQ;�٩�&�p?1F�d�ұ��,΀+Gg^�q���]�9�̱[!�� W��BS,�����'���`I�2�Q�B�\=:����el΁^�$i#��)�X<{J>a��(�^0k�
�>a�%�|A�X�Q�J��F�K G�Z����YZ�����@�l��r�J	h��59O�@���D�V��&�\������o���Q.�6���c�=F�(ٔ��{R���O�] �) ~���U�Z�U�|����\"��~���e��&;��E��&ہw��E�%/�bh�	^(m�9x�g�:yS@}�B��9��#=�4Áb��U�|�z$H���[v$4���XP�!���%Xm���
n�%��X�}�p8�T_|.$�����W8p $~���Б�T-R�ܸB��a@Q�x 6�Z�|�����m?��*$VR�㪏;|>R�PR�)Z1 �2�E�3������E�'"���#S� \\�2ú���@qC		g�lɨĪ
=;�S�Gќ��Ȅ��x��9���	����VE�GG �T��yI��:8z&њ�f�FD�QbE��1�z��㇒,:m����|B�V;<s2��s&�
BB��	{v�� "��GS��k�DC� Q��Y�!jٺ'I8y�Q�ys��0ҟ�5a�Ȁf����s�H-5=&t��Y��&�2ro�7w��z�Â6HD���a�C)%��;,�(O��R��\b�D})V��m�j��@��*Qo�mp�h��gO*h��
����
�Ɯ�b�@u!�$n�j���Ț�Wc�M8(�.w�D�� �����*1���Jw�ʤ�(O�@�p��%����q*Ԟ2���z'�Q^��)��E��*NP�̻"�y��+oP�₴�`NL�&�]�����̒��@`�Ĉc��c�ЕK�I3Ө��˞���G,?�V�e7�	�'-$q�9�Rc:kd��t��p��.0Js	=�6hKGŗ>��rS�!6*����˃�vV�d�	.2O
0Z�B��9�8|�'7d�ۥ��=�6d@	A�c��Ā��׻X�@ ����06�N���'�(��?7l�ȕN�'*�4���޾K\�zBJY+6s�Y����#;���T�"$���B���8�� ��Z�O*Eه@S�����OQ�L���jV?c�$���/T� %�į\��d�i�|B�`ҿs�d���/�'Jj$H�"bTs2�P3�@A.]�)�) B�lZ=h ��!HH�J��ɹ�H�ɐ��$�8U����N�v��knYp6�
�7���MӰl���v@W�a_�p@C(Q�]�:�&KQ�ij]x�'7���E�s�f1z�	�vSj9+��Z4�2M�f��6��	9e�h��)K5V��$EŹ,���S��� xYRoM(�VyA�cR�S��1�ׅ ��t�iT�C0<u��e��rA /�.��F(�'>�$�r�����3l��a��0$ͺ4�r$]�D���	��@�!fk�̋�)Aܕ
L|�Y��S�(�8o��Js���������k��U���M,4���JZ��*����5Y{��bC.hݡ�VFƷ����Xhb���=~�Z����.�B	�,M(r7j��'�*�*D�"��:�ƨJ��}�v@����	p���_�[�\
0�#g�̹���.�Ⴕ�@��J�L��y�a_/�P��#`�ȥ�����w6�B�LV'V	����A�7h�>p�"�S��rE:5 J�)|u�޴_�i֧W���ҡ6l�*X��'.C�l�t�ם"]�D��I�Z8��QD��y��.��ȅ!�M�t�T퓺r���9s.�P�;�F�Tkl7�1b��9A��)y����'*�/p�ey�F]3(����+z���ΧYY؁��P�Z5xuR���:^ @�E�*4] 	��kⵣ�BAG�ӧo�םvyQG��o	��3�O� xp�X��ܝj�`�e��[ Ǉ&������W���S�O��I/'��p%�QΑ�E�2j�Y�a�\X���/U�m-=(:��`���s��O�)�,
 9 U�r�.�1SEV$�<����UN!qǪ�5X~�"+�*ϓBK֩��&̔�u�+��/�2����b�<�Bģ6��)B�j�0���aaƍs,N,r�+�<ͧ4̹PQ�L�~��c5;xL���D�!_!���.J(J�^��%��I��A骐����l!q���:�~�}���Y!M�XY$��K,r�JB?���"Y�Pq���Q0N[p�C�$m�4�E��
�#�6�۴_P�,z�JԆkz��{iB[$�E��T�>D�s�?�s�<@�S�MC C�'e3ک;�g߰z.��C�E=�U����'r���> S2x�|��º>���S�Y�T�Ġ�box�q��K"
��$�u�M
0�9֦7LOՒ��W�
a��@e��6u��GD�,m[j����Q߸pkG`��@���.OFu��] �O{��f`�u�� ��\U�6aÓ�漫V'X:������H*?��t��,���P�'ɁHw�z���/)����+�*�+�0|�7	۹&�P��B��T�a�n	d���!H�>d��"ܐK�.m#��
TP��ր�68�v$Y��>+w}�V��0oqO�h���Y��Ɂf�>>��!�&��h����*�n����c͜2j��#�Ry�}&����N 0.h	)!!��t�d�Gi)$�`����mjp�աX�|��9��K�&�x��F�_����ɫv:Q�W9ܠM(�B��0�@����8ߦA0�@4����J�P��bo�z��TXF�ӗu/!��v�8���l5~��2��-qOxs&Ȕ��0|��-�+%��5i���&Ѥi
�PG�<)!F��p���@�1�n�%��<1�%k�xP����3��-K�aFw�<�$�)Q'<�Ȥ&	7�X���Y�<���*r.�p��� yO���`�V�<��T��V9� eЀ`x��)�	�I�<����v���f̂J�ᒐm�<��BG
5�][*^#TD�od�<鷁L���[�O�C@L��c�<)�A�&t ��B�H����Y�<ѷ�R�V	:�.̡[�\Ձ��QQ�<�����0)wC�6�⑙f��`�<��
G&z��'�J7f`�"c�^�<id��Z~�k��	�/8�3q�UZ�<�G��Y�d��6$��3h�iю�O�<�v��c.��ƀۮmE��YĪ�\�<�� 2�d#���&K�*�s���^�<!�Ƅ;� Qbǅ��(|�C��Kc�<������`��G�l��Sюp�<9���'Ȏ�#��?��=1��D�<9UD[�8������%[8���@�<���%P~dx���v��!B�HD�<1�'�@��іO��c���G�<����7�<сdσ��M�4�O}�<����"C~��P�C� d�&|���]�<9�G�&-�-�ս�����K\�<9�� :��]�q�S����{G�W]�<��[`d���ft� '�8*�t���A��R�;'�Q?-����ȓ&�2�r���]�� 3���#�����C�|�x��٘0�*�P�,�ȓE�z|��OP��(�7�Ư��Ԅ�l�v=3�Z�W�����̈�R��Ԅȓ�������֍�OZƉ�ȓ2юY妒8^<���K/D|����S�? ��S��<��ULF�z�1�"O
Qj�%�#�b�� �/�IѴ"O.��3H�~�"�l�7*��a�D"O��2U,K�t-\���59��K"OY��ܟq��@ �D�	s��9rA"O�)з���K��0q��8�.�C�"O0�7��1�n�B�퓌ܨ�J�"O���j Y4`���B�9���5�O̲!�����h�&`��!	=�����D#�\��r"O��!B�^f1xC�4$��ҳY��	�͉Aі�&�'� u��e�n���S�O�D��4��GNV%L\�P�O�N��H��v/fձ�-���Px�䟨>���j"�OO���!�(O�Z�D)=���Bbg�ϘOy�PU�V)$(���e 65PJ]X�'�Z�k��&IKh����?,l�z���$�M�4�ת
y�#��֮�(��ɕw(\�Rf�����c7��&ZnC�ɫKQ8���6��D����4�S/_I�\���$&R$S�����O���nϾ.E� �JT#$NObX�p9B ��$5����hA��- ��L�h�*I��GVn�RF�F�`��p���'���H�`��QV�y�X6��M�t��L�k(�wj2����˶m��'>��-�28�lDP�T$�b5��� D�0�c�)��ls#�J�R��Qo�?�n���h�1���-U��V�>]��JŎ�~��O)�-BR�H�/j����V<�~�N��CEhy���
A,4��V�+Bm���3ɳJC �h��OkNF�rD��:X�ÄDu�����D�<!LӒL3�9�s�z��i��d�#�N���cS�~��la�'�%0����T�suD��e����Q�'��� ��G�2E$��*1�e@2�X�?ytm�Aqҹ:#+&�����IZ<fД�X�۝��u�Gʖ/���6:0ջ��+Ta�gL��*H���>,��L�O�,�I�&�"]��)�%ל$X&0:�n�Gj�0�U��B\p�Y��#¸��76��02��*���i��I�<�d�	���
%���¯��QǄ��skǜ��W̐����74����J�+:p� ��wN,-�-^|����
�^�H��RB��S���lv:-�C�P�N �&�Y-%���g8�Q  �n���:�i}"��+ё^�h��&�-��G��D���ɣo���*�Bb� +ό�E2G�?n^j�P����SvgХ",q{4E 2/�$������@�b6��B;^(��z���+�c/ic4#eݱ����B��FC�`�@�磐u~R��!�l���n�#n؆)� ��$��Dx�lW�y����Fm1+��.����0)Q
�����˕�u�vy�2��:
��`��>�����*.(�$�B�6�j�سL[�4J1�R���O� H+��;êi)�C���'=ȾIa��((��Ӝ�p��b�ēUb���oZ�(�(�Ya�F�+KVŁ��O���'S�"f4�B	�L8Y��P�2C�&£(|�T�Ta�'o������'o* �b��H Q�f��,	K���m�VyI���%�F|c�/�2������ ً���~����%�4Y�m�a�I�A͈̺3I�y$r�;���,"�lȮ>�^���b�9�e����"A��O�M�)ܨ%�z�����bNJpJT5��I#NƔ���H�)i)>����p�N-�L�	O���~������?S��U�@	�
ix��'oN
|�Z�#��4�T��A&�򌐇��P��M'������aJ2������h{�aZ�~ƽ�d=~�zݘ�I��4�����\���+��Lq�����܌9���*'H6r�pDB��?c���e�t��EcG
F&P�����'��)D�P#9�j-A�E�������2B�!�SV�7Z��B7`��@�h["@|�2RF��D&Ti+v�M�f��Z$L��fy�T'��CN(���p<������H�:.w�	[䆴���iQ�,��4�J\���R����!�h�*��\��텷L�"UC�O���e�bm�';�NX�Ď���Q�Rg� ����D�/N�
��WK1?Q�g�!\�=����	\�ī������~�Il<e{��S�CA�x3!K�*xuظq���=F� yԄʴ����'gMdz��{d���FL�O�C���(7�ZP�Я�/k�NtI�DQ?! J�Zs��O���E��D)4�\X��/��m�Fda�D? p��(* ���f��f���!�@�+�(�R��0m�azR@��E�(xp$��(�P�����Y��s�n��E�Ҕ��o~H�%�VL�����4'��b�[ަɮ���y�0H��x@�8��Џ��9�����@�ax§IK�j��m��P=�r�' ��#1B�!]}-��n2}��I{T�?,~	�էУY�2	���4�uw�	Z�f�at��9M��=��O"͓�
�P^0D8��ٻ:�t�Y4��h� �ձr~��Z(O&��l*�J�>�b�1�GS>}����K.���9�˙�y�x��6]Ͳ�1+K���i��G��p<Q�+DSҙ6�)"v	��1S���T�])�?)Rб:�,3u�O(BY2�)#q����1Q�젊� ҈#_Fu���%�H��P�ia2�%�l\{eH�g�>��v���K��H��(��W���S&	�=mc< ��(
)�rd��\>b�6��f֟�\y��[)��ᲅ�#B'�QKm,ф㉚S��Wf��B: ��d3O*���M�~� �D���m@aR�� |���!'�H�l|�����&�n�5{Jܡ3dү��+�����a�@��+��^�2��O�����֩(�X}'EP��)����B+Ԅv_A1�h��d�~|� h�9j$@����>���o���)w�	Caz�;��`;'
��brl�ȑf��`E����kʶr���Iʟ���9��xJ���XS!�� ~k� �[�+LP&u����-H|6O|��v��*@�����MT�����<kЄ�DO��J��01O�ɫF�*B����͔�ē5CX���5\~����K�4t\�݄��k<��bR��r2� q�/o�N��^2:J�4x�̥"Ʋ���Ě.��1��dO6��6�X�M#��+�i�-C��X�j����`b�s���H�a4�I�T�F8��j09�vE���O̡�fBPȔ�!�珜iV
�:��P��m�Ox�ęv5Ox1�>���!X$��r��ܴ7�q�@oC�`Ezݔ`�S��5K�IhrB�I���0Gn<|�~݅h6��*M}�e����߱i5�
�<�r��5e�~��rέ�TX�!�B��=���UWX�����N@�F�K嘼V��|�,�R���i���@N	�b�n������~R��qK�oZ��$0�$�S )e
dQ6�M@'"����ɣKs�x�%��4i��p/�"� ��d�Mo���R�D\3Y򀀀L<�Ȅ���O/L����d��'qx1X,s`��ߝX��O��  ���IBDJ"�I���i��
#�@�I�'|.A!iC.�tJ�hO>�<X�-R�4�nZ�B��7��O�M�RB��Y�`��џ}1��#�l9 !�i�F�1��';<{��׀vtіʄ�?р� r���5T+�0�����		uˁ�4��*�o@�!�x�ЀO�c�����-��J��O����-O����)B�q04+W�&���p�X�CJ�r���G�h� �Ȋ���xT+�?a�K��'��l�2�<��U�(p.!�mU�c( �����_f��$٘o�|<����I�kL�8Q�\H�/�\��*���atڤ�å��R�B�����O8 fG�=]�` eo*_���	�csʌ��;v�4�ʐ7,OVkBFăs�~��=1bA8U��H��F��V��c?�q ���[H�@(���\����O��bv�Ĩ�Dl��P!g+���r������d�w��ͣ៟Dp���F>��S�����*W�5H�1X��9?7��W������H�BÁz�&��E��w��r3OW�7�4+�(�|�qp��7�~=83R�T��嫡�ڇ��O��S���#��,���$�Z<��j?T�:�B�3�V\�A���n�B��ӟ ��E$�T��4{��i��B�u+�t*Ҁ��8���
]�Y-�TG~�擑�V�ȕ�V�&�bٴ(�nSi�)�, dƛ<(�˒�34���*�耂@d�I����>�y҉(�
��=$�ϻA�6H��A۸~+4���DQ�Y���OT`R#	#�r�_��h��=r��K�i�yx�Ckn X	�녣ﾸ�޴~��S���*"x�hԂݖU�8�à@G:9���'=p�5�d�կߵ4�ȘP��T6ȽK�'���wD�F��.��:�t��M�!92�04@�8E^5�B Q�+�L�#�N�$;�x�{���.Ւl��0�L@��y�'�}I�,>\TK�H�J���B6� &�2��S��pI���	��g�TH�L;N`#��H���Zv��%�<��c��/A����f��0
�XE�����+"��
D�XJ�'������T��Nm�0c�	*#b� c�r�C� ����
`��#.�(��W<4����I�HH�Z�g�`�k������" d��y�)	ix��U�����'ե���D�u"
q#c�)N�$9��~"�|sTQ��i	�ku�
��N< ���)�ŋ%P���G�,G����隙G�T�(^�}s�Z�>���9���!Y�9�'�'ӎ�A��)\Y��`1Ǧ.��M�A�ڵ�'�v|BQ�Q|ք�a��P(_Q��8��.5�g-��@e�]#P�;/*�e�Pd��Y���7m��"bߴI���e ��do�m{���M;o";[`ip�Q���]��䕌C�:!S�i� � �)��Z*FD�p�+��4�2=qp�љ��u���TG�(;��H1Z�q�i�9A��TB♀'W�dф��E�Ҝ�>!��Q�0����I�c�Pq����|�1����ċg�IJ@Aa �Ks"�3 ��}��<�������Xɑ?���ɁOXu�Hʖi�L@��P</�hp�%'XY� �'_��@K>3��AB�)Q������^ �q:0�F�4��A����UB' |�a�	B�,��1L#X-�]j�`��:���቞��6퐳c��KF��'h�%�oEH{&(�8eV�2�J̡�dQ�f���c&��%c�Y�G %{���1~�hz���WZ0�Y�-�k�w!J�#;��+�R�0Ә��q�3x�L�?i&/����=��k�|�x�QGDm6�Xp��[)�X��
�xPD��cI����R˅�x�n�a��h:�Pp�([�5J�HѦ��RfX�8š�'J��00sD
i���i�'�d�5&E	Q"p���O��ԬO1	�Z�	@݂n��7~�<5�s�0T}PG �zD��̓��?I��P�u�e���z�,)�b��*j	�!�95����w��C�94����G�)7���	���9lN?m`��%U�v�8`"�/٢%[�9��F܍h����%&�-�e�"�N�[��Ө�	�rM�4Qd���������G+U�d�X��؈>ք�b�yz�>v�ISA���"�(�J\,x3�c�4V�`���-?��s҅�E�fP�T�z������$YD�t-G�^TI����)8��[���ߛ�6E !��DD���R �"wV�i�M�H��h��/fp)b'E��*uPф��GA���" �&xF�A��ҙ3��HG��?Uժ�Bs�G"O6�iCO��vw��Gyb�	?WР�j#k�"N��k���hV˕$;�~�Y��Q#
���.g�V]��,��&*iy�I�l���PK���F	
F\� 8"�;@��q� �Fy+2�́Qxp��Oz��� ���z'a�7ÈOn�afoo�޽`@ƉYˎH�Mb�2���M݊b��UL�W��Im�Ι0�FH\`�'��@����H@���C�dX��e�#�M�ʄ�.=:|x�%�*W��T(�^D��A�,�N�"u'C�Y�������>\�iK�Ȏ(f��l�e�{܌ģeе"���2^:�*�I�sEV�Q����z�`�i�L�,��`�S:\��

4���餌���:�)���{�hө�M�<Ւ���Z(@�����:K��1�p�:ŉS6M-"x����7:O��y���u�(�e⓷N+(x��'ݶr��m�p�%�΁��,P�^~�u7
Z$nq��\�k�Y�G\��?� ������t�QfL�)p�QX:-z$�h~r�����X2$���T��Za��8jc?��t�B6tS�QR�AB�G}@�'�O@>Hץ�&5>����}&��¶uW�MSëBah�O -:R(êl7��	�+�8d��A�鑡%�&����
�e�,�[0���O� �kXw{hb�	#P�ay�oR z^��Ҵh 8e��He�ܖ&�.�w��.I���&_�?a¯�~V��'�*��
� ��G,���i��iQK������{ɘܙѪ�5���tϝ�L)�˧r�2H2d<vt2� �D�2Y�<,+�BH�1�4���K5I1��������FT�t�6Y�{a$S�UR�%�[��L�:d��72ojx���U��hA����:xs�%?DٙK��!.@+�H��1j`l�á��
a�5�66m�>�9�Ë�K4�LP~��e�S��H� ��d��ۅ,��űE�����O�"����f�ʽbĆ�%��=�
vh� �H('Kt`r�Z2r�.��!'Ǝ�M�dɎA�US����@�Ԉ/���0�+WD�쀥bE"K"yk8�0Ҭ
�P@��A��$d�)�����#1U�T��'O� #E$<�t-H��!�	Z��p�d��N�*ș@�S����w/�����R�	v 	��_����gÃ ���i��ȇCƔ��b�8q$X�i�u[�h4�ɍl'������dàaNhp��	�	h����	�s�LA bEd�s����A)�2<-z��d�P WE�����d"MOZe$r�R��M��8�H����,;$ �2���EӐT�c�U�Ѫc�ig��Ӈ9�@��� �-8,�bCDEҤ��R,� b>�I(�B�@��|��Z/��Xp(��Y�N����rl;ڧ~%�)�jL�>���Q��{dX0l��3�V��B玷7?�hʷ�\�Q�
��*s�xK����x�θh�O���!��E��\��b��t܊���:H��BD�'/�lpG�/��/,�t��c�L�+ �S���B�	� ���� Y�{� �x��#R�n�kr
K��9�N����'#0�&8)���L�u6���P�Δ n�r�A��ܠ3��H
2�@i�4Ul0k�#R�w�|Q!a����Jkܥva>/l�e�,��&�N�1�Ie�Ыb�$|ͨ<0핞a?��I=+c�m�w����3%���$`2�6� :尰Ȥ#֝n�J@��C
��A^��0!X4��*'&���'�Vx���S=��m�6I�aط*b����!A�Lpӄ쐄x�R}�ʎO�O��B��G���̩�L�:O)�Y@�'=����N�`��I2aO��s�	 Dc��~h��H�,�g��� �2e nAQ;�Z3C���*rgه/U���'Ҝ	��$VS����d�?cT�G-z�"�&Y�S��)t-�. =\	(T�/Ve�Y
�I\3B߶�j���)�s}"j#8�|�ҭS8F<�p�ȜU����Ѓ�/�61�S��`��d��[�������X@�P���w�e�0n�R���F��1�gW�L14fVQ;�^�(�摿����	U����@�'��=��Eע}�\�µ'ՅP�X�Z�h�2|*��H� 'bE{��K/H���' J̒ƨM_�a�T�-��MKŢo�>�B��Y���	
D��a�LH�b��	����HBb�?}��J&IB�Zk������)�I{�+QT���� .��L��^�6߲���rDВ��c۴@�i	2."�3��T��NYU$��)36�Πo�!�D�;���Q�*7 �A�QHX6���s O��`�j#�?�O�`R�Q3G��M�Vf��|ڰ��'��E�fT}޴�')r 3`�Bx2U��B�3�1)�'���˂�ߤ 8�B���8�{��]����)�)|a�w�Ñg��y�1
 �m�!�J�KTr�kAb�W�jQ�)X1}�!�ą�X��@9S�I�Rx DJR�ɜ �!�Ĉ�WF�`��Q�9O�#�Ӻ'�!�D�3��q&$W2&��F��2I�!�D�/�F��q�.$T���D�!�Ć�	��ِ'�+�6y$�-�!�D�{�D���ڔf��a�eR�~!��ѷpK(I�`��JP�F�C]!�u"�RPH�4����W#��A!򤎽D�� ��Áx� �w�]�!�� �����_��*�`Cv�!��-e��0�ʥ>����cL�p�!򤏉~z&�` �!�Z���"h�!�D��lvŒ@Х7+�)"a�ǫLp!��t�بȓ�õ���c��6n!�D���H�sG[�ҝ� �9#!�dSOl,(�M��n<!�Pz�!��0e�u��޽R��Ie�־ !�� $�i�e ��m��l�DO�(�!��
6���CR��5CDa���!򄌧`7n	Z�h�]C�HrMʙ�Q�|f�� %�D��% �iD��=+����еK'�߬#D�R ̐3�.�Y.D����5J٫��Ԏ'|�t��[<�YXӀ4?�@7 y
���
lc��+�"��Q-�վ�E ��')��~���7�;A�Y ]�,PCU�Ur?1 �xB�Ur>i��o(
$I�(LZ)n�k�e�v̓Z(����*�	óO����Oذ4KP	�Q�D�Y��	�a���	I�)�'W��ѐ�C��輈bC�����'>�*�)�'���B�&�4N�Լ !'P�M����<�}���	�%�C�Nq^\+�$�<[=�(T��O:��=��3� �0[�BA5t8yJ�jR�s�`1Qt�L3ո'����)�|rgl׊8|j�Y6aA�dB�8��h�~�<��<%>��feO�g���$N�%M�z��U�>�dܲ�(O��f��k=T\�#�	����HfT��J��)�'_���v�80�8"!�)6	&�l���$�G%���|�V&.���4�&Q��Ւ����Q9�<��=��\Ga�$��!!�U �k��ٲ��@H%�o��6lhK3?E�d��'I�@�*#�G.}�SE\ h�x��+b0 ��a���B�a],O�t�A �
-xY�Q��)T��P�S�O�`��)D89�$�p������#��N��6�٤�1�83N��|���"��Y�,�e\���ў��'X����^>� IP�/-� ��2\��iX!O!}lG�e���ۈy��� b{���r(�(VA��e�~�C(@��y���JtJ�d�g��EY~AC-����PI��
�|��c��k������i$\U���":0�b�!`��['g.y��#�>9�n��\���|�<ѷ�ˁfH��9���-m.ȑ#OGX�<m-�4N�m���o\ش��CNU�<q%@ΌY%.�R�ÐM���gIv�<i����<�{�e�m �QfNQr�<)�)_>w�U�`��LET�(�`En�<���*�4��Ā&UE捀r��k�<Iq�3#s�ѱ5�!eu���A�{�<9���L���:ae��O�mⲊ�w�<�`�%$Q9��]r/��c�.�u�<Y0'���ɣF�?�l���z�<�`k1\|8��hT�u���"���u�<	�`Ðc��)��T���u���5T�����Q�D?2���P�g��}�so=D�����aN�)y��� ����E�:D�����V5q����=E ���&5D�@��ǋ�L�x�/�S��k��'D� X�� $9���b�. �m�� ��%D�h+��4y�������epA��"D�����g�н*v�#"L�F�;D��z�H�)s�t�Q��� li�KP%D�|�RK�0B�
���=�$@�%?D��z�7�6��V�U�(9i�(D�@����@�ۓ��$)�Viq��'D����A�`D�����;e3�<Q�A!D����B=]Aƹ3w��HL ���J D����aȩ{�'G7i��b	9D�����E�p��lP0!ڄa7D�����ɥ#٪x��J�0*�� D���7
��<#$jI�m-���FB?D�,�W��hB�(T�u>��/1D��b� ���t
�o�zSt���`0D�`8�T2>J�ө�W�.}+�I1D��C1��;cF�h�Հ@�?t`�)��-D��q�W1r��c��<X��9D�ђhN�G����4l�0If\�;D��ا%H�D�'CҾV���(�-;D�<�$�!-G�xJ�	۱&|$`��b<D��`lV�Ho>\z�A�ps,�m:D����K�>[�(I`a/H�t�ea-D�4q��ҖD�\����S�x�!�e7D��UB�$"��,��~��c5�4D�`8���+R�<�aM
"{�-yb&2D��D�ٹF�d1�EʙO�|�(�/0D�XKa�0�� �tȉV�"I ¬)D��A��!Y�:k.9aQ ��fjFB�əQ��So�7l�l��AMa|C�I�2j��C�H�|)�qq�IA;-LC�I�2S<Ћ`a�h�9p����B�	�c�((��eC9�lp16��R3.C�)� `l��ĥqa�xѴ����"O���a��_sNt�����?��Y��"O
Q����:(�"������2"O�zB ���h����1���J�"OD]��M�0lX�b�E .{�-
'"O,����%!��H@3��6A]e�`"O�Ur���9ԥ�CJ8Au��b"O`�9b�������~�\t��"O~T	$�#4��E��t�bX��"O�t�ʕ&Q��(�iK�B�ڶ"Oإ��O���}��ӥc��c�"O�A����{���efY�"�|8(4"O�y��E���a�1�PUR""O>��	;/��)`�i̥H����"O�# <|L{��<v�F"O��
@NY4~�MRe�)B�ae"O���	��ۦ��ǘtS6"O����[$ڤk $]�i�:�)�"O~(���Bn,n��p	��f�t�s�"O�IR3nY��(M(ɀ;�p��"O�i�Ī�)�ㅩ�9�� �"OН�֦ܝ-g �Ɂ+�X�t�j�"O��yR#�\�����[w�ġD"O$�bԭ;q�2q��	~s�!�"ODyI�Y�{��*Q�2{I<��q"O�U�T�a��ŰK96P0Q"O�9A��0=�j�Ɓ׫.��`a"O���b=y��)z7ぶk(bD��"O"iE�ޅ,pR�6�	T��T�"O�-���+� Y���L�f�\��v"O�l
���._��X� �=��h��"OPx��<;�6PIBD[�{�I�"O�����ιr��5�D��W��d��"OM�6�M}��@$"�>�ԙD"O*��G
a?ĭYr�vO�I�"Ol}[$�ƭWȸ�2�ҫ�0��"O�u�����6��R뒣a�rЋ�"O������J#�5뵨���́�"O@]�ևV������
J���h�"OT���#��Q�ƸB#)�=3z�� 1"O�(Ӣ^�c��8J�n�. lD�� "OVq���R��A�c��g
�5"O
I;��N�M4��@d�QbUr�b�"O ��cI
�9�Ѝ����Uks"O�|JaU5Bǒ쒑�NA����`"O������s��ɲ�j��K���J�"O����Ȏ?`C����	����u�D"Oz8���W6����	KI��"O�ɘbC�dלmR�%I�F�p "O̝	��& �Nh!@��͎��"O�l���M8��P�3�0W`-Z�"OL��Rs�[Մ��8�^� 6"Oj��7�H&X���0"䊤x�V"OH�j�͟�,��521�B��
�"OX��ca�8��a�[�^���q�"O��f�'6�P�"� O�V�0�"O^0�	ԁ/@�cO�#F
b�#"O����&�� �d�7n�?�<A&"O��6�5M�T�;!���9Ь���"OB!'��e �(�}��b"O�}u�І :�� #�:T����"O�m����DtX�1C9�ʴ�!"O2ة0�?Ȁ�y �W�2{��'"O0Ճ�м7�n��������"O� H]��;f�a�*Ԉ��<�g"O`�@�K��E2�U�

F�r�"O����_v�}!w�[-{�kP"OH$�J% �X�����date*C"O���6@2R��m�&ɞ#Kܸ�"O��$@�Q�p����Y<ұ�U"OTyZ�h�*0M�1��F� L6��)�"O�9���!Ш�2e��}-���S"O@D���bP��`Q�S�|,���"O�}��d.����Bإz� "O���f��0_�v�JAaN�M����"O�$Q�M��P��CJ�x= "O���։<��ń�>V�\2�"O�uZ��@�fն�`�a�C0���"Ot��!H��}�t�r�.T��"O�<HD�#����@�?!~�J�"O\z��؂ "Y'^���1d ��!�D��c>��1����-�: {���M!���a���J���'M�"�!�ʄdJ��)�j�:! ����!���j~xB�����D��8|!�D��k�W�G��P��F= n!�DL\p 4���M"�JMIR��pe!򤔿y�J�Յ]�b�"Y˅�ܓ.&!��)6����CNS���U�A�|!�Di��L �I�ph���V`���!�$�S�����`�v��ʣ�P�!��dy9��J���"s��.L^!�9y��7�܂b�0l��&��D!������@�_rD}�a��)6!�˂n��'��>E=aעX62!�D�uL����&�	bF�u�!�D����TH����$����&>�!��e����!/]Z�(�0�P2�!�ğ?x)��9��**���7FS'[!�$އN�סF�w�N��e�� }F!�dɂ<F\�b�`�9Zln�a�܋{9!���>i;@صjؿ"B~M��J3+.!�D��Z��{�d�E5�h���m*!�DI	Sq�dZ�L��"���b���7c!���(l�0�E�!~��Q���l!�Ӽ1��z�I�e�L�#L���!�$[�L�n䒔3b��둅�6Y�!�d��NY�a��7t->�B�b�C�!�d�����Cә`�0�kC+^�'�!�dL�ZԜ�8�Wz���Q���!���?@u;��0Q�x���I�!�?d�r���N:��p��q!��_#d��Ę��DP��
PH�!�N��R,٣L�\4`ad�3�!�$ԍ<O(8��.J�e"9�d�'f!��)f�ތC@X\��qBK�=�!��J-�ʂ��"8�����*���!�$��R���A���7�$L�u� �Q�!�$V�o. �#ŮIV���Q�/U�[�!��C	z�FQ��D=�ڸVO	�S�!�P�Y2�p�i��s��a�틹�!��R+k"y�ʥF���G
G�J�!��;n8A�#!�o���!��/2�!�D\=n��蟱�R�eH*(	!�9H���x�#��ڱ���U�!�DR�I�^��S�D�}�������Ay!���40 Go�~x�=�4GY�!�R>x��W �!m��Y�]�"x!�� ���s����:�JǇ5}|T�!"O�I{R�
;;���#�Ș'6u�Q`"O<q����)�t���'�7�UpV"O,d"%�Į6�
B��d�2Ed"Oܥ�S@�@�`��ӆG'@i��F"O@��e�C�^�<���Ɩ'&L@�2&"O(�J�!ӬX�|���<��u��"O4Q�"/
�4�^�@NW�o0�t"O�
VM�:Jy�YT͔�{I�tj�"O���f隵1`h;�!Ȭ)�Z�b1"Ot9��1H2�X��`� rR
�c�"O���>`~h��(�c�ސ�2"O�9P▄E�@�$N�����"O��87B٩-R�#W�˔r&��a�"O*�0o��=�l�R�Ge�0U��"O2���Z7-�H!�J��u	Z�G"O.����8��H��g	.|v"Op���Q?]���B'{�u�F"O���]������-9݌�CC"O84�   �T   �  �  i"  N-  �7  C  �L  �R  2Y  v_  �j  Uv  w~  ��   �  D�  ��  ��  e�  ��   `� u�	����Zv)C�'ll\�0bKz+�D�����b�����y� ��y��%+�9�I��nI�'�2��\Ȕ�
R�~�a"�h(L(c�I6p	�X�v���IU4���i�`�^��n�ZL��&�!� A� H��G�$�H@�]'�nE� ,Bc��;fMr�@�'�?��*\'DY��l�
N�����3��IVIN�2�[�D��"B;j�6�1��d�O8�d�O���ա����fÃ�Ij��KFU����O�haS)���ɔ'�r͔�3z�4�'��¹&SP�A !�x2#d����B�'�	ǟ���̟�3(`Ӕ!�PHV
q�9��H]�DIXh��ɲ6v���K�o��uJ��'8�,c�'.�Q3�Ӣ��';��jgH�&g��}S%�ǿFp�]�/­$����<�2�ǽF3b����-���-Ce6��"��"e��4g�2V���'�2�j���O`�d�O�ʧ�y�N

��T3��̈́r��7B��?�A�if7������4�?G�i�U��ek���H��c��Ї�ݮ7��1"_�J�tp��O�O�'c~���N�y@J����t;��Ol��P4����[������pfL	s�
+je�9��&�I:�i�j6��٦��o�1%֍-�h��E�J�Qj�*��8
� �qVkQ̦��e�K!\L��g��4�j���i�D���<b�m���l;"kF��D�F���0c%FW#ڈ!���7SR�c� ٕ�M���iz�6�+)5b�엙)1��2�FZ~.� �#�6j:bԢ�,ɓ���ciB�A0�m;�#S�C�b8mڥ�M[ �i�����aq�w�K���9c��Xh��F,a�~(�7���\�7�DC���L�-���QG�6:�X�$-�	*��P�2 O'�p0c��*!Vn͠A
9+����	�,ڴ����3Nl:eN(�&䞮�?��+��M�(���㊾'�:�-��ٺ���?��c���?���?�. N�`�-��/p��O[y��L����G��`��Ĺ�j�axIϹaL�U�@g��0.�&n�i� @�Bl	5e�q��׾8�����'O�)�*O�͔'��4˖�^(�p�9�(C�y�\�����?a����?������O����H׻#�,���F�?Z$�1���O�A�n1 T�2���n5lz>m2�oC|��S!��Z?.���"y��M��Iy�o��p��7��OP�?}ͻ@�ɚ� �T�0�PA��>�"1����4�Gfº	z�8q��^��M�e�
��O�.!�K�1�|��C�]��%�ҙ�0�7m�B�<�rG^<tv�]�1�J�t��%?ٛ�g�4�2�ᐠ��	���<?	T���8޴YG�>��'+z�S6ޛ_�t�s��!n���'���I⟰�I}yB�)�$#�����R�R�
T��(^7a�ў���
�Mk��i���w��瓱?����"A��e�&�y�o�ßؔ'\�03�Or�'�BP�Rj_l�tT��J^*H ��I%)�(�d����I�x���&D�T�R1�O���{��G%cɠ����tr�]rJC�F���3�F�*l&MH�Ě��&PF��>Y��Q�N�s�u���"J�$s�P�'i�8^}R|�ajަ��(O���S�'3���?�O���&(Hr(|�Z%$�/�hس�B�O��d�<�������I�F"n A@Ss�` �e"{Z�$�OʸmZ��M�I>�'��-O��gڃ  �<�%���/���,1�PT�P��y��'B�'���ןT��ߟ���_)O��HC�C�	;$&�س��M}��ۗmJ�Q5�}F8���.Ԟ��doΜ���DIE>��QTj�~���pb��V`J�P���r����¯V�V�����d������F+h�$�ߦɨ��%'{>Hb�H�!l�����m

2�5��my��'����{�+�C����Ɩ�('���?1@�i��{��Um�d���?O�7-�O~���9'�!gٔR����� �����O���o�O��d�O�m����X�b2���5�eYXc=ء�7ْ<�Hw�R�2��u��I��rF�7���'`H5I��Ӥ��aP@c�14*n�@3��9@��MZ�JR�7P��J@d�Q�	7P:�D�O@`o���P:sAӎ\6|
ҡ+m� xcK�ty�(H�.�җ|Zw��V�aJ�.�r��	L�)�"�y���;��|B�i��)1v�W&@eX4���Z����t�����̦��dC .�M���$�L�i�O-cq%�1��u)��8�B�����O@��^�g�R��0L� >�n�	P���
U@̄gn�1p肯Hi�P��(����X�k�4(�#+[�	����Ɍj�]���S7H�L��ȡ0^� �᜘$��Cc�\���M+֟���)�	c�D-0�MFj��<X�O��'�қ|��I�Ƥ)�U��Z�J5�Dº:��=1�m��v	o�N�OM��o;s��tA�+g���&j�����I���I=N��%�AA�����Iȟ��I�SE��� �0����rA���m4o���S�@�KDdE�Ra��ĖOM��{2ؔCF\�aĊB��q҅��3�Xɘcb �/fb,(�CF\��.T�90�/4@�@r�h�%��'a"�@��J�/580%��
Ԧ� \��B���Ohb>���O��dF�l����A�"T%���po��W�|�O ��4LOر E
[4Tz��*]�*`�S�'�"�u��Ml���4�ߴ�?q�'��-����ό�!솭�B����*ФV�lB��O��d�O"�����O���0a�>�vN�]��3"DZ�&�8h�KBV�j����Q�Bvy+&Ǚ!�Q�46��Fj8z
ְ0F�y�7�ȓF-�=�bF�w좵`dTO�V���	".f���pE�SF��E���q`�	��?���hO�#<Y�K��8�B�ECS�+�'v�<1�m�5����ň,tԨ�pAn�I��M[������!H[�X�O��cԆr��D�0��qNn�Kmӛ5/r�'7��s'�'��4�|�
���&g,�P��_�&��m:� p�ȡ �9N��u��*mvͣ"�'����(�%G[�I��=^��x3�L� "ᙳ�Ȩo���yw��'}2$�x�Bx��d�O�n�&1�%L�,-�|(�L��P�f�'�|��v��hHs�/i.��VN����)��<��v������O��Y���2mq��@*.��YT�'剨x���	����	I�$��C�b�I�T�� 2�m�jو�ɲ#Db�r�'�&�k��<U�DI�m�T�D��6J�	����?I�) �:4�1@f'ڔq{�2�G)?�rJ .����f��
^]0���H�2�"�>�+S�S8z�(��X;+ǘ�9a%?�a*����IF�O-�dѸZ��H0S�>}����aLF�L0!�D�pN���ʟ�`�L�9�k�o�џ�Ê��(>�$�WG5����dZ�c���',剧v�]��l�̟�����8���|:�J��hܐ1V��3҆�S'�ǶP�.l��� cQ� �2�
;v����|����B�>��L��1���	�'��qJ��_�E������R�QL]*d�ƭRTN6�3S�.	+��O��c�Kr�r�mL:L��1:r�'��	u����Or�=�E ��kvک�F�:E��!�
�y�RGg�B'�[�4��=�5���B�����'x�I�҄T��F�y>���!K�"{�ٲ�G�N>���ȟ���۟F����v>�x� ���U��)r����$�ه�
�?H�R6��"EZ��a�O�GQp�Fy��2,�\��+J��qP�ڟ(���"I6N����R��5�B�ф1CL�FyB�ĭ]4��{����RR�ȷK��K���?1�� g�$��b�L&��#|���J߂U��OD�n�r���h��s:�&�42ش�?�O ndq�� �	�FP��;�n�
�T�90#�h��'�)��'>�?�
�vJ܋��dQ��Q�h���a�#�&Vb��a$�L+`�2���ce�$�(Op����Kx�CrE*��ub�G�,����'���(� s%��k�I�B���N2��j>�dF�N��'e�ɾ\�܃Pψ&G� h��ʞ�1 �O���Y��6mp��M�|�j�˂,U���O�=ͧ>3���2��-!A��DAb��EC�?�+On�[��O��O>ʧI��@`�4%�9rw�S���#�6'������?��+Ңv�V�ajX,K@9:�^.� aΧ��	��+̅ #$r4a� �ЃC�I�r6Գ��˸�AH�$X��	�q���b0g�
��R/� ,�	�Z���OT�}�'���rcUO�(�Y׎I%q�\�	�'?V��D�.����)�z�pl���$�z�O��8@U�9 �|�K�G[.Sƕ ���?a��?Y� @3B ��?I���?��w�hBu�%>]�'ځ]���ϵd��Q���]=KˢQ�&�D���O�~ͥO��xG!V�~�25JR����]��ĖQu���7�_���]Ñ�P�:%1�p��J��Y��F9mLQ Їz)>EB���O�;�R���ß�D{bC[��|8���?=�hu1�k
-!�D���ūg��5#�
�ɦJQ2��I.�HO�)�Of˓oT�ܡ�U)T�&�.^��$��m���@fx#"�'���'�>�c��]�6�)[I�G�0�Kb��Mas��u�4x���NXF�1�-���Q��aӉB����@R$=�Y�&�W�0$�8)�.6)L�����5PKx1yP��	u�Q��Hwȗ�gm��C"V�'�����ßM�@�d�O
�=��$ΙJW�kQC"R���� l�!��9g��(D��ft)
��D�<�'��6��OJʓl�|MIT����[�\��h�1�ѯI	2ĳ����?I�n������?Y�O�*�� ��xor��'��'R�e`�0���%KP�FLz�dE�c�����e�'���S֍]q*:��c�.cr���U�ja1�V��E�`G�	�f$��N�}�'��+���?Y�O�| �LI&6�%2u�U*M�|B�|�'��u8£_�/*�9�'j�x6�@��R+�	b�*�³OĲqS��W-��?�.OZ�Jc�O��?=�"����$���	)bA��p�ȏ+�d�b/���	?���OB*��u���	(b56�Xb���O@|�ۀ@	��T��#��H޾��O����Q�p�K��ŷz��� �!aO?-�$�q�j�;�a�&a+���/?�G�՟(�IS�Oy��	d���Bk	0xb\�u�A(vH!�d^ �3�/ -�pD�ΉGџ�{���^���2T�à	p0�)��P����'\�	{ ���#D��D�	ğ@�	�|21��U����"I��(Y��. �Ҙ F���>��):թΕ��T�|6��"�~�	M�~(!	�/t��je�΢_<�����"�X��kA!V��4�%�,�8a�8����Of�� ZV 1���/�F��3�'���^b�$�O��=�H�;BY*��-P5\#Lu�����yr�Sv��x���g:��BF^����H�����'C�ɣ>�d(���/�(S�J�?����Pσ�������ɟhE��D��c�Ձ�+S�u�>�;%	F$GpѸS܎�r�Rt�_�a����!�Z�UEy�\�� z]�D�ߘn�$��d��B�k�i�hK4���5L�`h���$v����_l	f�řl�L]�(�vob��'B�d�'�0�g �߶��2��!+�NA��'n��8��
a$5�� o�
PcM>�A�i�R[��`ǉ��'�bP���_�O�� 
�LF5}�U�	џ���,L�`�I�|Z"J�>���;��O.*�E��	�<�dɑe��a �j4>�|���F(6�<�%ϗ)�����O,2_��ⰠI8bU�p��qF �s. |�\����\(=���<�	�ݟ���Z~Ʌ�=��!�5j�5)c�h �@����0>q%-^��9ze�Q����Y��l��S�DXإ(J)I�9��	K�(y��Cy�D60�����g���d�1k�ԥ�V͙�u�%)πh���D�O�� t(���Ҡ��P�[�ܥ(��ۇB�H�P�~�����0>�HH�]. >�SS��Z~��'ho���Ġ�88zxFI	L�%j�N|���.a�Sv�ݛ�X5a�����:6�d�Oj�}
�'�B�ۅ�V�B�����{D~��
�'g��s�
X1P����Ȁ
�(	3��$�T�O��uIP���<E����k��p���?+O �pn�EP
���O:���O���n�dXqC
�3���1!G� 9�@HZ0B�%7l ���ߕgN���)擌$���@�O�	��ĝ�z��Zt���3�(�Y"�� ��ަu���3�)�6@��|"ūt�����}�YQn߮?ۢ�k'�Q+��9?��N����I~�'�4@�e�P0$��g�_1D��Ss"O�}RP:1v��ThR#~�8@�Q�$z��4��D�<I@,A�~>�- 5@EA��Q+��X�
6k���?9��?������F(50df��աY ؅ٕr�~�x1�^5�5��gXP���I'�<����Y5b���2EHl�p�e�IR9@�*K�
<H��dΚ�^2�薣�~�`hۋ��F�= |�F��><�� E�O$� ��'S��O�'rp�"∨8� ���E�7�~]��'{��vI�%��00*Ĝa�*�(I>�ǵi��S�̐��O:��}���m�.���4c��}�B���ʟ\�����|���|�#�?|�H�7���J�B��Gf�M�<�V���r��0� oS,�b���,]��<QW��E������b=�W��wN�dX���ʐAx�F���8|S�A�R�<)!)�ԟ��	K~�%2�1��ʴk���e�ˡ�䓔0>�#�uQ$�0�"J?��9�D�l��4Q��0��s%�(Sm��ۤ�V�b0��	yyR�C=r�) �=�T��P�b��%I�-2���d�W�Z6�$�O��a� |��m�E�
`�j�K#"�SPȇ�~J����jPٳ�9cVNLC w~b��F�p�W�D�^����U�C4{�>���*GR��;:�V����/����Z#��	*^����O��}�'2�I��!ǃ	�9�*p���'O��  ��z�5E/+��1�����OU��Z&Aִu�"����=V�v1���?�/O>�jBO������O����O\��"Aa�×�:����7�y���� v�|���C�~j ����5��I�D�r�O��UƒJf��!�/;@���`�!��3:�@�ט.Sᡌ���:�Y�?=<h2���1,Ϙ�	V`ޟ��'��]����?��DS'!I��s6`B$r`b��l
9Rh�B� E�VO���6��s�$���P�h��4�4���<��f��N]�,v�^	`�SC�;�P�
턑�?9��?�����SF�GX|�IÓ�o�m��/��mr��7A��86T�V�ۛ��a��� �(O �!��N�L�j�y�U�\^�U�� E�� �Fh�y��ʥ#\0���Y�	Û�(O>��5
�-�� ��`Q11X�l{E�V��B�':ў�DxR#^#?v�y�T\�6I)���yb�M�"��h:��\&��͛T��	��Y,�&�'�剥H�V�bI~ʢ#�0�z9a�Ҍ8�J|���]� ��� :�����ϧ̒-pçW�����ӥ]�,N a�Q-�\=a�L
;5���� L#q�+�8ʓ
�h�RJ�6-��&L
#(3���l&��d�-^����b��QfL ��D,ʓ[JĀ����|�'E2t�EH�"����5��Q��*O>��>��}9�Q�SJt����>%$����ɳ�?i�� g$d��牓bl�����ğh�'􊵀��'�"l����OIq�J��{�
 +@�	��^ ����OT��$5�Lܙc���x�x�ʉ�A�*�ZSiG9��'e�0�&*Ֆ-�h�K¾��'zc�$�<��I:@��٬A��W�K����Ҭ��iLrbx�P�J����<�A�Or��#ڧ�y�,JOmb���Y1��ك'�ѻ�y��]�'԰��)S�tH�P�^7��O`�D�m�<f�B��f(ʙgq����?i����D�:~~tt��O����Od��b>�V=/�xG+� �8�EMp�i��B�M�ru rI�-
b>�qa�L8q�$߼3� xb㡚�>��a�f�߿�>MS!��?6z�� ��X�`;��K��I�-PO"E:觀 v���*S���yhph�BD�!@�'��	��J���O^�=I����]��85�@��e�C�ō�y��B
X*�������(�&��cC���dt����'m�I1
������@Z��y���3������$J���џ��I���\wx��'\��F�9�-YEΒ#S;Ӱ�$EX��Ն��r�๪���):,8imZd�24˱�"+�މxW� 3jb��3u�D�j�=Ѓ��y�֨�㖦aل���45Eѩ2��Z�Ԧ�!V�0���cA��(���;���2�O���ώS���7�� ���k""O�ը��;��\x-�f��a�|��m�"�O�Ȳ�[�S3xl*K��f��Y{�Ũ[����O41��OJ�$w>E2稍d�N�z1�H34[�5#T�B/X�U�`�Vx�y�IX�3
a���?<HQ������(v�	xbm��a#�R��Rii/�n&>��*��2��*��1�Q�����OZ�d0?D��CjL�!jׯ��uZ��l�In���qB��T :%eQ?'a�T���3�O�H��c2`���)pm� )��U����<!�gO�?���DEV�@�Ba��
�,���ϡs�$P�` �G�"�'ZZ����5e�0�Ǻ
��j�C:*6�!I?I𠄒�xz�8�E�ͿU����#I6?�bBH�~�:��4>��3Ph��5�
`�D,>���G�N8�a$�2@��?���
C�'�>�̓A~P���0k�@Y�Oܯ'����`�>7m�6�(�4�_��A���GJ�O��Ax����=*�Ċ#��Xp��?�)O�H�FFJ���O����O<��s߸;�������Ӌȑh �;&�+=6��Π?����"擹�Z���O(hP���<4d\C�f�0;|(�QO��3�$E�Eƨk�F�!:�1�v�PaO:�~b�Ʈ9�F���m�-���9C���?	�Ob���'�R����}k&J��WQ�АJ�H��ȓU\���f��0�P�a��	M��'<#=�'�?Y,O9�f�+_�%@��K"%���U L�}h^y�f�O����O��d�c��|@� 2j�fx�#jIHnEy�Ϩ92��di���HLx���.�:��&�z���<�eIG�{]�A�j�uKD<xJ#l�����\�Y�T�� ��N��1��oO�k2��1��O�� w��RD��@M�"Vi��g�w�B�e�X�oZX����(E��4�jx���ODz���'?1O>��V%�!8|�}I�c%V��`{ԝ|r�'�"[��Cë�5��I�O�(��c�4@�,#B��N�0 ���O��D/(�d�O��Ӡw��� �@�4�)�
�8du@ �G4��E�f�sP��S�KN\�']x��#�%qj�u�!iѯq��I�n�25�Y�����^�J�oL+�&�"�hя���s9����'{�	�B��0:SG6M�YQ�Z�Z\��O���$țf�z�x7��)Y�\�f���O��=�'���J��h�0#�u�p�	��]�?a,O��!]�I�i#��U>u�R��ԟ|��!*kةFȅ4J�V���E� ��I�آtkA�S��@�P��X�@��~����O����q��j&�`�����V8a�O�p���Y8B\�-0��X"-V@�4jH�<�L�S6���ɖ'M�2�:��";�����!�3#��I�GvZ�d�N�)§)���Ǟ�RC����C�D�vX��l�\��b�,fP�ۿ?�F�E{�'(�"=��a�"v�DJ�ϊstj�B�a�2H�f�'�B�'�ָ�G�4C�2�'���'���҃S�8P�4@ȸ+���(ƪ��#��x���ymJ��!�ȖTȺ�;��I$��N�I�J���b�R@�g�S�$��F��,E`�M��N�8ui���-���:|��A�� 5VT�wTQ��OD��'�1�1Opؠַ
����ⓨd��;�"O�<k�@x���c��-�6�h&W����4��O\m�Rf�!a�m�O	!
{���W��	q H�@�O����O����q��V0P�H���,y�u���<�4끣\?Z���ڳi۟mn�(iмiX�J�M�d�'�<틆��Rl����6 �����f�x��x&.?�d���p���S()�?�v�UU≝SJ�,31���E��ҠfE"9�L�*�d�OʔlZ��HO�#<�.�(E`D���p-j��3']T�<	����PCziA'�Q�Z�f,��c�N��MS����$B;}��,m��������Ɓ!������(
J��	ߟ�:��������|�4	�c��Q��W3?? �sK_��%���ûz?��ɖ�Y����׿arQ����aQ�(< ����)C������7$p�CX x��Ԯ��t
r�� �����]̓5!�ɿ��Y,�y�s��6�La���;�:%�ȓ��Q:�hS9V��	�/�I*�h�?���4�J����M�0pp�7
�5"�OJ[��O��)R�Ȧ�	֟ĔOD���"�'�%������~�q�h0����'���'S u�`��IY`��6��2/��SZ�$`�4f~e��� ���� �(ӫ���TOVUZ�`].qlب����35�>����F�3[d@��A<J��,���=?����J>E�� ��"��%O�����R�u���J�"O���@[1�Tc�@Y�|�N�4�ɽ�h��MP�L͍c�ܸ#���k5���pӚ�O��٢�� <'���O|�$�O���Y��`�2�h��-	T(A!ME�-�v8�+ڵ'�6ٙٴ0#v�ؒ"u̧DvI�⿟�Ark�s5�$Z$��.y�@��TK�4�T=sdEK��M��ϖ-p��e��#�(c���?O��:W�u�u(np\4`7遧FN� ���æ�(O29r"�'����?�O��C�`��0�R@���a��6D��C�ՔgԀu�P6#�(o>�|ʑ���`�'%�D(ӏ��of����'Dfȝx2+K/:�����'���'�"�xݝ����'�:(Re˖�60��ĆɄ0}|�B*^��u�f�*��x1� )��G~bտ]B�rP$PA���1P��a��E�Ecʥ0#BGo�PhYYu�3�P.��ח��ը��>5L����I��\�4[&���Fx�J�PF����슼y�xi�C���y�B�?�h1�T/�eް[s����x����'���Z�R���4�?a���e��$���`�&�+vq���?�ӥ���?������	 ]�XH� �.A���@	]�~����3����p@�ͯe1~m�c���4Gyү��:�����'^Y�ݨ`/�0@M��G�n���R"D�`7������1
�V-A���'���W6�'�^�#i5LYp�B�h-�~��'qxĨg�[fx��5�ǈV4X ���i>}r��vƂ)�!܋h���rF��;Kl�$��Bq�]8�M�&!�O�O �	T=i�"����ٱ#�M/l�	U�-"`�Q�N��`tk�'.Q>�����2F 1�#��"��9"�3?I�nJ�!7�!(q�Ⱦ%/x��'ʧ*�%kb�V5YjD�b���/�6��'m�Ԩ�oL���(�'���bީ=�����`C�/-L�A�	�'��P�7G\5�@M����B�X����� c�O˼�b��b��5j!��Vy�8��i���8Y�d� �Gy����7�U��k�u(��Ca�ЇI�1Oq""�'s�a�H��@���D���d���y2a���0=���)	�0��`�.���@���-���	j�g�9���E�<V�b-�v�́0�4���Y�i1��Ǟ"-� *���!urE�'�t#=E�47|)>e��k�xd�)�G��8d�C�%-��G7g��K����f��k��?��._�b��rW��dFف�㚣V��
жqy��'^�(��X���v��B*�]�w��l� ���´&'0��$Ğ:5�D�vD�"o�����&�Z@�

x�\t�jܟ^*N���i��4rl�R��	=1�4��a�.�0�2��	���|�3�ڍLl株�n�s*�,PENUy��'u�����\/�Qc��}��+
�3�I�b3�\�ҿ@ۊ	A+B�H@��+�u���?����)M2%�:��OV���"u��1��D%O��uAׅ�O^l+�f�$����o֌D]��Z�!�8B|�$�5q9\���D�-2��h�B�*C��9�dSp�fg�;3�B,EM�l��� x���Pd�Nh���G�(E<�扉D�����O*�S�Sh~B��?0F��25)ȴiE2��G��y�?(� ���'
:i�nXg+]!�hO��F��Ň0
|�{3�B�vd4�0��ǉREb�'�R��%a�d1A��'2�'���OD2�9r��q����[��M���tF�"���8*BJ�~�BŲP�$:�b8�I �ޱ٢��,�e��Q�*��T�Ђ.�=�C���")ԏ>2�+�ɔ8�ܱ2��A/|s������%L�]����I��HF{B9O6�ra�C�&9�@H�+4�P���"O��3��?9 N$���2���B�ğ0���4��$�<��aA�1w4ܠ�i�������=QZ=+�/���?����?Q������?�O����΅S�EbCT�K���!�;<��0aW#�&^��WG�&q�!F}�� �BZ^���G�X� �+C.t�)���%�.lh�B��EjBmCw�J@�'��A`��?nI�A�7���!dP�)� �c��hO">a���6\)�����"�4��s�u�<!E��c�N})��2�,�A�XuyJsӾ�$�<)4��4X��Sݟ�ϧW9��Д�Ԣ&���뇉�\IBT�	��V������I�Vd���lQ��`�����o!��2v%��T$╫��,:�0F0��F|��pӮ5����%���s`P�bfr5I��+A���Y�@>Ĭ��fǣ��O��`U�'���3�|�@/Y����dNL"F7��B��,���N�TƖ	�(]�AT�  �-#�Oݗ'���Q��#fF�nD-,NZ�(O�a�`D�O��d�O�'m�����?�"+H�Wd�s���>_�b2�g;�?�5���3�`m�V.��#���T-E�hz�ΧߘO��,j"�8/mμ��
�	kj��'2pX�! �h͐�S���[��� Ga�O�l�d��"�� ��F0)��'X���?��O�O�)� �!*��2d����C��7"O.��sj_���m޶m�D��6�ȟL�p�I\%W2<��L��v����q��O��D�ObY"�K.(Zv���O��$�O����O��w'��^>�����."C.�AwP��&$lnm8��_� �@�|���aq�ڸ�ʉ�')ۉ&�P�A�+ً&�|�iѶ}�`!��H$�P�'Y���,�UǮ1#��g/Z���`�5?��D����If�'��1Z��d�K�,��9���J�m�!�d�� �v=�wNN6"�X���L�"�(��|2�����1O1�3�U�hmX��DaB8��E��U �D���O��d�O���O2�e>b�Iݘ	��u�0d��&��Ig��6%����ΎT`bb��@���"��(z+2P���.�:H+�B� v��]�E���#�/b/&�!���&�Q������O�� �M�.�`H��U..�w��O��=���dϧ&�ba�G�\�,���	�E-2C!�Dٚ~v^�H��BVD�A���!"/��M+����oj�o�ӟ��	�|2�L�Ku�(2g��U��	��a�ǟ���a������<�ѕl��d��l�V3'�ic@:�#�3L���+�kֽ�X�Y��V��Fy!E3~� hS�m�*��`�h�f� ��ų&� E!"�'%\�Z�瞻n�����$���;��M�*5s�+Zݣ��� ?"B�4�X`�A��^:@%�v�_J��d�ty���g�p� hE�p}��cr��!����O����O����)���\h�r�)�)T+t|ұ�C"z?���w�'Y�\k�GH�9G$���=�D�5�'���m��c� �N<3萄%,ƨ��Y))v�6-�O���e�#%�O��$��N�]����		�8]��֍dY2��b��l���Q Q���������3w�De��Pm�(`���5(����$!y��'��@��2O.֝���I�?��	�<��� IT�dH�4�N�#d��m]��şXJȗ؟����!OT����2:�$H�Z����'0cp���G��&YF��N J�2�'sT��e�~r��?��'�?a&�c�\���([�r��p A )2+��?)�. ps�a��%����ܴ )ZA3&���*p��0A&f0�95Fه_�5O2@���'�K�����Ov�������#��� ���QP/�Y��%b�6>��I� �<�D�OXi���?��'+Jd��Ms���Bt�}��������.^�g�0�Qd�i���B6<z7����Wl���O�������D ��<���&��xy"7�X�+��	� o�
�MC�'�?y�'����c�O/�t��K̄]����"1����%�ip|�!�K|Ӥ@��榅��'�M�%�OT�S�?��;0���X�	� �<�A��2�y"���>ɠUA3(T(*���1!.ج�M����?�-O��O��?��^�9PT�рC
#�4�)aj�2�M���?9���?q��?1����I�?�ዀ�?y��
�a�8?�T��|�b�$�<�.O����<1.OJ�R��G�9ЩQ'$J8G���1�I�&���?a�'纥�k?O\��R0�Ø� ,�O��<����	���͚�&��ik��#`��n�Ox���O��OF�O0�p����J$yǣϽ2*8hfM[����ICyR�'���'A�	ȟD��U���,D�n֠����ZH����)`�pZ򏈥�+��b�~t��,Zd��DMlU����s4��ȓ  fm��Ђ+R�PCtjO',����{��i�P(F����´�� ��@��q
f�&a�Mk��
�&Ѡz�)�?�7�=\����$:�d���:h�2��͕b�)��'ۺeBiڅA�(]�Gћ4e��$�0vN^��Ӥ[6R<�`!"��LW�O!��l
6G���N�Z,`C��D�
�Xt"�hװ,�9j��>dm<�F L�^]�@&���Y
V�\_B��o͋H����C�k�Huk��I �>H�B�Þ9��층��.|� �I�<<�)�&[(��y�O�OZ2�K
a��y��X,m�n9�B�)e�L$�#��~!�MY�|ґ��>���תi4}��7t�<C�d�(1�\�D�O@9Z@ (3i�n۱_5n�a��|��&a��$�'�R�*wn�8l�SV�xRѻE��PqŪR�@�����S�&�/ix��E��Ldq�ӡԪTb:|a�̴A��jb�x�b�����R�Oۛ�✰<Zj��.L��� ��jF �y�f�%���3?c����e@�ml��=�' EQ�8�GĐ*]Eh�g���:���*r�����ɾ9�b"��Ο���러��� ��"!�<-|�t;���\x�"ac�`�ȳ�m=l�Y�R��s^>q�ӣ&.�9b�O�Q�V�8:"�)�I��)K`@�pL�Qz�9�R�����3�đ�v́e�VC��=h�Q і�Ԗ-�Z�+rA!U�N�a�iӌ7��O�IP��Oq��Iצ�˅�#�
B@I��w_��j��O=�?����>�f��5,/�p"�@E.T''�e?���z3��`����[��Q�I�?��B��낒9@�rU��($�;��N���@���$o�H���O����O� �;�?���?��'уT=���U~�8��A�� �aVA�#h�e�i���i
�,�� Z�{��q�l|��f�&�"m��T�P���)��Jd&��h�'��Qzv�#�g�@U1�Orx`�vo�OPu{��۟���M{�����O4b���&��U?$�9��=--�����D��=�J<���2���m�T��C�E�1�'487-��a�'p�Qڵ�sӦ�d������ܨ`[�|�F�S�T���	�O����ɸ
 )��ޟ��'C4n,Ϻ�z�N@�s�j$����'Y��Y�%A?���+t�G��3VN�'��Q9�%�/#�`*�)�pl$��C`d��:E�ՍEmlM�#�9e��d�����S��e7 :�D�.k��"}2H QW�u[�-�l�N��f���yRKS>NT�2n��|��x��j�(Oʢ=ͧb�L�@'	Mu\��a,�;5�h݃�ٝ��E���i	�'u�r�� l A� �T��=Jl1X�)g���?!%��MC�$�:cwZH �
�'A��`k��?%���e_B��#I��]�@1*�'Q�5�~OB=O*m�y˳ƱL½����4F�"�����2>�b�� ՒsL( jʮt7*����i�	�_�b�D�W�)�S�?��h�t�
���A�K!,�tC�	�=��T��Ė&�J}!���=��+��4���Fy2�&���aE _x|��-J7@�
mn�ޟ ��ߟT0�i�Ygک�	؟p�I���N�	)�^ȣ�O�g���^+%�4 �Q/�!|�t�p�,;h +I�I�g�	�_�` �P�)��#␶{t��c��Z�5��+ݖ;8u�Dg-56tء%P>�A��ӆ�y'��Z����`7�����';�TH#��O��L�4��#=�WjF9@��T���gtM{a��l�<9��O(^��ʃ@�	@�z��]f?���{E�����|�'���i��$XN��C�%Ҍa����n�C�\�
6��Ol��O��DZ�{��?A�O#��b�D�h�4�b!o@��B5/�i�$�N�,��İ�&x8�� ��B#D�0bF�p�� .��p1B��b�(E��]�����$�1�HQ�I�%%�a�d�7XLp�R��ǜ�P�'�r�	l� p�C'FH�jD"�	��*wc�	��O�	"
|��sL�,�ԍZ$ӄw*����4�?!*O�%J1�w}Ҳi�Ȁc����G�^4b34fD�'�x��!�'nR�'q�	��6$��C�'$�v�>�uq�hл��EW�#��<q�	\�E���7�T�u�a�a,u��!c�bڏe���K�ƍt��QS�V+�hO~����'��DyӬ7͝v6�	����Cn6��ꗳN����'G������b>	Z!��==5Z�CJ�w�b	`ca2�P�q��ik��I^N2L8J5*��zU`޴���.|�l�ǟ���D��a�:X�6�1N����4E,@�D˛�63$�d�O@\*�F$d�|IA0�˩z�&����|�������O��eԇ�p���) �xrL"x����R�:���_!�\��(]�lf�s�3a���f͊>\���r��	��O(�)��'Ɗ�O�������vD@�A��8��\8w"OvЫ� h�"���7M���1e�|���T�?ʓX��sp/�:WzA��̾��ʧ�y�����O��d�"�Z( 4��O��d�O���w�T��gX�1�]�DJ�A�a���ȳ���A�<:H��[�~�Vb>�c�I��">bU�uy��k�ޕ��n�9*C�`�uB�c��u�P$Z�b�� �I\7@����;P�J`�7��S
�H����5T���&�D��5R��L<9v���N
�Tu%�%�����o�<��2hO���c-�'�X)�p�$�U���D�x��S�!ach�9��dXbM���?9%J0�O��iᰠ�nظ��L�=z�� �:��0<��nE�|+��>%Ҵ9���q�<AB���x�U� f��a��r�<YD��=�Fu����X�򵸦i�<A񏌩>fX��
�xt%��Y�<�CnȠ_�����G�p-�W�q�<	�U�� �9v�h�*̀�w�<��ȉ7���mY
�1ʀ��r�<Q��XCN<�h�c!v��@l�u�<����..�Tq�b�5_�����p�<	����F� ���BF ��c�<�C >?�
8괦�7u��U2vh^`�<��"��L�2u.X�^B<ZɟX�<)���?5��m�3!�8��
%&ZP�<9�x$���!�L#>����N�<�ql��5グ��L�N�b0��+�J�<Q�+��V���K!FE+��e�%ǍI�<��E^`\^�C*G5s�ȃG�<AcA�$;��&��<���PH�<� R%a#�^%4fXT�BJ^
Qe�ɓ�"O��h��C+*,˕��'���"O( �.Ǐ*r��ş�2nR�P#"OHóh��^YRӂ�M94Mae"O&"�O�813�y���ϴ4Mh��"O���E��U�	����jW8�(�"OPڒE�
�؍�CDY72T��c�"O��S��<����K�3-8"O
|�C*K6�¬Y��ی0(��2�"O8*u�D�L*ʍY��P4R�{U"OH@jJ)S
��G��R?�4j�"O������Z,��h�J
/f�lI�2"O��`�29�,áJ�l8���"Op�{@$]F�.�s̙�h"� �`"O��)S!� ��R� 6���3"O�]��+Ào���"�J�J�1"O�c��Ď��̋b�ܗ-x,8&"O`,�fE�;���� �1a�NT�G"O��9g
P��LP�ٰ\��1�"O|D+vR����ē&�ࡁ"Ot��G�<`�=��Fρ1�h+�"O|y��Kge�8��~�"|3'�P�<�ת[�N4��r��E@`��D��K�<���
-����I�$9� �s�@P�<�0h_�a ���ɸ;|��H�<3(X�s��zF��u���Έ^�<Aa��>1��d���T)Ov�;2��R�<9SG)( "a�*<����I�<�׏QB�����%�{��	`�B�<I� I.H��B��&vjVl��EWr�<��)F2q��ɛT���@��qBWg�l�<�B�c�Ƭ�G�g�0A� .Vj�<9��� ���Q�^�z�4]SDDj�<A�M-x����A�"s���&$�d�<a�)��dV��9W�2Dfc�<G���pB9�&E&$x����z�<AR"�~�z�1Ԍ�)Z������Q�<��-P;}���C� 9,,YY�
�d�<���$$ir�	aj�������|�<qq�]�M��Ρb���pJUv�<�# ť%�� yw���Bt�p�<�6�dk!h430���ר]F�<���A�a�(PZd��QIdT�� @�<�〥���Ԧ�-F�⍨G��`�<�c�}��k�53���s�<!��7 ���c�ާM�,��φw�<�BょH�^Qk'k���v�	u�TK�<y�/�U��ؔ��8N��肤�`�<�3���D9	�g�zu�$�E�[�<��c� h���������z��|�<�B��|s4<��^dHI�S�n�<�&��"9�e��	� !�d�w-�k�<	V+S�A��I1�a��8�:�����o�<Y��N0���z,ǔR͂�xA�b�<����ND�@�$M��u� а��s�<��ݲa�����
�S��l0��o�<�0��O�5s��מL�Xq&@s�<ٴEġ��@+�mAt�rC��V�<!c.Gr=�s�O=��AB��T�<Ĉ@�x�Y	ҩ�Ill%�1l�G�<Q��_�ļ��bl�\0�i�����<)1�� d�NH#��
]`a��Αz�<1҂$0#���E�V��o�<Q`���9�
����z�J�mi�<� Ph���=�����M'y �yq"Od\+!�0=��R�B@�cd�Sd"O
�ٳ��b�� ҅o_�}�\��4"O��QA�ÖtK��Cu�E:�mQC"O \ a�	/6�b@�@m@��ybc"O<��/U�v����*�$<�Q�"Ohذ����Cxő��@!��G"OΜ�͊�M��=��h�wq \�F"O̥�����2͒G&E\��yQ"O�y	��]'BF1��T�\�0;�"O���$A,���BM�(߈ਸ਼"O�25l��=͞:c�F�@ƈl+U"O��j�M��3�U���I:6"O>(s���@�r/�&B��퐵"OV]4o�G��)�F-�X�p"OTY���3f�L��`�N�]�,m��"OxpSK_�҉{1���Lڎ��"OҕP��C�f�0�����r L���"OP��/P�N���+��ЉY�"��t"Op�3�4u�N)!��Y�b���"O��z2N7-YDXQHf٣�"O��˒�9�­{������c"O����G�}̨���C�5hZPX2"O8="�����s㙲$]H���"O�< � �,e���SC��\G��S"O��z&$�0P�R�����,4}p"O )�`T��i�5~���!%"O�)��������!�n�p"O�@
U��/r5�
���:�Čp�"O�u� O��6A؁zBA;�X�i�"O�T"��6E����P�:�x$Z�"OU�q�	8�,Y�O�e�2���"Oj$Cum��8�����Tܺ�b#"OPj�7h���Ȃ
��M�F"O`�cQ��"Hp~PiũT���)T"O�p�����l�d��
1���w"O����+�!�b ��U*JD�p"O�  0�L�y�t��c)Kad/�y"OU�X���V� kH��qa,F6�y �;K4�������\�P�J����y"A�ҕ!DC(B��d�8cPB�	�}�hЖ^;X����0HB�V`\��Z$~�Q�op;FB�	�XŤ�[I�G�Uۓ��
r(>B�	,>����ČS:i('a�qg.B�	2��q���!iv�3�ş>b�C�	�;��(���[j�'j/^��B� j�`��`B	�2w0]hU�;�B�I�rE�� 'Ó3']18�iE�l]�B�I�:��e�a C�g�8����WBVC䉳{764�Am�J�f��g�՟�$C�	)�
ip j˹,�l���E�6BB�	�hc>5 `&V:~�t!c��^�.�B�J�rqX�H�5U��I��$p��B䉗[�2���H¬$�^���%ޣ.��B�I�4rnQ�q�Za�үƹ:dC䉥!V�'��(��K�D	��B�I�U)�p�p���ڱ�b×{HPB�I��X!�B �\Ũ�+`��L��B�	1Ж����3Tb]�t#���PB�ɕv=*�D��Y6�Y��^�T;DB䉡"�<Mۀc��u\�L����p�fB�<I���/�$��a�9��B�I.����c�lx G�����B�)� f��f��mo�iQ� '<j�9�w"O"�ñ!ɍ��A� 8`4���"O x�`�v���Ɗ��rG��R"O���kݥzf���I�7oU4�(�"O�� 3�E
fAĐ��'�,%X�lJ�"O��X�)؊�H�#�a��$;v��"O�p��%]%�QA��Z�/&L�r�"O���ׯ�.;
��Sf��'�.ʱ"O�	2���(�#^w~ xc"O� ��N�@�pã�E�AI��!�"O|8��q�kPjϊ>�bM��"OL�k慌�,T^������]+�"OQ��A�j��@��OYB�d8�"OȽ�p�U)Vj���hZ%R(�9�"O
�ҥ�<�1��?t�y��"O��#�e���kT�8:e��s#"O��i�˒.%�0��1F'��r�"O�$��A�($`�����1�ݙw"O;�`[�=�� �!���B崩j"O*���=S�H$����)��Xu"O֡:W�޵hM�-欛)g �Eq"O���
����K��=3^�Pb"OUa��Ga����S�9�9�"O�{��$8������% �i%"O�=��)��Jv���R����"O�u���^w��P��a���Y�$"O�������v����W�<Ж��"O�����T
�|%hs��7��M�"O8T#1���@�<����r\���r"O�XS��[�=�`�JB�O
W��"OD�z$
�-���
��.,@}St"O�[��W%y���oV�m�8��"O�(k3k.>% ��NK�j)ct"OfQ���Z ���c���,{@����"O�"̤W���7����A"O�t����:� 	`R/��İ�"O�4�� W�W<�����Da�a�"O���=}��P"�]�&W^��""O�m��bxa�	X�B��P3��	,G!��Q�R�����}��}д�ͺ,!��n��|�4�	A"z�8t�V !�$�- �	��߬_���ɐn�!�ʵ}t�@['!T��j�*���!�$D�/��C���$%8�j�u�!�䇎<���e*�8rd)�H��.!��?	q���ĸcc( T�J;p!��va��p󎚿0d���ςc�!�Č�"4E�ƥ��tjͪ�'I(�!�ĈUT�aZ��q��\)�dy!�$�r���F�+a�X����7{�!�D��PlM ���b���C�q��C�	oO�T�qkZ�0k��`cGѦ,�C�Ɍi� ����eȘ��QD��y� �5|r�S�D�*a��1���y��K�WO|��������16O�y��k.%Q�ƅ1�q W��7�y��
�ft�6!�E`�����y���rnV���<x&H[��7�y�ٜ��<B���p5��c�ˌ�y�IL%l>4M��K%|��H��y��ؠQ����AO�Q�V�.�y��8�f\��m�zt����Ȗ�y�R�x�z&��kx��{��!�yr/�>&��T�j6&�eEŔ�y
� ,����|�:1��?�5�q"O��Hr$
&�"���.�%,�$��U"O|UzV�"	�l�j���_�H���"Oʝ���ҕe́{q����3 "O����l�_0�Z`�C =?�E�a�pEK4d�?+X�-��%��?��6=�ҩR��ݘ\�$<����%i8�a�"O�z�h
[��Re˽lW�MI��i���A�e�!�m��嚫	���t��5F���^���E� �z�s�c��yb��D�������"tgF�҆�1V�!J��a��P[��ĸ4P�!&Z?������)��`��@	[������Owa}2ω%�n��!i�,,H�9�L�))�1F��j��� ŊԩS
��#�&3�O��C�	�� "�t���A�u���@�8t��IK Q�:LQ�ʊa�7=�X�x�-�<D�hI�$8ʅ�`"OZdɇ	��~4���J̘�3W�i���q�ɟ��x�D�	4fʵ��t��5�`R�2���5� �g�j�#�y��Yw�>�� 9��{B[=���sS�{Ә�"EƐ)Bo@i	�_?����Yik��EE
`F�Xȅ����T��s#�G$���%?$h1����Y5��[���I�B�Aֈ3O��L��?��(d��*�p�cd]�l+��'���%�a����zl�)f_>YB�+�:��Ą/Q�P`ɔE�M������4�p>aC &St1c�C����h�a!_W6-�eF�>vs7-���l"��%7����f����F�\c��Ձ�ڽ�б1���p�4�J�����i�ĩΕ;�>�?e�T�L}6�IE�R1b���� �J4��o����'n�y��������iQ��DO�B5x�`�eL;|�����P�	tԜ���Ou��c�m|>!�r*��Қ���l��v]>��"��j'¸9$�٫���d�qu���.Ƣu�4�q"ߤ]ZRoHkb-X��P�\��Lاi�3��O{4�S5A8�#��r�ȀC�SM�D��D4Y��y(���*��)���m�j��C&�?u���խK�>XӠ�~�b �W� Zܬ�O֑>}�P�P�~e���jV"�q����'����X	��P
�	ʚJ�q��%R�# �*a"��SV-52��MQ.8T�
B�8�bѪAS����O�}�")ۻfp:�+����y�ɗl��i�C�"�p�8��w���δ�q�?]�a��/ eF�E#�wJ��C׵X��� TnT=�2���݂)
����׫����� �A��6M�3r"��x�j��{E9&��eq�"d?��q`���msf=0F�X�8���'F��(6a��9�É�z����QMC �@qeF�~����G�9<�et7��L��/�Z�?�;��[�c���]~ul�x�+E�O|�H����"GT���N|ꓟB�Q%�'\���Ղç64�\Q�/+5��p1���9~�}iGk�5|���Ob�9��A��y"uL�!@��$�a|Q�'�G4 ��O���E1@��x���q@I�=�����
Gd2�1��KG$��#�*jpU��>����i����1�M�Q%���p]�X�q�ŧXQ&Ѫ���$��"|�\wK�;fiF #���$��'o�8J���<�1O� �'��9R�S/��55�'K���p�n]*`�<�!&P�qp|��'�.�~�OA�Oi֤ R�CB�ց����4T�4`sj����@�a+o�'��rRP�P�݉U���!ݷU�,��H㚱�b�
�X�Ru��>ӄ��Ę����?��B��c�L>�яav^����1��$�F�9��y�2DKv��#SbB9�7�|ʟ�Ke��8$��òm IP�L@�8a�Gj�l[�=�O�2�'i�����H�U9���釚Y�8���dIk�Z�3�i>�D��4@����2��6�^h�t���a��$�h�p���!v� ��^�3񤔅* "��2"I� Eޕ�,qF�I�o���V�I�o�i ��\�(a��6����m�F�ё��Y&�i�F��+ZfHb�'N�1k��x�� =	��i��@�G��,I����F���O���Q�1?���O���U�$?�ɐ��;����`�#[;i"�,�7t~`h�`�^�K�:�'h�����4���擉q*vT�?� ��&![6^��P�jWp�t�j�S�4ER�,<���\�M�f'�;=4mْ��h2�f�A")���чHöm)qO��|�0�D݃4��C��@w�]2c�hf�>��怛$F��*&Ě�;��q���O�%Rg�&k���ʕIϙ?'�t �V�09�#G}��I�`��h�*O��j�	�;�?1�)ڢZ�Z��iS�[�,(Ђ��,����>X� B��9�{~���M�}���:f��-8��4�r	�����I�#݀G������X�����#��a*c�5_8r�sS�C�	�j0�ő����@����~�O)l���ؑ�*�h�kT�r{>��˓c�T���ǈde�}ZA/�O��*ĬG�:Y�V-G�$["L�&���A!B�xࠃu�D|����*��$�i�y7LUH�9Vn]:<��bv�Q���Q���`r�A�oCTd���i�|�q7A��]��)��
#@x���'SDI�!#I�i��2���_,|�s3M$ړ?�Hc�f��")�gQ6�d�'���f��'����?aj�P���*2,k>� u� +@�V��A� Iк�;n@�M2�j�!�O.8��@Ȁ7�J��v��J�z����z��	/7
@s����9��L�~���	ЂP9!�l�Jp�J�g�a{2K�R��@�'Y���Ꮼ(t����:X�0����ȏXX~ȋ@���ɪ��Oh`���O��P�I�����JH� &����dӄt�#�T�S�h���R��?X�E���|U<����>����7iY><@�S�#�� ���ȩ=|
��. M��M��ɉ}����&?m� M��J!L�J%��ě�Wgҁ�`�"G�L��6�\b<�7��)�\�3���.����{̓He�����>�(��B���a�|z%��
2�ks*���Bzg��{�<YwB	�LFh ����8EL�9��(f�qO?�	���Ca�"6�z���]�K�����>@��TR2�ao��i�tp��H@��̓^vv�+��Yg�R@�zI �i�2���2�n�{ױOL�Y��Ε��,+�i>�9֊(��n��HM^p���t�<q���zk��	a w5(��E�-�,ѫ�.*�S�b�h� �� C��uV�%�4k\]B:B㉂0�Hl2�
�"W�2X��������$�d���>	'��S* (p���f*~@��2�v��Ã
!�y�?rnv��ǋG���DUQ�@m"�#�&���0�B0Y��e��2�|c6�(ð=Q��G���at`�4 �t��CQs��>)� ��o��&
�A`�P?�O��W	<���O8�8+V/P!#!�dB�!�8��b��34�}�S,�&�օ�/k����w��?;A�֧���A�eJ���	�ab�{���Ye��,ܤ�B�A� 8f61����E���������Ɲ:�~4�u!?��{���i&�Z�H���F=���nz�ɸ�'�7|W�\ku��'w��Lp*P�60�� �'�ĸ7mЉ u~���g cW�6e\�3^&-��Ľ���P���F�9M�Iår��L�㜷	˸�)u���|"�O�y[��
S谒tH�q'4�I>a!�(PcNi����/�v�[�4���|bp`RH��}���t� �<�M��ڑ��9���S��A����t�'޶ ;�IJe�4g!�%Q	�$�e���S��]�1��i�7ݟ\4e%'�	޺W���b��!ȴ���I Vcହu�Q
��>�q�A;M&�s凔%�J��`_�4{�m��9.����LB	Q�)�s�쩓nߣ6LY��"��M���y4�M={��c��<<O��{0�];g�a�l�d�'�2TdX���� W���q��R�?)G�i�8�"<�M�^w�bѬ;Y�����~�����*.~���kb'@v4ݢN>if/( �4ܠ���!��)�)A�r k3oA)J$x�2��;Xb1T �vs��pI�nN!��-�O���c�d8��WI�,yx��Af�
�:����>�&�m�	��
:f��ϟ�P���V�]�$1�C�hMV��Pd%�j$��� ��s�F�-��ySr��1�m�����'g���N�`��)�6M�(;��~�䢗Ss<؋f�6���"�`�j��l�3�I}�O�4F�*���`�6APd �GK�l�8H`����Z��hI�tDȰ�sQ[T�E�&�4	� �/z�e��'s��u�N,�TXDRJ�R@˓6�0��"��6`ƀ`��T㠄<Xr�3��W�jy\ē�DRʸ��!oHS?~���U	�$T��$J*�*���B�8)l�Zf��wщ'1��+���X/"Dn�J�s�2]I�~J,�s	ޛ(�k��yd@"G�ri^=bU�:�1�C.� d��~��ߣL$�Mʇ��#>h. Sm��A	|=�B�ǔN=��
 P�M��σ��Lȃ��~�.QiȤ�yg�'E`M	�e��;^���q�H��x��~d��*��K���F�\����!M��!�B��e�L�JE#���^R���&��+�v��@�D"��H�_4���$R9'���b7�ɟ}�qOֱ���.j���s#�J9h�!�~�b(�z���@�K��r=3�O��:yhy���9T ��XE%�z䉪����Wzx�F}B%^z�0�śb���vm�[b����SڼX"��L��f�R�R���g"P�w��9���qv��)�kϵ?��r��?;R�8F��Y��]��1�p?��n���IGF�
F�"���!J2�MӤꉂqi��Q� H�~��DH���,m�(���uL�l��k5CS�4� P6{�Z�'<
�������
"�Q�F ��8�

Zx�G! �l��#Nʝj\.��¤�7[T�����"`�ݫ���j��y�A-�}�I1 �Q��bŦQ��� �6-<��htA�> B��4k����C�6 �4h��(�(`$ �Z%��ZK��n�d�(���P�5RZh��\ [a��Cb�R�KZ��Y��䍋X�.���hQ�_�*� �IPa&^����Z:Ζe�Ǯp؄�bꕻ8y����dI�,*��A@8�޹��C��|1�y�bK��fnZ��PH^:x9�(�'�'�0>ɥLQ�x�Эi�`J�*M|��Sɞ.QF�HC�i�MW��V�*��#�Ъ`�(�[�l٤P��8+����jE�=����I��nv��.O;0�0�F~bN��vu1���P9Z�P�-�C6`Iy�D&	�m���Ǡ.*d��`c��g�`��-y���N��l�67-� lR�$�$��̓+bbI�F���j/:5�(X9mn�͓)$ؘ��C�|A�����"�I�D���Jo�5�,P	|�$*�4j��= �(�"�jl�s�^�a�x����㦅�V,]�m��Յ�)� :H���0���B�|��h&���x|�= �g�>���ʁf�֦u���G���� ��� HN�����MD;B(В���]X��)�#<�O��+�+��;��y� �	 �̄*��_!Y�(�K�쟘��\�"]�`���d�y�� �L�+��W1&n�D��W���Yp��D�N������LBrl(ғ#��-�E@�?'T����X�!84@ƒ;�,@�wFB�N;8����f`Mڄ�
^'�%貏�m��c �Ȕ-�axro��>�T���̵�
$��N�W�VI�7 Q�9��]IԤX"�h�ywk��ÐT���ąd�$ޛ��zu���	VBLzeǃ	���1�ջ7gX���\p�ڂ���g }z2�^����	�����v
ȗG�����'��lB�Gŗ�M{6�:#��;DU^�+���=Q���
�,�3$ 5��	�pO|�� A�j�	�g��F�6<"��q���C���4P����y�r�����X3u[�������$Ao��I��c�p�`��!د)�Q����%Q7/	�H��k�-l�a��%п	��t𔬏�(�\�௟�V�n��,@4�z��@C�%O~�XiA�F

�D2��'�42��1fi*,a"˖�wA��P�`c�a���2f2�8Jw+I T��4
0��!F)�,` �i��%�&���c�.B ;0��[�z�3o�mp�C�	�;3��
�`����P�FD*)��1��0������Y;�ĥA��i����'����]��y�lF��,�E��C�H�1�_���>�5�O�YHfuY5,.&�2U��9�&��@cT
fC��`�'
�̂Q�ߖME�`Á9$}ȉ�$�"3`��mC1b��c>�3��2��%�qL�7����ĥ$D�<i���%�RA���+��8q&�w�`YV!Yk�a���>E��#��'���0�*, �q�%��y2-�>>y0�p�O�dZuJ����ē�ȵ��7<Ov�4��/1������G�/����'�v�0GA?t��BS/2|��%ʠ�E2q�!�$��_t �VȾ���[梉-�!�$у:������6u�L�c�2�!�d�`�� xa-�i ��b�.O2�!�d�0��@�*
,q�S�*�2�!�]X�Ԕ(�.Y�,b�́p*��!��K��Q�%uj�����z�!�$ɬe��}���C�Z~������!�ɬ"6���3�ͤ~L� o��!�d�/�T��Fo@��8��Ŗ:�!��8Q �31�(>	��a�!��[T:"$A�)xm�]�&��
!�ŃA*����"F�a��k 
��$Y!�d$*�p����&Wk.�)c&]&�!�dЮY�E�n��Y&y ��!�dԾ]ar��A���C�xd�A(Y�!�$�{[u��� f�StC�<N�!�,��a�����7V:�C5aZ"�!�Xx�d�bFg�'6R��3���\�!��=m��� ��1C\u��RM!�D�:���1oüI�X�c���BD!��AaZ�c���-�hha1NG(a[!�d��'��a�D�GP��a�MC�"�!��W9>b>ܢ�k-%���aEl�S�!��ή��I�c�5�m�ĀH wj!��?D���r���B�I�g��{!���v�" h��)4��x�GU~T!�D�XT�1;Q�G,S�t�-ԲL)�"O���[� R�n�:z%�,�"O�� ��?d�z}��Q�(o:�R�"O��{���C���z���1j�)�"O�͓0�G(����N�6J"Ez�l04�ē���M<��W�V�G�>�!$G,D�8�h�a�di��֢[�¡�u�/D�d�VZ��iua�r���/D��X"ǒ!K�d�֥7�v9B� D��%�и��ŀP�_}��S�<D�$�SI�-^����)||����9D��VN
aXh����!$��}9w
7D���s�F5mZ>9'k#�y��4D�P�0��+����u���T:\쀐�0D�� � ���@�}����k!��K�"O&�{��`P�5��o��Y�T�A"O��{�,΃pܴ�b1eZ�A�d*#"O 5���	�\����4��ɡ�"O,��j�q(�X��<�H��"O���L��l��ё�1d��Ez#"OJ�#d��
i�Lxp�BF�����"O@�Gk���hq�O�-V��pK�"O��� �^�O�	�Q� �x@ �"O�!1�I�`�i�Q�º?�5��"ObpЖ�Y!H�>���fғNn0`s"OD%2��,Q.��؀U����"O����m^�W��{1��[�D)9"O�8���=�qbaM�m��ܳ"O0����iY���`�\�l��"Obh���0�.�I��S*ey�dZd"O�	`�/9�P��ƒ!����"O��kui<D���ᕄ�	J8�5"O�h�.��G��4)�B�G��ؗ"OP͸aM��HszD҆�·h,�"OF8!1�ۑR��bPD����"O�YvC��tv8I�@G�1�2"O�A�ޓd�ô	G�yP"O��0��?�8��#�{����S"Ot���+A#�F�w��]И=��"OL����1Y)-"D����D"O�x��̍�&���za$T�Y�ia�"OTu����l�|� ���//�ά!"OHy	6钞&AB�@&B�^8X-"�"O�4	è����b�S�@P�R�"O��c��V$dX0P�Bcd���"O~���G��Ϛ��NL��B�"OԬ��h�	
C������'S��L"O�p����D<3���n���J�"OJi� ��
��`�ˈgy -J�"Or|w���x��� ��!mr ���"O���Ħ��-�n�q��Y�wQ4e	�"O�����/c���:ጲ3F�0"O|�`͊"��P��#Z���r$"O�8���,Q��%x���[4"O��s��'�)�bg�-<��v"O���R��(�6�Z���v�Ja��"O:Ph�`��n��	c�O�� ���Xv"O�dHG�B�J`D#go�:&��!�"O4�X�@�m�4 Bm���{d"O����@2C.�2�MB.x�0�u"Oy�f�����푄]؀��"OE0d�%VRݒ��R�|S�I#r"O�h�1�h1$KT#t�j�d"O�0�ǆG1�|����$�6�х"O 8D�
%%�S�G���bp"O�ͺ���t�����D|�:%"OH�J��y܂)���2m"l�b"OD�p�
(��q:���$`���"O����B2͐���@׳z,�\ b"O���K \q�P�E!V��"O�e#$�	U�d�M��c��$"O -D����6݁e�]�L ��"O�$ w����[PEFb���
�"O�p�E�<%�a�]�w���P"O�d�Q�.Nɼ�2�S�}80S$"O��yt�G��aX�m��X�2"O�� F�Q<E2���@
�.�M�"O�4��K�M)2��_�I�"O� �1ZP�L$L�r��͞,���Pf"Oh$�!��?�p��/E��R���"O"��J_�b%f��`���g�F "Or�A�!{�8��ħ�?N{�eb�"O�R��7�А�D��IFR��"O��z6(�?D���A'��3u���v"O,Cc'�h���k_�/��Y�"O�Т�
?`~�z�+A*~M��"@"Of)�%%I;p����j�%<��A!"O�$9 ��6�l8K�K�~����"O�с��^�aʶ �A�<��"O����O�:@ `�M�[ײ�+�"OJY�cU3v�4`P�"�2e�Q�r"O~�qb�"�J21#ǆ<��"O�(�k�/���A�#�����"Oh��Q�L�i0�%��`��t�\չ�"O�A0W�X�tŒ�ɣd��7�褨�"O��p�*F�pBv�$�#vC\��d"O�;sl�U����v��ީ"Od�Q�g��@1�u��>P�(0"O�	ٶ�9h� �Ԍ��J�$�3r"O*����%?��$L��z��|-�y�,KE�2���]�Zt�[6.�y�LW3b�VQ	5еX�&��`���y�G[X�wӀMȾM( �¬�yR��]�� �pg?A2�H'I��yb�P�e�2��b�D�Q,	b���yL�1���{ bL0,���[bY�y���$8+W�V'+ L�4L�y©�XX��Q(�$j�� �֭�yҧ���,�"l�F���	��yb���Xpkv���aF�P�2� �y�K�0l��|�Po
�X�@��6�y[$C�$|sF+w��\	4H�y�<T�4�넩W�/!ŉ#˒�yҋݪz�)����%���!�Ļ�yr"U�"8,U�oW!ch��p�M�y���D��T蠃I'洛`+۰�yb@#P�tM	�'T���������y2����!��L/6y�S��
�yBH�:Y<t��U*� ht����I���Oԣ~�e�>ik���%pxpY�Rd�Z�<���Y�)����ˁ~��1P�DS�<��*J�M����w�$՘#�{�<��ɓ�Y���a��t�~�86�R�<d��A�B,	�h�;w/�T���EO�<aW�Ĵ,7��9��ʋS�R���+�L�<1e&T.dkF�J#Ή-�z��Ǉq�<9�,W�9r����_B����7a�G�<���_��T�t�L�$���֤�C�<�U��,x�9ЫP�w3V�(�N@�<cnŧd�\}Ca����B�H�|�<Q�o|�>%"ǫ�2X��ԡX|�<iqJ�!�z��Qɇ�9 q	¤�a�<Qu��. &��u�['~�@���[�<�vƙ�'���r� &�P A��EW�<!u.f�ܱӔI:0����l�<i�M�@��C�O��O)��б$�k�<!���y�j� �L˪M��ĭ8(�!򤌾K(�B��@9t}ؒ�C�^?!���2&�NAB  N/_�&��7�	�(�!�H������Y-X���PQaѬVh!��
�U�����$��l t�S RO!��ͩ8\��9`�RZh<���2gF!�� `tH%fP$�l i%K*a�l��Q"O������/��zB�7L�VA��"Ot���)Q��t���J���YE"O��mծ
h�dRk8���"O�i3d��'	j�ۅ�6 �d!YG"O椸��'�nmp0�&f�xh6"O����Ծ�R�P&�޽�\�;�"OP����)��ݒtI��q94"OX����C�ʪ�c��[�P��v"O�1т$`lL㥩�7G��YS�"O�	�`��6����"Oѧ�xI�A"Ob����ئ)��p����oըM�V"OF������RQ �Jج/qpAA�"O@ّp�\:6��a�5�Mpa���"O�)1�W�">�}9ԯ�.xc���"O�bi��c�hj�%C�4T��Sd"O<�Sk! �:��R�>H:8M �"Od�hr��9]�B���#ǆ.#�e	�"O��@Ө[�30]`�!��*���"O����ő�F����4�F�{z���"O�4�r�B��2���O�j�"O�P��.	��vNƊQ;i!"O���"��Gq^��� !j���"O���8K�r- 2�� �L3C"O$8��,�6�<k� #HI0{b"O�q��m�"�y�����Ӽh��"O��ŨKp,"=y�A�/%ѫ�"O\4�TJ��6�d]PW�¥v��3"O8�ka.
�O����s#�~L�I�"O`��Ԅ�f�T�2��oI��0"Ojաӄ�E$na�5kΓGR���"O�m��+�)c(�$
�J�,:;R��d"O��K��)	�(թ�%�$�"O�ѱ�/e_P��Qbגv6�г�"O6�	��K�P�R屗!��� 4"O�����l�����K*�R�"O�XÃA�TK�)޿Kp""O�m� v�<�rB݅%�:��"O
p+��b=�a��gѢd���"Oh�"�E�h����.76ne	r"O��á�^��)*�g�(���w"O����?ʨ�+W�;F��*T"O���#Ot��* �W�:�T��"O<R)E0.T0���!��U�p"O�ræي_*B}�e����U"O�s��Q����w	��f�rف�"O�d�1�[�_�2�2�Cf1LY�"O�����]8~5
�c
"&�ph�"O�i�`N��~%�UVK5��@@"O�<�TbND��uAW�����"O$)a�ݱ^��d���G��\�A"O��s�(پ]�L��2�Z�J�<@�"O~�9�.��b�s!�T�1��4"ON	��Eՠ1d��P'Ǫn�� "O}�P
[0on�)$ ۣV�jU!`"OD�*�*�h�p�#��,<��I(b"O�҂�2T|�5��3@��q�"O�%R�䏔㐘
�"� �Q��"O��S�T<O��J��߷k�J��"O��C�zI򵢉<�f�����yR���:����B*{vݒG��y�d�Vz�(c� 9x�-ѵԯ�yB@��e��as�%K&�$P��^��yR�A	eP�C�Kρ�؈�2���y
� ��0 m	�3|�l gl̆%�$y��"Ol�rB
�y��
$�z��V"O��e�"Q"�Pw�L�P����t"OWc]�;Ҷвǅ"����"Or�RØ�:���E�<K#
Ȕ"O��X�ғ_����$��:��ye"O|��%��'��8r�ՇX}�t"Oؙ���H�.�ĸ( � a�a�"OܼYd��7�F`Ig!¤^�,�#�"Ob1�pA�Q��l��E��d2 A "OBh �W�[��-�Q�D.y'����"Oni�A锐QZN��c�5.��P�"O���CG�T��a�I*�2b"O��ZD��_V2)P@V�b 	�"Oڕ�(�	�l�b)�m��i�v"O�-�e��,���i�G���!)D"O�H�ԿC|l@Q��L��va�""O�}�.�c�t�
��K;	�.��Q"O`Qs�f�ER��KqL_��H�"O�I�6mQ'Q�f�'�*��
�"O�	�q�4X�4��'��Dk�"O���_6hצ|��吰u�:�@�"O��RЬ��8�Z�Q�$(N�-
�"O�}{��C(P��p�<մ`C�"O�ȑ���'	1���Abj�J�"On���88C��Un
 v�pH0"O�A��^�N�$��s��f�Ұ�C"O�T�aAڶL��iq���J��q�"Oj��FJ�/�bͫ���15RH3�"O�Sȿ>����� �)SF�$��"O�(�3}���)Tl� xYG"O��ҍ��ัH0[jZ�v"O�-`��[�H��zE� bm�"O��Z��Pւa:��	�H�z�"O�4�'F0fRX��$��Dl��"O2r�MȬ;5,��l����d	f"O�݃a�I����e�S�j�h\�"O8����q�EzA
L�`"T,Ȣ"O����G<o��ّ)
�z�It"Od���F�En�Gh��A��"O*��#�=)<f�o
!K��	j��5D��b��.b�2���N�n��$?D����� � ���L�u�@+G�'D���	
Ah���`�:@��G2D��Q6j��z8����V�W (0g 3D���t YJ���d#T��7�;D�@�DI5AfI!풵t��Q+�+$D���6쌔e�b�s��ϼ��=�eD#D�`�Xy�a�c�;p^A��G!�yb/�1/�*�i�,�1�4�P�yBF�mX��ZWA M�1S'��!�y�ב`CU��M�*�`V$��y�Aݸ9%j��e(G�Q �m�Ń&�y���W���y��(H�~�0�Z(�y���N4�qc׏;M d ]�yb�Hd����-
%��B�KJ��yRm�G�X��^�rn5Zv%G�y�-�!V���cA�.j6�I)��[��y�݀{R���	�\7�h�Ł��yI�
X
&-0�M��R�����
�yR��_��b�@�? �
�@�4�yb��32c~��,ďc�U�Fȍ��y2�cm��B�j����V͋��y�k��А�7�P3�v-qVNM7�y
� "hz���Ѝ�F�<�p�'"O�:P���/�t"�Q�L�����"O @�S�DP?�������1;�"O8�iè�?_<�;�ư�@��@"OLMؕK�0;6^�`�ڭSor�z�"OL�+�$�G�x�"b�Hg���Q"OJ�k��:c�
�ہ@')r�j"O~l"0-�	9���9<{ �y�"OJ��O!��<�Gd]	Pi�Ȣ�"O�(���^��@�bcU!fV=�f"O��ցзb�Ц�R/���s"Ovt)��O�e!��ݬJ{��t"O�dQ��͗ �|:��
dZ�hD"O\�zv%��7{hԮ0g�lZ��߷�yr*L#F;�	K�7,6�x0����yB䜺1N��F�ք?�̓7��yr���
�{��1#������y��ܷF�>�@��[�x�����y���P5'ѝY��8{KS<�y�FB\��u*&oY�%�~��e�3�yb��y
����^Hr5���y�A=(](�����e:��ٱ�yB�\
� �ƳT��($�y2$	,{�dA
��W�L2RUT�
�y�N@�F��hJ��̞yfl,r���y�ɍ�G8���k���Ѡ��y�J0|���k�,&Ł�욑�y(�P0��G�Hچ�hWS��yB�,��&Bɝw�j1�ǂ��yR臸x�xh �2q��'�y��0d�Bdd`ߍu�D:���y¬�jMӉ�"n�PO*�y�%�"+H,X�Ë v��1h /��y���[Q��C�Ӧn�0����y�mɈ$�h&�_Ǭ3�
\��y�)d�.}q�޵[r���@��yld���.��Y����C� �yR�]�Bۤ�S�oK��M��l�yb`V4G�����SY�%K �Q�yb�Ǽ4`0�
���KtA���yr�	N+.�1@dH�ȹ���y��ԳL+�P��BZ�(�V} SO��k2a|R)2w����7�[#
[�*���ʰ?��'D@�[�C�)*LFx�PAǐ��A1	�'ur�ǉ��AE����F�l�����p�O�f{��/8�35@B�a�,y��'�����Կ#��,���u�B�'�X�0���S=���4�U���eR'育n*NC�)a�2�t�_2�v�&h�=S0�c�4��	�Kp�j�H�;�z= $�#f�B�I-E��`�"�X5�J~|B�I�O!
�&���Ax���$v�xB�I�_���8������q��Y[J.C�	?@��ibj` �$��w��B䉬6�4��Qb�Z0�S0D� k�*B�	�po��[�擌Hl��U�|| B�I0	����dF�*4�>��c�S(G�C䉪5�4�7�<Ѳ�4��C�	�v0�����M���Q\6�C䉁V"�2��S(=N���a��)��C�4q�|����	QXT�xQM�_XC�G|���
�8��(�h�2�NC��h�j��[Q�}�!G
m�HC�I( j��&V=F(�MA����BO<C�)� x�x$OD�!�~e��N�]�vAɡ"OL�w
@}�%!��ݎẌ́��u"O�xb慭~�y�NݬL�4 �G"O�)(f�%6��)��쒺y�����"O��h���#��hJ�+�b܀ �u"Op9�Vb�� Xy��D�T�"OHy�V>����G��Q��U��"O�C
M#���'�M���T��"O0my�Oԉj	���7!Yf�ԝC�"O� �e�ot�˲�C�l��pk�"OZ���߻hd*鍞b�,CC"O�T�A���A_�,q3�eKI�<��R�*���q0G�*�|���C�<	7-ܚt�Ai �΁^��1 ���{�<ѱ(�DC��A��j/����{�<���F�XͲ3Ŧ�Q֤xj"{�<yŨ�5SV��â�y����N�a�<�ACW3�Ţ�熀Pa���2"OT���FQ���ۄ�
5
A��@"O�I�قO��Q�􅈷--쑃"OH=a�,]�6\d�`E	(}!z(�C"O���E�C�s�إjڝ1��cs"OШ�̧;��z�
b�6��"O�٩p��=�|9
�)��J;�ND�<�  ێ'ʈE9�Q�4�C��<���^��K����^V�ڲGC�<��)�*I�.� �?��N�I�<Y���2�@�s��82V�
� �[�<rm�8	�e�z��Y��V�<���/��ɣǆP?4c�(���V�<��F�w�&p��<;���20!D~�<a&���L�r7�I9+C؄��XD�<I��	�x�Vx`C��8K�j��B�<q��&�T LY6^�$�3��W�<)�G�S�Z93�H�笐I�L~�<� �^�+ܸ`ÇKO�Z�t�hc�y�<���
&B�!��)Ȏ�@WO�m�<��jԊ:�Z�JT�Xe�y@�Oj�<Y��3��x��f_�Fņ�@Q�]c�<���[�8:V��Z��*@j�b�<�2ϐOU���G>%��a��G�<��R�1�$���:n�p)j�
~�<	��_}�Ƽ8��56�*�i�m�{�<�w���F�:�(����#G�d�C�v�<���=O��1JgƂ��6�p$'Bs�<��Ο^���BS�HޒyPq��o�<1�$\�A���/=�>�z�fD�<G��3S�й3����r��CBY�<qV.��杀c�:�y`NT�<9�MJE�>�҇'�!:�܅���	I�<Q �O� ���Ğx�+0%C\�<���ƕ�� �7j/a�A��M�s�<f&\����d!��-�쵑�h�<��!q$2]i1�؍9�<�g,g�<I� D%�49@�X�H*�(��f�<��
*��]W��=X�&�v�c�<��F
5�e���/v�]�Fg�`�<Y@'F=G������)W�&�x� ]�<����k�l�����&`�$�T�<I���RP���'
��cM�ɚ#k�x�<a!A�{���7mP�6$�J�MPx�<)�ö"���V��hR`Rq��u�<�e��#=�����l�*e�-��EX1Z���'��Q#�NӘa�.-���t�	�<b\wZ��W?~䋶E�zXL#t��?	�˶%
�R3��;��\��ܙ���W>���U�Co�̻N>� H"���//��a�5m$K�6�x��E.�-�㋓1]���ďS	&��S�m�bU�%Ο�E��!�:�/ِZW�Q`@� *Q����'Ȃ���?��xB�'"^���F�ԖQ��u��%V�g�X�X��� �I����'̑>��;'S.�Sf�Y^x����{��Dr�q�J(m�֟���4�?��'��(�!I���'=z�h`l�5C)��3eGZ�����O(���O��DR�vz����Ol�d��4h�A���DYV���;,nԐ�؝:/�IJ��>`�R��Ѧ��!(ʓ/hX��J9.}���X�Cm0�HF�����t�%R3e�r'��]�´�Љ�W;��ꢠ4}b��?)�E?o�dl�@`Uq����8.�@�x��'$��T>a�`K_� ��z��gi�`�`�%�K�N�H��,@s�mL���q� ���	_k?9F�i:l6�<�7,��f̛��'�2]?�(�� ^��(����<4.XKg���<P����?��|�H5Y���,,Ή㧒8@�X˯�@4"��T���A�(L)6��3�IWZ-00g��r�`�1#�@�O��dbɱ5�8��$��`����D͏o�BIx���lZ��<�O�h��7f�@D�������F�tl�Ox�b>�$��iv �ݑa/ߕh�8R��.�O\o���M;ݴ1���#���؝�0'�AE������E.\��?����)E����Ov7�?*|��N@�hء&�$������Sˢ0��
�j~X��L��D�pQE�Y�\�uǷ��Q��HT`�J��A��Yh�r�ĝ�F��@g]61�ԫD���6m�P�r*@+u�y��5f&��T����c�]�#!ޜ�M�W�A��	����OS>7�0i��e����.9���хh�2t�$�O4���[?!q�ܨ&^i��@+Qj*)�PC�m��?QV�i3�7!�����]+e,��U V�G�V�!���n[V����?��
+Bh�X���?����?�!���dp�$���.�0m��;�gԈ0��r��o���'�:'_P	�k�1G�$���0I}:�8�DS�9j��pG�Q$I�4`I�/�1OP聘�aΓd�}��Mh��H��S?�2��[u|����>�ŉ�1N����+xl5���V}�H$�?qը��wp�'�b�q��'f	��@6l��K� 9+\U��'���X�\��5Yc��?��+�NuZ~�l'�MCN>ͧ��/O�A��[�\�d��1�E�
�����sb�.r+��''��'K�DK��'�b�'�*,�pbJ�BZ�s5�8Y�:���"�'�ɲ���GN�%�v_�s^�tyQ�W7�(O��ʧmПp(�����E�/X�����.�å"_�`D\`�f��%��z}X]#���+5L�O���6�'���5��&|ˈ鳅k�!D��LB��߱\��O����O���'#
n}�k�"'�llA�d�� ��]0���c�' �l{CC��(�q�e�\2G��m��'�7�D�&���	ɟ�'�<3d�   �$   �  �  !  �*  1  [7  �=  ?>   Ĵ���	����Zv)̜��P��@Xx����W������K;G� �$��=� ����8�҆�
zn��;W�Ԏh`Pr�-QF:��A (P�J����9%Y
QT�*"���KEʺ[L�"%B�0鲲��nE��[5F�>*FJ�Ae��#1�2p�GϰOW<]ã&��	gXC�m�(^Wd�:�b��ݶʲ$t��K`W,W!��#Q��8>� �֨H�k T��!��Ȍ0R�xa�-y�qR���zF,Ԫd�*'�8zT���vV���vcC�p�����	3�uG�'�hY����a�`�~�C�%K�B�l���0���2T��;�#�x��3�i���!(Z�MR�Q�0D�9���UJW9)�M Te%�P�q�|�ԇ��Y���{���^����_��M#�"<�X�r����J?!��hO��I�K��A!!�J�.ִI�G�=M��B�I=r+JM���Ъ"p���h�(SFPq�4vi����X�'H�����OݒP6B_�D����㩞!W,���'"�'�2�~����?�t�OYD�4[ebY�p�&�{��Ï>���QqI	Nr5�蟲>\�(Yp�G/��)Ey"K|=�W�M����>3־��b@�4n�9d�@ Lz<0r0�Oc�L��@Bzv�b�H����O�E敻aGȤ���p�T��A�禙��4�?Y-O>�$�Od�d6�S1W��<����/趤�@J9Y���$*�L_r��"�8{0l8c��˖#�Иnϟ�2�4Yޛ&�'0H7Or&o�����ß�؈�DU�0��X��e�6�&�"7-�r����O��7!l8���]��P�n�:�8�'sB�L���#(|�����P�8�G{"�P3~���nIh����aد:����gڇ�
����ލ~-�uQ&}�`�Ey.��?���<���'��I��q	��Je��9+��"��ӑ5s�6�'��O�}�1SjYj�jI/NH�$���$J�֘%��E{�O� 7m�ڦɲ��b,�ձ��˭� �������MPXlZ��If��Iڨ�R�'��)yQ���e̡p�PL���PEaӊ�s�l�D�Ȥ�\[�lxB�0uT�yt��Q̧t�1�)Ӥ���K��g3Z�;����ݫ1	 %0��U��$*�Ax�.�9.�Z�Q�PT���5E��F�{$��S猫D"P]��*S�l�D�K�)�'V�V9��۳���*���cf�L;�'!�}Ba�285��3�n��a�a{�}��''�#=�'O��Te �9Q�V���%[�fa�E+��i��'������#n���'���'B�����X�a��ӿS�p����2�Ā��<hx�S�*J����˭|�iY���J<I����W�V�[4�;��ՐG)ۉG��v
�K��1l��s� �p��j�{�O��V��L��i�ͺ���2py�IH��^��ȼuK�<Qf!�� ��d����
�s!�8��t��ē8���%��L��q�%�@&>YzLᡶi�L#=�'��<�Q���ɝ�.Ti����D���UF�?\z�)���?Y���?D��h���O��S�r��mqE�6)Jt`��#����
M0#�4��J 괵c��'1\Y �C�x��0 �	�@���(� .;��#�X��Ι�Z�z��B���A�8� �|2嵟�{)��x�9�ԋ�]���;A#S!�M����"�㪄"V@�:�L� ��oT,��A�'�����iЖ8�Ty�D��:��59�OH9n���'��Y�&�~����d���l���e��B�~Y��E6�M�OѢ�?��?Af"�I�ȭ:b�O��}�W�4����ޡV2��:3×�1{@h�����hOX�N2�L����@N��oF�B��	),P�?�(�$L.��}ځN�B��A���,���I?���O��a�ø=Lfu2�`�pf���O������z�y���R�E�lkA�ʊ��''ў擴���.�T���n�j(auOз6��	)4<���O���|�"���?��"�8��/�.�BI�	�zl 㒺i�XE���^�`V��']X>����dC�Y�`H���E�:��'�3a{�H�>���#P�Ig�0����k��Ԓ��i$g�P1ß`����n	U���$O	sB;O�6��O�O�Ox ��@N���*��-�7`1��U���Iy8�t�B�	�@����@ܳ@4��s>�TʛFjӐ�O����r�|�Ð��o?J����=t~t}oZݟT�ɤ�Ll�1h����ݟ�ə�u�'L�ݪ�jن�0W �dVA�7$�o�X�@�C�DizL�dG�Ocع��(O��AG�����e��d�6�jq�gNLGp
�;$R��
���3Nu�,y2JǱl=�=ܰ�*'�� oJ�HQϏ*"�1�'m���{�azr�]�,�Q������=�Ǎӥ��x�*KS~Ω(eE6]��diF��8ZV6-F���t�|2b5we���F�Y*°{R��=Ue�� ��a��''R�'4�םڟ@���|"��z�X��J!x�PqSOײQ����� �t=b���'���2�PXḅ<��@�t���ug�LӜ�����tV8Y�gI\bH٧�G7I����c��<�׏�ןhC�A׃�\W�:6h҆��<	���#����D<SL=����"#NR��ȓ�`0(�H�`�I��G�S��'>x7-6��S����
^�$���:�(�+֛M^�0��@��մ<ޠ5���y'"nx��bL�(_��xW�B,�y
� |U+�Oѡ�v��*3<�)�"O�<�4��Jvs� ӳ:�P�"O@��dHI�mm�P��m�0t8�"O๵��{�����d�U�"O� q�	ڃ1ަ���E�=�.�`�"O���,�-�xՉ���Ǫ8ۢ"O&9)dhA,z���F�ɔ~<H�"�"O
�P��,B��C�/O� ��G"OrZu��v���m={��3�"O�� IY*�Q)��Ȏ�Papb"O u�F	�<	�4�	�</� ��"O�1���6 �DD��hݣR1Nx�d"O��#�_*R�:�v�-� ���"O�H e)	@������)�%��"O �e&V`��3���0pzs"OfP�b�;�3`��?ln�D�t"Oz@�&)M(9� ��z�B��$J�R��!��A��4cp\�?	
/O��Z�d�D�p��ۨv�8 �O�81�Y����:!Ѹ[8(1҇��3�E�r소S�����3]*�E�H��q�p|{��	n�J$��Cފ��<y��N��$��OƺvI�Y�%�~z\h���[M橐A	Db]��'� �!�X�<���F�9-�H>��
N�6y�-�6P Z����K�ȸ*�曪8�血I�.2�´"O6x�a�Ɲ#A��T�	�Hb��Ud��>�j�;l��*5���4�
�?!�/OZ೵��X��ڡox|��sO6��i�#4&e0ǁ�.r;�a�.\!_�V9�BgZ&3��� �k�!BGBC�?V�D�%j�;,  ���Γ	��<�'n�+`����ƃ)	�d��/�zt�d��"6֔9
q �Aqb�8��'�KI	<ܸibvC �܊����M)|\�,�E���R⢁�=9����KM�^l���	1�0�ʄ���0=�焔8r�'�r�#�	���h�Y�a����(�*2����DЮ`����*��O�~˓ua�C7�	X0��Ѧc���Q%�Й�E׊O������S�JJ%��J�3�0A�Aޚ�8�K��\2 ��4k3���ԇ���Ob,`+J��sL5JK��re�QaFrQ�'T(,�q����;��P&>m3G���W�\a*F&ɼB'v�[C��3��(��i���UC��R�����.�mH�ֹ�4���'8o�C�����`�%>ڃ�����Q��� P%��� $D��0<	�(�6F*@��@&`���� jܰɧ)C��Bt��ɖ�Z����<2e��'T�XlH�c	1��=�򄜄��p�#Aϵ|�=8�mH��$}W�Y��ؗM� � #�SK�O�&TA�jR�J,�ǥ)MK��)�jB%4/�"���28��а,ݽ"k��?11��*G0
���f���p�͝x�LM�����Zw)4�`w/�R��b���Od��Ь�2[Ԍ���Z��+B��a�a}R���	1t�[a<��+GF��SDp	�f$׾��˚�2��8G�0/Ƃ��H(u������>���gK��%��d�����O�i�VN�ar�Q��EZ��8��p�
]$G)�H5��f��5	\)w.�Dp�ꋡ4�a�cl>�S���-�lmc�%O�hnV��䘠c����Eq��O�dG��k��$6�>%��)Z�\��|��aV�N^�q�0"L�~�"D���o�f���m	�k�B�����-x�r!X$Θ�T�`��x��ـ3'�b���	��!�#T>�2�dĬ�'3��s��U7,�]�2�)�9���
7	Z��d��Dhq��"���Ż#�
r�\���*��+��@�[�(� 5ĝ���LF�G�b�>qw�N.f�`E3��_r�T{ m-O� ���+�|�kW呔u��6���
���L�
,�`����D�8�^���� �9KT�¶����U���	͙*1�dOpw�1q���3���p2�[h�䉪�~2�K�}���{�\?=xB�Kp?w��!��+U���@��*y�y/��EZ�b$�$<�\������O�	N9�������y�Dl ��C�*e�6-�2��5R3g��-��q�R��oy�� �����]: ��ʢZq���.N^?ؤ�}����9�M3�i�f�qDۅ��-�C�V�s�Zl��f>��F�3��l�����M�T����m�0tS�$ŵD����d�]�`.�S%�R]I�#�*����?Oq�
��7����NC+,ԓ!(L�	�м#$�[*qO��ĘUڨXe��,�Mz�>���&߮A��AS�"�?T@ 1I�a��I�8L�'yv(���?��L>��(X,~X���tc~քre\EyBKíE��X6��1��,�=�OAbL�O�
q��I�EU=ĀJ5��>Y��]�X�z��%��I]�w)�I����bq�9�Ώ���Tz�J,��+��$	��; �0�4b��\���`M�=h�sF��M�vb����n#�	-7������ $L��"V"x����n�5,��`��i7T�H �L�]��̰�-E5l�����#IS�ͪ/�+�	E�Q��a�GյF�ڭ8�J.�Dŕ��M��J���+��dY<Mr͒����Yu������9A>��U�_����Y��(��5pd/Ft����EM'��,I�.G#vb�y���,1��|z�;�,��#��y���p�+g���H�_�d��j�p/��(�+5�|ڛ'\����&��q�Dy��YQEF�9��ɼC\����.��V�E{��Ic���<Ա ��C����^9
�^�[�{R����䩞%hvh��%����ěP��Eص��=aH�c�%ܺA^��O��J���6�¬�S�,Ox� 
��eP&u�&�S�|XB�"d�D�{���[mB'*:�Ƀ-6L���e>O��S�]3!r:���
�J��{3,�<�Nh *,�3�ݐdhT`A�H�����̟¦�1/f��£	���V}�D�Q2$������$�k̈�c�J��sbL�;�h\� �
R��:B����%�e�Υ;A�!'�J��=��O�F)��O�}?\pK ��
�����d��	y$8����ĘOe��Q�OӅ�h�k��ͽ4��PT"P=uz4\j�'^^�J������	8��Od��Hdq�	�'@�f;��2gS��s#L�@�qO�Ӯb8�ؓ�0[&\���*l��CƮT4:d�g��zh����$lJ���K1�W&�.^�\1YGiў1O\0[Caa�(}+�K۰"�J���ϐF+�,�w��u���#t"�Y+�RW�IK	�=�y�,��\�>p���:���׆Π�y���*hL�����P-h;�(��|��>�X��)t;��cC�6�u	 /"D��D�?np\yg ���,d�ɰQ�0��υ7��L�� ����' ��+Z�r9r��0(5�P(�'[��{A�U<&���x� U� �5�VG�W�\ą��R��q/�?" ę`��-L޽�'�DA�7�$N �OPH���^֌�A�_&
��� b"OD��'ʟj�)(%K��W�FI�p�>QTR�H&�֝="^()O��1�(�*��S��C�*�"��'%�i����yr�an���}e��_>�mZ���_�~��gNb�'=�!ӵD�7eD�JCLNg(M���W$:���X� �� ��	�f>�̡cl�(�[tؔg��c�K�|����HB�z�J��� m�9�&�j���#�T_n�Վ�ӦY�G�!�)��ƛ�V����� I�a ��2���y�錸%\$;�N�3�U�&�S�f���Y�IS�t&��'�0��EH��~��ϓ;T�z�+-�*@���6��>���,�<�{voߊ9���c��.|kש�O4�&I�x}ƌ@B�ڇ]jl�BoǺY-m���\�ҦC�Mh�Y5�m�ɋ���@r�\��� �9`#=��3L����[ y�\�O��@q"�.x��4.l6���F �Z�r4+ڴ6���	��X�X�N��g蟼l�<ѳD�C�~t �B׽9QX'�Y�i1f@ͯN`\��(� Jk�9m�r��|rTO�M��hu�̷;^�E�ܸON��2eC�7�}���ѡx�N����'��-ۑ`}ښJ�D1P��9�g�Ҧ�&�\q���I�;���M3��IM������\'h��Y�D.wX�|��L&.f�4�e�-\@��gbK����aEE��\�^�p�^�6��'���'N��fj[�\,��cA��r��N��`#]�}46a����5�`�=�E�C�. �JSb��f��ڟD{� Cy�S�� �cj@02��L�N0u��o��7M(���K�a1�D�0�	�=j�|��!�p�5�(=���N��G��΀�'ʛ^�M�OH�PۧN ] ������.��i��T=k& �*�;/�^���a��Z���dR-��I��؏t�ܠԥG}-&�'i��E�[�pzZם[V�m��T×�9����eF�+j����GQ0<�X��	�~^���Ľ(r4�� �$1���A�r%H7�q��$��Y�puDaw�L)w�1�ՀVR�O������)
;r`q�RZ�J��$�V&(#|����
|$�Ui�&� `B"���^@��O���`Vdr�<'>�ٍy�gPO�5��k���ԉ�����u��A9! �@T�J�&��rC�(���o23d�b��!�<!㓇xI0H�4K�!i�,�C��3r�>x�ӓe.��ZUA��?�(qKҎ�p������uUY�A��dmȼ�׾En2�XQI��(p�v,q�E�P7T����ޡ6����7 �g�B�I	[��cte �B脎u��Hs�A]9z�V�bva�B蜾�^Hr�EU)Z���apm$���YU�w�T��>��L�3B��.ޜ(���&f�����6F�Q�a�<>���BY�dd�)R���'�2���W���iGJƾb���{�$�=\�x�DA�6$dc�$	���B7.�A�&֙`�����c,ړ	B���؝+�Х�s*@�d��,L��T�����J�^�z�d;��IÅP5(�ډ�����'�fq�	ӓw&� N܅'�>���i�!"�<1hrc��D]y��8{& f��f���F̥g\����e�B&�0ktoҟo�2H+% ��e�$�����������'|��e�$�4@
n=�2iIE�⥳��T�B��H��ƃHSP"'F
k��%+&� ���ݴ��ɋ�ʊ�3I��%	X�bD4��iW�<�jlV ��B#?!��l����Vg۠"p\��&Xݦ� H��ru�9H`�%=�Ks��
�@!Q�)��D0Y��+_�t�Ƚ�t 2�8Kf�m��*�t0�e���I�pi ����Y�n�Y�A�&T�j
�Һj���4��5ܔiA#)D/.�PW�č,�t�jׅ!R��W�B�)V�V�kz쵆鉈.�.��FbƎ���)��N⬈��*Kd����⟾2���� ƚ�N.��Bj֮Ln~�*��,.",�#�f"�f&+~8��`��6e����)gF��K�!�
35Ύ�/�rT�D�d�Bp�ը� 3#l��4 1gE�I�]?�eCχa��8)V�X�/ḡ�B߂�|!IC��6?�&&�BB��B�� �%{��C��B�M>�9#"DT��ђl����֯B*Zi�Q:^�-��8l�(����m�Ġ�ɢ@����Ο��'X��Kq�ڧQ6ػ��&m����-J�TG�|{a���l�T��("�Js�ҷg��ٸ���*���KA�R�*�0��)1f����.H�j�u+��)#�}��Ӫb��L!3�K;}�̤���L�=���)0%�$RC8�ѓ�\���؇�����6�O-te0��N�v �����5 ��BC�kVP*bM��g���k���@֓kC,� ��Kp>�p��N03h-{R���=μ%��S/w���3�΂U�����CP^��q��f���[�����QqT)�G�؛b�!���%�1O�#���e�1K�_��(#bXx��[�� Ӧ=;S�(
H��F	��[�<K�@ߣS���A���T���ɓ$	�<D"��AC���G-�/"�๒L��K"�00l�	��� F�K	Ĉ�"��a&�;O�4ẐH��k��D��\�Vo�#^UjA�C���x���ZX����� ,���x��̪?Ȱૃ�T-@����'�V�C�O=�M��� lcb�{��ĺ�0ઁ��L�n�) �F�J��P�e��&w��J�B�륮�.+�n���˽V�`�pƆɇ6+<l�#)K=[?�Dj�-'�7m��-��d�a矣(�|����/-�O��Ӱ���>�8�����o$�}���x�/�1f_H��-C<<�v4q��78�`����o����43Bc3hצ9�N�)EIƁBɚ12%��VC�l������=yu���>Ph�+@��)�P`��7��R���6�����j�&�zw��ej>Qj� A�)�������!�D�!����RH<�G C�[�����5�qR����Æ��MNyo3.�5��X������'U8�pT�'D0����
nf��s�F�!��y�$&�6�y�V�aR�x� .�6V�Z��d�
�'%EuKǤp[~u�G��.p+��i�6�놋�= �U���H����?���P�D��9ۦ	�	�r��� �x�I#r���(�]�DH��i<D���@��(a<��Ծg�!�D�� ��S�b0:�ۜ>����R1:о�,���D��O� 8T$O[��i��!!���"O��+c�404�Z	�F�
Vb^�r����P#�a|ύ4M��x� �� و��*��=���!,q�e�(�dm�<Ypl<�!��r��Ņȓh���8��8݌X��|wB�Ex��^�wQ�?��Fc_:f�� c	ޤ"G 8j�*'D�P�P��V�n���E�(��@��%D��``m�h�L��$d�3*�೫9D��I�哳xJʔ��J��x�\��8D���ńP��F#ah��ՐX�i8D�$�&+�"��Ax�@)!4|�s�&D��a!j��8�@8 ^P�c&�/D�t3i�^0��jD���r�<�iA�9D� p��e��x2'ά*⩪Q�$D��y��7d�]B��Jt����� D�\90�פ���"�+Ҡ��m,D��Yd üwE��)��3G~�ZՋ5D��,�/9��]#׫�4�q'/!D�$�GL.�e�WE�8LH��c,D�|��"��N	8��t�l�^�6M+D�$��Q���9ѩ� b�$���(D��7G9R��)9W����!D��)֦t>�l�V��wi��bU/D�� �@�������R��ɸ��!D�3���|��yUr�P���.D��#%��S��#	�%Zxl��+D��Q`�L���M�'�RA ��'M&D�%M@�U[�D15��wS@�B-7D��h�!Ȇ\8Y�r�����JC/7D���V#�V�D"O˪�p�2D� s�E@&��	!Ck�aD��X�C�I�G��1f��?J]x�{dH�U2C�ɂ֦ݙ�N�/o��x�W@Ծ@�C�	<A�x��*\���I��Q�u��B�)� �q�e
�H��z��d��}��"O�`�����ZqB"$�$���	-5�5��.��0�! %��f7�6�P�HW�R�I0�@�Փa!�=8�$����ڸ"�j���Ȕ�n!����iw��f��q�
�he!���%��@㏒'V��25�̸D5!���1i �щ\<gΜ��ŰP�!��T���X9�,�4��C O� �!�d@��4����:*���K�_!��;$�:�I5/áY�Yj�m��%J!�$ą$- �2�=���&�=!�D[�:��tb��[��!�5��%.!�$ЖfQ=c��4�P�'��!�$�4;	�A��#L��3եÃ�!���VLA�`��0���E�,N�!�䛹7���x���r���Г�]�V�!��5F�`�9Q
U�9r���m�(5�!���v&a)���-�<�Sfcύt�!�O(T�|� CW���b�!�$�
1���R����!$�LAD0!�Dߚ:>٫�/̱`�A�,\�(!�$G�C����d1SP� ��/@!��z R�
� 1�:�h&h]�q!�$M�#�2�c��ߔK��gײ�!�Ĕ�p���A�G@�Q=^ ���`�!�,O|f}`b�L�9��E��!�D��6N´��G.f�g�p�!��_�P��2�Z�W�~C���[�!�D��E(`(4 )�U�Ilm!���S���ɍ5��Y�A� 
$�!��l���ŕ�Ж�bF���~!�$ӫ)p��2H��P,�}�qm�;|�!��~(R�N� \�X�b"K!�ƱI���UF@�Fsx�"E�F9@!�Dׅc�2=���#[p���aN�_$!�d��L�
#���XĜɅAW1!��:|W<AW�C<&�p-C��n�!�D�	��$�d.�	[=��qO��/F!��R+bT H�堖3<�R���(z5!򤐯X/�I
�ߵ7$N׎XL!���7�S�z�Z(˂z��ȣ�'ӎL�v�X�+�=�Ƹl5(]#�'�Z	C��5&�͐����bɮd��'1l�ǆ@�}2DM�o��S��pq�'?�� HǄ8A�.��E��)y
�'�=�զM�,<q	#H�!A���P
�'� �)�aZ,d�A�bg�0@�v$y	�'�z ���5IV�
�E�(9	,@��'�0-Sb�_>Ӥ�8@' 5p<��'.�jHO�rV��B��+D����'o���	}~��q� Q�kq<���'�i	��7:��IXR���_��u��'*�<��H�7I�b�@�e�p�Նȓ�Za���9;4ib�@'l+f�ȓw��AJ��pT�O$(56(�ȓ9���hf�Գ:?��� 2�|��"�����	��b��a�q���RY�ȓq���g��H�2���a4���o,@�̓/t�8��6�ȩHE���r� �ځɜ�'4����k���ȓ=�~0Cel�"%p!B2S ��ȓ@������2~���D�� A!�%��vVs�e��YvN�	҇��90��G��8��&8��m���F"�f	��S�? �Hs1�-!_P���3� !�E"O����i�5Zz��r �4��X�"Ohlűs�,�Cў����"O4d)Q>��V�F�b�"ON`rA��b����B'7X!��"O��*q.�?7|��圜~��"O��@�mD��,H��ؚ`F�3"O����(~T����-�( "Oh%1�єS@5�s�Ø�⁓�"O����-1֔hd���q�>�ʑ*O����#(z�m��O�B��I�'��1�E�\�J�23CC�I���'�P{�KI#M�\��2胪L:���'�ՠЩ=j~X��2fJI�"D��'�azQ��� �Xz'�1<��Y�	�'d���R��jR���� ��4k^�R�'B�ȺN£YW��{��+rhXz�'�F��D.�H���+�C�"�TQ8
�'�p0#� YL=2"��h�
�

�'�8�ZD�>>��0��-i�>HK�'��Pa1�DZt��V7����';,aRg�����25*�5�����'? m���>��I@ѪҸ.�"�B�'!����)�]*�u"�K �#����'򖬹�`3	F���' �5`d�	�'�RL���9��m�Sk�aF���'� 0���,u� <HB�8����'Y�dx�㘭�R�j��F�UK�-Z�'���#$���}�v�p2��:S9��
�'�@]��BQ��"�S���x
�'w���(Ѽz�^ ����C���K
�'؈���G�&S��{Q_�$�8�y�'R�""�;x���	ҮP�Z��p�'N�q��`O	��Х� x�,H�'�� $�
^��쒗L��s�53	�'@���e�P�1��7@3(lP�'��#�eՓ,0�LK�ᝌ>�$ �'�8�x��*dR��2`�L�8�*
�'�:�P���L3�H�G'CI�d��'��ݚ�C \2PU�.i���'`~]�4� 1Ry�-T'(��a��'Y^xpE*�%Z�ɻ���p�,a��'��8c2��(�x@�\�����'�ې��6 �"��+j4����'�����+o2����%+&����'���v�@�`��iͪ7̠�'QX�AÖ)�tM)�k�C�*]P�'k�<�!�/KP��0��/.��H0
�'&���VgJ�f�%yBϩ'Ȯ�x�'�'� e���Z�S[���A���H��'��1�#15�p- �/"Us���)����h	`l�hʃ�ڤk��ڹ�y��Ё$���C�N�J}�q��(O�]���/.0mRǇC�j�l��n<��C�9���Xׯ�3b�2!�r��v߈6�!�a����9� @D�.@[��ӹ�p>L<ل�U$P~�0�$(���S�ADc�<��@P�t����# k��Õ�U�<�͂ W�x����*7Z�E�Bh�O�<)���0�x8��A?�|�@�G�<)��Y�S�a��J:e�t�X��C�<!�-�$~pE�v��8X�,T�ÜT�<Q�g��{r ����=!���FH�N�<Y���)y�����80����˓O�<� L�V�P4#-��Z3l��<X���"O��b2%E��R�`f�I�G>��r"O�"���87RLi��aڪ\�#"Oz��A�H�^�1�@�}���	�"O���̽Ag8(9��[X�~�h�"O�iA4*D�X\JP�ͪe�,��"O�P�ө�@�+�T�8�֑��"O\)��Y"?�PzB�L�VDxF"O(ِDg-HIP@��o�.S���"O~5p��!����2%�s�"OƕB��#v�~A#���&���"O=�0��K���c@���
���"OP��B,�Rm�5i�O]�ⅆ�E*!�$-<����	���`��֥~ !���Tn2 ��<d����ǁD!�T)t��=H�뉙s�T�y��}
!�$K��@"P�FB?�T �י!�Ă�"`�����V1n9�������
!�$A�l�t`��L:O��i��ɚ5�!�ϼ z�T)�T~��3nL��!�䚮4=��z6h֟vkV[�fY��!�$�2��*�kO`�tLJ�D��E�!�DC>U�>L{���4áB��e�!�C�gU��q�?/�8�`��˦
�!�DҾj�>L�W׸sK�H�vk"d!򤋲a���!tC@�d1�KMʥ^ !�d�9Z��X���

^La�U�!����*�Ja #�*�Ig���J�!�W#<�~�T�٭���P�!�� m�Qۤ�C��H1e�U�P�!��1����N%g�"�	SA���!�D8_x��U#�����Ů
 [�!��PmFe�Q&͹w|��[�D��!����2q���̱3✦^�!�$ �H��9RQ���|	�9k�/_*�!�X}
��唍�EqO�4
�!��]�\���B�S>�<|�0� z�!�,4	�a�2l��h��\�s,��!���8
F@��,�n�p�s� /k!���7Lގ)��$����(ڡ��C!�d�{8�ةU�Q��J݁�@�%2!�d�|�т&�|�a�N�!�$�91fM2Q�^��{����!�F�
�@!���;�l�+2���
�'��1��f���z�׭$p���
�'�f5{��ٜ'nD�3��!J���'5����٣Ҁ��F��A�46"Ol\�DȜ$���1�ҕCjrɡ%"O���,<3�05�G��V^ �"O̒&Ņwe|`�#'F&�,e �"OV�r�C8�8����(0M�(x�'gHԹP+�9:�c^��R
�'`,�*��ޫ"�a��'�">�P�'�)�p
�o9ƅ
��5	Y� �'���b7�Z|�09A���r���'����#�]=}�~0��̸z5�K�'�\��ŌLBN��%˧t[<8�
�'~����PLPr��w%�>h��J�'e`��E\�T�|���#�5[�.���'�HP��h�4k!����#��Q8��C�'��1���
"u\tٴ��F|zWP�<q`�_�\�-�4d�!kd�t��̄]�<�
ܵUleHf��� 2�sf�W�<iejۨ}6��z`H׉/��RE��V�<� m��D̀n�"�Z!!C�gLxqG"Oh8e��JU����4��6"Oڨ��/�~~���K� ��"O��5l�~����@92r*�g"O��!wjʢ"8��9�+�cmHc6"O,[��L���P�d��Ai�aJ�"OT�g�
  ��#�\�B�	�6s0$�1*��5=���O�(��B䉣1�HL!h�8|�(}B�)M4[�B��q��@�j�0�ɪ���;nz�B�J��)*���]�+�n�5R�C�ɋm����ƯƬ��<�FѴzHB�ɿu�D�:b1YYhh�C$5>�BB�I��L��r�o�@�	�V���ڍ�4��%)�A� ��,��}s���bE�5�,�'B�4#����f��XE&�6:����F�h'�4�ȓU�ჵE��RtFˁ,/���h��р%�0��0ӥ�7/�܆�w�^͚�����5A�L��&m ���x����D�ƒ|8��9!u���ȓV*��%�Gp^x��ʵH>����\
��_hA8�T�՗x$�ȓV�j�;�� �g,��,��ȓ\SblQ�"��:��T���ȓH4��b(� ~%�|jV#�������9����)�Ѐ�c˙f��Ʉ��ta����=Q���E�;�ȅ�ȓH�p!�	��p�(���|��7"ti{ ��#2���'�U�e�^<�ȓ7��K��b��M+�G�Bx�هȓcl�4A�����`��-�p��%�ȓ	W�@� �$bM�q@ōGh0� ��sl�؅'�.nA�P�/5$]��S�? �ɗn��Q�%Xp 'H�j�"O�����l���DVY�Ja� "O��'���D�2�#ƅ�J�u"Ob�B7���b�<[g�
*�p��E"O&�b� g��0Xv��5���p�"O��!2b)-� d��~�$aa�"O��Ӱn5J��	q�M�y��"O
�P/V�e�,푳� �"O�U30��9!��aÈ��oj�i�"O*��QN�v��@�֞F�xd��"O.�ɒ�OS��Ic��E�T�FD�"O�]�0��c�书���[��3E"O�PSv���'0R)����2XX|xD"OXT88kN<LhGG@DJ���"O\�1*ʧ]x.Հu�ښp�(�"O
�*��=�P���JE�>�ܹa�"Od�U��:5H�[�Y˞���"Ov���@]B&q�dVjgp�5"O���^A���cÝ7HݣQ"O���2#I>~jh��Sc�U;���"O<8`�����93�azSN��&D�����0 ��ȢA �L��T;p�>D���Ǭ�� �R����`�`��.<D��Se�:S�D!��E�_��d�V�?D��XG-ޝf�t�Q��RR�@�6�"D���܍T-H�؄�i:���$�4D��$gI�A�l�Z�
�=gV�T+�N7D��䤀��}�����#�r I�0D��i�Nֱ���1M�!G �c �8D�h� �-)����4�Q?}����$�6D�0���U2Lk�e��&�!��XQ��6D�H0�Ժ|���@2��N��8�n3D�@���Ф	�a�KF�Q��-D��{�f�qx�� �,�
��u�v?D�\ l�R����N'`E���bo;D�d)��   �`��<�*ū��'���7�>NALJR�$#����s:JآG�Z�&��Q�'��H�G��Y��4������G|���I���S�O�0h�'C�(n
Ԫ�/κ`���"O6��!���h��x����s ���$�O��Gz�O?$����:-t���QK� ����yӠ���O�6iO����O����O����?��od��R\�^�U��Q�!m@�س`K'�M$���J� ��3FE���剠L�0ɑ�h͊O@*��� �|x��-Ǧ� 2�D��B�᫁{���$v������h��%���Ȉ#��	������V��\�dˁ@�T�:f��&=(�@�p�8D�`��GC;y.�{��LcV�x�"z��Gz�Ox�'Ƕ��gC?�$GP�B�GL�XL�ť��&B�'P"�'��םş��	�|Z��d���$�Y�f�t<�dNV;7�h a�7\�Q`�lJ���<���.\�H�Q�I�	M}�	"���".ò䐵`�N�D����<��`؟(C���
+3�iP#��`�T�UmC0�y�e^���#B�]�p ���y�aU�T����c�
]�W�������5&�X��H ��M;��?��OD�11��G<X��{���-p��h��4x�
�����?��eVT�$k�J��MCTq}9z�a��m�Q�"�h��f̔z[}�a��)�Q�`�q",���Gi�@-�Ŋ"�� ��cB�>m�!��P�n&�m�B�U�
H�Va H����	*��hH��� *(�`�^� ֞!q"O� �r�G3��CSk_74������xb�i>]��O��C卉�!�,����г$��hk�^� ��)ۆ�M��?a/�X�S'L�ON����Vx���-V]�x�I�#�uoڎlr�m�%��#�="0�S�YjZI�7�Ղn�f��|��	���
ȼ<.�ych��?��灵q��p�� T��Z��@Q�>|�ST�e��t�?I���[�x;�APF/�`A��K��ퟘ��C�O��%�"~
Cc��&�v帀�?1�xe��c�/�y2��pH���G��4�|��v�����'O#��|z�J,Ӡ���Ǩ^|3l�.Iכv�' ߽^2j�5�'RB�'�(x�a�i�ݚt�&CAr��@#�'7r�u�Ё��r��哇"B,9P"�sҡW x��'?��O<L�+���8c-��]�Z�:1
՚��! ʻ�ڱ��	����˧��
�lӻe����u���4FF+5΄ؕ�˼	@PI�'��8#�j�az��̐e�����B�a���vc�
��x�g��� ���M�(�5�WB��!��7m�k���Ğ|r�A� �T#nY{(,DB��<�d�L9#������?	��?�������O�S�<��C ��	���& ��=af,@�x�&��#�ͼ"������O$y:uϞjLt��Zu���a�P*E�Z٫�	PXҔI�V'�:*C�mSt��'X��q�V�D�&X��#[��z%�� D�:5��(7I[%m#HB䉃f�mh5�feJ=p)G	E{���?�.�Dd[bMJK�͠D���'�T7M8��T��@�n��IR���)�d�$Ș�'s�`#-Ԧ�z�CS�0������УA��=��3;#��b�ԇ< 3��5���!�M�-( eBD��
'W��<I��5<F(�iA�D`-k�f_�9T��aǔ5�u���'gq���p��<qA�J՟T���I�2m!B�5b�J���D�OJB�,	��m0�� z�8�aab)	�"��$i~k�+;�UsaP�1�������d�o�2�mZ�����i�������'���X1@C��AА!�N@�M(0E]xk�)R"�R/ΚA�&�K�RΥɤ�Sy�'!H��24��<�l<�w-��"�rL���`�p����M�N�K*C�h"\1��#���>ba�8@������;	�&-Ku�쟐#�o�O��'�"~Ga��&������];gmjԛecB�y
� ��q� eTڭ�B�m9�����ȟdBc���Ow�ш�*��Z�rAR�!�	柘{��:4h�Iޟ�������_w�ZcZ1�(�J�� ;�dB�G T�������=���D�� Q����u��Oc�#<�ba�}�@ �EK�~ڠ�c+A�s���Ǌ	/o�T��)�0��ĕO��8 �� >�`祉���iŪ�<٣	ɟ� ޴Rc�'/�'���EFD�P��)N?�Y�D!r�O��=%>�:��M�w��Y��ȟz{��Qíh�DnZ��McJ>����"(O��8��F�z�ǆU�A{�9rv���X��H�W�O����O8��˺���?y�O��B2)#�`kP-��.O��{��Š�j����K�>���a#Q#�0<�g�<13rI�F`A�f96d�4$6�v���"�($�D�EO�w3���		>�$X�6��gT���1��O$K�D�lڐ�Mۍb%.�禩�$"��9����gc6IL��zVB:D�H9��H����NM�$d�4�FŬ>鑸i��P�Lc��ƌ�M3���?��O?�$����!`��63�~���4|��A���?����A"N�RAå�h�6m��-9��ܪ��U�4�I��X��%B|jў�@t,�5Gsx�9��lQ�D'Ϝ�,�!FFN ��5��5���	����K��˸t@n/�'Ns�A� �;!�L1�ЪY�>0��ȓ^N[��--��(�҉l6�y&��E{�Oo��4�ع@΅~��]���`�N��'Pq��r���O"ʧ&c��c���?�a���k�����1�LkPB�"X��v�^E�� �Mh�8��M���8$��c1�fY�W*P�vȁp�ԅ*�0ɱb�O����h�Ȇ��0�(E�X04�܉>��t�sʚ�*��S n� �)b��$w"�bA'8 �p��	� 6b�$�l�)�;}8�P��K���ש��W��-��' �!T���vT�X��&A�&����}��'�"=ͧD��H6k�XjYr1�i���U�i��'�ȭB3*t�B�'�b�'� ����U�hU84#�*Đ:��  �|Pt��s2T���T)2��	0p-l�)�3�]�L�;ueSbe�c�E�#4���V�J�j4��x��<4C�0CC�AV�����P�,�2=*�D�� `�!�Lr��$�ď�����O�$��I�L��!���	�`B����x�)I�sd��>���D�<�Ƨɢ9-`�3��%[JM��>盖g��nZ��hݴ=����?�O�z-�ć�	R
�4&̮n�Vŉ6�����%I��'P��'�Fp���֟0�'q�� ����3�X�����2J��SUD�BΪ����_2/�p��J�b+� cj7ʓUή1���[/�&��_���C1;��h+K"kպ���d��M`Ұ��̉+v�8 ��kr̓u�88�	A�|!j�o��Dp8���/r�Dr�'J��:7��&?��X�[��}�˓�(Or%���&�¹�U�I�Z��9�Q��M�M>	a`U)c_���'��ݟ���!�R 	#��*�>x��i�l,��'kb�'�N�0D�F� �̐�� 4n#��Q��Q	u���
'�;'�	ۆbB*���1S���(O��g ^"7y���e��X��o��G2er⍙�w>�a��?�땣�=�^�
��D�<��<�'�uA����@$�3D���fI��ȓ9ch�A�F�7}��\ȓ+ɺS�*&��E{�O�(�)��1����a�� 5[�SY���'H�8�f`Ӥ���O��'nv�y����?Q�`I\ؗ�Eq�\{蘒Z� !2�4�����\�@����b'JP)��c>qAag�*��"�G��e"˟�+���!E����R=6=1ra1?�Ҡ��)w(��O��)�g�(P�tȃ��F46�$L�V�'w��2�l�ɧ���L �%�0J��a�7JX'0�nuJ#�;D������3(�yr��B`b�qsE9��ٟ����4��������2��0�-]v��iG�����`c�@Υyp.���џ��	�8\w1Zc�bA�5BΪ_�̭�uA�x�j�I����?�WJ�#\�P�4�_���	@Ade9���,�<�aLR:Җ H��ZDѦ�郤J(���qK�|Fyb�Y�#V��؇nKsT��fJʇ���ybn9LOj�;$��!(�PZ�
X:]���+�"O��#퍜jXV��Aˑ�B�^E!��i�Z"=�'��:y�3킙�H��CG�>RL��ǋ�e=���?����?����v���O6��&&$!���7 ��a�H0E[��s '�=�p�Q銀"��'*���H�wX
iJV�PK0`(�k`{���*��TЬ���N�r�џ�)cH�OB�֨�x��g�� d�����Af�<�"فi�����Dµ34��zU. WX��Gy%.2nb�bfєa��H���½����̦I%��#�"N�9ƐMtn��\O��z!y�"0��#��5�H���莪p�`œ�"O�8�K�5�|��1�H�ѐ�"O��Q�MɣD~��`IP�|��"O���2nſyh�bƏ��il�,r�"O����DN7d	xT�c��#�"O� �!h@ ��I��!QM�o[���A"O"��jN�l�R�e�D�N^\H�"Ob��@n��MM��O��b���1F"O��:��;W�Xݚ�!X��� "O�����F�lh�<�sl�j��� V"OL�JƯ�P�:�k���:O�x�q"Ox�"଒�{�z��!� {ƺY��'TE�QDG32%��h돂O��MS�'���pU�� 'a\�h$ǹe\Q��'�D �e� �(���l�}��@	�'5d�$a��Q��9�Z�x�6}	�'>�|��jD� z�`�6-ɚ J�!��'�|iy�C5p�x�g��\�He(�'���.��a�L�
�HN/s���:7��A��x��̺p�d�o.|��Lɖ'M���'F�
$��ZE�Ά:�P�)
�'���wˇ���R�0F}�/�_����c�1h�pm ae�7�b�?�Po��O<PI;�0(<�Q�Onx�H:� _��R�W�k5���v�J*|`��X���h�`�Ng,����j��Y;0@ۻ"�b�I�I�7�"a%��H�M�ˢa�����C�4�(�(~��OXP�e�E�if�ũ�7�0�
�'\L1��
O2DO�+ek<Xx(�#���h*�%A���2v��n5W����'��M��LW����cB�u.S�'�}�"�y�б�u� .OnP���їjaR`�;�* ����Y˞�?��O�XƔq!tj�&�v-�w��Kx�p vn���-�s���_zdw/��s-���,�:)Ӏ\X��07�]9�.Dq���DYc���u��BL�Q����E���:u` w��n1Vؓ�6����#C~J�!�A6`~P�H��'���ˤP�D�&/�&�г�^�
��TC��%�dl��i,}�B^D��[���qy����,p��[�Gt�	��F�ē(�=j΋�tx�#�S/��Z�X��!�HQ,�0&�F;5�)���M!��|��)#�lųW��H�`U����l�������V�z� F5��d �.NZH�-�L�@Cǋ��'	K@0��"�\�yYp(�b�Y I�@1����}�cOv�t�rbi
�|�^]ʒ�ٗ{vt@bCBGg�&��a�Ņlٚ�,LcI~�g��j�8�;ԉfAt���Fy�TI��΁D�1	֨�=���M)�fȸ���2E�-_(_Iޕ��f��{�`�*u#C�Y���	R^y�LϺ�)���,c)�xd-����
3���C聕T�("#�'l{�%c5�?T1ԐI5�0:Ii��'C��AK�c@��L��z�џD��DA�Q���k� ��*���� �Y4[�%���O�ɪ��Z�M��ʧO��!�}.[J��3��7K�5P�ޜD]�V Eф��|�)���:f��t�%J5N4n���j�)N^�a�g_?ѢU�B�,-���N?E�ĉ.�I�?o�mQj�s���E�Rgџ�óMI�E���BGWMJ�ϧ&�~@���,a�]*&��c��kv�G!D�Q��ʅ"2�6͜��O�˓@A�hbLݩ�
4��4\)V(�''�$�*Sp�Z�$@���>����MQ���2�MX�0�2��)m^%��^���`3Lì ����ߡx���AĎ��LG�Ȁqאi����?����aSt�'V�e;�I|�#�5B�z ��b�.)�ԮH���p���>@a��V�G��H�L<��?G9l�x���<�5��JS1a|�p�ߟ���Φ����FY� f���$�$=b��g�'��٫dY	�*�ҫOb�(�&�2W��Yˣ*߉c亘9W&��)q`��|�r�9�4�J�?��(O<Lc��� ^�[�&O�4
�:1�x��]�.�h�qj�g�Om��J�!cTtcg��-t��un�� �T�3BU6���@�V�Ո��Z�R6z=Iǫ�>+IV��N� �(�{�K�����i*��bfF�_2�y�V#��)0�C�I�0e�����	���_�<8��W�����?�`ɂ�d.�ҕZ��0�sc~�<a��w�p��*���"N�y�<��!Řc���l[ zЙ��'Py�<�r�L�Q�ᕃN�:�ޝh�Fw�<Qя�7�ZlIB�O%l�p�J�t�<��O��X��(H��
T����O�j�<�R�c����!��%1v.�K�<��L ��%���-���ذ��[�<���&i�܈���@!<�����ƃB�<ɳ�Q�,�y&C%�^,����Z�<� ��`���qP�s�Y�8a��p"O�ܸ��O�8��Ɋ��D�D�a"OV@�lv��M���	�3�U��"O��r�l��t�\QW,��s;
�zP"O��sӄH#�`ɸ!,�#!�Q"OF�3<Ē2!	�XjU�C"O�P��C���N���IPyf �7"O�@���ގ{,�)ɂ���R`E"Oؕ;छ)|8���ڮI�(xr"O��&aD(����*ĺ"�Lzv"O�,"���r����C��<~t��"O�e�1/�*����'�v���5"ObAj�oҎK[�X!e�%���0"OP��E�b�6��1�ۙ6���"O6-1qOC�"(q���4a���"O��S�9vn,�WlN��D��'z`�)���-1����K�2l�fɣ�'Ӱqqꑮw]�A�d�4wd�h�'\�T�5 �z^ʐC��h+
�'9d����"XXN��V��)��"
�'��IBE�#e�E�A��+L@I)�'� Ӂj��l�Xۡ,�Fˈ��'���ȶ@��r��9Z�-�)D���'&�Ts�Y�{Đ`�a�%�"$��'>��B�]�2˦)e���tY�	�'�H�#�MĮt`���O�(��M�	�'ڄ0���&6U8�&	�2vX�	�'[���pi�~����C�7���
�'* i��ņd�JX�3f$�T@�
�'|�EY"�^7�Iif��-��+�'��XɃ�/�b y1�_�vtD���'m���ԬGbQ�g�bl�5R�'��#L��4�<���k����'Z����+˼g�u�s%�*5�`�'L��Y��W�6]���g�T�d��r�'^�(���(v��#��'S>��
�'{�dQ�[�L����/;D3�h	�'h�����7<h��Y`�[�M-� ��'sn1�g��7��x�V�ձH�`�p�'*���"N}��p��ܳpt����'Z]�g+
MtU��W_}��h
�'@��L�]� �SG`a��'��e(ugH,'���m"B��	�'F@51J��-*(u��	�'"�^�Gn�hvkιk����'Fa�b�*`�v�qq�3h�1��'�l��gR=u��L� ��6���'��dX��](Un��VB�/51����'T���o[�1?�kV�B�1Tn���'ʎT��d�*)��NA�:v@d��'H��!"��&�����&J�,���'�����F�'�fm��}����'*(�R���1 �i�t��`�,Y�	�'31h`\Z��tA_�K�Vu��'��L���D6&%�M;�$��AgR]�
�'�*S`�T`8�!�V�F���
�'mҙ���N�h+��3)�T8\}��'�����1�b\��Ȃ-]\����'�x���V>-��f��)e� ��	�'�����F'D�M��#�4���'�%�&�B'J��P: �(]��'�2d���L�=_�k�A_'\�E
�'3�A�(uT��<g��	�'���� �<E�ʌ�T�\�cdB����� ��)���$�~9{d��!.���r"On �G+N.�6)��_69-\l�A"O��a�e�< ҥ蒀ѷV*���T"Op�&�Ӌ$5<t*Qe��{�;'�� g��F�m
%��r7���z@�A��y���	 �t�
<�"���`̣lmޜ"i0�IV��~2lZ����� ˈeA�qR�lZ(�y��L>y�@c0	��G?�|%���8������Fy�:�x��� <*X��9��-���'԰rqiݼE�p�V�':�80@�f�)���*KIF���^x�"bj2l�4 ��f$r&2��a7
S���' q�O;� �6��4;��w��H�@P�
�'��� 1�|�IpF�lmH��U*�|�`���D���8(R�?�'zd����>X����i�bI�Y��'�*�ç�ܳ4J "$��Y���P!�<��<I�,
�* ���'�L�
'HʩC�Q���vĸ˓��E�6�4�&�u����LS
_"���TOO(T{S"Or���j�F���,�O��[��x�Iy��3�NA�n>��W�!��=���8KF����-��B�I5Ow�DB[�BRh߼Q������ Hi	R��O��Q��o�g�<>�,�Є	���P��˸{� B�	�e�üBn�qp�e_�����d)J6|�0�)��'7��d�뉥M�,Ys��1��4X��؁�"����q&�5Z��ȡ_{"X��43��t�5�W�z�D�r᧘�c� ��ʓ���@C��4���+��B\�4b��)��R++4��u�m�Oh
h#�)���L]���͎<��h�'cn˴�2����ϝ*f*�*4����0(�Q��� � �g~�Ĉ�k��UR��� LD������y�a�d�viI�܇S��z$E��-��B2`����|:	�S����-�(y S�V�S����'r�l8�R�x����|�q�?Y�q;b�:D��;��Z#J5`��pHN�s)�m��&9-��%)�'y��iłI���X�_1�C�I=2#���Wh
�_�|Q�"#C�gC\��oR�Nr�hr��9Z:C�ɏy� y	D�	<G@�T9�䈬Y\(C�	�)k����*��?��x�'��ygC�	:�J�"q#�+\�̰4o,A�B��:,"�8�aC�?%�$1�)L"m2DB�I�/�8��3cO>D��r�L=ɡ��_�q��`��b�nG
)�ƫ� �!�dM�Ob��"Ĥ4a��:t
�H�!��ǪMK
%j��B�7E^0i4�_0J5!�ȃQ�ZŪFAՎ`�D�h�*M�!�d׹Ld^܀s�}�a��d�!��r�@Ac��۶9��"����3�!�_�=�]��eUil8����9M�!�ݕ,�>ܩ��Ͱ`:Vt�2-�,k!�Ĝ�JA:1�FN�e.p �e��.�!��](`�P��d��2��Q�D
$6!�Go��cG�YL�*����:�!� �Ҩ�sG� V�D@�E��!��N�;�����Q�Z����2(̕a�!�6*��'��b�dy��)J>�!�$�8$�Ε�!��3�����'!�� fv(���ah��Q�O�9!��!4r������Ą��n6Jb!��>G@���d ���>��c��9p[!��ح=�(a�B	i��u�fi�
X!��C�:)�Ј|a0�	R����e"O�;���G�$��@� k��@0"Ov����.��a�(;�!��"O��!V�DkŞ����؎V2�"?��%^�d+�Ń�K������#�Ȧ�q3nE�l�(#F-;4�r�'D�� FĪ�`}(7�_1"^~]�"OB����$�t�`Ħ�L�.
P"Ou���>?����R����%"O�<�Wk�5��c]�@�
d��"O0�0DH�0<^��iDE&���"O�0�V�É2Lpi��g@��Dr"O�P�V���{eh�����<��"Oذ�l�?)bn!��Y'/�d� Q"Oz���◳�fX�����"Oj8 �!w�z��)r(!�"O�4�H��6>@�r��MVD@�"Op�¶��j��՛�P�Eʸ���"OR9Y��O?	� |�3*O-\莰��"Ot�a�IΆ+����)�+K�T�Y!"O��J"ᐩU��t�b�ɖ#>�8"O$h#Gۈ~�F$2�E�Z�����"O�aǎ�F
��$��F
��c"O@��łф+��$��������"O(�i��[�q�Z"��>3�
x��"O�)G�Z?�ls�Lҧ��Y"O�T9���Pz�$3EЫqل 7"O�a�A�tX*hJ \9 K"O�A1�Y�1��Q02퀧 9bX2�"O��Jv@�R�� Q �؈t.�`��"O��3���6R���b�^�9(uk�"OD��0�B�������yu|ܹ�"O�@	�h�Dl�B�%hshK�"O  ��ۗf\z� G��)]�Ԝ�#"O~8�2J�Fv�� #t2��7"O��N�{]b� Q� J�NM�"Op4s�D�N��8Q�FT���[�"O�)�Td�U�\2�j�#�,D�"O8d�!�#�ֹ�lV%��A��"O`�Y�@�:m2�5�CD��S�Dd!�"Oj��@z2��@�O2��L��"OA�� �^h	�%O�'n� �"Oؔ��;Z���fF�"kH��S"O���ևˁABr�Ӧ�ҪY`1"O�Hy�+X-�B	�J 6A���#"Oґ�! ��|���H	a$F@�"OB�X��܀(j����i	�h�*�z�"Ov�'�t�DQQ�n� �J��s"O�(�A�@9s���{�-� p�R4J3"O"�y��D�a���!�G:Y��u"O�y�Q�6y���A�ێO���SG"Orp(���:�Æ��9���J�"O�=pGb�H�8�3͐�W_B��G*O�t��G@c*��@���%�2e�'04�P��A7G���c#�<Uؤ��'k恓B�͉LbU;IX0Uᰙ��'��L)��]S�F�����JY�9�'�:��=$��E���#Z�bp0�'v�#�1��a獃(�기
�'T@��D
�:Y�0!�5J�p��A�	�'��S��ٕ��8	 �k=�m�	�'�~i�a�j� hq�X�4��[	�'��J�<`�d��6l��50�z�'����#W,D����v�M�<r8�:�'�����V
ߊ!wlՁ::l�'�|ԣ�@R.^w23���#/�2�
�'|���,�:���Q�R
�'�eW�nV�1`���8F�J�*�'�*L���tI|�YщE8��1��'E�<y"��<#�Ђ�j5����� �]+[�i"P��
� Q3�p�"O�lbA�A7?�4��5w1�T �"O�=�tB�Z�µH�I�;11ɣ"O���� �`�)��-W�5� "O���a���ey������'"O�%U�Q"/���B.J�����"O�!�m���t�)% ����1r�"O��J���'�^�zw>$����"O\�Pu�87#�4�-ɦ$u2Q"OB4Y��k���/.��"Ov-!�j�-7Z�H��L�>pZ�${�"O�AY��ȁ;d6쳒�$GpB�"O��	@�
]g��
ϒ#"O��۰�ݗ���#sH�;3����"O4m2W�ɍm���j�O�HF��8�"O��)��{� ��E��ps�"O�u���P)9�����$X9yh�٫�"O 
�#��b݋��C�hL��{�"O�A��N��S�4aT^թ�"ON�X��+S8v �oP
Q�}Z�"O�:7�K�@������ߴH����"O@�j/@ �`�4kW��]�d"OX��g"R�P8�y$���Pl�S"O��8A⑗L��Oʢ%�r�"Oة�r�M�`�,�$��/ ��b"O��׊��_�@�F��@����"O�p�7�Ñp.���C��Zl�a!"O��i�*:��"3e�)B�&���"Ov�sW��+<��⋃���"O� �B�@+M�V�y6C��h� R"O<��F[�~|�V �z#�l1#"O��b�B�nH(���@~���"Onl��l�E����ϝ'`|!"Oz4�J�ak �hϓ�v[�!j�"OR�2���	*��rFMGDu|��"O, s�h��
=�њ%f�>����"OD�dX�$��4�7VuF-��"O,$3�"_�+��Z�#���H�"O�X*�`#���BTʠQ��p!'"O�m+�Mݘ�V0yr�I 5I�m�"O�hIw)��.Il ��	t:6i˕"O���Ӏɏv�v@QP�U�^��=��"O�Y�4/I�:��pbP IY@��5"O2�j���3gk�I�8*���$"O܋cdٓw����u�W(pɪ����i ��	:� }�^�*Mv�
zT"���v�X�xc��q.�u0��0In*��a�N�@��#z�hm�ː�9H���>	׾i�,��	K�geD�� ��}`�(D�d�!�ߡ������&25$�ר�%\}�a��i��'��E�,O.� *6�91�$�	aob�B"O�ŎR�R`��mL�!l��S/��l�Ƒ�F��qX��bS <w������($d�U�U =\Ov5I�4�*\�'p�x�n��FJ2a�E�ߜH�Y�'�PMx����>�b�x���;By�I0�����0&n�G�4��<�T}�U ςI�M[����y%]�����3�4��F��U��KM�sđ>�%i��dm8~���T&�=�\��ȓ,TBkN�H� �Ef��mڙ(�(�Ory:EF~��ٶ�͍��4`�"O���iT�_<�9���T���b"O�ZuC
����)i��t��$��$x胏�) 7�Q)p
�-��D�t�	0n!��'5Y�\ �A*M"�It�G���	Vܓ�h��� ,h�ǌ0�~��*��\��Qz$"O�%��Y��pʲ�G�~Z��"O��BGH� )R��$�T�q� �I5"O����`��$����fH��v��e"O
(��\8*�^P��H]�u^��"Oj��wX�,��rV&[>z�U"O&t�U�C;�Z�u�pp�"O��ڴ��&��*�>vi�EzR"O�5�c�S!��Ы�B$H�V C"O�ZG�Nl��D�֨�5>e��"O�P�e,=���ڕ��5��"O����FsR��![�ҷ"O�tCDg,E�Ttst��E�}��"O�	s!�&G�"=���)c�j�"O�J���:9ґRtcT��萖"O�����i`(2��²V��MXA"O��p�,	�nٸ@bP&��E�"Ot�����D�V��!'�	��a�#"O�y
!,��%� ��G׶QA����"O�ᴋV�	��S2���C���y�"O@�Jr��#��"��?~��<��"O�QqiA�*��:��Y%T�HMT"O��5��1����$4x� ICA"O�,��a_�g��ѡ��S�\8"OZ�&��;)\	k1��W�zX:"O$)#��׻'`��r#o�Hx0t��"OT�B-�)%�$��t��2	\n�"O(�F*�4]"�)S�=k\n�Yw"O�`2�΁%v\����F�,ɥ"O*�����,�|b� L��6"O�1���:8�����O]�i�ȡ� "O��C�̗2q��U�7�*v�L�"O0)���D0�H��4+�hT"O���슶T����m")G�+6"O��s) 8![�]PdN�^+��1r"O���s��RO�@���O��e"1"OD5J�GT{�(p����)��2"ON����� 
�֤��-�'��1f"O´k&!3Z����l�
��0"Ov�5'�E�ny�ĪLT�)�"OB�{#LN�lh�SCILB#�!��"OT�1�OG ~�|����g)��(�"O\q�a5C�9�V�-�L�#"O8����B<AG̠�@-TQW��"O
��U%;i��[ヤz@�H�Q"O��h'�@�C�DB�g�9UÒd�"OLh@�G�F��:C):(ش�d"Otl�e�@8f�N,�4��j�4"O�8���D9�M��	%GlY;4"O"�
S��Wu���� �,���"O��nW�Nt���]
6/ԃT"O�D�
�q�l��B�W���"OFٻ��=�Ni��]�q�`�r"O��a�iޑa����R�R !>�!"O(�d!Ç�D5��j��
���"O�5�6�;- <�j�G��S.!�%"O�����a!�q2�߁F��"Oθ��+ �0�q���B��ȁ�"OLLd���{����9[�6� `"O� ��;"��f��Lq�=�"O��&F�%Q @M�DJ�[��X!�"Ol�`'̂
��(p��B
7��e"O�ժՄU�"C�5� d�V���Ã"OD�Q�L�RЄ��fi:2h8��"O� ���AM�;g��'�7=�*y�"O"����3��m�R'A	���Js"OԬz�֛r�>���6f,��h�"O\@��
�
  �fAT��'&�4���D'F9�R�H.Yg�@�'TH��p�O��zu�ǞNC�x��'b\2SR4)�Є��
�E8���
�'ӀKC�q�l��lG�<��m*	��� �U�u��`#����E	Ϙ��F"O�I����U��-���+% �jw"On��6�� D���	D̽��=²"O8X��NE������^g�*��"O��F¦>B& ���72� Yqc"O����mRd,� �E�i��E�"O�d�"z�:Y���#RX�Q"O���%(�#6��r$��7���y"O���ֺa�֨��b[-S���Ѐ"O4�0���[٘����]�l3�0�"ORyuOɟO!x�J��Q�)���"OP}�T����� h�!($XZ�"Ob�����9Z��q�G�z:`��5"O��s�Β	�0��Q�H�+M�yK�"O>ub7�B�j�.��lҴxE�D�a"OB��"�_J.�z�dK0���"O
�u✭�j�`u�˻5@bp��"O(��p��w#T�bCZ�#Tj���*O:pk�� *�Qadd+d���'�hSb���;9Z���㇢$�j�'��8��׎SPZH#���'H�h}2�'D�t�q�N�s��F:���'N^쉴�#-�"%vA
#u����'Lr :��Ƨ~��S�҃2Ht��'���$�:�0ԣ�/Jx��'���(��\�w����3N�	6�x��'�4��E=s�����.D��'5�	ƃ	7��2��@�Pv���
�'����+]�n��ALѴ4HB�9
�'!Ԭ��E8Y�&u�V�'��h��.ݑ\�t� F�!u��-��'^�$�$m
)fHA�0�g���i�'�m��&[7;�D���B�Z_� r�(EP�
n��-�GdӼH���cV�T�T�ȓL�~�p�%��J}>dS�8U��-�ȓV:�K ��6~�JIK5�W[����ȓ�j8�ݷ^���ӍX�:����?�>U��K�|B�8�# f�ҕ�ȓb�xT`^�-J��A�7�T�ȓzO�!Y�"�3q���ѦBf��ȇ�Q@<�s'th��rN�$�����es:9:ր�Q��ZTo�l��W�����H�`�
�qb��$�Іȓ�\�g<SH�&4�ި��D�8$B�L���"��ʉp�6��ȓT�5��(��]�2�!K�����QO ���.L�vݺ}Іh�?m��ȓK�
�%��9��h�'o�<}W8��ȓKs||AE'�oB��Aa��J!�)��?X})$
]�r������*��ȓN��m���XPP��HE�`��ȓml��05m/r�r�#��C�l ����m9� Ӥ�6sr�Ӂ�рD���|E."7
#+00|+���7x�y��e ���#Ԣrg%���h�jm�O�Z��_
e�T���'X�< �D��37G ZC��=�ti��`�~���4�F%��<�6 V��J���$I�����a0���cӠ��樑�I|-+Ri�`�y��H~)ϓb��f�7zA��M�9�<��dZ(6�h�G��+ޢ�k	��b��cՕ&[6b�m�Mn���O�d*��o��L	� �,Zj����K'@+������O��G�r���B���-�%ʒ����y��>��ˣ��z�aRI� �@��P��>,�щ0��$3��up���i���R�X%�yW��?��X��,���c�W6��?�v�3=*:@��a���x���d�b���������!#PXh�"!�{:��� �Г䙓F�(`�p�W P1���fJq� ��'[PX�̟�A2��G�/L�\B��&2����D~߬�RqĊ'�m*�Gf�U*�aظ&\�I�t�+6�'��%ɂN�.eHU�aF��2�$5����(�q�B��dH0��K,����3wJL��ѫ{�NC䉡u)"Uj�7u��C�I/q�p1"�GУS��Y�A�1���"�*�#p!��N̹���V�S��.\(u�����O�;�0�'#�aBD9S�l)`D�,̸�#B�Z�`��)b0H���� !��[fIء'M*i����)Ķ��?��2��l�3.Y�5���bf
�b�'Mʄ1$wƨ��U�ֲP���S��8X�8`�)�7	���郧Q��Z�!Eʀr�T\��IY_���$��fa2>|�'R��/�(�E��	���Ot��5�ݪ��x���D �V��)[�ޭ�Ǫ�GP�H�'`a��@BΦ$k-Q��_
/WD`��p2)ISH��=�Vt�"#}���4x���O4��A�\&-��(0�o��v��#X~�A�R�ɀ�j)@��2�������+ �5J����ak���c�5:9X����
���9�^���D��Wx"��"G8�Y�L�c����������1J�
"����� -��@+��N?���bhɬ>	���'�������BHn�i�Ɩ�9m���{��c3�X�P�Z��&��M<������ &E�@�#d�d�x��f�I�6l��$0�vMї�Ҍ1|\R�*.ACujc���!��~2h��"�,���<�v�ѣ"B?	ħ�R ��"���2N%�c E[��򤐷^�2�`0o�h�����
g�}��	�@ٮ��Q	�ɘ�8h�Ÿ&�قuA�J�i�<	{pGL6��0K`�I�]o����'v�t��O�� ��֟�pk�mչHv��H��xH��qtˊ5#�L���猑=�R���	E��O�У��4�vQ�Vě.���b$Fm�y�0#�*Zu�J˫ D���&;@�0a�ԅ/��3�ċ*/N 5�'���BV1��_\�}��d�|�� ���4�6���LF���KFC3/Þ^^�u����y��������T��a��I�/S�(�J�
_2��q�k����'�~e�D'�Y��!0&�Գ�j�i�N�A_�Y٤T+8I41:m�b��jE�IJ���$�#r�l�q&,�#EW�e�d���=C>):'�îK2�T9?�~�iW!øL���s�8�ɦXHԑ`�,����呥����7͉�#�[@�">�؄�I�p�lC����V�n�BANb��ZWH��g��H*헾"07�S��&L��O�����<-P�q����9T豹��B;9A����Tqg����e��)h(��c��	>(X�i�&:S�ėsx�C��+8u��NB�?��Y6"��%� qp�P%]�"�nڹ*�J�$V#$v4���':n��q�ؙiW �{r�E�5x�C�)֖���;!ծQ�	�"3z�����ڦ!ZW�۷$�.B��L����� ��iG4 L4�P�.N)s }ذb�5u�IGz�Z%Z�G�<�, ;�Dƨv�>�ʧOZ�{���pa_�tJb��{��A����!ׄ��w�>�ڗ/&|�����Ol��Qmϴ/]�T��$�rƍ�c�?���P}�ÛoR�d�%	�=5��K5��7<�ɱ+�o�L��P�)a$H�c��8�ʬ�������b�B>B@������ J(b!@�s�Q?�󕉌�{�I*��7Mȁo_�^�����_�dgp�30���ཫ5��=x�eJf�G�>Y��ϟ9]�̜�C��0H����+�*1�Ȼ�≻9����O�Y���'G̓��^�D���eH$Gβ50'��6P�$��d�-�h*4�� txY�qeO8L�L�ҁȤFͰ1G�V�]��dO�/�Hj���(up�s`/��^=��e�	<�@h�"���4��-Oj��a����� ���\��۷�ͬ&�6d+#�8BH:�P��ӹ{���"��µ4n8��B�C5&���M�.#�*Hk�&C;CD(�0�O�љ ៚`����d���B�e�_���9�	L� �8���m>��р�d�����
G�Q��ޜ�ls�C�e*���͛�o�Y@b4!5 �Ƃ	�Q۸�ψ�&��'�q��#�A X�v|j]2I���;�(�c_��$p�����N=7��$s&�¦ѐ$n��d�2��W�q�I����l�iBH�0HRTd:U�q�qO0�:`�i�$+/>�r�K:pp��g偃`� #&%O�m�Ha�+}^P� 1d_��(��ex��G���a�0v�i�p��馵�r�	�|��"������-{P�)��K �Hq��D�.2ܩ��tS�$���-c�.U#�$�Kf��!��C�;��b��S7@�}�䦋6�*l����/g����'6^Ҽ�g!K�M���m��ys�bG�� 8�g`T�xyv|���޴'`<���B�McO�ި�vD��]H�/ �"��̨pKI�uf�*L�I���JgY���(9W��/��ֺ
�(����8�
�<�֯��O$�Y�KN�l2��vb��?�T������ ӈm)�ȆO��K4�q���h,���n��D�fED��P��#�Z�%,�褮��jSH���ž<A�aE|r�����{���8,t���'K%�,��ЈZntX���X{����ý7��(`��$z��g�'�"�S#j�W|�{|"�s���k�0�3�@9/�@�Fx�_	_��l�'�ޟ=ޜu�eןD욷'S�'�ԸQT�=!a�v�C�h�(��A��P)�c�P%j�Z�8�"����?$A�։�F�z����2:,B�ԎZ��T�ʢ�A �C��w�Z���߉B��$�Ӻ#���9V1|�'"ѯ.� 
t���vE�$��J��š\�[B(Y���N�!�$a�O��E���P�ba�T�K����"��=��i�-�!l���H7�ߟ�KP.݅V���O�
sn���bW� ��i��#h�xg�ڟ.�r�Y@F�(c��Q����p�0�HV� on�ZƎ�X�,�E{�4��Ň�;��C�I���e ��Lw޹�#�<G��h
�އ��\���\)E3��[�h	'��QxP�vąJ�'I��;ԥ� �T+p����Y��=#�����H
�G�-�f��~J�ĝ?@sl���@*p��5�B��Vt:�������"w��*x i)ŧ�sr�ñ�'��=�GSTq0����g��d��%@j|q�._�4�W�B����IQ�YѼ��W�ǲLqZwW�P"��6j��-��,q�,�]:C��3���r�t�jgEZG�k��Z29JT�3��'W�@T@�:3@��#T>c���A��?c_��P�I3<�8$��Jɟ�+��ʊ��!�㭃Ѧ���ܝ~ǰPi!B�4ar�UR�U=��)����h � �*Ȏ��J�<f����6ԉ��8ړc:�ыRd���x��4H��)p���:Jm� �«� ��X�o߃>ƨ�����*��$HQkO�H��9@�Í�Lb��"�K�?	����F_
U��&ڨ=J���`EE|�'TR�;犑�BWI��FZh?���޹P��� � ���Ђ�(�B��dnh�Nx����S�#���H��Y���G�i;zu�Sd2����T�\"��QNN+Fe����fh��&+����т��Bϲ<��N���0wG���<"v%�s9�|��T�wz@��BK�30���Y��0"��@Bb�)�L(;S�'J>e sBH�&!L��2��2���A��ӆ��	�]&��`I=5*n�@�=4c@��L�)�#Yf'��q��\��v�	0�i't0�`���7gL��%��G��r�Η�����EvDh��"�!v`�Rǋ��u7F�q4�D6+�O��6��A��z�F\��Tŉ(&���R�!��|0�!DHN��bb�)�x�J���CH̸!�Ⱥ��K��M�'�C:a���9�*�F�zBь4�0��*�v�U	cJ1}"C�1�)�6��LqX��7I3�01�0n�Dq�D'@4^R#�u�v$���u�L�@R4N?�y���k�VQ�� խUK\�s�B�~Vt��Dg�'T�r��T:"Z:���喃F�Y�7@�/":�A�BK��v�9wo�^.��Abc�A#��l.6���%��8NbpYR��n�*�߉�H�.���K�$ȉ"$!�@�+����'CHIP	��BJ�H���{@�hb�œ�]j ��WJ�@�G��ur �s3�FP}�+�$�!{fU	�Q;3�|4AE��G�8�����O�����$�R�Y�gQz`\�:�jN��	��&vYෆT.2��ĠaO��!�F�B'Ѕ}l@�*��i2�Q�bA&��,H�¨∖�,޼Q�ZܴTPcju��-"���(�x
���L�|Pi��A�x�2�
%A�>�𔪇v��%*�AI�)�`J4�J�h`��I3sS�8 ��))`�郯˭�0<���#�Pd�K�yW~az�Y��ݩ&�NҼ�tl֕%+��A�j�l�����2�ĂS;R	���)	خ.@L�5Y�h�nW��fxh!�8�@e�O������%zԱ�
�H��:��
g6K�G�*Hb��I�O�=�j|�T)N�~ ��(F@�,��C	�H��л�`Ѝ$�r�)t�2�	�A;��G��#��uU#>���;��y�2Ab�-ܕTm�$�c��?a��5�w뒤'��U9%��;���c�(�~�,EnZ8*�&�A�LY{IjbТ��=�Eh��Vʖc�@x�R�TϜQ���V`�'W0�Y�̯O�XX�F�D̔д`�?�4�j�V��0��J*��'q-*��GdO|j��o��"nJ�7]<!;��:M�(���A-`�(B�S�!����S�Ĩ�M͂�:֎#Hr�yF��*1{J�V¡j��,*F.)tpֈZ#�=h�F�T�E��eSU��Ta���wM�@�F�a��]�T���I�~���6�	- �KA.��	6 J��  H��X�>B��߉>�@t+��̎�$��'}���3�Ac� ���k܏?��s��*Fx �A�kш����#I93Y��"�� �e���"sb��[ը9�`i���2���ac��O�0u��'��)8�^�5Qv0�$KR#�l�;s����挖@,yЂ��9�.�z�,]��Uj���B�(�Bʮb�J��\�GY�I�)���b1+�4w�EA���w���.[�F�Jf��*D`V�ˣ�I�u��| F�E.bk��rtF�:;���JW�L��?Y���@oH���))p��d8��D,fTF4��Q8:������nT��`�]�Wޅ%��X{���՟��W�E��p"/��A��C�Gle�2ŏ$#��a0F�c��ɑ/*]�D2r�[m��yv����H�B��1qd-�3���`lO�xi �$�%V�ι�RO"�z�+5�*h�F��\++�B M��P��6��H�P�3�%�E��hWJVS�j������}��؉v#ȫZ%��7"Ҳ2�b���h	l=������|/8C#j~����'�����LL*[a�R	�z~A���\�h8��/�������t��-;���%@Ker���k�9e���C��}^X�TFǌ'MV��G탗SO�Q�A�@�w�X�y�4t)-O�E[ AI��a�@�U�h�t�Ӄ
G���� A�_��"��T�c�*��֏
x��I��b�@=J�Fɣon�Б�A7_��J�!g�<Za�׍D��↓M � ����v@(���=,h,�@A�V'B���Gs|ZwL08�CU�P}H(��A��\��1�Ҹ0���2&C�/c�(�P��*T�c��)c4��"(�>x$���E�5���Z��K-f�&�p��3+Z��ɇ��ՙ��WQ�������%j\nt���tqy�+�LrL�e������ O֔P������G%mQdh0�+�7Ip C�B�#�&�S���|��`�d��!2*pKC�&P��w	��H|�qN�c��S�i�<�ЁjŐMn�4��f�*9�dhݚ�L�fH�Dz =6HM�ر�q*E�Nl�44� `�,%�d��Cq��o�< ��mϢH�m�����p��&l�i��ʓ~/����JZ�ϲ]�ӈ�����oT�RЖM�o�{̱8�'ޡ1����FY��!AP���@z�5B��1�|X�Oy���H�?DmX�q&�ڌ��'�K����*Wc�a$�y�႐p���K�*t8�UP6"Y�?��/G&���ݏ`��X��G@�ղ�D0F�k��̲=��!�����)�3F 
u!��Iv��4n ��f�8h�8�b�g8[w�(�y n�:��dT/��	�� ?%�0AT��OB��"˟�%��s�i��x*�!�)1Rt�#B��?DwT0y�
�?]�1L%\�.ݹ�nV�m���B�*ۧ�b|�%��~�t囶�_-B��Y�a����d4g�z9B�m��f>8��'�E�48$i�t��D �N ��M�hC�0��u�Q��X0���?qy0Ȓ�]��᠈܀ ��L��Bo=B�¬��\hJ��A*��N#6���Y��O���,J) ���E�*�\M�O�>��p/ɻ2ؼ��)S1~��h�� ٪����!+;�4�g���j����3���C�R�{��X�q���#�E�q���	^j@�!�,���D�����K��,��'��!�:���S�Ff�:��a�iD`,h:Q�ݏa�8��LZv<	y'���t�X)B�i����ŧ�q/�q3���f�,(�V��M���C.Λ֮Îf̠q�B�	�6Ҍq�/�~"��)H���1&�2�~�z���2b�(Y�R��	f�(����$X� ����w�י8b�%c��"k�� 2O�8~on��[^@����1�\�7\������]H��;4X��䚄�h�i�,R+H��c��ոXB�Q8p͗�p�6���Lݱ�?�'�`�QG�)M��1[���:U��t�D��9����n�/J*�X	K3�������6�R�(�l֝iq�F�x���H����0&�+��Y7��uJ���+f�A�bJY�q�^�(KȘ���&_�-��qK�=�6���C
N���V�4�3P�'�jQ)��!~Yd%�O����֩�2Y
J%��K�p��Yz��Rct`�^
b�Z.�(j�R|�D���h�.s���09:}��D�nū�D�)-���)�\ĦO&��+.2��X��EyB�
�Li��~r��[92l�4>�މ��,$-��уÀ�J.����Mݩ���bښX�'�
��ť�F�n�PjM,N�V}b�Q�Y9��rC 3<�i�a����0�"9HcC�(�l�(ŦO�s����+WS���&iSo�*��'1���LM e�l��ނrT�2#?}�IV�� Pp�Ǽy���A3��L�d�C`�J  \�� ���� /u���eg���Vp+�
Op�A��R�TLj@�/M�p�C����pe
���4��'�\q�a�QҘ��d`
HY��Vt�da#�C�!�dK g��Pd�g�����mZ�M��j��� My0��[n�az�#�*#선��CI��aȀ�p=��P3tY R��iR��"aV-F����@H�4��"�+D��B�"	70�|�I��]�qN�@`�f&��>���Ѫ��&��HG�n+w0ZD��k�~|뵪͒�y�O�?*�IJ��U�i��HB�^ D�����NX�u�Z�'��>�I"/<��1o�/
�)�B�F.lJB�ɱi��1�@ �=h�*��>����  ��P�'�r3ԭA�{��UI���־�y��50�zA��=�"�x��ȩ�yB%ʶBW�mc!`.3@���kA��yB�J.>�B�r`��7�B؁�$ڋ�yF���Ȫ�(S�<�X���,R��y"�\�_����I�7"��w���yB�aE���Ǉ�2�> �&^��y�F\6HR��eb6vƔ��,R9�yRnDi�8��C>(1�����yR��jPA h�3(hJ�H���y�#S�Iz�	k�N�Uv�i�i��yr�߬+����H���dYw.S��y�����X��6K�-�zW���yB��~�h��k�:� Y�d��y҂û#�8TsF�� 6�!�eG^��y���&'��M��B�*r�E�e͍��yB�B�{2\�QM��-�1h�HH�y�+W%"U���R�ĥ/"^Q��oY(�y�ʃ
G_"UNZy۰�M�y���(���PB $0��٪�y��ߐ7ɨ�NP��4�K
��y�*�9�	i�d�+3�j �i�>�ybgMw��=I�!R�!9v���I��y���$Tr>�j�&��!�>]s����y�.��P(�8�rꋿ"M��CR����yb�I�&��|Qta%I�L�ys,��yb� S�:���W7tax}�S��8�y���\>�8�ɜb�	�agҟ�yr��=���ՄY�\>��#�H.�y��G,��P�b�ӕ^y�4B�M���y�/2n�`E*`�&ِDS�ܦ�y¥Y�8�R	X�	ג�����y���+l�#�(�� ���yr��:X��K�O�RΥ�
S�y���~���g�1}t"䍂��y��еO�+�&�X�%�(���yҩV*/���E�ޮ]�9)EFn�<	GH)���"�Z"β��7��F�<��%^��<9�U����SG B�<���ߏJY�0%�_x̘�z�i_P�<1Gg�99,��)Sg=toJ�R/F�<����#m�V��1�baZC��D�<r ���Q��9\�qrLTF�<�6͞
�^�s�f�0�A���Qu�<��J�:y@ ��,�3!�<�`��[�<qt��d3��N.|�բ$�L�<�eK�.�؅� �C�#���*�*�L�<m�d���oI�v�~͐�a��<����iC�?a�t�S7z@a�u��r�S�ԵH9RB��-~q�A�@�&4� ��g��7l��'����~�M�b$��8P���{r�/raY�d�N����sj[���<Q�$��O���	�_Tx�QF$�Jm���p�Zy����M�j@iB��ns~m��Ɋ 0� S �>S�С�Q�<J�'��['È�y���XaBĦe�*ѻw6�`����� ���Ra޶>���-8KCP"O��S�I���j�{G�\�<A�!s�Ú�D�6aq�iֺs,�]���_�A?���?������f�p�!n Ib�ח?u��e�Ǔ6�0��$��o*�8�C̤_��Yy���	�x��S%	e1�Hn�*�:l!"�-1t��rG�J�й��҈��b�p�p0'G���da ��O�9�"� 4�<��NRd� j��5�@DGW,j�^l�0���%���� �E~f咦��F���8���HN�!!(�. ����>�P�N�Bd�P�-ɒO�p����&���HD�V�ې���矂|Xs��{C<����KɆ�"f"O�$�X �숱�EH�N���� %y��(���mW��ɤjб*�88��?]�rdO�S��e��w�\yp֏�r��ЫA-Z�M�ZY��
���@,�2�l`Ks	 ��IW���g>�өF52�.z��@qx��"�AB4�zH�"�	�zLP���C�
��-H�`L25�V"?q� � za���0d��YՂ?# �s���!l�݋'}:qj�b2"p&�Xb� �R�xG$|9�K�	\vay KEO�Z}�%�Q����Y)�d�t�Z�?�����.���b
�H����Cȏ�z�B��Ʋx������8$�N)� �½:�d��%�tjY8���I��[��2s�1WA�Uc���A�J�vD��3�`8;���7��H"Ʌ�fG��"C��0UB��'L&Fcr�V�t>���[�T��,���h��i�-&���Ai�<����'{����N~�'_Bl���;�����<}���!�:/=��K;xK���� ������Ѹ�����Ğ��~��]��Ν��%�5'�6:fg�e�
��E���AK����aur�=��IP19����'*(PpŎ����P:c�tKF��^���a@ 0��S�藱fW����a��WH]1E���"�.}E���Ag� S#��,&gH�Y@�1�$˓c���	e��(e�2��d�>��*�	�Sc�zf��~�s�Z8����@&4��-˳��U�@��"5Oh-؄F5bt�x����(B�$�Ia�ys�'Mf�j�P�Є1ŪY"?���z�-��X���35�͙Q��-�ë�)D�*�$>1S�V��a���2w����b�
5��@u�V�Q~|̩�n��) ����URf%RE�������9@>X�rC��$|�� �E�%���鴮I5-4� r��	(N�hRL�M�x��cˀ%fā��č'�����	�.<��˗�0��i����Pm����a8z��-�@���⟘�S|��x��B�s�5��Pkd�S�.C�#��X� �%���`u��=B� ����!
�Q���O�Rmv�#t�B�%��p)� \��Q	��%G@|�cሒ!��<��b���ا%IE&S62�Pȉ,v$A"D�\@J�㒊rO��u'	e��)�nN�P� 7��Rr�L��f[ ��؈��	v+��1�i4�x���<��jaޟ� ����=i��S�L�ٖ��u㌲>$�\�3f?a�̴��I�_7����?l��k޴7;��a+��dy\,���"a*�H�d��2G�$T��0]j�	"�rӔ��0�ɕa���pf�|�>�Bo�iB�aZ��M�F�ٖ ^(���ۥ"�� YA��j�I��o�j�޴Qf��`�m	7�0֝5��L"�%��h���A��+�V��J��$Q�Ɇ�
��HOBՈ0+A~�P�1�A�jyi�C�Q�F�JQ:y*��V�q1ҩհ���b�3E�`aAǃ/Q�@-��P�~%�=���r��`�!^T$� �A�B4��?�qF� �pII�`�G��`VC��|q"�V�&���U�?~ I" ��X��X+ ��X_�1��g$^���uK�7�Չ��<x.U`%΍Y���'^�D���"��f�Z?���ץ�MZ��⎃ks�|�e<yU�`�t�A�z.�$��片X:��ۧe�p�,���K�4,��spOk���K�/B\� �	z>,D��l^x��O.L����zbT{eg�cV��%��:2NPa�k�7R}=I��_�^ᦩ#�`��HkUQcQ�5ѕ.��4ZpY���5Vu�E�Ȕ��J�'Æ�W�Ca4��k�j�8I�bp)O���*3���0c��Q���<r�HIrA��?Z��a�،X�$X���E$)^��Ce�@͚��C7?�FhB8:T��!���Y�6|��OhP	�ȅ+�nUga �@�ÀF�Q�T�R���r�b�*D�>	fpAU���`A0a���Z8�c�ǔT�@A�d�ԃ	̖ #�&s
j'DՖImXؠ��2l&-�� �w@V�'q�\akW���aI��J0�R)?{��Õ6wq�BVD]�L4���gP
X9DM;ǧ@ꦭ�� H�Rq�<�Kfޝ.]i�	�HóQJ��Dޣ49J�:�{2�њ��O$^xBϐ��F=
�S
i+�����Թ ����#ғ`� ����y�V����Y
m3"9�LSh*��؇i8�����c�07M�mQ`��_�+�q8��f���+�l��NѴ<��F��5P��`J�<Ƞ����
���� ���-7�b%�p�E�S���Ѭ�#!�2����F�qU�����8�'��l��L+fh�l�"K 2$���S�-�0%j7�I
GR�$�T�C0|�$�BHR u���l��D�hhv��% Q
IT����,	ԩP`.<�P@�78z���g�/�t@�à
@x�'JpX!C�5Y �	%/���#EC�;h��h�����Y�	!?V<�æ��59��;��^�-��9��E�8n��(c�?��Q����Lܒ4af$E^]��SuOK
 ����͉�e@X����;�r��u	��X����"I�5���q��8?ɰY��d:/���i3kO�ⴳSL�zGڜ�R�4���+��9ưm�gT���� �	US(`�d�ju&T2�>�*C�;�����t�`i�.����?�	��6����o��@�8#Ҍ �TR�Y��oAI�|!�	���IU�������o׳E�sB��VQ��*�C12�"\��3L��Y�E�c�4cjC'%'@%���՟֝<�ƀ���ɈR�$��7������@L%u&8@�(/N7����KG*��X"��õ�bc�f��l�v#0H��D�^�0�"�@�6Vp;d�Ș0��$��)whzá�@䊰a3���\�<���� %0FP{��I2�,��j�-�$���cä6�&�A&�?	�)�B��93&PB�."ړ	i�U�B/CgǶ��RfʽQ6�0�P9g� E�(>/j��+U ��e�k�NR7<��ɻ"�
�Q<�&��b�6M���Z��?YԪJ�V  Pb�M��Dz���W�RB�'�lLr0�T6�Z0�D�ۑv���D���q���-"�3&B�Y4)��Ô;2��țR�K�c#�*a���4R�sS�L��?)ި\>=�CT;3���-{O�$�Ug��;�V�S���1|*Ԛ��ΐYx���jĿg+�����5�Ӥ�B%���~�V�	�o��c��!���H��U�ԅ��E^�-Ib*U��,�xW�݃2� ��3�)� ����D!n�����%3^z�s�E�OL�f̏�W{�P"�EvӾx �	Bێ�)�*��Nm���@�����`EÔ@b k���%u�v���	_ dy�$�1�XF{r	]9k��+�/��&��E��& ����´9`p#�+�~\�=@RB	|&`�� �G�,ѧX�$&�Ġ� ô>	|T{T�'e�]�#��%s��k�Ԕd��3����;ac�}ң�&u��{�'����� *5� �R9%��!p&#��ɚX�B!H8�r��f0�����/8n�'vC*��d5́��Y ,<"b,O 7������5(���� "��R��˸���a�N?!��P�RR�5l��f\:vL�fs�� .]�>�	*��C��F�2苺��Eɓ��O0�#��.����PΝ�=�2�`=���4A�1SD��FgX>&�P��>��B��^7?��1U
� R���yӐ�Ö'�>%�X��� �E�6�w��9s��fY��i��S��g߸Re�{�hY��`-�;�hQ�#���/f��P��0��m�u�o}�I	' �ؠls#	�6\#�a�v��p�<��MK�2��M��]֦��R����.��"��)Z3��
��3V��4�p�	f
UH1�>��,��8�2LaPGцN	��S���4Db!�SC�w}�䠟;�?y���8;fu1�7O��3B%��2Hv��� ~ e�FDB���oy�-8F1�@nL�dM4�b]���k M[dFE�y#d�f�X;|��fWWZt���2gl�7G�mZ��:��-�\�b��L�.�d0�֥�2��Cp��9�+T�X��I�¢&m#^�\�2�z�OC�(]c!B#<Wր��R�R�>D1a�R�%D(�Å_�@+���b�J�X���sg����
a`&�E@@�'�_�'
��w��1���i����jT� <w|ޡ#�iٜ0Nؠ+�58��K�睺4���)1�D��t\��4x�:M�7�q.�58���<Q�҆}&����I�J����.%Q���@Ľx((Sj	=��M
��ءOD��g"@�1����Sn��Q���$�E�{/J�
�8��yr���%˚��B?��U[aI[�(I�Ę	�Ա�@Ԭ�%�V� �P�� �ְ��lֽ@��E@5�L�
d$6��7����稘>����M�G; �!��X.~��ɓO�"�AET�x�d�"7+λ+T�'�Z͢NW�r\�*b�م0���҂��\�p����#��m𥈙�!�p8dJ�QpdÅ˘�X��M���O�E�&a��eƴX���u�D�,Y��",%i�D��b L�1�l_(f�}����l-,B��_�s���
���l�X�&"âA�`���i�7�_D(�4�� ;�m(�-�_�X��1$� M�1OZ��q���O����n0�S D���`�&�s��`���7jD�h4��͟Kg�b��	CfU�@����k��Ԁ��7�t,�w䇅[�j09D�2a��jw-�&G6VX���A��4+��� w����~ʂ,�:r��As�i�h���Kל?2�A�GN�@� %��Dȗ�f��_�M�6h���0�2W.8|lг@�O�i�(
���(�D��ʱ��.�m�,P�q��Ֆ5�~�8.��a�`�+p�N�{�VyqcnG�,����8��ɓ
|7pdJV��{�l֤�!{�.���CF�`�f��W��$eE�<�Gi҉���ҁKτ1��S&�.����1T�e�ʗ��\��o»���1%^�S�l��j̄j�,�?b|�t�W�U�/W.�3�Z��6����H#dR��2�Y;O
%��O��z��zv��������q"�h���TA��|�w�I�F+!$J"K��%�_ J�I�!�3A�<.���KߠJ�u��0O� �ďށ1��)��^5L+���	PJHQ�b��	��Q*����s_�@���C#�p��Nܥ�?��	QI \a��M�
��]
�H�0vV������IR�$\0w�fA���M�0���G�eJ�%;��W'Q�z�t*
u�a�1u�j]RE���?ёb׎ u��k��'8����?`GN>S.Y�3�~u��u�ǋY2���U�L�� �*��Y%~���cE#q�2��䂆5|�q��C�J4Wn�dF6DS�3�͑����r�"�yUzШ�'�ܱ[@͞&[�΁0sꞰj$���*���q�eꝊ6��5Ӷ�i�̅A�m��X�ȑ#jޱl+��
����Qr�	HuTT�S�����8�eC�!�F��$���Č���KU�R����?i�eܪ��F��";��c��h!b����(:i2� �Y<a|0�V"V�-뮁��F
$2��{�fo,v�BN�<>��o.H�IQS�	U�ӛ3Fn<	 FC�{��(e�u�f�L����&@5BEx�(Ig�t��b�s
Rf*%� պC͐7X/�e�QG!d�(|,�8�]�E"�~1��C�$�"ݢ-���l��Mh�t��CH )E(I��)M�|��̇�:�
�R�a�%N��x"e�Ll�l���@(F*A�4���PO����ңl���Q 靠4�$�I��=-�&�&	� ��)rI� f���R.2?AԦR6���7�ݦ �c3�O2j.u���[�������5F�h�58�����9 �S�O3i e�����̘�1A�<����/y�, %s��]��(�h˴�W��<�G_�+��6k���O�q �MX5t�8A����Q6|iQd˒�^Z<\[WR��(#�@�2)��4w�:7m���pĪBHW'`��d�6�ݥS؝X�̺�6��@�e)R�; %�Q�֘��+X_J�ӺkW�ջ3�d`��* ���hUo r/��abf�4E��c�Wa6�C��'l0d3��G:D!�&º0���!��F��:4#�ֺ����4;~��e�!�Hp�����������e\r�Dn��	�	��M�ƬK5G ��BMT�.(51���hʾ�ɖ=���"��+7VQZ�`�		�|��@k]3.	�"�a'0�Ȱ�V���1�'�>0 )�[��Q�5�ޝt�PI櫏�H���8���mZ�(�lѡ�I�u�$�C�<8=����m���A�B;7x��s���a�1a�'�%���d�:f��ѡf�~�T�'���L�0�����fR	Y��S�49ܸ��/�'�4y7`R,NP�1��ƨj���A��v(墄%�1I�d��Fo��.�� �,O\�	�TL�*i����J9A�X�4��=����m
Ŧ�уd�Ij�������Ӝ!c�i��Td�U�F��f[V��E̠P�`P��zo���TD.kT���'���G��?NcN��6�rH1�ɟ�m2C�w�R��v��ZI�A	B OgX\BB�Obt@��J�NQ�B�3+JXi��R�����Ѥ1(&7=�\���ջEl�2�ќ;C��*씬|�T�����))��H,�\���,zy���� �P4Kջ�1�j�YB�� 8n�:�����h��'!
� ��+AY�4��QbB@ɂ{2z�r$%�.��3��-!�p�Q���$g��ԥC8<��:�O�\~r鋇r}>l�]w9�,�}g-��! H��cJ�U7>���*�s�*���,9�@h�c���a�mӫ%h���U9$ũ@
ҼS���Q!���%�2aCQ�ȟty0� �sH�KB�>�~:r�N䨘k�Ԙ4��P��ur�=`2B���T����/�|MiW��%%^�+!�T�6���OL�p���N�!Ql� F�j�B2��2w� )�O^�ȥ$@��~B���*Z�J/'n�π �y��"ad��3��k���g�d.�r���:��4���\x�Q���	,���2 Kٌ�3󆕥'۞�X�`�`��5�*5�.O�.��!j�h�^|�e�|rVxi O> �%)	�W�P�'�p?�r�Mp�
�+��6A�ř`�*�l�$<��a�<+Z8�a�n�zg���(�29��w��\�&F#��4c	>b�<�	�'U,���ƈ"Y�ƌˣZ3��1���d��L�:?o��9���֘����b�g~�*�D�@J$腡tڈ8�E��y"��V����)ڐ�GC�p���=Q~�١�0=vE�W����
S�

���w���ҤEŭ�Lq��l^%���͚���1��]wY��"O�`�5��7�����	X )S>�j'�dJN���֥rޢ|�T�w��鉕��`E��)��Q~�<1D���874)X��<b���d���e���$�N�XG��'��!�J�Xp��✠#/�P��'r�d��h�0h�qzG��'u\�M��'��QS��{������/
TU�Ӥ�Dev�ؕ!D�l,��9��#�!^�d�B蘳;�!��͉V�6�ۃ�%l>�t�1�!�Du�(02����6<0P􊎪y!�D��'���y�ქ3�(3���xR!���0D�9lN=`rh��*Y(P1!�d	���M��Þ.F��жJʔ?$!�A��H ��w?	�@ۖ�!��DXN���HH�d9�Qhb�$$�!�$�-j�ިq���d��(ElC�E�!�PRT�s��B3��a1���5�!�,_D�j�/}�V�놆�:�!��2 £��D��WdѺ.�!�] �:�ï���!���]�!򄇴/�*����5mM}���"O}��؝R�2������u"OJ���O�N�ʠ
gн: ��G"Ob����;��`� č��"OV���E�|;G#��O���"O�l�`AҮ?�(��A�o�Q��"O,�لbQ�,�8h%?�N��!"O@��Z��trao�g��9��"OZq�&��*�"�yС� %�pс"Ou���0��`K��P&9�Be��"ORAs��#;L���AX2P���J"O�x`�s�"�OÐ}��g�'��KAD�,bH��Kկ�~� kŬJ/�u��ą1N�Ɣ�3��*_>q�L�M͈T�o�9d��]�3Mn[��s�p��GFZ>�0���G�3�W�Oβ��@'?�w�O.x��a+�	�N>U!���J8�|D"șP'BA8d�f������A%��e4?�~:D���܊�a�&�	Xl�ٶ"�;@��=a0�D�q���Ӯ}���y��ƙ8�0�9��Q 4rV�O2��<q��3M��i`���k��I0�gL=��1��:O�,�<���[c���0� c��XQ�F�"&:�Ӻ#EAZ���c>��#!�\h�ah� �j���*A
@9�ɕ�?�$ ����\ib�p!X� �Q�!i���M>	�4�0|�p�N+���B�%�`�>�Pĉq�I-`�<�XԩXq���OԺu�@&,i,}���Hb`$��-O���?)�'g�]�>)�e�$XF�8�OҔ~'X\�pIFYdI�u��OD$`�Fg�_~2��1G��8�T�0Ud"�I�5N���?CM p��E�3bR�5�4'��^�1O�1�$�d�S�'}Wb�Id.޳qg�q���Iu����'���낣%�)§r�z��BˁQ2XLi�^5	� �.�5�%�)�'dVͲ�E�)�\�q��2]%d�o�*Y֠� $� K2L���uw�O��9P�
:\����H�T�%-�����Hy"j:�&|�t@�-�������%�I�r�i����R�� �O�?�;�燡5���`C��R�4(`��S=s{�I����g>�C �x����6�V-M�
�G�>Q���0�"��ȟ �iԝ KZ<����f�����j��D	Rr9{�" ٟx��g�? �����*#� y��nX.:��,���Iέ:�(p��	�UR����O>@���֑P3��:F�G	>��'�D��Qj�?t�`��$��)=� ���'�j�RP�ڜYN�a��ޯ.ŉ�'�J�@�/�d��to~��'}2h�'М+@�m�aǄ�|�́�'�"h�����Mzʘ���{2��a�'���I���RB�� �\nE���'{28qP�V��HY@�J��*!+�' 6Ձ��ֺU�����10��
�'b"\�p��.�҆&ۛ�v|2	�'0�k���{j�pӊ 8	Ӑ-!	�'�z��e
3zBL���{5��Z�'��Ag@�K�@�+�  h����'����2�Ɩ0pPX ��0�4���'��P��*E;#�R�h��8#���'�48�R��z:���l��b��T
	�'͔����ܑ�b� ��
��Y�'�2E�`ս8\��D��*h 
�'����ɉ�]+.��``z��%D��b�"�%7��@lE.S�@���%D�DS���^��l@��C�E���{�)/D��k��!f��AL����%��i.D�HӲ���^4]��342����*D�L9��^�1���r�F2^���5D���D���^�J1#gi��x��`Rb	5D�䢁���%��p�B�s5��Q��3D�`�pe�S��Uaj�E�h�a��2D����  }������&�`K�b0D����-ɂ �����o�"�9D�@�(��Z��iZƤ��d����4D����)]jv�㐏ِO�p���5D�Di�c([��`kT�hy�렡.D�ȲA돾">X�%��&�na�e?D�@"�K$Y�(��GF�&�p�8�a=D�D0�=�p�x����u�1�;D�<�t#�"gK�e�l�n�&q��&8D�T2�H�'�꼨$�D�{a�H�G0D����f��`UFκ�0JA-0D�d�4�.T}��b�L:qϊٱb)D��I�g�*n7$���ɶ�@�TM+D�qS���Il!҆���6� 6D�0+�F�4h��pz&����RF&3D�\�e&6�cψ�1�Ԃ��5D�p2�ʷ	�*)b�ɓ�Jp�`�'2T��pvW��,��N	5��0u"Oę��d`��+�K�"k8� �"O�m@�eH~��A�jc ��8�"Oyr�o]�VmAwC�e�T�a"O��R��^�[X�a�"�*���"O��Ch��g�(�(#!���%����y/�\S��+�|x�S@H �y�Ƌ�4Z��e�()'`�a�=�y��T�DQk��W���RU��yr�.h� ܂L���BP��y��)���`��B/��ڕÀ�y�L �F!��d ���A(d�`��w�L1�-D	v��0$>�x�ȓL1�ըc�ڜ{i��kC�`���ȓ'Dt5��=��=*0/\2O\��D��d�Ђ����� O��uN�t�ȓy͎(A��ŋ�����H$����(���F�m����ۻ�<<�ȓg�b���*Ӎ"Pb�C���v�����S�? |u�q�U�q���	��̀�$"O�2cX��P1,��Ҹ��"O&��cP��hMu+��i%(kG"O���h�q@��(��T"O� N��l�A��wK�( �"O4P*vGG�r ��, f�L��b"Onu@!&��-�ra٤�V>d�V�ٴ"O�u�͈R��!���G¨���"O%H6�W�5MJpp&�� �dr"OJ%���� $j�8�I��&���"O�8����-er�h���P��X"O��hq�*~�ۢ��[��)[P"O��3lô�9[AIߐ��Q"O�Dc�k�7`�R��5H��(րxx�"OVdpTޢV��:A�&d�2"O�P!�N#B��*��?�]��"Ov�k�����<}'�:5"O*�X��$Y�:�ÏhXk�"O�IBW�52�%��'Z���"O~<�u�W� �2�kҶ�$���"O
�z��,1~�lP��Rd�0W"OT��7��"�i[�\CT"O��h��SM�vH1��:���2c"Or�㡆F��I���	^<!�G"OH�{v��&.� �@\���r "O6�	��	&�NmZGS�*�ŀq"O���E ��]SqD�0_4�m�1"O�,0��Q�;���ren<����"O�$Y�MG�4���m&W�lc"O�5�En� �+-S=�ah�"Ov��UJ� �O���p3#E?/!�Άu6��%S<:,�ba�Y�!�E<���s�hG�~*N�x��!��ɏz�̽��l��F|�+��;v!��ʟb��[�g�0��)��	X�d�!��/=Y��Rw�i#��"�\'�Py��'f�����A�#$��ShP�y"� &M�욇�x�lIq�\��y���<e�HmS�On*�0"�@;�y`^k����[�Z6a��H֬�y2�@<9��K�}gb�A�!@"�y"JC 7 h�Q6�J�b1 ���4�y���p_���ƋH@�D��@"�yr������=H�t:,Ҏ�y�B�>@Y�G�:�@SuD��yBH*%~�#��N�2��M���(�y�$؉8��ۖ���ܱ��.���ybꅤy����ʺ|�I����y���2�x�#���_�4sU��yb��q�@X9�F�*PZ�Dr"�Z*�y2��/6�(ᒅ��L��*���u�<ᢡ�(~.
�U�#�z�(u�L�<�'얇f]���Є޶=G8EH��p�<�$�I�wjp0��:Y�Є�gWT�<I�dQ�C�ɣ���-W�����L�<W�״�V�* �G�+����I�<���Q�{_¹1tFE�[�
09��D�<Q�!Y�([� 1�F�hW�p���
I�<�3Ǆ�q��i�ua�@�P颴��D�<�)^n���u↖V�"�E�F�<Ѷ�D�-�i�@	�:||�!`�K�<��H
��F�9a�T �6=��n�n�<!��?K��ъ)�*|�d��P�<9�̀9L�pu� (�<R}�0	BL\d�<� 0ܒ�jJ!	8�yI?��9�G"O�X ��Z.g9��y!��-t��  �"ONܘ�鎩~�\�8�/a����"O~:�"��j�&YIǌxN�T��"O�|P.كdv��f꒰8I�j�"Oz�"��<���0��	�FP2���"Oj�8M��M�ല��Yz��k�"O`���^�h�P��"����s"O�Y)���Q~��	�].���qe"Of����&|�~d�Qi�?m���"O�Q'�M�7x��;ph@= Ʈ��W"O:0+���N�4�Ӳf�9!���"O�P��� 8�U"reGT�+�"OfP����֍�i�ka���"O��s�*~`��n[.b>�I�"O��6a̶P��T@�lO�},%�5"Oj=8P�Z

֠ �5�1H �3"O����x�-�!����B�"OXhW)�
����#	���Y�"O��2�)Ƚ⦄����H�L���"O��v*ɖq���b�Q�9�<l0"OƸ���p�����-.��a�"O
 ��	���D��#eZ�Q���[�"OT�2���/g���A�Ǎ�<�R�"O�QkEd�!p���b!�L�<��"O�:�CFw�(`G!Wrݨ$"O���&,ֲp���=id���"O�����Gn�,��d��{���"O���Wž�`)D�L���52"OB���@Q>HlĊ)͢)ǌ(��"OT�2�$i0�Q�+M7eϊ�K�"O����A�;����)��(Ȥ@k�"O&D���Մ4>^)��O2W�M��"O�pb΄�6Y��c���C�qS"OZ��jc�����ϝFgX���"O�]Cu�
�#I8�Y�`I�w��D"O0�@��@$E��pt)-8�h���"O�i��ES�<L�mՠk�H�a�"O��aC��7�NpAҢ=5֬� E"O�m��f��uJ7���6���z�"O�`��א'vP�B"�$�h�Ѳ"O�0�s`~���C�K{�P�"O�P�³G��R�ѓ��<'&!�շ!Z�����̙Y� ��=!�D.
g�"`ӡC�d�����x�!�$N�+!��(�هzp�]��M9�!򤓙 �<�������>=x&+��!��O�h���!7�Վ'2ࢩR�x�!��B�lr\��D܈V)�)V璳h�!�D�uKY��〨4��a8�.W�!���|�K!�	�Ŭ�7�*[{!�$��b�����3t�@U��'��D!��@f��[7HW%%�f���F��!򄍅Yl��D@�M��XS�	/�!�֠�2"�֖hd�³��c�!�DR�J��YHƊ�5H�|�cA�W�!����B�` �X��rx��oP�4�!��_$1�H��G����n)K�!�DY�:#lm��Ǝ:n��hydM��!�Dۏjr�*S����ˈ�?!�D$z�͒4ϐ14<�8��i��`!��	�5N�hwC�#u.ǈ%�!�DT G��ّp*˿B"�@	�M«l�!�υ0-���홨b~t�Xp�8Z�!��  Cb�߮dXHt`�力#�H`1�"O��ɝ?.��z�/ܽbf�Ж"O^�pW�_5M��)���%h��`r�"Of�:A�DG��@t-���a�a"Ox�Y��['F���*g���x�"O���g�ǂ}&|���+e{,�D"O�x�   �   .   Ĵ���	��Z(3VɆ	>_�����@}"�ײK*<ac�ʄ��	ڤ�Z�x��	?	n6�΅9� �r�j�0k́#�I
EG���K)v���F ��-!H�=�u�Ŕ�QpYom(|���������m���+D� 6F��:�f^�7(0�[� ���w��U�H�بBR9t`гp�SHxv�8��R>dT<D�W�]�4��	�Mq�A��)i��ʓ1V�k���=�h%�'@��fFĚ\K��j�͟�]��if��?O%N���x�(Q
k�h�R3���ğ�/j�[�
R�9(�iM G���Ө�e�b�z� �)��9��ɀ��tHb����'t�pǋҿ2�`��R �w�Q6��OrAB��	��P�Op8+'��tR�'^dЙBGN%؎$�F_%�l����(v
Tj�,�OJ�I�d�$X�b�|ΓI{���3�����i�#��5x�L��
d����<���r�8�EFayRgF�7]�1#pH��p�E�e+�N��ʠm̖11"��O�(�v��?HX�d�<��<!fA��7�ᢋ2;H���Η _���JK�\�!����8��'}���`Hy}�he>)��B�5�m�L�\80��U;NRh����d�>���Hv�|���p���L��ӳ@�')�
�H���"^L5K�8	�L�P��>���OJu��ǆ��i���p�A6%cJ��2�ҏaa|�� B�),�Rԑ �,$��	(o6�j�fIT�Ƀ'&�BD���? `�%Re��!�P�x |�P�<1�HY�E���	�B�N�ɏ�r������(��pب�	���D"�xҀ��fx4�N�7������F�K_�=QeF+y��PP���{�f���EE<_�����N�A[::��ƪI����E�oZ�A�i�P�On���qM´
�"�F- ��Vr�1Rb�P�5�$�%V?�@��%�¨��O�%{�-a�E�7m��'����ͱ�'{�H[Ɠ�8���aTޚ'�&�7/Go!��L� �  ��-��!ӂv!�$O'��=`g�o���G�^(i!�dY;*�� ��,�U�r���'��!�dE;�r�!��tzܒ¦Y�]r!�d�+>��ex�g��{��4��DڍCw!�D�NV6�x��X�B�d���2U�!�d�!Fpj8�i�(l�>}�`,2�!��
L��� o��N��hx���" $!�DO=@���n�b�bӴ��!�ċ�2�hxtk�&��   G  -  �  B   �+  87  �B  LM  dV  /c  �l  �r  by  �  ��  8�  {�  ��  �  E�  ��  ͱ  �  S�  ��  ��  �  ��  ��  �  ��  ��  ��  � x C 6 x# �) �+  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!����s�\bV��^� �Z1/O:"�]9�.?D���dd�R����7�˟&�������<IE�)§0n�a���5�F�p��9 @����I��E0HSgjMC�p�X�E�|�A�p�.}��'���D̎g:�Y)0��;j�^�."�S����[�c��=X�M%R��჌R�<W�񤒇?�X�G���iW�%�6yZ��I]؟���Z:* Т��ݞ2429�2�:LO.�0�]���+�//2Yu��P�!�<���,Q�}��J�!�dF4x����)hp��y��F�R��Є��4M�TeS�%�i��8RHH�FNC�I�L�!��F{��¯n�z�ȓ+~���j�}3��{�mǋ�X�'�ў��B��`X2�9��Ԭ勰�	$�y�L�(�ޝlQ�{�IA�I	��?�,Od�O?�h��Χ(
n�o����H""u�<	V�Л:!����OVXB�`�UR}�H�a�Z�<��@Λu�m9-��'� �ԉ%�IC�'��I��qQ����
�u!�o��!�C�IB��3cT�=,4X���"ړ�0|RB�A�(��3@��+֤� 
�C�<��)ݔ z�����T�[A��2�JX?�M��O�>�f�ϛ7M��b�]�$�E���5D�P���+L�m�L��X��`3D�ܺT�u�q3��S��|��4D���@��
t�`�e�4C¬��D?�O��'z-PT�M�����,�R��?�S��MKgLh��IT�R�X|�g�:�hOD��)I:+�!�O��w��%����-AZ�Gz��9O��KU�A%M>����
���DR��E{��� 2���̚{���,K/��4�iz��̞L��xb�.P�k=���CCW���)�"%?i���2�I~�� �T�ի Ԍs�+_�2F2B��-Xo�
eg�!����� d�����9��mg�q1c(P�(!���J��y�C�K|��f�:{����@�U	6LC��J=R�y5/��m��P�h��5�T�I��HO?�g�ҽָ��3�Ԙf'25Q��#D�dʆ�@�Ld�(��!=`$E#��/�O&M��-�ae�4��K���-���'��	#�R@�cDG/P��[e@��kC�I?D"D5H#��'�������"?1"=�'��	�K��"A,MA���l����<���q�ʝ�L�R���E�1��h�'zў"|z%��5�F�Q,R�]��	!��}�<y��5Uiz�ђ �&�t�aAzܓ��=a"M�
e����Px���x�<A�ԋS HI �U8T�0���x�<aG�3�x��-Y�>�B��r�s�'51Orc>Y��͙5 ����E�̐Q�`QG�5D�0���k1f�#� ����[�+ D�\0����k.q���J�NJiTh1D� �G�ӧԹ�ң�6�LE (���>��3�L�Z��?�R�iP/���C�5��RR�	�@�9Q���m���$\F�$�n�|�؇b$a�XMA�-P�ў���Ӏg��u�,�v��ڕ&�5�@#<A�n0��,{n!e/�Y�0�B�n�ʵ*�"Oz|�֧��PMУȋ���%����6�HO?�$J HI 	Ѣ�ڢh[N$I�Á�k�!��̌n��m�
;OF٘������Iux��#w�+�ҩ�&�࠱H��3D���`�W�{�ʨ��H1+
�(�/D��y�A��-��h�%A	^T�4kb+D�p1G+��y�H\�fˉ�2�Z  &f*��p<�Vb�r^lEq�Gb��m���V�<��	�lJ.xheEM�r�M�vf��<у�'��iq��	h���S$�J��X	���M�p�s�dχ`��T��b�@�*����>1���AT���s�I�x=괣Z�<f��=h\�T�E��q�VU�'���G�Ԉ��`JH�da���e@3�HO����(?z"���U O֍��%�?!�Ā0C�l��ŌJ7�$	eD݂A��IF���;��Q�v�� �]�.#fh��e<� ��17�`�B`�,Hp�u�A�ݼC�	���驕���R �*�!8�C�	��aP� �fT�C��	v+�O����d�]��G�?9������.��G{���'b, �-��sHִ ��׊N>B�:�O�����=�\����jM�9�rH�-l�!?YۓC��ӆ��*)��x�uoڥ["��ȓ>�Z	�7�A*�HH�̓!��}�ȓ~��|���B� p�0d��C� ,F}��i��>�fO�hj�j�h�L&�̒eOː�M[����bep�n9(�7��%��
�O�c��O�$$Jr^)[@�=��`(	!.����_S�<ѐE���<��2!#+U^�"�(�O쓅��N�O9&%j���n
�,��-�	�jk	�'� ���T�4��e�	�f��I<�	�B)�	ŨT	4�����W!.��ȓW�,b7��.T������4� �����d+�~&��2/RK����d[�kft�R�
n�<�����>j��L�q��q�Z�CW�%^��~`a}
� p!��( �+jRQ{��@=l8˰�'QԬ�?	�GX�~��n�_4De�rJ�[�<�sEL0����+�0W��#A���7�(�L 0��5+B�@y��>~ƺu�U�'�Q���&뉄=��i%��H^-(�A#t%<���I�3�2���R)2F��;��  k�bB�	�L>xa���b�)ȋz|Epش]����=�B��>`,�x9��WQ�T���h�Io�'a�m�	r�$8H/��+T�F�:��4�3�K��!�G#|�TX"���2�%�,�$�!��͓6���c���R~�\�'��T���2O&���K�dQ�����V!S�v���Oޣ=E���ԃ{#.���~�)d�G�y��Ӹ5q�)zE�s���P
Y���	OX�H��ʩ ���a��κu�" ��D4�O���JB}������hH�)�xC�ɾN�J9�!Gy>Xpѩ�&B�ZC�ɖ�0��HŻ[�NЙ��L��P�ȓgĔ(VoD>/:Ԁ@�C�E/6цȓrPz@Xt�nŀF	I�-��)��k����D.$THR��7p=@���A���2 ��)��ܫ!��0f�(5��l���蚸zD*؋���Sxl��u�~�Q���e�U*V��-E}��Ӝm4ebe�W�lY����D��hB�	)
�B�`f�]�@Z���'	1E*��hO�>�b�MRP��|�0ĳR�*D��;��ː']���# �a3�(D� @��$s��-�aY�c!�4��`9D��L����  &4nh�i2D���&�X9V&�Ykc,��&���cJ,D�T�AŖ!J����!U���{�+%D��v�S�'�6�����vz)(%`$D�<�!�W�M�S`�+u�FY���'D��k��X$p5*�j�' `��9D��rPh��&�xp��iB7��]JdG6D���#] V	�E96�ߚ1>`0��5D�4i�锡��D��N�<N l=�i0D��+bm��(��EJ#l�W�|p�֡+D�����ɧnR�C���e� m	�&+D�(H�UG���#�8��Y�")D��A�F<Z��4O�2�t�J�.1D��0��
%�L�i��T�}Pjmq��0D�|z�hl�����рA�XQ�q0D��l��~��0@`[E��/D�L�(�
\�(A���<�-�k.D� p7�
�wn�c!)p��h�@?D��+�&�4������=ڬ�Dn<D��y�c����;�NE
^�xKE8D�p�W�Ͷf.*�[1��#A�d�
 7D��i��Q %��5��+Y�����5D�\{�@ףH�<0*��КC��Q��b2D��qo��9ph��e�'e���S�$2D������m��p���ٻo߬���1D�4��f_0Q�)G$�.���U�.D�0��M1�ur�Թ7&L
u�,D�����^�����ŗ5lx�[�d.D��Ȗ�A�"�p�i���8�I"@9D�@�"]�\� �z4dZ�2E����7D�ī�*�#�\M�D%�t��,S�(4D�t��&Q��th�@Ź.���!�0D���DJ%o&l���nD(�L9��,D��#&��w��z�IB�I�j֡(D�d�aJ:%X�� �I<
{���O&D�� RE�%�F%<��y�r�M<}��!"O���t��*~�,��X�d�H��"O��	����tLjG�ӫ��3�"O�A`bH/E����#��Y����"O&�
SG�b	���C��W��U*2�'��'��'"�'���'���'>���Fӻu^P9`UM�.��`�3�'br�'�b�'q"�'&�'�"�'	fQ��b��Cj�� KZ�G���p�' b�'���'�2�'"�'���'-���4-�d����#��<K�\���'��'�b�'�2�'�2�'���'�4uy��Ǚw��]B!�((܉��'~b�'�2�'���'���'/��'r0Pj�o���I�4��BQ�'�r�'���'F��'�2�'�R�'�̍�iĥJ��ㅮDÒ(x�'�B�'�"�'���'0r�'r�'�nЉ2c�'�v,X�M�j�+C�'G"�'�B�'���'���'4r�'s�-�Cg��w���ka��O 
�2�'��'4��'L��'���'�"e���`(3��`��i1
�2X���'��'a�'��'��'�B �<T���#D+K��e�Gb^2#[��'���'!��'�"�'!��'QrɎ��e��$�~��8d~y����?���?i��?���?���?���h�Td@q�z+
\�-�.g�%B���?I��?Y���?���?��i��'�XM(�@� d#]�a� �S��<������t�4 X�%dg�6->MuE� &ؐ̓���r~B�mӚ��s���ڴe���m\�hP(�0G��;w�iG�ib2K.5~���� �6�K*,����~:��� *��RW(OS%�����F̓�?�+O��}�Ç�Ǣ�2�hcX�n��$L��؊ژ'y�,hoz�a� 	N�G��MpT.��t����&�M+�i�>�|J�
��M[�' ڈ�W��yF\J�
�Y�Ь�'/h�s E�xZ�T���i>�I?E�v��S,N��!�r��f��qy��|r�u�q���D�=c���2�� =�p�Y$�	����Y�O�l�Mk�')�	�<]��{#��M�4� �Ǔ'U�`�*�$TJTL�>����|��� �uW��O���c��"*�j�(4�/;��1tM�<�-O���s�H� �D�B���j�ǚ#r\�:�~�d�ݴGMP�'�L6+�i>9�7��gkRt{�����m3s�y��{޴�V�'֕T�i��ɟ/��r���|���Q`f1l�H�)��8�`YÒ��_��gy���y�fI�.1�	�AH%)H��FL���ąܦe A�G۟��	ϟ`�:҅(��ÊNG��V&ω8f����MsB�i��O������5&�d��L�,I4��Ô7-b�JF��S���BN\�0�j&��=�M>9)O��`�oZ�D`��+0v���'��7m<N���$ެv�J�Q�N]�PJe��(*����֦��?A1V��ܴ[��Ov�*�⣤��YV�R���*�`�N�9E��51O�dʡY���"csV�ʓ����#�>�Q�@�f@�(#p��5ϓ�?���?!���?y���'�?���0{��X�嘢K:�<	��ճW�����?a��i�|@[��'�¯k�L�O���a�!~0*���*;����{Au*�ئe�ɫ]1<�l�<i��?���asb�-p��O��+��4�b��w)�9S`T*����"��(�l�SpN�93N0-:���� %j#<Y�i�tH��'�b�'�哩c���;!��!b8�L�CL��h�X��I �M3�i�LO��{�I[���,66~<
�*Iܔp���0�HZ3F�qy�OU�8�����na��K+0�'W W�ȰS��=8��b�#�2���
6/P�m���.l!�`ˣR
C�xВA�++PP#U%�v�Q��2�ȸE�D�yS�!�J� 
ȉ�Q�jfZ�
3��>-�MaE�����05(INB��A6e�	O��ɀ��M��dAegr��P�X���p�*Lb^���`�{�xE���q��p��.3,!y��Y�hG-�	�&)��As@�A��E(6҅>��=2��ɋi<Q�W
UX%̽!��м�X�J�> A�v�0<_�@��%�5[� ��?���?L>����?yŤ�[1K�gҠv����MԊ`c&��F*�L~B�'�R�'h��'w�ٹ1�'�H}��VP���i )
r}��-}ӈ�d�O��D#�D�O��d�4�LX 3�i�6Jp��,+����(�!�}K�O��$�O����O���?��ʧ�~҃�;�"M��M�^Q��b��6�M�����?�?�1�&��n�I�r�r��F�~�%�`o[��47�O���O����D�*�'�?���:'�; �r��R��`��*܌s��'�"�'�Ji�������i:E5�Q8 ��U�ڄ�PC:���X�y��ԟ ������?͕�5F�ğG2Jx0�MF�SvFA��E��M����?)�g�+����O�������:Y1�![E�pqٴ4����?����?��'���O�����!��� �mO
D�X	 6�`��Ulڇ����?E�t�'�fL2 !
��HdkU��3�Y���P�D�O`�4AW˓�?����?A�'��h��^��R�se�݁Gl���}o�%x��'���'�b�ѭc�P�9D�LiD5!֏�p7m�O�\�TH�<���?�����+�����!4�D���o}�K )'�'���'"V�p"��6��E�k�2AM>�Q��j� �'�"�'�2�|2�'��i;� ��z���yX�hg�.'�$}��ՠ���?)��?q(O$��3�?!�A�
��a  '��`�3GuӨ�d�O���>�D�O���];Cm��Ƀ���B�O�/Tҥ�T�	{�r��?9��?�,O�9�4�|�����X�E����g�4+7���M#���䓖?)��	r�2�{"��Zg���,���o�Ms��?)*O�E3 �|
���?A�'f����qE�Q����#ǒ+EP W�x�'V�D��<�O��
��k�(� B��3bA,/��7��<��ؚG��'��'��td�>��0��`���lR���-À_L�o������6�pi�?Q��D%R#T�ͣ������;�'^(�M���$�?����?!����,O���Ox���@�v;�l����Q�H�F���d�T�S�O(��O(��0��A2��x�P�<�7��O<�d�O��
R��<����?a���~�
�/r�`���`�9�i�f�(�MN>1DK�(T �O��'���aQ��� ��#7���cDMEj6��O� ҳ��<��?�����r"��2�����8�||��jVK}��h��'�R�'��S��Q&�J2�$�҃���x�*,L��hI<���?�����O��Ӭm�x!b/M+P�t��M�`X�7��O��O����O���t�u<��Т�K2eՎJ��B��Z�P�I��,��UyR�'���ޟ��"�O�+�2L�"�7r�S��ٲ���O2���O��"ꁡ���J�0a�ū`��F���c-�#�l6�O(�ľ<�����)�O�˧�����Ys�  � �����D�i��'��*8���O|�����1sΒ@�`-Y�a��
1YӸ�lRy��'W��'gb����5�� o��)�P,ݎt����E�>�M�)Oe���Z��q����D�z��' �3#+�"��4�&K�^�,��4�?1���?��r��yRS>7MFQ�� b�	ύ��ReJ��`V���#J�2�'�R�'��D_��Q���s$	��a%@�0�
�B,��]�����9�S�O�$� �C�#ZQRlS:�DER��z� ��O���3&���S�ě>A�J�2,������%��tj�+S�pX����'2�d�� =�k�_�4*����X�v�'j��cR��b���� �qB��q�Tl�4��{��ђlY��ē���<)�����O�4� o��,���`�7{����Cw!�N�<I��?ُ��'��ĉ�z^2���@hۖ�P���m��� �9��'��S�D���[�h�'uJN]�C�������oZ�8�IO���?�)O�8�P�i����Vc�U�	� L�!2��O<������O�s�o�|���=�pL�4�����RMz��gIi���d�O��-��H&�x06�*�t�%N�KN���Lm���d�<��[�i�*�����O��������_��zY+�b�D�����xB�'��ɣ1�#<��]�8�#��́Q��mx�c�2�nZGy�f�:.7��h���'��$�2?qp���j�t`�Ẁ+5��\����1��Ο�Iן$�L|Γ��iǖي0+ݑ
C�A�C��;%t���4 a�ԓe�i��'�B�OZ*O�V�o�@��w��-G����Xo��n�ȟl�	���IQyRW>�OzH�����8����%��5���u r���O��dȏ]��S�$�>��� �4�1C�@� `��([��yFx�.���OP���O�i�����U ��L�6�3h�֦m�I�2צ�xL<�'�?����$)g�ީ�W%|�n�Q�0	E��l�{y��'[�i>e�IwyR�'���q�	�U؄��P�uy��sF,I��	ğ��IM���?��'�"�1��V,<��&X�i�x�p�4߅�|~��'u2�'{�I�Q?@dk�O[���A�C�:p8V��#^��c�O���O�Ľ<)��?�r+ӛ�?�2�ʧ]�d����(K6y����w��'��'��I PBD�BJ|µ�D��v̓q���9<��{�jɢ'�&�'0"W�8��؟���l�ן����qC�K��u�Mr�!�7�,�3C�i!��'o�	4J��M|R����X'����]�|D|��R�D$���o�Qy��'&�c�=;i����5�^k�h�Q��͵I���*��@?�M���?	3�O����'[��'��$�O����b�.�A���=�7AP�1E���?����3�?a��?!-�$�O�&�h���
s������@��L��4R�P%AT�i�"�'[�Op��'�"�'�x�6�*"Z�ƩǼ(}m��e�&�2�b�<�+O��Sܟ�;cB�EV�x(1�&�1�����MS��?��Nd����'���'y���u獌�6�d·.��q#G��M3���D8��?��ʟl�ɨ��ʠ�P�Jb�ը ��;@�L��4�?I��f���'���'��͢~��'h���D] ~f"@E>x����OzՈ�?O����O����O.��OL�i�L�ReR�f�,�S3BH�U�0������E�	��,�I��8��>��?!�K 7�0Q�IO�M�1j��I�y���ϓ�?����?A��?q,�¬�n�覽�ŀ�l��\�b����BJ]�M����?a���?������Ol�b8�X`�#
�4����ԱB��@�%����	��l�	͟ ������s 	����̚�O^& ��`U'X�D5���M���?����$�O�l9�3�Z����� f�hSJ�3]I=��iZ7;:V��!�iQ��'Xr�'��E�Q�t�v��O������2�-I5*�x�'(��9�����B�Ʀ!�	ny��'�8��O��]��s�`(�7^\.9X7�N(B=Ѥ�i���'fpQʲoeӼ���Oh�D�����O��G�3j�I�Q �%Hx���N�U}B�'���9��'TU��So�	ޮ3���hçR�"���x�����4uF\����i*B�'%��OG���'���'_:U8B(U�fɒԹ4 �(F{ t#4ef�,���O�$�<�'��'�?��j=!���D$��>(@�!��'�&�'�R�'�Ҽ�эd�����O��D�O����>U��%�m��m� /Α��,p�ir�]��b�$k��'�?i���?����c����U�I�y�h��s�ެ����'i<�j��|���$�O���O6��O&��M��ӧ��w�1�ßG��	�T���<��̟������O�.T�3F[�.m��e_�/�~��u��5��7-�OT���O��dQv�TU��ɔ�֨	n��>��9鶇B�L!h��e�H��ӟ���ϟ`��d���C]�\7mM�5ζ�1"��IZ�Y�T���,��m������P��ԟD�'������4�#o�����Jb��5���?����?a��?!��A"E��'B�гs�B-��w����+Q�3��6m�OR�d�O���?)p.�|
J�0`R��=�j�@�^?�e�e�b���d�O����Ov8s�����I��t���?U!֤A�i�q9�D�3I�*TXS�M��M������O���S7�B��<��u�dB��+�.�S�48���@�z�N���O����٦]�	˟����?1����dӡ���q�����(�����������O��2f��OƒO��,���T�&�R3�QPk.=�b�A��M�$��:i���'G��'M��H�>y*OX��d��}�` q/�VOL��4�D⦹��x���	ɟ��	V�'�?����
�Ah��Z�y��ys��fs��'e"�'��p�Q�>i+O��Ĥ�<J�����%㜔[k�5����=I=���|� ʜ�yʟ���Od��1�@��@R�6�*|��J
�"��lZȟQ��V;���<9�����Ok���6��9T�l��My�e�#W����E���	JyB�'�r�')�I6j��=*�$�3�� 7O��,Td*����ĥ<������O��$�Or�)�@��^��-��8Y�ؘ�g�&��ΟT�	��H�Iy����3;��ӱr�Ԅ�&��Cp�s1�T6&��6��<����O��d�O����0O���ƌ{vxaf���;����R}��'�B�'��	8d�M|Cּ MB��e�����IX<��4�?�I>q���?��Ȗ��?�H����؞OV�%�eV����i���D�O&�ø�E���'����=:�D�Yu���TO"��cDN�V~O����ONИ�6O��O�������ȴ5����1�n6M�<�tEBOÛ&�~����2��i�*P�g��TM�x��XDGc�R���O��ɣ6O��O��T�0�!�"AE���S?z��Hy��i?,���h����O��d��H%������R�	�+ɕ�t�8"I�ZW���4v#l԰����S�O�#H;_�D�	ǉ!RzD����q97��O:���OH��/X`��ԟ�It?�D�&��"����C\c�ަy$�D��(�;�ħ�?9��?���-6غ�x`AYq섡H�ʛ�?y���*���x��'R��|Zc�<�aM����1�S�K�V��O��`':OP��?�����)�B4�p�?ip�RI%R�Z�*"�_uĉ'�B�'��'�R�']�y���2P�����^�ƽ��d���y�_�T��Ɵ��	~yr���1� �j�:U��;5$m�D�,[Ѿ��?)����?!�T_̨���A�ح�A�W�(�0T��� qk����V�\�	ݟH�	WyR�@�$���r9�lה;�Z(�옷�*yI`�[��i�	O����l��2(��	d����.���Ĵ�H4S��F,���'��P�h�FɊ0��'�?��'�쌲c��1}����^3LHP�x"�'!��vtb�|��Z5�u *0��h���W�4Ta��i��ɛ/�)ݴX���؟l� ��d� U*�vNN
x�>�����'����s��|�����(#�@�PvO��[V[���@�MSb� Bɛ��'��'���F9�4�.YT�@�`����J�A�"$*/����H����'P�#}����0,ZE̐���k�D�p���i���'����YI��',�Sʟd��;�p�����&�Y�tA4�
�W���&>!�I۟H�INN���U�Z �i�&l�/�f��ܴ�?	�L^2ډ���'2R�>�,J��� ҆�c�Tp9�I�_}bF�,��'��'S��'�Rf��E�pT�'A�
�`!�c:B=(8��_����̟p��z��̟t�	.C2H���ǋ6�vĈ�R�&�`�r@�B;V���?Q���?q)O�H��BH�|
��|YC�kA�	B}��'���|��'���'��D�xmp%�k]�K�4�%�U�q�����t��ꟈ�'��Ȉ�)�I^����3�r���ʗ,t�X�o�� &������[B?��6�dC��-k��ণS�8�7��O�D�<�bb �5��O9��O�d�EM�Q'V���]�5��0�'1�$�OH��]�[���8��R�
�Nl�Q����f��n�ty�jAK��6-O`�4�'����,?�1��EbbR1@[�N��� �,�Ǧ��	��r�<�S�g�? (-���!�l�˗��3H��;��i�n|�'�'���'�R�O�D-�&����EKĿ_� |Y�i�4c6M�"W��t ��ʟ�j'��>a�A��敉|v��KP�İ�M����?��^������xr�'���Oα���A�\]����MKLMZ���D1P�1O��$�O �Ď�;��HK�d��o�jĪ���[�jnܟ\
` R3�ē�?������[3�<������V�<�,����g}¡����'�2�'�"�'\��� �8�Y"��;jޭ�T���>���s�����OX���O�|�Oc��d�W����Z���q;t��AҸp������������	Ο��ޟ�����M��BZ�r]��
�*��	�]�qo�ğ,�	͟��I����'5r����D���P8������ F�*�ArH7M�O<���O��D�Ov���h�dXlZğ$�	�g�� w��$���@��߸�rܴ�?����?I+O����1b��-}��d�^�X3��>x�NTK�B�M���?���?��=<ʛ��'���'�(Y{��a�.��jK�t�s���]�d7�O*��?y� ����D�<��Šv�u�h�5nʀ~��q�tӬ���O� 
.�ݦ)��ן����?����P`�qn�Bc$��%�R��HF�����O�h�E�O̓O�I(��k�[n�h8���W��Rd��M;ֆq;ě��'rb�'�T�OHB�'/"��*"�L�����%J$��M|u�6�X4���D�Ov��|JO~b�U& r$�&*ܔ{ֆG�y�؅���i�B�'�r�>��6m�Od���O����O뮎-�����2��B�H�	^y�
���4�P���O����/�,��Ѕ%t<�BԯW�r��m�ǟPa�
��M���?����?�CZ?E� jFT�!�;_�>���l9?���'*J �'��'R�'�X>����*NeT�����R�T�Im|`j�j�b���?y���?�Y?��'^b�4�t��i�^�ZL�U@(�қ'���'(����#1ɤy�vU'a�Lj(��l��(x]0�n��f�dl�.P64C��f��ȂO�
�xU��.�#b���j7��C�p��nA�z�h��P�|G2q�t�4p�^��5,߄_\��p���tva�.S��=�M=����GF�[c�Ӷ*Ҟk40t�`��4iL�[�g�4g�t8�ƅ�'f( kpE�� ������� n@`��1F�j4�t���ܘ>����<8 �h��W��d$��,`��E��E�ח\yl$�g�'�C%~����tJ�\Ȕ�0���O�^��IM�h��I1B!�A6�0��M���q����b����1`0J�d�O�ٻ��Q
��P��;X�mN�Z���O�d8ڧ�?��+�Zz��0�LN�!��/��x����$
b����]�0<���I;q�dA�� TY$�}Y������ߴ�?����?��E��dG<����?����?i��fX�1�O+��5�՞$*�U��K�"��a#F�a��	Q�Q1xdb>�$��sH	r20M�ŊP~F��+;�<��׀mޠ��d���Z�&�>�'������Kvl�u�R?x�`=!�� �����GVΟ�>˓�?a�*��E�x�g&�!"|NU�����xR
WO0L �r��:hL@Te9���@����<����e�}��&��F� Iad�w�йQ6���?���?��g��N�O.�Dm>�[�a�5ps 8���k��A�^��8�b4�
��� 5g#��<I�.��sE�,X�F��-�Z���*����Z���6O:L�!)���ay�H�a�d�'쒘e��0�m� !�z ��!����q�V��a��DŃe�T��AN���8\aF��2�y2Q D~�����Su�1�����'�r���Q�Y�'���� � ����\0Li�����'��P��'j"9��hs�.��JO��H� �/��7�U�Q�c��<,�Ʃ�r�@���xB���
�l�bĈ�+1p�\32�io"�I�����b�/r�
�b�}�f��	Ɵ|�'`��+4��	s�Ȳz,��y��'����ˑ�l�fU������m��'
7���X�d]i6��"7k�#cͮ��D�<����5;�I��$�O6ġU�'�0Y���!\�t��=^::e�"�'�RO���i�De_����e+�O��N��+ӳ�8pq�ꝿ�xЏ˱��ɯHI�pR�B��s'��%��^�OYB�!֨ͼk��̊�)S��N%iK�����O�d-�'�?-~H s�c��:�"*L߬'�C�I�;�X�cᑲ{����f�(����'&#=���Xkqƛ!X�D%��.A��'�b�4�0ds�'8�'�w<-������c��$,��4z#e�:?ԸŚ����vy�+M�'=1���SQ͡>��bO�l�U���F 3�@�xJ�x�� ܻO9���ŴC��$�}*DW����V�%!vQ����|q��ٳ��ge��lZ���W�O�����0a�\�
c�;^S�ˆ)\�A�!�D��e��{%dž`�X��(���	5�HOV`�'��	6]]��V�P�앀#+
��4�)��R�t���̟�Iڟ�
��|��d>��vC0`蹠��	h�:�ˠ��wy���CB
0Ş�'�啣ge��c���sf��2g�)4uå`�g����B� \,�Ecҵt7^����Ɲg������O�Po��M�����d�O�"<��V�+Bޱ�S��,V0��*<D���Z*�����U�<<"<
��9�	3���<1�ϝ.}����'r����5FeڇxobyȗfQ�y��'����7�'d�1�.��E�P LBĥ�d�]�)p���P6#`F�����&fmd�"� Ϲ�p<	7 @�S�P5	�m��0A7�H�1���؇ñl)��J�	q&5X�kEM�ؼFx���?%�i��7m�O�Y�DJg�<��WhD5��C&�<��������,�3`�D�����Y�.�D��tOl�mZ�H��Ѡ:��Oٱ'�x�IGyrCR�`�6��O����|��/X�?�!�'E�H��IM���9Q�]��?Q�"���2���#��͡R^��'���,f��4�u�K�h�IP��,$��{_d2�O>`h�:����I:q��Q�8Vz�����p�`�	��Mּi�R���[Ңa*!0a�\ y�n�:�1Ov��3<OP�(�e��k�J+U.P$o�!��'��#=Ϛ������h>B �ف�X�R� )2��?��J�0�*a��!�?y��?)��P��Y�`��8䩒=1�|�ˣ��,Tصr5�`+/�������52�c>�O�L��Ą.
R(p(�퉵e��0�͆#�h����nP:5&TC�q��'t���ũF�ҭ�&�&��z��`��l�h�������>��?9���&�<A���.��� g�A���x2.�=��a�T/�Ը���t�'
�"=a
��d�'���e�P9\��m��:��s�.��R�fU��'�2�'�"��~J����$E˱!3n� ���^ 9 C#R��A�a喇5m��i��	�4G0���Ik|��X'0N� z���k4��f�#Mk�I
�O%g1F��@��Pe���$�> �'���dW�%����1l��b�LS�,���$�O�iH"Y����m�!6��h
�+���#��'�����IY��#\ԅH�X�Cl�8)Ƭ� )$b����4�?�)O����<i�;VV���H�5 �����}�@�����?�e�@�?���?��I�O^�Lّ��
R���b��E����=I�ȹ�.�nvm��	�J���%֤N�f���Kէ}윉
d���^r��R��a_`������F�B?o>6��<�R�������M��kM��+���0 ���7��E�
�3.O��D�<a��	R�|��`�	�=M�`�I��H�"���E{�O���	m&� O�=S�h��&_�6��<�ǊT���F�'}r\>�2DoVß�SX�,���QA��MB�J��$�ɤ=J$X�L��߆��C�L�O��4"����ߴJ(f5[�L�2��'؎%@T7P6��EdϷ-�Vm�u.ʬ_R!�W�9R7��Bn�V�"�Z�*1�X7'��DdI�	:�M��i���i�!dB�.��i >�Q�	Ydb1O�<<O(��DX���⦎������ F2��|��ɉ#�>���悥o��(1Y.:�0�4�?����?�瓑 �I���?����?��;$_�9�f��&�N� *�ho�0���R�Aʈ���p�����O�,�'̞�B�]Α�@�p�؋1*'=�8�#Q15=h$`�!���O[��'�D|S���(R �[�9'�9S0���9#��L>�� IrE��$��$�)�JSV�<u�A3����&��4���vɜS~"(2�S�O#�-S�FO�]a����>$�5�BvD�ղ��'�2�'��fo݉�����ͧ*Y
��V��d���5�e PLf�$����^���� .,O �kr��K�b3E��*UE�Y�)�/�M{a��r�i*�E���<i��6�	T(�*`��+��E--�*��I/�MK�i��[���IR��u�4����R��\�%&Y.�8��[/�m���Ӯ+JJ�('*�5+���<a�U� �'dtQ��'m"�'������ CC��#�n��AعR�'�_�$���'��Ɔ�w��kaL0%#���<��F[J�vU0úNzZ!��	Y�	�D��;�:yh� I�x��x�T�΀_t��K7�S�/��}V�' z�����?��Y�8
d���/�l��a	V H�<�C|���	ڟ��?E���;�6Y֣
�I���0�-̊���&|On�oZ;O�Ty"��Ȓb(�@j��jH�e��4��ǷEE�PoƟ8��U��l�d���4]u�a K3N��y �W�VR�'�����.䦽KN�ʧ��I�3-dpZ��9�x��a��)u��[RuS0�T6d�,��i�`i�xC&!T�T�腓�Q<C4�`�%����Mk�iJ��)>y�6L!��ҫX�DN�D�1O4�.<Od�)��"V���SU"^�Q��h(��'��"=Q���	 �#g��2��y�� $3;�I���ɞ���&CEß@�	������ߩI3*ӈE\xl�V��_U�`*�+���	)׃"XL�QBdc���"��|bO<�ĭ߾��-L�� 4�n ȧ��-5q2IѶ
�8�(�;`iJܧ�ēwΒ����{�zĉR;kC�i���iȊ���]�i>���S�? �	p��A&I�6-Q�,�{/�T��"OrLu��x��v��r������Ȏ��?a�'�!���L�
�İ)h�A�Ҭבa�x�@���?���?��g��O*��i>B��� ������_��Nt	�
1(�U �j1< �X�I���<1B�ى+s�p2�k��~Y&��4..�1%�>�i!�'�6y�ay2CJ^ׂ��b=d^v�"#���=E����?&���'}��'�r�'�"�'w��0%�|��D�T21�EO��y>�C�I�8Hhb��x>Lc�h W�c��8�Oh�0א�q!�i��'���;o]�:�Z�Z�k�^���ce�'�B�_;���'��)�㸁:���h�Ԭ�f�&�Hsf�3B��ĚU��'r�n)��'��q����e�Ċ��	 Pa,�.�e�)T�t�[����0<��/ɟ��ش79�	�:�
i+ ǒ�-f2� W�B	4y��I���	B�S�OQ��Ѐ��֦(p�'��i9�'��6�D>ap6�Q7�����A@�$�H���< ND�'���O��[>=��ʟ��&nc�a�.�+Ɗ�:o�̟��	�O�VAѡ�ܱP�X��H���?�O�哺rG�=�SAJ>36��d��k$�'/���2�ŸV�thyDh�p*�����,� *�pʧ�⬸�lۭ��	����O��}���O�PCE�
4�>i�TaR(O����'rvy���B�ZQ�iA�ጁC;l�	�*鑞�C���b�bE ��,#Y�=�i�(��Qx��#��E�@z�d��bv(pE�E�:D�P �؈Q�!���X�n�ZE�9D�ZdL�[��i� �*��UЁ6D�|Б"Μo],\�0�� ��5�T�1D����=3h-*6K��]������=D�$J5-ˉ#�4��ր�j"����0D�Hh���o����Í�m&@}�$�<D��:�ð[Z �P���k:�s�;D��%�2��Y[�i޾>|���2o.D����E֣}�F�ȧ ��,�P�q��1D�l��.�2�81K�w���0�;D�l��Ɂ�-�0q��H��z8�8D�\ S-B=簅���X5]�C�9D���)(m���QH��\��"D�̡u�	n��P�uFC-�qr#D<D�Yf,�S��+u�[�F3���A�8D�ؚ��JCD
�{�k�nj��Ԫ5D���w�Ӈ%n� �F0�^I��m2D�+�ȓtm8����-;�p�k׭/D�`�J�I6�Y��cS�Nw�H��.+D���^4x=���Q�=|��T��)D�|�V���CT"l�#�P#w��t�h5D�<	�-F)U3v܉#*J��>D��`�ϟjKHce�s��$�E
0D�`3qs��ZE�ԫ�~��F D�,ђb�O�E�#G��jw>!sRE4D�h�m8)|�8qd-Y��!�u�2D������| �h�v��9��[��2��0!k�Y�'�4l�U�	�93q�A/�����҂+�2�@�aM�{�G�M���i���2�#�I���ev�޶QN�w��)_�����OF?q�g�#LN�j2��,O|�ze���%�C�j"���7d��SΞ�2>5�"J�;`0JA{ϓ�!j�������'QT����iM�1���
?�����^@��<ni
� ����B7�1r��ᒮ�	@�쁊����7h�\3B&��y\k=
�B���ؕGU\�
���N���3Ȯ=��D���>q�%&�8��'X��h�w��;��'%�D��Ŝd��3������O&��)�rD(� ��0"W��%&��1��D}B��)B� !vm���7����T��B}�h�%�ߥ/�b���f��
Uz#�ϝ���\��$	x�V�Н?˓���P[��<�B: va��Ǆ���*qh ځ�?S�R�9P��cτ�<!��R��R!m�nF��N�4br>%1�N
�y�X��%?�O�(��:t`�q��qඡb�ĝnK��G>�hO�aGg�-(X=s���H���L�4C=.���M�nS����O�9n�(nP�a�6�|R��*jX�S$R�&!�P똊Iq*�X�/IP�\��w�g@)��%S�#��V��
 xH�f�
�u�'p
�tO�y*P�`Tn��V���N>!�n��^�����w���
U)m6(����
h�
�0c��E�V@J�5�=�$✞����E�O"��u��Q����1���f��tyrFO�]�p�� �tJ��ڤb��Y��h�#���eK� ��C�8Fq86i�yٶU�ʄ�(O4�0Q/@�B}��Y�/G�ʕ �C�Su�*�Oμ|r�'�L�KP�Q=�F�'��S�� rpD�H��̡�a�1u�H"O��!�=�)Sa�h�i�-r�&J�)���vf � ��x�7b��L+�Lϒw�8$a'�|RLΐs��Ӵ��E��ƪ|�����ăx �cA.�o�zeX����X+n���&��R���� 1��7O0�㑻[��Q��9�䐹_���"9O.q�p	ӹ������<a� 3���^���%���m��֕���X�͎����j�Eφ{�j\[�"*泟,j�Ⱥ�����.��8+��PqH!�ly��2�� {�(^(L0,��d���(OR������@҆`�@޾?�ԈS2)	9�()	 e?�����G}���S�'�5Vo��q��IC�D�E[beCu��S%� N4#>�����(ˬm
&8�����G)6��ᅅ#"K�]�`�~�	.o�[F�����O��,�Sj�Ez}��
�ɻOP�5�tM�|�"�&\0��6%���c�"�/do>��l�π�C��`NR�|4����Nq�:`	�(&a$T�O�O�l�j!a�Y�4/��N����5j�_dfȢ쑵
s�x��Bɯ#���An�*@"}�Ӻ��+ʽ;���BL�9�UR�Ŋ`yR+O(q�b�SAQ7k���v'�.�(O~�P��V?��#Z�Bi�X�1��E},b�KQ�<��$+��%]�~�S��5��Y5���)�BϏ�*`!�蘹U<�T�Daʿb���F{�c�J��08bf������`ORӁ)�f����c�/k�08�'Њ@��NI�Y6�X�� �0ā�CqBz�� *���V�֒~��Ms
n�Rb�\���T�=ڢ�K1���`2��T��9`�V��DY��h[��&D-�Abe�)�yb���(@T��Y�'M�  ̻u��:���Ǫ⡠F*ia:Ys#N�SYx�+t�� ^�j���Sq��<	��O��r��ܩB4���
@���Q.�-3�ڽʱ(U!
p�H8Ea��07�͋�(Ol�A�)E21nՐl����R�'�5y��AScV��7Om��'�2�X7jI4{BxPi�O�fA�1���m�R��/9ھ��fb_C�AK)�V�'?�i��k�IX�gS�Dq��3f�W���(ۣ×�5�6�I�O2�R�N�<Y64��79����#C*1����K��н:�Cā/O|-�p��h�y( �I!h^�%�зg>�.�{��B)���@Z M�j�"�ӜSP:D�F��H4��в�)�pi�+l�2I㘧�T��2�y�'֮����{�4�st��$�M� ��w�0��u�"}J|�����u$�ɡsyr�{!�Yx��9�E8'z'ƿs����~���w�Ё7�b�9��-v�T��R�˶CXz�mQ�2���:ܶ�N�3,�c�������4��@�?�͟_?�a���'$Њ�&M0pX�8��6��O I�D#���c
m�t��#�w�>�Áo�8���Ԏ�<��1k�˧
��s��C\x֍͓Tw�����Ǝ5Y�1y �սB� (�=���N3�����G��L�v����#���u JXY MҕyB
ђ�͢�^�����e�\�!��1����/0%,�'��-���~zӉߚ?r�M��ꂶA��A�'�Յw���'��$).i�cğ\Χ_�8L��暆!zv@�-���*����%�O�^.�� �?a��w�D�y���(���O&�6�7�>1��Ḡ>�Ѫs�'�P�{��5Tl�A��G�������ԏ��M(#d֧z
���F�/:�����J�}����:p����������B�/_��]/@���ĨYr�p��Q�\�p��nU�h���!�@W;�䉣N +�����<!�/�r?��;���h��$g|��MG[�G�|�� EW;k{� ���&[�L�'�v` taH`̸Q&VI�uq�O�2�Uʔ+U��Db-O�}YP�>Iv��^�����0���@��S9�-�P�!����,t�>�e��OE��I(���w��:D�x+ i�@����T���`�j��A��Ļ�E�:�?AY7���:X##ˣ�����՝}��9!�膡���db�>~����fw��1�L�57�t�z��&�䆁�����Ž=�����b�1����ưI�6͒�߾�F���A1Yj���!8l�!'v���e�,))��P"�	kϜC�� N6���0��Xz�h8ZG�q��M�t��� 4�� ���V�@��RD[�V��$�R$�/�4c�$�V,�"oP4�i���iŴ�k���<Ѣ�pQD�v�ɮr/ �<f������H&J/�+�y�I$N'�)�
��P�a�ራ��E�p��IB��(�BV9!�V� �c�L׸� 슪r�d��a.��D�u���)!h�:|��	�)><��THжd�k��s�D�	)I�M�D���V�0�9C�i�<���@�T��}T���N׸:d�x�U���Eވ�'5H�p�D�i�<�O��W���'r4���P�a�f�bQ��;E�̑!#H�8� $Rg�����T��2̐�;-w~�0�̀��8��e��&���҈{�F�Y�䓟zȰᅶ���E���AP/=� QkR�*n1O� UcB�j��҅	$���p՛|��X�Ii>ib.���p�W,� Z�
E���|R$� f�D�039�j ��\?)mJ�
�T�!#��\Z>��gW�	2�Ш�EU=r�*m¡��P�v��I�t�^�{�⁗5\�	�RmO�N㤵I�䥟��vDP�*��t۴�M��#��'�~�I�lAK� �8N�9�.��	�'j�8$����m#���$B].qX��� 2
��D��i�O����.pZ�wE�P�Љ��<�H��S@� DCt��'�(Q��֧oVy3��;2�P����z�r��Q�����A�n|�h����<�GK�<�9��Ȕh� q�&�T8�����H�cӢ ��
�t��P�V(��K7,��5m��}_�������ͻp˒;S����Y�azR�ߌ�Z�n/��P��	�d]^)"v/H�F*y����6��� ~�`�J�_:�i�އ �t�Z"O�j!�2S����掚!֨8�P�Vx 1!eN9/������C�֩:8� a���Y��qq��T���]�o}"�Ln��������>}����۱-����
�7��(�
���'l�)���h[b!Eɐ)�1y�t��'�F9�%n	"��sr�(n�>��g�<)#��@�'1�I�4gW\����?9�1��0�� ǂAV)�	� ��lü��-0��c�J��M3�5��O���B�Ƥj�l�".g(���be\�d\�&��-�v��ޟ *R΅�P���I$4�̹C���OrF�84��V_VE�'|ў�>�af��@L
P�F�ȏ3�2��0�����+$��:����±ͻ�x�$\.�> s�3 ���ɲ09�'�Z��E,�"�B���M�P<pdT%n��p�G*%�h`�Bg�+�90��>Y�`�LUlt�6mS�>����w�dʆ��s�����'�Xt��)#.K�8��-��P����h�~�agؘ�M{�m
9J��Yb��C��7�P�'&�Ex�dD,J����Ε��5S.O(�`�K�ڟ���D��+��-�ɘ�PhӁ"T�dT��`E��>���U���>��rkl���G�{R���W�	0�z#��V�X�Tи#�I�G��]�w�6��t�X+Wl|1s���8�69��"Ŭ�O(I؀*�%tt�4�Ʋm]�a���ۧ^�ўXȴK=�̲�dK�?��1��g�v��Y�]���6dޝQ�0Wd�	�1O�';ٗe؜{��):e���B<�ٴ8��X`�Y @��	��
����m�5K,�!	 �!�V��QkE�|�&\�3�Ke�1�GG�H�,��#I/�TBR��:��͂�°I���p��'�t��QD�H�Z��2 <{)�P#DW?Y�$q��5�S�'Y�t9��"��#��!����'X��${�����0>!�.�+$\�Ty�oM�?p�qbЊ�?%`�T��l��@C�'��U'�P"P�����d�� ������+vt�6k��8�
	1#�7c����A5{��l��KW�5����ī>I@���0k\Y�RK�1�"Ț�,Mr����1jzD�1II�$�h�2n��j�X'�&�� y�&�QF�V=Y�`Bv �<�&g�rJܨ#c�t?I��@�	$� a�'�6�z��
=\h4�xr-U2^B���d�7����NC�gWB�e-5,O�����0�\��$!
=:�𒧲i�u3�>��C��&�ў�SLD�m��Y���J�,�:�D[�RBT�ē]y��Ѐ�`�^��R�ș5;*�ڑ��*̘'��	YH���ᭆ�s�vU��w�Z�%X�kGB8�3d��8AxMr�=�����K�]� P:^;*���nP2'6<|k��E�$̀$�ly��p�� 
��g��?4�G):dn	bE�� s��@�'��4�W-i�`f3"ž�/�M�5,�)��!����_���\�H�����{�H�&�RE��@^��Ș-Y1�	�)"�q$'�.��\��~�'	���-�lh���+�"����y���?z(d�6�٧���2s��HO�hd�*�h�쀻�b¸J2D xAK,Y½��"O"qҒ+:X"P)�:K9���U�i�r�CCc�S��M��gՌ(�>5@���i�>HK�ȅg�<���7�	�甩d�T�d}D �}'Lt��	|1~D2"E�sF̳�*��Sp8���E�3'�q���p�ڕ	����gFFt��R7�T����	�s��4�� �SN[��Ez2�(!f�G��͋�o	B%���)�)`n�1�y"͎�m�\��maWd���ȉy�4[��:A<�)��=R���
�0�b�G7]2I'D�,��7a��rS�
DPa��>	筅�B԰��D�4(�T��0�Ɗm��/M [a}�EO�@6����fal���F�6���{t�^��B�I�&C�yr�ӼlO�Q#�32\"=��Y�aڊ�}
�eĞ
�L0��jWg��(�oE�<y$�˦9n&���E9"i0ĩ�¦y�0��$VqO?7�9jarC�&�y�n���aޕ'!�ؠ*OLL����<->�xhr��1�I�D��h��'oX`�UÄ�v$QsE�rz�8�2��:�'���i���T�UH�"l�~�A�'BJ��:G6W�/.����
r�<i6��)W���k�C	�T��vKo�<a������ ��YXYp5�l�<Q�+קd��Y�6�_CR!Xc��e�<���?&s*�3bi  �d,HP�F�<�P�ΩQ��I@aݿl����d�B�<� ,��b|.4�:TN�θ9�"O򑣰͈�9V���κ@��� �"O�U���R�R�0�k2������f"O�Y�WJY&�`YƧ]�t�f�iu"O����Y�UV��XF�Ҳj`A{�"Ov9���� ~}��d@�O���,�!�$�A���Ǣ�^D��(ը�W�!�����w��!gL�41���E�!�$Q4<�Ia�!UY��M)Gc!�Dː?�x�y��_%m���w���Sm!�D�W���Ҫ�Me��{`�
.P!��@�HVHD���� fS�r��ƅx6!�Ě�z���C�^6{7�Ѧǁ/)!�I�J��C��14)�(��;L"!���2���F"O�0ʅ�
{!�$QB�p)���<O�`z'�
o(!��0_c� Y��,Yvx2 X��!�D^)"`Ez�Ʊ= ���Ve��P�!�d',�0$RA-ٌE��ܑUD�+t�!���.�^�їR���:QF�= �!�$�;�`y+"���J�f$\%y�!���I���1p���FÂE23��;�!�T�sjd�PϜ*�H:p��y!�
V��Is��ۋ6,ĕڧ	Vn!�$�i�z��]�v*��aҝB!�DL&l^nL��'�U*��!̲p�!�$	$}\��R���H��H�ď�!�$�V
��d�*�:��"�	_g!�D�w�H`����F��aph͇;!�d_�Za �8����g�?l"!�MQ7���2��{[\�3G֞1�!�"g������p��̻f�_�R�!�dV�_�:@��*Ǜ����#D8/�!�d�*�[6�VB����#D�Z�!�_#zz��͓9r�8�YP�� 2!��Β#�ڹ)�OL��[���+\w!��-�����6+H�g�Jf!�$A}�VD�$��t��5��a�!��T����*�~�tx�%YP!�$ИTĆ���A�� 05D�7(4!�D��?�QN�(b��@�A-G�u�!�1X>NX��I�$c���E�]�J!�$ˁ@ѹ�%����QdHǒ
�'�)�M_/Gn�,A�'3r����'����u��X��fp��'��,Zdw���")5Eff�
	�'ՌD�0ʯ7��(���B����'/4 a�%ˌq�\�1V�Q+=�����'��0��k�T:)*�h�'bF���'�����ײ,Rб(D`�!^�H�x�'��$��k�0r6@�AVj��PUz
�'����R=/��EZ�jV�v��'����懐�M�����
o$�h8�'�dڴ'8�d��T�:��'���`ባD�05`S��6#N�
�'����4o����ʳ-ɚ��s�'ݲD�f T��6�P�@�%XH��'�&1pf�l)� E�=� m1�'��M]�Y����
H�,�
�'�m��E�p�(K!Z);}t1"
�'v�z�B�/q0mХm�1>�1	�':�@�-��	r����K�!i�K���"O��@�"s�[�*&��c�"Ov�;�%��B�^�[��
�k�D��"O� DH@���.?b1����7j4��"O<������ksH�{��[�3�n��Q"O� �V�#n��)qb�Ǖ�j����D=LO��Y2���[��J�c�5�!�"O�q�3���n~���Շ^�h����Cx�dذ�0���c�'
QNع���.D��qĀ>"���%�/�j�Տ-D�{$�Q�*'�k�GE�9�V��a�0������j�9i�P1Oϥb�����"O<�s6MJ�H:��WĞ���Q��d+�S⓾hq����K�9�%�t�K 1��B�-_�� �K�P���I#	j���p?�䡐#��Q �H�&"�2�zu�r��=�"넌��H¦�k�&�H ��W�<a E<znPAA�P8 ���E�O�<Y�$<�)`�Cߞ9�pj��I�<���0:lUz��֠6\���q�<�Gǔ�0�
ذp
�kQ�7i�k�<��
���Bm�0s����s�<�1d,|JN��C^� b�dF �m�<ɰ�F���+PT�>����k�e�<��˖�;)��)���`.��%"QM��hO�O�,Kf�ίU��ؠOZ�_(���	�'d���D�}��|�L� @��	�'�ۢD��C��ppj�p%n��
�'W�+�'	�n+����"f�jz
�'3HUǌ��}~|��"X��)�
ד��'#�� ��`�&��M
PI@��'AU��f�5��Q���	L6�A 	�'�:|a�a�U`
	�2�����	�'�\��`ѝc�`y+b����q	�'`�ٰ#G�qX��( �n�BI<	����ކ\"!��Al���P��%5!��P;SH<�aŁ2A[P��q�]*!��\j����	�U*��@��y!򤌭T ����CĊyl�p��(V�.�!�D�4��H�D�D H�y�\:&!�$�Pxms4�H�Z	6}��P
O4!��T>�.Mi�Ӎ  j���ո\�!�D��_�Vi���[�E�5#!�$I"C~�m�g�\�X�|°�G�=f��>�O:U!�*�4]Ԍ�P쒚[Ǯ�"O�)�2	����TP�k��'�|qG"O4�"ܴs�j���Y��.���"O�M��8�ܑ2D���n����"OT)�-\$X448P��ڌ+t�TZQ"O"�������r(ϸF���"O��h�3/��qi��U�"��p"O��)�l�;�쁑u����?Ol���!�D@f����!�E����!�щZ����-@�!�bH{Ռь1�!�$�r-�������X���%G�L�!�$K[��� S��I����@��/�!�d�J����w��B����P ז'�!�D��%~��iD" �>�B����Oy�f�P>`�\����\�;�|TA�"O�0B�㓶`��dYg��j�P�Y�"O\��h��rX|�v��>�eb%�d*�S�1MI�1�#��^��Y#�_%5[!�d֜J�tyt̏�)�0����-Xw��=E��'�(��re@(�b1��h��S���p�'��ԫ��B2_`����/JV���s��0�
Eb�0���G�4)�ȓѳ,ȈE]8"��,�T���S�? ����CqH�ES�� 3=~��f"Ox�0rA��x��]0 E�- d�1W"O��f.N�D��
T@8P�p�"O<���O^�a�T��l��ɭ٩D"O�H�cFF�	1(�%kŉ�D@��"OH$��ޕ8��x�j�76��|	D"O�]�o�;^n�x �'��4��Pq"O�Q�p	H�g�h��I	�G�,��"O(L��C�,���S�ƶ���H�"ON8q�+#S��r�R�����a*O���\�Hyi⊃�9�0�'WJ�`fF�x���� �0~8qY�'<�K��QP}��"Fp�{�''�ٓ��X?��}�R&�M��q��'_F9J�Iĕ:�4�)!R�G>�,��$g��#~d+�<�Θz��چ^���U�VU�<�ĈI�p"��>5����6�JL�<��e�{���`P�t�Zl��)�_�<���A�����ϼm@��7��Y�<Ɇ-T�[�Q�E�\d��o�<���R �(���~�e�BA�@�'Q?��։�$e~��eNQ3"�����=����|#d�Y�P=p��.
��%��d.\O�����L�\$dd{���((�:�"Oj���L��>'���P̔�[��Y�d"O�;o؇�&�Δ N����"O�%���1F-\���^�_~Z�y�"OHT�B�E�{�dyۃ��o� �Z�"O6�I%���@�F^�	��&"D��A� 
3>lY�w�R�!ڵY�>ғ�p<	�ǒd�r�"KM�KQ�M%Nx�<ie*�UN�՘�	�n����]�!�d��|�b=H5�T�[TF@�p�R	!�D�-Ӕ�yC�M��$3'�Ĥi�!���|������NN�Ms�T9�!��RP<����E &�.�{��F�a�!�?M[.� ���~�T9P�_�	�!�Y��:�PQ�M3�F=�!��!,�~�
��3C� ��2�!�
�abri;t��h<����ǝ	V!�d�	�hb�@�t(���E!��48!��G;�X@vm׸f7��X!�/} !�d�8�!����<*2R�6I��!���]�^=����S��qH�
a3!�M�t(��q��@�k�4�S�$@8!�D�4K&�l9�!��a�����>
!�dG\�MZv��x�V�A��\�!���aZ،�2JC=&제]�e�!��ܭAw��A$2�"Œ���5v!�D�C�ءsF-e���ԤX!�D��(&��
G F���S�!TL�!��?�����C �f�j5�ÞN�!�d�=eU`X{�O6��0��hW�)�!��$��5�cLA�m� ke��@�!����x�E�D�������)v�!�d%p�a �tl2�#���q!�D\��b�O�/J����ۄ!�ܨ&R@9�c�=e7~�"m�Q�!��XI�F�����(?O�1BVΎ�}�!�d�*
�a[1j �5:0}+T��f�!�d�"H[�����00��s��H�!��Z�@Bp�R�Ү&ni�¤�N�!�D�R�H�z�mǊbFp%D���!�D��f�J���-��Vdd��!�� �ѫSbT��t`��&�2X���a"O`��	��4���{�DW���8S"O���Ѯf���R�d�j�0�"Ot� 4m�n�9�Wf�������"OXDȃ.]�j��c��8S�t�"OԔ3pK��#����gje!�"O�$�@>'���K7t����f"O�z��Q�
H!p��<Q7"O`� t�]�RPB��e�^)͚|�"OR�aS(T���3	î��d�"O

ČЏxQ6 �D�FU����"O(se)�
1rpA٪4Q�TYU"O(TYG�W?����&�%CC"O:U� ��/{���%O6 ��`!"OX�YChE1%셢�P�a`���1"OTd�� �H��įZ�"r���"O�uX�F��&���R�˴5��d�"Ox @���~���K�ʃ��F�#q"O���5�E�Z�m����+�JX"O�M��1~��  E�8:� ( �"O��XA&�pX�GNS�d�F͚C"O�u��"�/a��@�A�@�rC"O�,�e�+_���-��t�4)"Oh�egI+[Ba��탨4ި�"O��pr��V�0�j�+�#`�p"OT[V#J9aZ��8���"�\Jw"O�����8<��2#�\�l	 �9�"OF8��
�0>ҝi2ŝY���p "O2�:weX�:���R&Yq����y� Q�
K���;&up���y��ҶolA�o�!�ʩ3&S�yr,ҡQ�����%P8���)3)ռ�y¤��"-b�	FEyӈ[,�y�Nudy�Х ?V( �"φ�y2�f��Z���H�`����D��y�k 5>/d��a�M�ȥڰh��yB�ɏN�}Kd̒8@�R$�v+ֱ�y��!F `���15(��Wg�.�yR ��~�
 �a�5"�U�6��ye�L�b��65r���y��H��|�Ҥ�<��#v�W��yB�O����Z�*;2l 1%Ӗ�y�W�:l�A����T�hdjE#�y�Iɣj�T�:��P��9�`) ��y��ى%� U�r�=31VYj�eZ��ybD� �蠸���(�� �kF��yҊ�}��L��S�7�32��yR�ǐY���
2��5uv�rbY2�y���[�����%�+,bxq�=�y"��j�1	`�T Vx�z#B��y��֏k�t)$�Ê)p�H��A
��y� �[����
� �"87�M��y�цޚ�P���|��j�ybF�	h 4I���4^*���Ӟ�y2#Y=B ����˔2.�>��@	�y�L\�1��$�c��v�p�����y�F�Z�\0��&D�s�a�MF��y[�ER�p�ٞp@�aWK���yb�R�<3�CM�?�
d#�-[��yaÇPJ6�ʖ�)3b�5
���:�yi�V��Q�'EM�0:=���/�y�����@�r�� '�R=�4I�<�y��;4h�I�6����`�׿�y��-86��P�*G�R$HbSN��y
� $!R"�"OXR�k���z��Y�"O��1���#�u�P%�3�p�{3"O,��T�ѣ�D]r��ׇ �d��"O$���A*0�ȓ�fC�Y��=�"Ox��h�X�ఫQKI�$X�!"O��0��۽(7P���ɮIDL�"OX��(��6�~��E��*%a)�'/dB��x�����A�8w ��'S�Ղ�j��_)t��e*1�M�
�'-�x����av ��W�&vl�l{
�'Q��@���	f(z]r��A#lE2T�	�'��\ �o�"s�p�3�XX�!	�'�4���[
uvn}3OO���'�JU�ENS@�T<�8�P�'�4��!њV$x}��
Z
3?�'լ���]�Z�n�J� N`.^m�
�'���0�z�.�Q%��M����'$�yQ�%S�i�` j��C�d�H�'H<A �G����?�D�
�'�� ;�˅�m^Y2S/*�
)r	�'�>ٚЊ§1��]��&ފ$T�x`	�'q9�&�L .�s�B�/L7B���'� qq*E�T�i��R=�U��'� �����V6�9�S��9'$���':�%(���9�A� *����'%�i(v�W�t�a�R��N�TT��g�4�t�%p��oԥcŨ@�ȓ$fq!k�0,74JQ�D(6���}�N��D]�Z-ltC��$^� Ѕ�]1��A$�3����ŞH4����s�f0�2�,=j�HS�b��h1D@��n`NP` �y�\�C��%솸��>[^[�+�o]4l��Q<u�6��UṔ���X���w�S"8��Ɇ�4����4����.�S�O�X݇�ZUF)05C�E�����-�@��ca����z�k�&�o���LwN�Y�& @�l���jە^Ｍ���QJ�^T�L�m�ʬ��z��\{����5(�ٓ˂ik�q�ȓS�vE�3�N��ͩR��aȌ��ȓ�T
4�^ʆ��!�F�"�d��'a��LU����  !�p���'K������(���+g�:/ ���'�(���'��M2��lޥ;�@���'ĎD�$@'B�����ΐ/Ca��'�TP�3��/�r8��-)$5�(p�'��i)p�6��8C�:q��'�
����uB&����t	�'o��J$jK3I�l���LV "�l��'��[��M��=�D�
���4!o6C����u��\?'@R�o0N�C�*A��0	 �F�?�>)��Y9(�C�o����7CH�W�i��.P�B�0 .��Z�c
.>�y�D`C(��C�I�y�)�J�$Ú4����*��C��M`@���C'+N�sD�X3��C�ɹ�N	���[�ɃPc�dKnC䉲)'��B�͓5���YuN��4=xC�ɘo�FPa����H��m��N�.D�B�:Rt�i�\Ӟ\��`M�}�&C䉭;0{CK�;OBd�#֏�?I�C�n�	p�&R��Dp�FI434�C��,c�2�s!�J�V?B�s��< ��B�)� ��Ra��Mw�y�� ��Ig�	&"O��"l�t\0���3�~uK "O.�bi��b�j9��H0L�P*�"O�xB�K&c�l[���e�U�0"O,���nə58`C%��}��c"O�PP'ς�PqP@CS�D'#�h4��"O�D���[�r�S�B�Zt�A"O�D��P?|����O�-Y���U"O��1H��nv��kW-��
�ȴ��"O.8)�J�2QD&N�SϠ�ٴ"O!h��O>Z@�1F�`�Y'"O��h0Dܓh+dQO]b�0�"O@Ԃ�(oHn����\�Y�B��$"O�t㦯�o��{!��+�(�)�"O��UJB�G�c`�_�в��""O,�R5E��z	�A�5�-dδtB!"O�4��+�\J�5�s�k��P+`"O���`�v@��s�k�*����"O��PJȅ(�9ƪ^!�p��#"O@�a� L�k�v(ʖ�����@�"O�I����9gzvq�o�$y�V4�"O�S @�S=$�����ET=�r"O�]�ؐ�X(�fR�[^���T"O���#GA�ig�=��G�/gF�Y0�"O6�.ʣO(M�'_�	lia�"O��S�B&CI&,���R0h��"O �%؊[30D���h�@��"O�$��8�̘����?�h�S�"O��1��ʲ:�����l2�*�p�"O�TYcl E�}����K����d"O�t��"/�`dXT�ݞS��xV"O@9y��'|0q@0$�eBfXQ"O��A��F�s͔��##ىz4dA�U"O�eiS�ߝ��8�KŊ8��I2 "O�pQ��_�KKz�G*��k�T��"Oz���cT��"�J�:�(U��'��-Z`�çvShXZԎ@�J�����'2��c�+�1=dx1R���!n�`0[	�'H*�ҵMX"1� 
f ϳb��T�	�'��%�%M;BBr����*�<��'�=�E�f!�C-2�.@��'(�B��Ȋ^���`͟���'�z��W�/4���KS�-��j�'���� hE;�.�6gȥ��m��'Gb��m��Y8M(0��)����'�t�����;p6�c`�ɤ�9��'мI�v��,)���ƢNѬ���'.�i���\�R0��2P�'Lt��#���z�s'�
^�D��';`�$3(��UpgG�Y��"�'s�u���v�6xcfǄ�U����'<T�#��0���A��9L<@��'q�h��4i ��@�Дlس�'��ݪR,ϡt�F���B��:u��'D��i[�|�X2` �,�t}�
�'l��xÃ��u�dj���e��'qbQ�gE%Dv�Q���^�.)��'���5,����a�O ����'Ē��b --�4���B�AG��
�'ap���	��U�ۦς5E���'2eP�
�4=���s��B>��B�'`(�gH�	�Z��EL�f���Q
�'#�t�7 ��@�ɀmC��juk�'O��xׄƁN� 	��Ț
?��x��� ��:UȱhC�Y�J%n%z��"OV� ��r��,"�I�D�[�"O�	X�`��d$�$��]t FI��"Oh�#���eՌl���Ǝ(�0т�"O|�X�,ޘwQ�A�=	�<��"Ot�&�ޟR���V�Ţl{FͲ�"O(�(�J�-/�Գ�BGAkd)�"O1B�*9�bl���N?Vbr�"�"O�q��ƅV/��á/Q��Dd�&"O"� ��CEx� �8Zwh�0�"O:k�@'\����ꆫ-�:��3"O���203l��I $�_Uv�j�"Opi�d�"2�QW�t�e��"Of�{�aN[�65���U:x2���"O~d�ц6$���)Q���g=� [G"O�`�s���%~F����Q.2Z�D"O��i�ۛ$(�:u��
0�ģ'"O����Ԅy��	c%��k"O@�Kqh$7GƴӓH��>�:d�r"O.l{��إyR�Tx�Ɋ$⢥ʖ"OX���hI>N���A�Gǎ�s0"O��%K��y����R�P~� �"O�Ĩ'�Xvb�UA�h�|:�"O�]{�-�3` I�s�]�$�x+�"O���k	W9�IYT�Z=K��3a"O.���Z���XËH�c�JxY�"O�t�%��.)�AqI�=_hh؂�"O�ԋ���7hW���.A�GiڀY'"O:]�ŋ�_"rUѣ �>}a�\�"O�]��eJ�⌨c%@HW����"O(�2�HɫC�ڰ�&E(^��H4"Od"@ȏ�`wn%�
�n� xB"OHi۶`W0w��&�2���a"O�����0_W��`�A[6O�x��"O�A�L����X��@D��"O�eZ_���I��
�`��L�1"O0�@f���@ܠE�ƨS�����"O,tq U'v�`��CO$;����$"O�]�ggےT4	dbVWd*Q[�"O��S�o�/Q
�`�)1 ȑ�"O��+kK�:�\ p�@�"2��+�"O�T!���6�X`����2~�h�"O^�k���%C؞ݣ#��%	��1"O�s�.M�Gj�[0�U@�JQ"O(���B[-���Љ��F8:�S�"Of}A��˨N������U�,(�b�"O.�蠬��p�z(���͓6(�*�"O^���h�_�4�ѱa�}���"OtY;��@ C���	�%b1"ON��m'�n������4 c�"OV���b�Q���q��|����"One�Qm,Mq���͓{����"OT�0!Ȃ��
��G�$mk$՘�"O=�%��GJ�(��U�X\ny��"O��#�GK�W(|aj���EI��Cf"O�H�c�ÿp��M*&��0"O:+k�-4��-:�q("O:бp�Vy�D��g�%K��u��"O�	p���*l���UGٿ$N^QS"O��� !�u�p�% K?[
�s"O�!�䅃�Zxu���űn���#�"O���d�%j�d�B�L_�C�8�"O���L�4A"�ˍ	��5@"O��`�d�-�m�* �,J�<�"O� .�� P�
6pF��!S��1�"O*��?EF\@�E�^�iR@�B�"OJl 0)�n��MY�Ǚ�(�
�"O2��Sh�=<z��K�F�?��A*�"OXx�qlO=a;� A�I���y�"O��8V�E��n�$����"O��kQ�J:#A����#Q,G����`"O�<s5�=U�t����38>m0�"Oޕ1�-�r:�-�GKҾ!j� g"O4�{ Kƪ8����+�_:D-"5"O �*CÐ���Q8B^�;���"O�a"CL��&�@���$3@���1"O�m	V�٫R�l�eY�lP���Q"O2DT��9dV`��T�PK~��"O]*t�\�N
�JҢ�d�iC�"O�,� fO#!� 27�˫�0"O(u�6�{T�"a�3%�&�z"O�4�%޿��Òe�5�.��"O��aB<��1���@#�"O�J��D,G(�d§cŬUkL�� "O`e
@o��-�69�#-Ⱦz�zDs�"O�90˄��>2�L�<{��=,�!򄍏b��aPBh��ĉ�L^1.u!�D|m(| PN�8�ܡ�G$u�!�GIN���Eů����lT�NI!���4 C�'�;�p蚷�ԩ,�!�U 9��x�\R�!��鄬U�!�dY `�;��RLN}Z�
؂�!�$�a^�! w��];j���&X!��T\dq�(ǀU,񒢆��.A!��-$V�2�مv�~1���#1!�d�{H!ۀ���!��J1ΗQ?!�M�Q:a#�dڂ��P��S!��CI�--f� k��A�L�Ԅȓ�D;cΗ� �
�5zH�E�������n u���7"�r��`��&�0�A�	�� "F$)Rf��iN���ȓR?�]J�2 ����0̬��ȓ�pԂ�A�+:]��1�ѯU����ȓNLt� T��abl
�  V��� RĪ�VZVȧ �,c�����D�MK�$�1���{�O�)x}���ȓuU�s�	D���[�MF$;�@݄�oX�e�VKF�F�esp`�'Cv�I�ȓ8oB-�Q�̠5_z%��hO &�U�ȓUq�rEn��X� ��ܤ=����+s��*��/�
�`@(J5bŅ�B��ă�Ý�p.~y�CI�[x"<�ȓ{�D���H=��pe���q$�م�1��=ځ"?m�@K��w�2=�ȓ_�~��BY�Q�����$V ����n��@�35���FjY�SH� ��s�R�"^.8���P"�8��ȓZ*��Z��-�&�hѡ��Ewn��ȓ }�aH��JxJ>Xr�$�0��ȓVﶸ!"��?��0�BǙ"� y�ȓ1��%�b�)��- ۷%b��+B$� �5��DA0B�"�Pp��|#ΰ�R�^:9�X�y0��!*�hX��%�P��Ʈ	���J�
57�nنȓ{F��%��=Z ��G�܌l�J��ȓ=,�՛q� "Bni�f$�	��`��Q���`#˗1 ��"�f��c}��H&X M�J
2fO�u�֥��S�? l��V�V-	x���a,G�{�)�"OP� ����d�V�ᳪG�H��]��"O��B��Iw�Fh20K��
��s"O�]P��)�!�"s�9S"O��@Uj�	,��0����Cf��8v"O��"��u��U��K�nah<��"Ov�'�3g
8��E�ݗ2�� �"Oz���߹$��XIw�
6�<5T"O�4�	`Ò9*g�ɒ#�@��'"O^<�"��_�\��b%:7�q�Q"O �Th�@�j���4��pp�"O��b��ƌ�C"_�k0�<jf"O��V!OI���A��9>V��*O,���҂A=��{G���<dP	�'� my���mz�����2xj�'G�aK�g�������G1'*�e��'�8`)�(����Pn�0�*���',r�I�->a���p��
3Q��<��'����H��Ip���)��E��u[�'*��f*����fD��gb�P�'2X0B&(��2W�֓_����'�~�AT��<n��IAv�.��l��''J��'j��Q`����ʜ�>"�'���p��D0.��)�S�
)ni��'�����6v�́ &��|f��R�'���gL�7�����M!ua�ţ�'s
�
�ĵ=���թ�d����'�@eD�!��D[T@�)�'�����Y�WO�L��8GF*���'q�l��5JƬ��y�%��'�D�c��"|i��!��r�]B�'8l�#��3
���⁊�fR>\��'�2)#��'b}�(��O�L����'@ ; ���A��� \��5��'3viRr.
ٰ�ym� J@��'�8̐���Ppt�p�k�2s�d���'EjY���(A"|��JC�!���']Z]S�[�py<<:)��f�h�'�p8��R�=d��xv�Բ�
�'���0�aʀfE�ԃ�ia�mA
�'""Y���_�:�
�+���0�,��'	���	�,X��Q��ۚU�D��'H��B�)44d�g�X�N�D|��'8��B胦f�DԲ�+� AJ��'�^q�$�
|:��"O�<3S(��'�fdHa�]�a,�|@"	�+$�����'�$q*������A�DHL�'vjE#��ʠ/�q¡�!O�=Q�'<"J:�H[1��A[�=��'���s�LAE�� !%\7����'�pɀ�S&��}Q.�W��@��'�������ty#ҫ�U,HŰ�'*���H�6E����Z$`�6i��'�0�!*6j�S��ʬ$�P��'��i���:�$PT�G�e��
�'O�l	�]�yylA��5HV��
�'�
0��$�O�VseT�r�
�'a���˝��|�`I-J���A�'�B�ibF��R���BVC��%b�'�F��!Ll���C8�d��'^!�ƮZ�7�*���IY0z�d�a�'Y���:D�M@�F�1��'s0(q��;f�X7�?➌��'��'`Z,)�$���B�%������ *-yp��I�|1��Цm�r�"O��C�F᪝C�����e�f"OxD��(KL#��w�	�|X�"O�[�b�@ӎ] �f��v
J<+v"OJ� F�L���%%N�q"O��Z@�Y�/������%l��e�"O�p`4�k�8�G�\�Zx(M9f"O�X�$�#`<}ڂC�omr��"O��I��Xp�\�db:c(��"Oԁ`5O��ya�-�}7\��f�l�ç
I5Z�	����&:R�)����qSU�>��bE$7B��Z|f��7nۗ
9 ��0h�%� Ї�5�i�)�x��RԇQgo҄��u&蚖C@�Blb�ש#�<I�ȓ}ੰ7���gZ��&��b�fx�ȓ_Ҳ��ƅ�I�E��OK(h䘆�k��j��C��ʬP��&�<��2�*Yh%�U�q�����(Y�� �ȓ&��ٓ0�ы�V	��!
"Ѕ�Cf�A`ġGz�i��,Y6��ȓx�B"K��;�0�+MU�A�ȓa.���+CRq#��C����ȓ��$���څaa2��w�S��E��}XE����vvLui��H�]���ȓF,���w�UI�dM�+���"O ��a"ͣu�v��R�\:<x`YF"ON�kq��W�\@	�$�4-_�5K"O��Y#�M�u5�@�لT�|C�"O�m���Q�<�lq����7��q��"Ob��.0F��3T땅�B9:Q"Of�i⣘9b��\("�K(:���;�"O��E�� $h�)T,JJt�G"O�LPw���t�N�*����9(��Q�"O�,Ѐ���P�T3�O�[�����"Oh�*ԠZ5r�4apg��Z��pj&"O�*rE��v��	BjB5c��hc"O4��c��f���G}6:�x&"Oޤ@��K�P�K�@�Q��"Op�� ��)��<P�)^���r"Of�"SB�F�<9�G%j���6"O0|��O��FRԌxa&W�{��	sb"O���X+,r��[ ��qg��3T"O09u�K-=?2%ӥ%�(0J	Ha"O���v�}�ЎI�kO$YB "On�P�SN�(Q���N�Ĺ�G"O6�IևU�f�R����@�=Δ��"O���N!�v��D�(p��Ȳ"OP������x�����4z��C"O����#sI ��$��o�V8�'"O����UB�,8�t�<3ΒY�f"O��c��Hr�{�9�"O�ѻE.��RAJ��I1�ΐ��"Ol`�"@�a���@(M1}�>�q�"O�ѰF�
�f�.��U�&;�|�w"O,�
� �\)���Q��x�*Ox���%�j'���gY8Z*�
�'{�(Z ��$�>�e�P�X}��'[�9*��Īq��؄�LA����'�ȡW�J�TkQ@�R�Yr}�'0��"���@V���o��P��H�'�V��f�̆MT�e�d�H�zfք
�'zQj��k[.�	��kx���	�'��|:��l�&u��(��[	:����� �u�6�^/n�X������z�"O�� ���g�bA���4;��x� ��2�S�IЖeL�Y:fY}���H_��!���3B�N�s����)6'J�9�!�D������G�#X
���s S^h!�$_�'��@��K9L�l���#Y!�$��5:�bW�ǌ6�DUn^�=!�Wbd�0W�&������3�!��#p ��r��I�C��!���;NG.�YWn͞c�N��
��}�!򄕻]��x��D�X܀���7a�!���usViZ�O�\1� Ɛ��!��\
�2�0�%�4a9QBQ
[d!�D��)
��K�@��3�T��!�$w�͒�1*�d��OΕ�!�a���x���+x�͛a肌{	!�$P9L��0���*hv&���dN��!�dX�~�����I�Xf�|Y�i���!�D��$��ڤ��VH�I�%��!�dDg1���S$C�{>(��HO!���A� �� �Y �d���G׀K�!�E�14�ԉpڲg��Ad���!�˰��"p�/&�BQr�dE�W!��]("��P����m��4�W�B!�d�7�=��;3n)zQ�_�P!�D�<"~��u)D�I
����A�ch!�D�y�΁؄W2Ag40�gb�g�!�d��h.F�p,��a_JI3"�كr�!�ܼ�­Q@A6"��i�����!�����c��CN䵲�:y�]�ȓ����3��0V �+��.Q�|���V.Z4�`�'ζc�R�V�y�ȓW"V�bSG�C�Y�Cj�$&�,���yRqω*4�E󌚣L���7�x�����34�Q�V�=�荅ȓ5�Fq��+�Eb�-ʃ!$x�H��������sl�)��n�V��"�D�3 ��'<�s�ퟘT,�\�ȓ:�bl���ַ4��!�Fn�x��L��e@R�PE�F�B���b2�@ 7AbC�I"lb�2�a�>ข��ߵO�LC�		L��ɹ���Nj�
���9
_�C��|�V��r@bȤ@ ��O�C�I1~3�-�7�
V)�����TpzC䉸�4��h�+wd5Aїn@C�"Y����c�'i�ȱP��fB�I�F�T
��H�5������2{�C�	1 ����aG�'"JPI��N�0�lC�ɺ0�N�ha�, �X�`jN+
�C�ɕbf�-��/�~���)��x C��*|��P+`�/GZ���
I�Pn�B�	;����#s~��cR�H�K~�B�=22��Y�#[9]�r��b�){؀B�ɥKWb����?~�|\;�fV�5|�C�	,6�ȝ)(��4SFxs֭��A�JB��3;�R-9!�UF��rn��B�I� ��+��xO�� ��͌?��C�	9}��+*R��1���˭C�B䉛��2�-�=&�:+�a*�C�ɕ}D�"f�]36��A�O27��C�	�Q��ac���'�v��&��BC�=�tI�=3Tvi�Wa�)�C�	�2��aiG_9�t)I3��3m��C�8��4�a�X+ULɉ���.FtB�)� �=�C�#^p%HB��xH
��"O��lS�}L0�r 	[� ��!��"O��+"���4�Uybm��j���"O���3���K��`�6�G5v|�A�"OP�Ұ�O�+b�ACAF�RY� SP"O\�(["%I&�Y�o�M>hB�"O���Pu��2jN��r"Ov��ٗj�$���lR:T�d��"O��& U�h	"�ꙬyAypa"OƩ9�\�?��x J!:f�6"O��uZظ�Mu(�x��"O�}���Z)2=�!o�#3'DL3T"OD�J�e��lM`�{�m
{<�G"O�� �k�6$%As̊�2y28*�"O5�&Ȗ�L�x�ڀ��@]�M��"OT��`ˬD�*����K�p$~�"O"��6x�9�X&,�=j�"O� �Rdъg���#d�!�L�s"Ox"�^;7F�p���P!�"O�����<�>�`cC��4,Z���"O�ܙ��I�==Ɓ))!Bt@ "O�lBQ�;B�Xl�/F�0�|��"O4�y7��4��3$����U"O|�� ��p��0�P��2���"Oz4��kO�?��P� ���tk��"Oj��eJ�W��� ��"R��b"O�����Z��{d���1U0h��"O�}�B��*q�十\S|!��"O�y`m(-~�*S�Z,�R�"O21��$h��P�mL�w�,�"O<H��)�1w��%�����r��p�1"O �q��%`p��Хo�E�� c"On\��@0��h�Oݝ�&1�E"O�K��*��AT�!E���"O �Kף=  �i7/ӫI�ܓ"Oz5�rk�;VƐX��_e�rY�"O
Q��\?���2�  \z(aQ"O�uJ�	�i��!x�+��]Ұ'"O�����J���p���3��� �!��W A�M5�E)zʖ�`�
H,�!�D�Y*��5ƅ+]��(z�(Z�A�!�D�n�d���ɜ0Ĳ�Q7��}�!�$X�8���г�E�|���E!T�B�!��Z&dUb�c��(�ȩ6�F�^!�ıY�����D'ZO�ae��-Q!�+���1#M
pfX�y���(;;!�DȘp� F��gR�q�@'O�!�d�?V�L�bϺZ8V�0�MB$Y|!򤜣)�V����;��LAq-�)b!�DN-S��� ���]Ȇ�Z&-a!�d�h��q7�����폂.O!�B�`T~p�qg�%^�,t8��>!򤒦sl�0v$��
���U��1s8!�$O/:t�pr�֊:�q�+L�M!�Y[$����)G���Y���G!�D�"Z I��U	B1�hC �!�Y�!\�d��-�L�X��RnP�`�!��]!�ք	�n&�x�ذN�!�گf��8i�J�+B=�Fy�!��M�y"0am�,?��u��S�:�!�䞚ig�	��k�m��%�.�O�!��́&@ �SS�M�(�����ʊn�!�D((��P;�
P{�Ҙ!��A��!�R�-��!�f�7�~́��h�!�� �0p�ϝ��0t�� CQ�૲"O��;�A�h[`��`���訡!"O�)x��Ő�D�S��9Pڼ؉a"O�!�6�T(a�@Z�����"Oj{�"//Z����C,_�%�#"Obl8��@m�T�q����P6���"O��s�^��� e�3�8�"O���ȏ�:���v)��_�hyS"O�Ĺ��C�s�ܕ�T(ħA���@@"O*5�Pȅ�%l������R��	�'��)r ��1�n��Ƈ��hԢ�'���� ͥ[�PU��&ʛNJ�h��'����n1|�XJ�i�-Ka*X�'�0���
	�
z\���C�>},���'P&P ��ΉI�8�WI�2L3b��'Vh	B�F�T�>�N0Qnx+�'��t�!A�e�zi`���Q��@��'��ԍ+9���$aP2<�ɢ�'���|m��QdL�5Ś�'���cBd�?zƸ�*GMR�1�D	����>B yZ� *GL�qB@Z5�yb���L�P�X��όx�!��1�y2��6I&���,z� uj1ݒ�y���.qO�=1T��v�$� �S��y�J�7%V�}ӧ�kaD�]�;�lU��'�V��Љ�P7V��2�W!k�5��'�\���C*T����9L)����'��ɳQ�l���r1#M|�l2�'֬X @�S�jg%J񏀑H��)��'�. ��"}�0ҍɅ
�
pi�'��QV��f�(Փb���z���'Ɋ���g�)S�.I*�m��+�4}:�'�؅��ǦS�>� B-ܖR���j
�'L()�ŢS�9��Qk�> �x	�'�:����6>��!R�A�E�΍q	�'�T�&�H��Č�Ԁ��Apv|��'��A��-I(n��(���8*)<��'�)kE�֬O�<�#�+�;�r\�'��y�CE�A�B��-�f8��1�'� $���2z� �t�9K4�U"�'���U���������-<ЌR�'�<�i1�I�e�f):d(B5+�����'7pJ�Ĉ�!��a��!hҨA�'A������{�űN�5uƭ1
�'�Y �C�)�I%��	�![
�'�x����*/Ԭ��P3j��{	�'|�!i�X )�@����đu<^Щ�'��l���ݞޞ����4X>n��
�'����F��!��9&��g��� �'Lp�ӳ�G�o��H��S)�����'Pj@��*y�h���. T�H8"�'hHKᩉ�O$�۴e�($P��
�'_�J$�Gc� F&�t��'6�a���;�d�:�'IA��8�'hv��T�ϰ����/�l�����'&�ۃ��=:z�l�d��0���R�'�� 1��x��5ɣd��0�R�	�'v�Trv�
W�r�����7#����'��DkDJԥK��#Ђ..�9a�'%T�Ȣko�`�PRCF�5ђt��'��Yu�,h\Y��� '���
�'���"畑���T*�`	�'*��w#�2�:(A�G�~�����'��
������p�.�B����� ���ի�y���O� ��%��"O�X����RF��ỏ��<2�"O������"�l�#ӎ	*�#P"O�L8������#J�n�y��"O���FsK� �� m'vQ0�"O��:�B�Wz��jB�ߴx8L��"O����\)`�fXcd�"r98�"O��	�B���Ĭ��/ڰ[Q̱"O:���B }H��LG�Q4J��S"O�TBv�#�TMsWL�%*�y""Opi�lF� ��iX@¸og<i� "O̜�����e�,�g�X�Ex~�S"O���
^f�,��F��U>�x�"O��#&�E�]���1@��L-Pl �"O:���F>0nT�wO�V�\ј�"O��"qG�/H(�����\�G�\)Q7"O��i��Xnn��Q�9�Ʃ�Q"O���f�=܈%���Sz�X��"O��I�1s�H�k�d�S�"O$�	F��(0T������2����s"O$��R�5�+5T�x��"O>�Qq+>��q�*�"Z�1�"O�Qx�-+=�0ʋ��X,��"OnѺ�䊸f��I�Y��"O�X�JV�=p��V֞�a�"O�a�#�;oL-�k�\�<X{�"O��3���3
�G��u0"O�����W���EHt����W"Oy�RgX3R��eK�Q���"OBhժȻ2��'C��h�̓/�ڸ[��T�0��/�E\���;\<�ӑNӶ(,6�i��x��ȓh1Ib��<�hX���Ȣe�Ѕ�Ͱ�	�F�6�h��O".��`���%�F>
���Pbc��NCՄ�R}�A�˶+k4A�'V=���ȓO�t5q��S�B���瀺��Ѕȓ=@Hr�#8R�JUP���=W�)��f����U�f!@𛶣�]H��ȓY�.t�a)˕>��H��Q%[����_L};Se�;�@!�m �q�p��/���1�Q%E��`M��C2�E�ȓQR���KP5+����`�=;�)�ȓh	I���L�_���@�(��R���'�:4!p��()�Ya�u�Ȱ�ȓt)��ف%ѲC��AP�!R	���,[`G�s��)Q��(�lՇ��2�ܥ`�H���[�6�݆ȓ$n� J�mǚk�f9�t�?,�8M�ȓj�̕K��
#5��<��g��)��ل�|c����jE�`��S�f�E����ȓ/8���>asn}�T��S��ņ�aN��K1 �	E"��Ï�kT�a�ȓH��Y�	6�ƱC��ԮL�e��*�}�r��]����1OD o�f�ȓ,d"i��LTC,t�)�������_]�Ā'go��L!�+ͭ$f����sF�ظ�H+dNn�a�C+�����_���B�酡c���Ȓ@+��ćȓ}�&�� cQ�y��Po�9*��ȓ��0��B�q4�B�\�z���J��]�� ђ&AH�d���zGj5D���#�K.�y�7�7b��:V'(D�lQ@"�+o&��%"{�,��+D�� �a@'�+�0D��B�
ig���"O81�O�>T"�X��Ԭ_Y)�"O�T�SG��x�`*W֬@�"O6�q%��j�L�A�</ܰ�"O�4[��6�� gɥXpr!1V"O�A�J����73�����"O��0�$�Y�>����.xl��&"Oa 3���~�N5�Gʴ/����"O-�S�ŔN�Q�d��(btP8G"O�����)omZ�!�f^$:E�i2@"O��
��1;�f�3��A�Z'^[�"O
k���?Y+̸A�dX�}�	��"O�-��NŘa�-��C�S�!�S"OT=j�b-H�*IQ�s_~qc�"O�i�'�Z�v�u�iۤX� ��!"O�	�Pe\�m޼��u�U�?�J���"O�u�7c �|o�B��xE�F"O���o�a��A�P7U.Vt�"O�]�v&(���ꆢK&1�"O��dcG�+��	#��	` �K"Ol��)A�3��:t��V �i0"O|Ep�NR#��ͣw���p+�eȥ"O6`x�G�e1dP��ǂl���!6"O4is�L�L`%{��ܣW��0�d"O���˘^�p�r�N�<�`"O���� �)�ȸ+'
^g���"O ����#f~���iR�N��"O��A��;X`��P+�p��hY�"O����mI;�h�X���%����"OzD� �|^<B��1�\�A"OL(u,W
V�v���ٍ]���"O��#,�� ��7Ş��<�G"OZѳ�-Y d�`#�dc��Y"O���t��z9��+�CT���@"Or1�t*�N|���9%[���p"O��7�
�"l\�t 
G$�Ih�"O*�4'������� u�s�"O
0�2�\���Zr-�G�*@R�"Oq����DH���J��X�[�"O<�Ȕ`�a��]�"�7|��Yb"O�%�E��6+B<��l��/t�qc"Oj�x����1�F�F`�mh�"Or}z��5ga��rG$��l��jW"Oz��޲�"1���g�2,��"O^p��J�aX��;"� �7B�A3�"O,4�ʕ)�PD3 ��5%��A�"O��S�f�&}zX��7DN82��-�"Oh�r�W|b��qD�g�"�"O$U���\*���r "O�p2C��m��k�LQ�p��9��"OT������\1�Q��8��"O�	�;J�(��OBn�Q�2"O^t�3��_'(Q�6���
-�a"O洓�OR�����Li*���p"O�5�-P�O����a�F�	�5"O�����I�x��,�#T	4�i��"OX�bځf��SEK�Fݔ��"O�в�E�gp=FEV�p�T���"O8���`�^�Ic�F�E��#�"OJ��ǌL?W������,7� �"O��p"�+�u��TƆ��"Or��gj6Ly�"��\ݨ��"Or��R"M~���qs��}�"��"O�D`к{��m��j8?�|	��"O� �t�1��uXX�e�_�U��9�"OP|�%'�1+~��oּ4�"O�B�U�B)��+���}��zQ"ON@�猙0>G����ϕ�@d(�"O6�A'e��\i8�^�J��p��"O!i@�@x֨��EȁLv����"O�ISn��?<�p��O��%�"OT�@�֣#V�8#R���V��!�"O�|R�J��((��M��{���"O~$k��+el�5��kˇ|�H��"O�ux�F\3$F�3�+_�R��x�P"Oha���8��[CkM�i����"O����\�@�W� p[:<Qg"O���B,��=��c�K�f?,� �"O�š�=���y���f���ʰ"ODq�B��0,�\{Q�P4����d"O2�A��T%fQ�h�Rŕ�s@�zV"O�e�p� 16�u����C���hG"O$q�$!?�Ĵ�%�H�P��Ia�"O��w(5V���{ҦP��hÕ"OpA�C�T+�Di�S�7�h%��"O��K�#�s��(��[a"Ox)�'țI�:� ����B�߼3!�ͳ+��y�p��(HZ��u��xY!�d�>;�\�Q�,�p)�h�&�E!�DI�}߲,{��@<6��(w�p�!��'X��+1�ީ�,B�aYv!� ^�z}1	K���̺��כ5!�H�v�U3���s�4��Х�M!�Ă�{��l��:%��I�1�* !���WIj��$P<`��Qb��?�!�D��r�*�b�c>��S ���BV!�D7u��K LN#��$	��]�U5!�ց[䘹��:��@s�!�(!�X8$X[��*x��Z!�ñQe!�t����Ő�Ka��I��H�RZ!򄄨�l0��BGORR<�h�64<!�u��P!�\A3�xKT�Ŵ
'!�����FW3���
0!��G�����/�.G(T���-7�!��R� �B0�ҋQe�-�����b�!��Ƣ}NH!��܉.�x�XgH�E!��Bg�o���$/�|�ԙ��"Oԑ�
#`THY#��8��H��'�
v#ς.x��8w*8l����'�p �V��*���
�+�j���'��E�������B!ˣ ��<
�'������x���h�N��Ձ�'���#R+�j5���)R9,+>)�'RP Pf.hs3 �X�^���'���qp׺W�ѡ�,
%NN�e�'exhP-^�xx4�b%X�J{f���'�h	��d=z]�MWŗ;z�d��'��5zr �A^.ݚ�'Ց|$���'�����QDy�uQ5h��w��0�' |���C��;Q��F&��t�j�a�'�>U� ��"S�t*E�0�ԁ�'�8�Vc��M��Y��=	�j��'&��'ƛ�n����֡����
�'����U!V	z�}�g�D�	���	�'��<�ԧ�N�v=c�n	��b�;�'�.E�l��B�27����t��'U� R�j��2M:�����z�n���'�t�;G/�7t̝� O.%Y�!��� bl��iJ�$�XhY��5#�4��c"OF<�q-��}<��dØ�]/  *�"OnPy�N�<l�HQ��!M�n5Fc"OD�d�M�dĴ�e��LEm<D���b��B�N<��E��>�4��A.D�@zQ��z��G�[Ǥp�%�9D���a�Es�qR��8�E2��8D�4`E(�:z��'NS�pgv�c��)D�lB�b��k�F��#Q]� \:��(D�pz�jӜeB��A��ΎT$�Q�!D�,Ra&�8�~��@j�2D+��q� �?�O��0-�17� �����q�`䑀�'��B��<Ā�d�n���nY�0D(T$O�r�<ٔ& �4��u��͌aq��l̓A͚�[Q?��t��55Xx�'jL�f���q�)D�h3�A� 5�1�� �8Q�d�@4�1����$�C�J] ��
�`���P�M���tD{ʟ.T3G��S.,A3��X�}�H�"Oj���#P�h�:ِ��
:BH�r"Ony!ա�C]H,!�IS7,lyxg"O��D�ڡ7���X0����Cr���q0�O̒O�&�S�Zv�h���߶mL�����R3�B�I�`ƈ��%��OK^��3���"<	ϓ7Ԏ�)΅{�`���Aj�d���'Zd�&���E��z��Χ�")Ȕ-�I8B�ɦ`܄�2有t���wc�(�"��D"��,2��M�n�4��"F߈ZB��/�6Xچ$_*Qg��q句��C�I�zb�1��E�c|�I���X��C�		vx�:�Oͫx��hXW�֞��C䉡2[�q*
Р1[z8jƩY�>��C�!2Z,`{���<�M�Fjʊ&��C�SsV��f�x�h�b����Kv���3�o'"�p�?{�U��B.��d��EI�o�S֠m$B�@���&�@C���I�0R��=�5��5�	;��PCI!��~�N��7���I���sp�һB�O�q�牘-���xRK�=hgb��j� ?�d)�S�O�^딠O�aD��pI	jQJ��"O�m�'�ؕdn~�P�����:R_�|��t��9< 08�a.��+���ʐ����':a}�.�uM�q�ů��a|y�悍���'�ў�O�
�+4��\��Hdd/f�|���'���R*^&��xP�2iS���'TT��U�ߍ!�PPPD��^[48�'G���E��2o,�Ā֤	ĸ���xRQp�d!�HDD��y��ă�y"ëm����n��7�3���y�;$�z:���eB ��u#�$��'����)�� �2y��r�%.�$�����y3>��X!�V�y
�фdI+�y��Y%G$D�wi��
-�|�SH�<�y2�ǀk&�m8���6��� 	A��y2m � n1�2�Ȕ�V��7���yb ^;W2������yr�Z��yR� >lF@�۪f\	��[�y��W몰�!g�:a��P�`�+�y@W,Z��1�Ë�U� �p@߱���8�Z�����n���W�Y�RYL��M��>�J���V
V���=ɓC��k9�I8�0D�P�3�N i"��e��u�9��9��蟰� ve��Z8XEc�&W��B<O���d��N�H ''Q�%.��jǩ�!�UP����,�x%�P
��:�a||
� l�9P���n�6�T,K	\ˌ����:\OrpyU	@��*Ī$nƍ'��Ё�'a�|�O"���'D�=P�kR�*�21��"O��u'�3b���I4&�8Y���<!���*BT�`��w�|���꒰6��B��(h�2u9��Ġ%�����Ϗ
!�6m8�S��M�ARh4d2'CT�UJSW�W�<��ɧ4�f��̙�;��򧄉z�<	u��A�vq�&�<~��:�vX��Gy��1L��B�Q20I쨫T�@��y��N�Q� �+�̕��љ�M�J��F{���K�j#*����U7T���`ր�6�p>�J<�7"��X,8j%�<�l<�g@Jb��D{�S#?L��G��?��D[1I3��'�&	EyJ?U�.U��ڰ2�lU�_�4l�fB�>9��:�S�O'����Æ2N�xUj�K3�&8҉��)�Ic�D,� CF*�-z`1�a ;ω'K�|R��)��"�c�83�p�ǐ�ژ'tўD�I<1&-�F�tB����X
��f�<���Os��*��Ȅw���1�W_�'��'��|��r��ZTeKD-�� .�^�<��I�&
�+�>4����s'��<�J>�4�0|:'�ب7Dpɚ�,P9j(�(�b�px���?��#�)mI���s&LӲ��y���6�V1x`%$~��E�҄Љ���hO�x}��B��	`Ǐ$"���s�I��y"�S�fQid���! �:2����y��)�'����蚂O�>ݢSCg��8�ȓ2�0���X�0�g U
s�чȓa�����+D�"o�����}��ȓ	�\�ĢR%-�*H2a�\�P<X��)�ʑ�F噻9�V
�-�S�2�=ѝ'�ў�'i�� b�!�2Yn�y���3i�Єȓ DM R�C�KJf�{R��^��ȓ�	!��S!%"i����8[B���I��k�+V�:�`ҁL6%P��H<��V��G{�w��<1���ym���R�.m��Ó��'��d�\x5*���|���)D�h$�9�O0P�0�M�x����a�	zi,�U��$�<�{D��*��@�]��֍� ���u��=�gB[?n6�p��F^��'�ў"}z1mP�`�D�O˱;���;�ZS�<A���+f�8kD��D�Z��Tj�<�w(B����-���d�����n�<�ԭCB`H�@�C1$��*��i���0=1���0vS�Q�$�ϿE�.��r�_eH<Y"��m�`� 5�X���2��8,!�Ԡu���)Esن�*���E)���'��>�aL˟-��csL� -vZ�1��!D��:CϰC����� S�&��a� }�C��O,��|�L���Q���ߝ%ذ�����yҧ[
�BeI���;���7�B(�y^�D{2�;LO�%b��,�(`��"��t��P���'I�	)HJY���[�Hȸ ʐ(g�C�!CΔQ�4c�W��%AM�1�ZB�I�(B��h�g�����̴B9�B��#	�4�q�A��DI�HJ8o�B�I:a=�ݣ�F�$mV�`��ܪ#�C�	�|
8��n�/��E&ܓ&�C�	!V�$�#ǎeP������m��B�	�`�N���L�93�"��go -��B�Ie�@�tF��6������$b�C�I<�������5����q�ŮpB&B䉁^���� *#Yݎ��
D�0B�)� �d[�@ذ|�B�X���*N@
���"O�es�cT!{�i�0�ކ{W����"OD� 0@W�R���ff��uEb�`A"OРQ�B��}�:ჲĐ�3`���"O���l��1c��fJ@(�"O��4�O�%�L�tER�mX��[�"O
8�sC���a��d� fM�	�V"O��A��YT>�(RdFI�P"O��h&�O�\L��AF�\��U��"O�M����) Q�YP��C�"OR���#w�@��%D0):�iU"ODlƊ�����#��,��q1"ON�Z'@���.�%D�s�,e1"O|e��E�(l�Ru��aJl�`F"O�t�h� X*�(bB OQxp"O2��CE�{#Z���`�]U����"O4�P5�E2R6�p�fO�%5�,lP!"O,��b���6�Q��	a�Ѳ"O�h%-�s���������z�"O̴�A�Y�?|��Cퟘ[���V"O��Ra@�oT��E�4�f�rU"O��I�LD"i����ư5يP�"O��*2NIZX���lK�<�X���"O�]����$D{r�W�V��"O���R�0Y����±C����"O�Q��$��y�z����|�n��"O�K¦����P���7�� �"O�	+��=c�2a0�B@�r��u"O�Ӑ�s�|��E-`��*0"O�J��)a(\i��@���CA"O�H@��;u�����T[zh��"OF%�ۭ)��W�&/t���"ON���E�R�j�s�`8 [�
q"OB��lR�`g��2�O_=?���s�"OP�+[))�Va��.��}�
�P"O��i ��(mja!����,�l9B"O��U�Us$�Q�KS,1���Q"O�<�%Z#ƍ�E
�#u�*���"O�u:����i��yWG 	� ��"OX�����S�DĈ?k(�AP"Ov\YFMy y�棕;~�tUB�"O��*M[�Bu:���ġk�"O��Cp�K�>�]/!���Ӣ�+�y�l]�F�̓@� ���jp,B��y�A�/A���6K�G�Z��F��yrG�X�^YI��I-="���5&�>�yr'�.�Q�H=xthxtC�:�yr��3A437�0��\b��]"HX$AI��tn-sè��0=��Ot���BM��%���b�<�PE��{ga6�q�P�	CXA�<1 �[(�P�ehJD�h�����`�<�c�[�7��]ç�܌O�h�F�b�<����10��Q��4�1�r��D�<��	 =	Fa�4�A�(i@��� _�<�˾^�PQ#��-z�h�P�<ɂ���c���+���DHY�3i�<�L��	O�cf�3�ư���O`�<aC*D����	@&W��IZ ��J�<qF$��'kZ�e��NVi�<����xf ��h����<�OR�<�ꑨ4���ꅖ*G|�y�a�<�F��$���0i[48�&�v�<!W��'�����K9]��Y�hA{�<q����[�h��R�
.~���ΜX�<� ~U�����/��$+Q.N�0��"O��0�_< �.�B�l�p���"O�zQ�ֽ7N��9@j��>����G"O�0�b͋�1��$��	�H8��"O2����./��i4�>X���{w"O�A1�(F9H��3AߪW�n�{C"O�1����1)ц\�<hk�"OtIä� `Cb�5U���"O�b�H rƱ��!�(%]>�$"O�Dꆂ(0}�XA�덞E-���"O�{e��!-�x{�$�[��P��V�q> \�g�	O�r�|:!DX|��d,�#Tڼ�Pm�p�<�%	Ί�줳beȵ��aU
2��'�HiQ�𙟈 &��1(m��c��U�c��"4����	ͳv<��U���4~�b�L$(��0��{)�Dz3AJ�%�n����ϲ*�PF}��ɤ6��J��&�S-Px1 ���o�0���2b��B�	�G(�h���Q�P6�C�lC�牉G���8��	g��S�O�0aō�o��ĸA���H1*�'�Z0�O<z������rhQH/O�*�B|sVЉe=Op���c�-�����7M����P�'�����M�M7�QJ2&������0c]�@|\�r�M��&a!��R�'���rT��*x�28�gk��yў��$�ȴt���ªļp�"�)��@3��bg�ѯG���ȓi1�,�b��u�4=��J/9�e�I-q>](�� +~�������TsW%��2~�x�p�ٹ
�\�HT�4D��C�j��`̶ɓ�O�h(����<�v��=c ��$Ǟ�0<a֦B�Jz�m��.�1}sR��R��jx���2�[(cg><���^� ���˖i���A��(��=��qڐP�D�GN��ӭ�1d���G{��7'S�i�#�1�b��%�V�X![���"x�P\�"O*�C��:tЄ����B�+q�5Y�1O<�cW�X9L ��ڴ'�>XH��	��X����R��&"��8��I�E�!��w�z����v��'ͮK���IO��Mk�B[�@���t���\��x�g�P%��Y1aV�4�!���|�iڞ.V�)s��7}"� ^���q�,��Q{���!YB�t0����8����(6V�y��OEU�.X	��B�K��]/�@U"O�ѡ���<�N���	ճ$rf����	�?�dśs��$�3���;J	���PCȦ|@JC�I5�tL�.����F�ܾR��\��I��}��E��O�yR
ck\@�Ҽ�ިSOH�Z#�9A�$rpN�X�8%���I�w5�Ź#d�"��>�/I6`*���l�K=�!�cRfX�P��M�u�vpS4\��*���O^�@�E�$
n�Pą3D�p�cCF�y��Ա�k՗'���X�3��׫,G`�y1�P&���j")��(�����"O�]Y�o~�>eW�

�M�� YF���'��B� �3��@�UPeaH��(h�D+!�A�%�xJ7E�����4I��%�w@"��R��Lx��r3�k��@��7%�(��Х;,O��!"�,i@�E:)ON=�b.��-Ԩ�S��5A�@u��"O�HI��Wj��$
	UkQ�B�xɔ8��,��VŞ<�����v>����?Cp<���d;��0��2$����B��kFP�	��d-��8R�@6E*�5�N<aQ$F m�P�c�{c��F-�!��(ר]�x�XDG�K�\�fD��0<	�k�;��T��" 1!&���.J��#�Z��xԹ1.����T�P	=1�E��]���"��A"�ذF�~�'Ј�/ׄ(�0�*��,WV�x.OL�X�$�+Bk�LAaCY�0f��S
5N����~bQ�K��lu!�#­��11
�Ǵ�2A��w62�� �'���#��)��P��7 �NI�P��A�V��QN }Zh3"	T����G�2�YM�'V�,�۴[F*�鳈�,�e����ܞ��I3}��H��������U(��W2|���h1.�0�Z�^�&�[%���=����cC�
���I*;�yg(�?�t��k����tf�B�4	�;�L5T$���Jm$���dJ�F��	�#ūR���ړ��4Lx��A8:~h�b�Mި;��Y��'��͡�+�i����)� ���3K�:����Y�Jqf�(q�O�Uڶ�0�jyڣ�ƋM��%i�'j�R�AK~B��G0c-P���/ �0#c'�BNr,S&���*���2�I3lOޅ�!��C�L�5Ä,0r� 3�\j��kDA�Z:V������6x�S�Vf�ha��Y=��i�i^��:��C73�]A&	]����m�8eick�Ia���4!�;�D���U'���Fn�lc�Ō%ߪ�Xg��D2���Z�$�6�F�=I=�'7j*�xW�R�4�P	�B��R��hF}��Rt:� C�T�^)�4u�%1f2Ѡa�
b���� ?Mk	2D(Fм8�+�Zy2�P�>|D���L��IQ�ƚ*BP[��4q�
�I�ͦ��HAB�8x������L�m3ʸ���L+���w��y{��	�,�(dɒ	�p���.J����%ɺ���΢r������"�$�B	��a6�0�a'�[4B2A-$���K����Z9@4%�'Ʊ{fGė);��ʦl� Fjl����66�#W�*H��J`�P�$���;ca
���,����8�H�u�ڤF� �I�Fj���|�p�,�]�XРS�4.� �E~���2d˨�*dbF�x��yag��=�`�;"M=b]���'n� �U��8!��4g峟��G�<]��Y	a'�jCC��<7���adl�*����c�;qW񟂝�A!�1DS�Ż�SdE��	"O���ׅt����g�^,�i��ک�M��.�t�JT�`D�<�X��Hb��r�C$� ���ţiD\��f5�OR�B�邹)�F)25�߿<\:\�d� �cd�ˢ��#��R'���Nv�)�)�e��C�	2TTH���/q�џ��6OD!�D%x��d�WPj��yt�s�DQ�IuE� ��dɣ�>�T���9�� $+����M����1�'�����/F4hmT��OQ>���oʶV��\��I����p�/|�DS�O
�O�2��$�9Ovr5�AMČ�,�`�҉!��O�ua�A��=L�'4p��b�B�J t�̓xUDA�$�,h�(����x�꽄�I�zSTiS��45G���2
F�P�e�8d�YsST�4h��E9+�ڭp��:?�|����}a���"G)a�������x�'.�q ������&>)1Щ�h�K���,(��C�t݂0���5n5�IL�#|�'uJ��#�ϢuB�%�5�F��|�@�O�dk�˔� ��O>���*J��	#�s�V����]�d�����b2�|r��P��<8�CY��� I%׸'y\I����k�� ����Y>q�����B�����g��U\�-Qe0D��9���(M�DE��K`���G�.r�`�9#����h�X�#�#���Q3�$P�40 �'����\��:I����N�^�q��^�wQq��nSh]��D�>���O�ȈE�S�)w�J	n6%Q՘��!NJ�&h&��|�5�:@f�${U��!Y�� ��l�O�3�FʰR�d��E�E
��^�(��!�w{��A��>I�O�(��!pK~Z毄�.��	H�(}Ӽ�ô�/oi^�� ��5Ox��'S�Ѓ"Q!dƂA���T�	N�� +�=��T�dY�U4l1��p�Ocl5���=��\;���:NHf�X��D�0q���\;��'��V.��+B��jġm��x�`@Kl�F��>���Op��DN1.Pq6���Oztt!WW��h�!٣6*���>E���Z����{0N֙5�8Pc=�?ɱO���p�ia>lO��5�N�Kޚ��+����s��O�DL�#\�A��.�i�!Z�]�񧎒�MkX(0�%d���1���L@��Ha�*8��Y��A�`��4��(N�=Г��l�'?�=R���<i�ɧ��Zm���1�$�b�*b��$	�џ�jB!`�`�����4i�:��P�R��8uW`I)��WM�$9��l������b��-WDD��.L�c�@��k����ݘj�P�p6���i�\�$>�`���3s��؁��J�:� 7�;D����CĊ3���c&"��|[�p9�	�~\��p+9��
)�x��'	R1�����w�]	�"O���ԅK��F@����DV�Z�H�<͸'�h�(����	Fώ����?�H@,D�� D�� x
�  b���p�Z��F/��C/�!���'�=���H��!C�� �rʈQ�	�Gㄍ`*}2g�7L.e��A�bOZ9[�,ɓ�y��F0{���$Լ_z�=4AT/�'x�!#D��o�Şu�B�*bL/(�X*���yS���2����t���)�.��قEo�q;C��?�(���L��'��v��I1u 3<GjC�I�\�T$�b/Mi�����(OB�C�ɑlq��FY�d���CXJC�)� ΁��KGYN���j�('[
y��"O�Y�צ��
*�S蟿(r݊A"OF����<�c��6 {�Qa�"O�}�$D�8G�mBH�j���r"O�t�'��b�4���w"O��JS�G�{�����<%�L
2"O@�C���ư�À ��t��"OjPK��<<�eɒ�P�^ �IY�"O�*�ᑯ�fqrBL�Yp�	"O�d	0��N�H��	چl
��C�"O�a���;O�Z�H�'=���"O�uf�B�&������ZI$D�#"O��T�&��逇�ˤr`I�"Oڑ�T�\�7���"�^5Q�\�"O���h�'�0|�F��F�H��"O�1
���~���)��Ɣ��i�"O��Ɇ��<:���br��8m<8���"O���t!Xx��y�����fI�E"O�e�1�,H���geܖ�䨪"O���Ɩa^��X��ǮvW$<�"O�� `��\J�)�ߐDjp�%;D�p����f�I@�ߡ% ����F�r�<a��E�_�<���M�)%D���C�V�<��J�~9~\�Ճ+a��M�i�<	Ī�3K�����)�v��!Gi�<Y���@[Z�0�$��k�p�k�/k�<9ǥۛY�����D�C�28�7&�a�<�@��N�~%hU�T+a�d��'{�<9 υ2s�.A�d��P]�H���j�<��EҠG�>�1*V'}�`$��C�<Y���#E�0�	V�X�$]e�<�3#�	D�j�R���&�h�f�z�<��A�
2ȕ�T�)��q��w�<����DN�Ȣ(	+Y��A$jUq�<y�R��L  ��-rF�y�  `�<qaJ�,EU�yI�
�(S�a�t�DX�<��Z�ꔩu	Ħٮ����GW�<I��	�hsn�p��' i�AJEK[�<QpOX?t��e1�����*��L�<!�%�ob�ȱ��:D:DSC�<a�� ;j0�bm
o��ic��`�<ɀaN(VJ�)�
F�`��@��^�<AUG0q�H)P:~���P�_�<��s��{�k�5�hX@G�S�<!���@Y�1h���1K=���)
c�<��g�(۴dHe	�:6d��3�IQ�<��.@ }0���6NX0r�޼{���M�<�,̩g~$�;�F\�X�����KI�<	ċ��
�HEiS�1m@&� ��A�<ai˻k�DXJr���)ԀAH0�Y�<ф�́�H��f$طZ%��c� P�<yS���3��<1�J܄j�ds��h�<�VG����LЁ@��A�DH�<q$AS/O&�������#:*m��E�E�<Yai�#�t�0�>��e	���G�<�Եm�R�I��Ay5ta*QkV@�<��U�'?�Ea��oǸ2�l�~�<�Ӎ5,�����e��\-�q��t�<����fj�7l\@�b����Z�<����R�jP:'"֐>Ŧ���x�<�G�V}��SS/Jr��� (�m�<�F��2pF�8#2�B�@�P���e�<�⑘_� ��ի�,X�0��c�<Q�	&>b!j�B03c�� �Z�<� ��WÆ�(`��A�+ؐu��`8Q"OL���.� (ISo݇N��<`"On��N�DJ
�Ju��i�$P"OB�����N�v�&��9^� p�"O���Ԫ�/W�z��$둖yv�Ҷ"O"�3��5Q7b�"@
C�?nޔ�"O�a�nE�j�ǹ�_&���"O��R�bT�sn03�(Q:�1r"O��!Dk�c[V@�'�U��]�"Ox\�%TN�$�1#^��½��"O`���B'5������R���"O��GJ�|4�B��p���R�"O�`)�G�p`T`��)X$e���r"Ox���CA>g�l���h�.�9��"O��RC%5� P�f�'�f��"Ol�N�6@`���I�rx1�"O��2�"�l�ȭ��RV\��4"On,���KT�t�$�G,�"��"O�IC�'�M\xJb��n��$ �"OJ4�'N^4�9�& G��6�	3x��90��Z�'M���І"ת?$Y��Ξ'a��|��e*p�/I����FK��z
��̓m�P�)ۏc��ӧ��f�i  �-�~�*�ZF,�
"O��@$ٖ�3����M�!AC^�`K��A(��DMy� !"D��e^���m�#9=p��<�O-@g��'H�r7�8	`Xf� �D\ ��`�],t�C�	*e~ș�ʈ ��`�/lV��=iҪY�~��R�B���O�|x�ԟc����SK��[��!k�'{�i�GY%N����F�^�<��z!�}�D�K3?�`�-O?�#�\
w$Y��� ~m��2ׯW\�<�d�/�=zT�>Lm�@	�]Zy�H�<�(���e�ukax�ė�oB�b�k�⁅ߙ��>��EߛQDh!� ���QS2N�>Z 5jP�	�y�	�'��j� ��_=0��d�N�s�D ���C*��5pW׎-8c>���!8	��$�e�@�����2D�| `d�B�J��B΁uY�ՊcJn��0�
s.�H��>E��J�+!p)"O]# *�1(@Ϛ��y�  s��!�f��3����n]���3=eБ�'ΝzX��8��V�0ͤ黅�Q80`��R�7D�L2��I �4�9wX�P#ی�!�䇃#��9*3�ԯt�QG� �!�DC!3�b|��k(jQ^���V�5�!�$֞W��j�J70n��Ȣ�[� �!��'v�(�d��� T^�)���:�!��ܮ�������/U� w�Y���{�쀇���Iغ�(�)�f���DA $�C�	-�B�y�"�:;	�(Q��R7�`9�r��e*֭��	�6��	SG�O�h��sf�����4���GL���\A���(�L�>.8�:0e�:&!�X<�B��&�׿2���ڣ�Z4Y�'g����l�,G��M���B�S���1SK�yҢ��IB�)bq�Hh�4�h�<!�>y��Q*���'���0���4b@��@=20��'4F�؀��-��L�e�-{gҰ0�Q�t�,�2�Odx� �w�&r߀Չ���<.�`��,,O����fKV���-O����KsCx2��$j�h5�"On؊���+�T�x�(�6�l����x���i0�e�GM̧m8�R%gg>1��@B�9Q�=Z��L+#O�:'- D�̊t���B��)�q'G�wn�� �Krh�O�Xdk� [����u�`�iąP�
<N�3ӯ[�e��6E>�O�i�kZ��?)�o�#̋�.�5X\�h��1}�� ��:�����;3`ȅ������8bs*l9�d_!K�FdɅ ɴ^J� ���	0s��P���C�p�؂�~z� Y�>5�db��t��D���O'�Q�3c�$3� )kw�'�5���:W� ����ےH������"~�[uJ�\ݼ��t���T�3��a��{��eo:� ����B�6UX�3s��'�Xp#�"O�yb l _�z�0��߾[���K��'�^���'���ӥ+\>a��I2pLa?a�ϟ,X��!��:�2�HtM�>j���W��'KM��	�{<r��9�<�0."D�PQ{�#+2�L%ϝ6�2"�J�4E>�$�z�D�!7)1��>���)^�,u�$nO=Z�L����|��h���GmеQ��q��ܟ��'S#�x���Q:X�Q`�L�+h,i�d�
�	���e�u� ��D	�B�$H�F�<�y'�%wx�\{�A�Z� t�Bu��W>}i���5	f�US1	���4��ّ�bB�+P�dz�i�/a��ȓg�(|Yg��z��ACާ�6�I�w@Z���O�3;�eڱ� e� |q�O����oR�P�4zЮ�a��qE�xjA�R�3����R���	� H��ȳ��-��"�\�t��3�K�)���+ƾ@���*��DJ�v���;bh*��>��c� R���#��9>b�3��K~��!wv��wn�<t��ċ�~t��)���f|#4@KT��pE��
�KR�67ބ�2�C�F�����4� ��N�;�N��Ѭ0&=��Z�H��?���m��dS��~jR�ک������5B�< ���Ʃ�/9,��I���Q�ڗ,jdMD����d����e�B�P�D�Tܡ笐,Jt��DǊV̀�ࣁO�� W�?Y�џPsn�� 2(=�"D	e�h=���:���Cד$̠�6F�^����OV9�B�/WB3�H���ӧY�T!u�U�J$&h�i��eb��*�����ֶ�`��Ԋ��0��I7"O(}�ǜ*"�!_	��$3"O�H���H�F���4N1%�P�%?��<�����Z�8y��=� �*��\������Y���;2M@�z���R�b�"B"D����!���`��x ��/��S��|m;6�=|F���6HN�?�$�?��X
q��1�V�:���g�޹�$o%rT�|��Hׄ��%Pv]�M��	.$#|�'�N�4�	DYKT�(:9�Ny��K�+%��(���N��S�h?�-�bi\�:�*Ưq~�VcZ *���5�#�O(1��F6`��Sa`�j���,�S����2>��3��9:R,ĂFoh�����<�qF�4�<A��
J/�m�EOv��h�� W:Z@���;|���퉟$�$�#��z�	�kE�!�!�+"��Ş�(��B��0�_�Fg����0��E��(�TC%|c������'j%"�܆S��rf��9d� �P��\㕌1�g~2�āy�M�#�ݜ`L)�b�;��d��;��r��>���:����M�)wxѱf��0��`�c��
�J�Z�'ے�bwfA, lh8�G�z�R%��{�OĽy�M%�` �_�y���6bX��`%��	�4�`A8i_�B�ɕ1�`4kQ�W6>Z���� �#<�5���bf��h�R�r���6E���a�/+|�Q�'�}���O̓?����"�Syʡ��ɐ$'6q�n߹,��+��>���O�(�"d�H��0���}\�����xD�F�/��p'�"|�`��+���p�(�?O
���ߟ����r����'�<  Ag�&^%Y���p;(a��#}�bK�8�xL �����=�`|P��ǦA�3Ƈ�H:�
����:����֭>�O�Q�����"�m p�I�Xy[���,+���z�/���[Q�[5$�5�h�&D+Q+&P4�T`QJB�`�����-Z�T�`������Om��zdM�%r萤��Ջ"���&H�A�|u�N)}"��A�Əh����#}�TPK��<Q��Zj���km)}��)��?`�	�@�ֆݮ�릀(D"f�xE�m�y؞���Fu�ܨ��mX4`jD��0��I0j���H�O�Y�0k�̤pҏ�b?��k�q}-�e瘆^�e:5c����?���t��a�L:q~�I�i��A�MA2^R�O�9���^�&��O�4D�x8�^���%��/�@)ڢ?I�AL�y��Ӷ�>�)U�di�t�!È�)��2EA�}R�Z��Η3qO?��9$yt��Q��	Z�my ��-Q�I��l5�b \�)�'I������
�Tƒ�ڠ���L�ȓX����� ��C�~���݉Y�ʩ�=�֮D,N������9X���0
�]S�J}v�!�"O�:���@�Z%q�.�@��U��"O�m�[=���KQ�,��@�w"O*5�u�	-��Z񦖳�@4s�"O|@Z%�W ��M+����"E��
3"OR�$l�_s�hW�S8@F�S"OƱ�w�$tZ�ڤ¦N�%(�"O� �Я"~A�7�\� W"O� ���V,ѱO��)[�.�;}f��"O`�J�A1kD�a��"�*yh$"O��)��W!,`�#ҡly�t��"O~|���R8B}^
EK�V�!""OR��'g���N�XEcҍq'��P�"O�40BD��Y��b�/��P`4"O���h�$�˵m�a�ߪZW!��Z��ԓ&�U�.���ҊH!�� Ffl�AS%g��T3`	�@A!��9�ά�" [�8X"V���8?!�D�6^���;5I�>-���d!�d�6c��S�Y�C�HT� ��	'!��P�� 3@M�z����3L�!�Պ.�Pa�#L��N&@A`�T,�!��%b��E`��,y���RVo��F�!��*$��P��8H�
=ʳH�`�!�d�7rZ��ȱ��)v�$i����X�!�d�D����#r>P+�&�h�!�$W�z�F��U�[�z���ː	�!��ܮ�Vx����4��qyp)�!���@�X���h���[v�����',�$�����l���ş� �pT�'(#��ųtd<�d& �`��*�'$dzGC�.E��-#3fJ�s:*�'	�hq��Г^0(}P��C�� ��
�'�F�:wd�o�La�i�}���Z�'R����)�S*�=�"O�js�;
�'.��[d�
�bx�S�m=�*�'�8S�	���1 �DB8dz&S�'5@�����(�Vu�$AZ�_:~��'�]aQ&J�o-��!��6XJ Q��'��l�t�ÉT!Q�M��'z���e�����QG�*Jr|uP�' ��&*Z�V�d݂��6�
�P�'�ȑ�J�Z{����^��%S
�'Z�r�EJx|swᔚ<ڔ,K�'��8���OH$��i�(�LA�'����Vg�a�J���H�X閱�'�j8��I0y�dE��lW�Q�0<(�'P~ԩGAN+Pv���"�
�b����'V�0�l^��`�b��"F���'ٰ��%�H�E�mS$Z���H�'�b�#dR�$[j�s�&̽Q�D�*�'��S��*9�J�+���+�'u��oY�i�vZCcT����0�'��MK��O��4Yz�.@!Iv�i�'�����+�$�"J^�N @D�'�RYY"]�W*E*1��:�Z���'�4�RE��6Z$$z�D .;�@h��'��p���~|8	p�Q�o���'Dj���5k�FaZ��ʎ�E�'�=�1�"���7b܇L�0���'X��S+�a�g�,�����'6��:�eN���d�&�ޱ}�B�i�'�"�FLc�p`#�'v����'�h	��H�/1r=��gI�X�i@pO�	�8����(s���{r+HԦ	��Od��	R�
��Q0�ē�����O�Q ߴ���b?I�!T�o����^�~���A�>��)ҧ=%$�B�JޘODzU`�J*RŸPn���T���ӎ&�����$Ӫi�@0 �ؠA��OD��Fwq�L)&X>�T��N�8��@� #t՚��<��C�
6��t��%<̐E���5Y:�/�5rP�$4?!.xQs1����_�4KF��|�����7�}CD&D�X��P�ǁ�M)O(��O��'����J�B���	Q�b�m�G�����T�i��I�>��4���0��g�? ��ъG=r
l��de�=3A�q�Z��[p�O%+r��k�'��'8��k�9X�؀�U��.`9nZ�W3b�'�n�Ӻ�O�2'8���Ҥ,0���à�'�$8&��G{��t	�P�1%�-n���q���$4�S�O���B���-@LEC�ǚ��8a����hOQ?�X��C�b�H�����9���'��0|*GX9
}Z�+�=���0��]J���hO�'n��p�$�%Ku I�@�?f$I$��2�.�S�'	�P�) �|�<�WC2$q�'A������E�j\�a�N6~ ���՘l�7mK6��?ah�/�⺻��F	+���U��#�.��dj;[��'�,��tJK{��6�S�][�4�&��4J�bظ��;P~ڑХ���?��������t��i�m3�#ɝL���%�Q�*g�6/��C8���4�Z��~b�x�!�?�O,#"��RY�=��)�=���Í}r�!q��O�OR�X��Î:���a�%�7z���#M<�ӈ�����O�00�J�t?��ӊ�&n�}c�OZ���(-�)ҧ`�d�cŃ�;�vY�M�)K̪Xo�ly�|���?g�*�	�r,lp#DC��`\hB�	�0_P0�����H2�abUtaRB�	g��+q�Q�@��j"F�)I.B�I~�l�� ӂ4�rՂ�|�$B�I�q�g��3*�U�@,F�0C�	�qA:X���d�p��A��wC�	�a}Z��)E-�
�x4��GuPC�ɘ}R�U�&�?��f!ϥ�lC�,$�h��bc��AJˑ��C�	$o���b�ՠD���
�lC��2F�Y3��V�'+� !��H�$؈C�ɟ�zT��LB�@�\KvbǑqOLC���h��r/��`	��1I��y�VB䉎C�d�A����`"����M�4B�8O���D/�$��`àRQ8C�	9�Fp����$	O�](�߰J( C�ɎJ�V�b�F�?��($�ɍ;(B䉿4�0�nݔ7%8e��*]�QNB�ɝ �ua���:�]����G�.B�	�}R��eF�=�0J׊��q�
B䉩^��R��	G��ӅI��C�I�P�IZa�mb,�3����C䉌3�l��cȸP��h� E��0�"B��'�>����-K:��Zh�
$,C䉉:�R�� �Ă@�Q�Ë�;KC�	�r*|Ɂ�)��������}�B�,U�L�^oȤm�F����C�I����!���д3�)Kx#�C��8X,��C��M�6��H>�~B�+;��1��y��*+ޟJMC�&WS�%0a�[N�<ЁE�ў\�B�ɝ2�~M�.ɽk����D9��B䉛uy��"q)yR LH"A�R�rC�ɉf�lM��lCy����3�rC�	:/�`�r5�A�.)��.��i�C䉣��e��&�e��#!L�0C�	2RȚ�Qc��?�6PR@���W�*C�	�_����d�ܣj`�Y��/�S�^C�x����р�E&�T��g���"C�	k�x�
��ٝ�0���	�bC�ɔ,��d���qɮ���#��5�B��h��� ��V�C�0Ac��f�B�	�*�Yt���N�Q��Ow`tB�ɧ[�HA�6�a���
��M�|C䉚-��թ�-A	zxx�����cf�B�IQ�����A3hPx	@I%�B�	�}���&W��ш��/�ZB�)� �"��*��e�p)G$���*O��[)��12�"� ��i�'�޵
1��3b� ����E.`C���
�'�%��j�4:"�E��ބ]V�0)
�'�X�AW���'@��r�X��	#�'Ś$���D�d3g`[�c�q��'�B$a�lؘ(���1�a�"��'��[G��B�d��Ѥ��V�ވ��'� �[E��^68�c��� "�KPm�<I����1�C �3�\d�/+�!�d�^^5���*b=.����6�!��B+:+ZTۇ.�]G��b���Ld!�JAF����8!7Z���ϑ2�!�$),�q�7;�P��G�d�!�ĉ�@X���M$���Y�w!�S$[x���K�M氬��k^9,�!�Ĕ�O��р����}��,��O !���6Gj5���4‑�e��<�!��ۗ�t)�d�<�6�%��w�!��M�`��G������E�j�!�4y���Tͅ�$=S�'�s�!��FT�a�ĸ32@���4�!�d�5�Q�@Sr����+W�!���8�Α�s
]�up$UѤ��7o!�è�� �*�#6gJ��e&��`b!�N?��0c� 9?N@�քȔ+!�D�9T7z=���i5�ݨ@��#v!�X��2  ���e��Q�\!���#x<�����eC�*�!��P(���@��4S�pIBt���!�ğ!'���2�JPS��x�R��!�dM�T�f��`�V���n��z�!�$ݘ8�`�!L^�oJ�� �Ǐd�!�dS�n �U�bJ�e��S"Ds!�dĤ ׌ih�(�,1����I3!�D�	6M��/J+Kl��#/�!��E�
ތ ��ȓDA�c�-��A�!���|tC��ܲPP��r�˝$Os!�č
Q�`��&&?l�\#�A�'�!�Q Z��e4�D�yo��д�>!���}R� ��3'A,`J���!�D=	D���%}(����V'7�!�䝡^�X�����9��R ^<@!�dA�a9D1; hN)�u@Q�B�x�!��ϓ_󆠻dZ�;꘱1ӎ۱R�!�D��I�s�Ml��Qc��
�!�H*�$��)(�>��$aݲ�!��Ȗ3S�iv�U��l+�Mć|�!�$qS�(����/C�x��&J]�Z�!�$ջ�(��@a�V�&C���!��~ffH�3�:��ۆ�ڿW!�DB�b��xP��N�m�hl�H?>�!��B!H�1Y&���C�@<d��K�!��V�Z�K�
+L��|[�O�!��ϝ.cJ�*��.*�8`�A�n�!�B3.�:�X�M���JQqr]%g�!���`.~PQ0� ����S�B!
�!��\$%8�����^^�T""�� �!�L.��E�g�T 0^&p!� ���!��H<��y��pJ�,{�`�6�!���	q���c�F-n��}㕎2!�).�l�kUDD�p����([�Z!�d�&P��u��]�<�v��ɝb�!��"u�b̐��t11P��X�!�� &����,��X`���ij�lJ�"OZ�R�`�'n�xT͒�XFa�&"Ob�X�E�=����D�T^�ц"OD��7O_�F�<���޿s[�b�"Oꉲ �K�*�l�Z�(Q�"O0�!p�V /����"��n�^���"O]r��5y����<^�h["O6%A�ݟnq<�S���O���"O�y�4���;�^��ݼe�*���"O�ɰp!�7�%��F��U�ny�W"O�k��ϊze�(��+ �\�,�86"O�ѐ�KrPD,)E���2�]!S"O����7{�R���N ��D�#"O��s�DfQ��A.b�����"O��1 D��W^���6�[+����"O�E`$�T�k�<���Kl��
3"OJ8��.3����̉	2R���"O���Օ�^�I�ɴx�d$6"O�$�n��o�$a)�C��k�v���"O�X1��P���I�@� �&(Ad"Ojb�DA!R��8��ƕI�&�j2"O��r
��e���Y���,v�H)"O��;��+p��͊S [�@�>�`"O�h�S��?�(����.a����"O@	��e.e���[p@گa�$q��"O�������$��I�s@@�"�X�"O�����Ԗv�������'�4H�"O"�	"[����T�ޢ|) p0d"O�8@��E"��U���F0\*�"O,���Ë>s���.�O�9��"O>�h�N���`�)���@"Od�Y5I��&�L\cbE�]!�]q�"O`����>]^�`��
��P��;D"O��#��F
�0�����F���ۂ"OH�ZGJAT� �P� +X�BX�"O`�������Q8bn���Щ�"O���"դN��A4��1Y�й "O@�����v1�E��W��(�"O��4f[�kϬ)��hC�)��E"O�|�p�9#�[ta��)|ȅi!"O��a�ڂi�P�qn]/pJ�{"Oʹ��A�Wb��
��Hn����"OB�:�F�=bԉc�
@�*�,	"O�����s�2���[�h��*d"OH���S�k��5���ʁ�hA�S"O^���eE�%2��w��c�}#"O��%�ש<&��v�U�e� p�"O%AdÝ ��E#s�!g��r�"Ob1�b��>[^�j�DL&b��(9�"O���E+�]X�HP3�@�&���Z�"O��)҉b`IX��!*�M�b"ORtp�/�#t����a��
����S"O $Ab�΀#\X��嘷�`-"�"Oh��ș�wwn�*G��3c�B�3 "O�z(�}�*��mR#k�dE:�"OYSjC�l�*ȃ��/5y��x�"O��+��[�o<��ҫADΜ�T"O�h��M�<�f	aA:-(�"O�}1��<.��iPV��N����"OP4i��
v|� �F�u����"O�����g�Թ��i%��bd"O��!H�wh��X�g��#D  �"O"�K��0S�,Y���_2|�:�"O��
��� ����g�A��p�&"O� �����=鈱*7d	@��"O�3�W�,}�����T��,���"OȄ�ceً%�` ��rbę3"O�yӐ�Ȭ��D��`ȍ
�2�#"O��K&	��;�� ��D�����"O��@�f�ô��dAX��,͠�"O��@�P Xʂ�t�2�W"O\8���\2\`��p��ĤZWd���"Of�br�K�|e ��'MT�)�"OZE��I,��5	�$0�Ba"Oip���0.�ج)�ڞ@�dAK"O��5�Ț;�{bf��|�z9�V"O��KFJ[-o_�4C�C�5dp�K&"Ov�C�A�8�Ш�0	U���tj$"O�e��� CZ��a��/�1*�"O�#������:&'�Z+rY�u"O��p�)J�Xr@�	$m�LJ�"O$} ���:3l@+�N^�Z���"O�@�I=:��(��m�z���"O܄�!�\*i?��@F -��� �"O� Z�.=
$.Wn)�&I�s"O��8$   ��   ?  P  h#  �.  �8  �C  P  �[  Zf  �o  4y  _�  ��  ٕ  ��  ۤ  (�  k�  ��  ��  K�  ��  ��  �  c�  ��  ��  4�  u�  ��  � @	 � � H # I) �/ K6 �< GH Q �W Bb {j �r 6y } �� _�  `� u�	����Zv�B�'lj\�0bKz+��D�/c�2T8���	#Ĵ�ƧИ�?Y�� ��y��%+�Y�b@9�J�G�V�A�̸U�$E�A��Oɴ#�t��MI?g��Na��	�0#���� ��1��R�E�6�@�]�$>`[l��0�5`�aKf(�P�R�%!�L��H� ���'u��6��+bXe�fN�X,|���$+���Sf�n���3^Z`�E���~�mN�A�I����Iҟ��I1@�9PcF
�=�&& �9a�=�SñJ���a��������?A��?
M���ٟ���Wi���ANP
2.$��k������Ɵ�$���IƟ���b=K`z�Ґ��EL��Id`_�3�^��&�<oP�x�� ��I�~ՠ����D�?n�}�E!�EvL��(��iA���rG�>��'��ON��H�&_2E�"�b��١���05 �����1���O0���O����Ob���O���|��w!���diU�/��IK���%5zhh�8����y��Yn3�M���
��f�[h(T7�˪�M�0�ޒZ�,k���a����p��$^�mZџ8����H�a���6*��Q�h�#����צ}y��w�z���GכHG�uِ/G?5v�0��
�N}���q�SZ����_��V�o�2�� �|����u7-�3z�~��G,ץ.uļc���gқF�۽F�śT��w:��wd�٦q���N�O�z�m�(�M{�iL�]#0���>��P$�
�>EB�� 𭘐̃�= 7M��1�޴q�HL��!D�j�^T��Ƀ2�: ��Ȝ�$�t|��/��]�� 	�(��a�p����\'/��1o�iI7m��o��|˔b��H�G-��hD��JM�Ӌ
02�Űa&U�NEd9���t�:PAF��,2<�*���,3�Δڳ��O��(S���@��P*��F1�P05�@�)��4$tR�'tN7m�D�It�`<��)�غ��'��m2���	\&⸲��Hp��=��'y"�]�=vr�'N���h����p�B�B�X7�D�{��xsbI�N��1fk�Rhb��d�)O2��s�K*h�NDk@mk�N�!O��[߶�5���Yj蘙�˓K����)p剩���Y��ha�F�R�"1�V	
����'=B�|b�'	�[�`�	�c�^�;`f�|��4f�:?�$�����0�&Q(=�(�'�8�S��M�'8b+̓KkN@�R�=|�����A��?�,OF�b�
Ǧ!��e���y��[�B%~��d "x��)���]�?!�ET☻�/�2�5�i��La���Q�\�@�JԀq��yJF�P�(kv�'��j�΀�m6�P3 �+�S�ܡ��'\O�z���Q�V�Q感W�\��'�����K��f/!�'���'��o]�-����	`�-{b�A9���?���?�.O�c>a�1��]��G�Կ]ц(���7ړ�?�ղin7��O�l��|ZQc��$�|9�t�&o �E;��/�M���D�{�D�I�O.�D�Ohʓc.�2�䗊]��U�3�B�85�$�W�F?1*�y�-S�?����PcG2��I��qOȽP�d�7 �Mit�
'���ґi��
3�VWb՘bˉ.^�9!��|����8A�;:���8���W �HGǄ%@�p%��4 �	�;&4�$�b�g�	
3�v��m���}�dj�3T�����$�'-��>�@ [l<�a��N��Å�����9�Mk��iTɧ�D�O��I�yz !�BS�A+ ݓ!"G�d��a!������O��$�<a)� �S�/@x�X` ��(؁JМ:6����? ��"*�Ʀ���A*O>XPc��2��E�6,��-�:�:�ND/�Nh���)\��������j��D�*I.�(O��PH��eMDuz��1\�Py�w�� '���.?�3��^W�}���?����V��ן���	~�Q������%��KE!Ƙoрq����M��'���{Ӏ�'kw
H�ֻio��'d�AK�$l��ે��(qd��)!�'����%|���'SR라]���W�µCj6m��:Uhe� !���[�jW^�Q�;O���#@G�<�dA�j�r�U��<m�Vq�T�~�IA!Y&Wɲ|�թؿ�(O����'�{Ӑ��ң$�^M"��.�$�:t�S8?Oz��?���ᓿ%f����Q%^�SB|�k���<��|2Ѿix-�D� �l�j5g�_߰�ӔvӠ�Qu�a��i�2]�����?���+�>0��	ѣDb�M5�I�Ԥ�I��xrրӎe@��Y��A��M+����O���m�(n*���䑈�0h☟bV��&Od Cb���P�ˈ)_UV�B�~�$il�B�C�L�!����שa~��ʙ�?if�i�f��b>骠 t��/4r�0��)�$�O��O<"<�d\�b�Q��v�t�X� �k�'�Ng�P�l]�I.�x 	���2�e� ��-�4���4�?Q��?�5�ѹy�6�`���?���?��wg�])s͞`6�!�r�
 u�B�7���>y	6��*aB�3�(�!��)��qO\��G�v�9ࣙ�>�  ��O �Bf7_�8h��0�Q �|�4� :j24�;(�}H�`�'y_� �D8b����ٴI��_BT���u����I��I�G��V<��莂y1� �Q��z�IٟP�鉼L1(ѵ�ͭ*�ıT��*T�x�D�OҐn�M���V�'5���O��
jJ@ar`o](P !�n�"�~���a��MK���?�����	�3>����Ȋ5�0q��Q���<Ag�x�r P��_�F���˓
��Y	�,�&Q��A:��[60@�V*�1�"Mj���(�R�2���	Z�D|i *=b�T�I>Q0*V=ao�PC�Z�.�|IzV��sR�Q��ҟ��e������K;,#�bB��N/p�R�'&1O���e���)"C%U�;��1�|��j�(�D�<Y����RV��Ο칠C�7;tQoU�ߊ}P}���O��c
�O�d>��"*�\M���1y�*�mZ^�? ��`�C2e���v*��s�B �3�T�'ML���&K>d�4���$��v�6�+b�\T*voR�|������3'g:y#��?P��7�3�I��D���O��U�v8CwC�&%RH��Iߵ/v��$�P��ɛ'D-� ���|�:e�&/؝b�b��G{�O� �dB&,暙�,\�D1�!k ��_������)�MH~�-���4HFP=J�JZ 2��MP��6��$�O�I@��>�Iib��-2B���J8�2Ltzue�k�ԝj���w�NE�'�0M���1_�dI��	z�\���S�R�Q>C���h��h�ܹ�"P������g� 0HL�'�����v�<ҧ��t�8(��aa���)w�贱��.��>��O@ʄR|qBggL�;�UH��ҟ�x۴g��V�|�c�5e�p��6�6l̓VQ\�C��i2\�S��Џ��D�Od��<�R'ZR��cD�Vt�E�aO�%8jm�B�'�cU��,S�#)����DG�K<�ţ�j,J��kң@�m5�0.��N��J���b�?Dr� ʇ$�|�!��0�PU�;RK�4�vd/R��yj
_?t��4~���Q�r�����g�I�)'~P�q�
�|����D"R�;�L�GBi'�'P�<�x�"��9 4	�k��:���Ο�`�4f��|�OL�4T��+�c�*1��E[r�m�&Б7L[�O[�zp^����ϟ��	�?A�Iʟ|ͧg4J5#d.:q�p\ksd*d���h�M�u���Pul0����%�ɮs�!؃��ec����oX�E�B�X�m�>4$#�Z�l Y�;S��\x�<c��z@�h�g\8�l��*���͟�D{b�		 3Θ1ţ^ (p#� KAp��D7�	#F��à��9�tLz�N�4�O��mZ���'<j}*�mӰ���Oj���"W�uH�À	I�\Ʀ�C�OR�d44�����Of��9A&A3PKłL�~H����3;_���7c.#��l*%gǗ�X|��)O蝠�]!Rb��4$�!I:���<(?,�|("4��.x�)8��'
x�������<Aq���h��8�C�#n
�2��J�Ip��O�X���W�腂�� ���Z��'n�}"Kj�"���g$~VD�i`'
>p�4��ڦ!��(�M[�" �?���?I���N���?	��X����p�մ"�H�	%'�"�?A�7��bH	�gR�G�T��p͟a���5e�t��s��u�@��P���k&����0��"o�m��\���!K�Χ��l�C�-it����Ɖ=n" �'��d;��?����h����+G�_Z}GK����%�1N;D�����9�8����^�+�����d!ړ�?�v鉋2�:tK7Ě���Um@�l/f� �4�?�,O����H埢���O��<�V�^L�	�@��g��a����=)A��i��X2�#{�x��$W>�3�,9��P��O(IXDѨ���-ќ��I�L�����e�U�q�-�^v��I�Wƌ�)�΄1q�@%��FS%7���o�����6��O��3�Ę�\O�M��><٤�/	2�=AÓsZ�4J3 O�`��y�KZ'̮����xش�&�|�O|��_�d�5�^�ޡ�˙�(��pb�2�f�E����Iӟ����?���؟��'�,b�B�77DJ�	@a�䩡�'���nhHp�	�� L)ݴ."?�nȜV�qـbZ>2�����-�/c�œ�Wa��S�	˓�MK�#��h��t���'̘'��t�"�[Αc`n�-XBfhF�?)��hO|"<�, U  |�2Ƌ�j�f��e�i����<aW��k;LH���XO���vcg�I��M������(I�=�O�r��3U�Hp�&��C��y�'OغQ�' r9���Hab���+��7��6׎���5隨� �i�i�XP����]�s��ő��C�k��� df�X�3���1�"DR��a_n��`	� *{��Q�m��!�c��I���Op��0?�"���3$Pt��(H��ݣ��F��b��D��p���Gé#~*�)#�"��j�����Oh}�&���;da�bE�d�a���'�剅R���������S�Ĕ�;�"�^*�RhQb�Ǚ!j�51��Ʋwr��'�� �1��S ��52��6ퟔ����?�iR�"r�,"P�˹d�Rj#�>ٶ&�D�!��& ,�9�ٴ���s	T�-�0�Oq�!0G ��'�ځbL �ȩ0�OR�u�'.B��<�5���W��@{��ވb�N(�6��s�<i� C�1Z��V�
�>�K��}�'��3ғ`��!��46����`n�i�|F�iN��'S�dʳ3j�����'��']b=�R�d��= ݳ�5Wi$�"�Y�~&)Q�$�ঝ�%���F%.b>c��p6�P�F�D��֫�2u����gAg���Mk�G�m{z\3�<��i��cju� ;�np�#�0|y"��Tk�8|B�19 �$���9|D2��$���Z�g	q�:,p�C�!�dI�6��}�IO�F�ҒR�k���'o
#=ͧ��6�(Y�C7G��H�TnU1>y
�̀� Z�d{��?i���?������O��ӧ4
2��4F]�u�t��d+_8b�
�{���xC
�Yf�Y�}�hR��'9<�� \�۠��<���`a��'Bp2�*X�"��Ъ��z�+�1h�\=�Qd�4:�\�OR-�1��rW��i䁚�4�e�e%n�=�OД�6Vovth���I�HH��j��'�1O^�~F<軠�Ik:�%�ǐ|Rv�v�O�81dl�T�'[���c�G���I7ˌC`5ɤ�'*�k�>r���'
�i̭}��T"���ej���D�wӦ��h��>�����f͈9�lb�� ���O�I�j�$�LI'�^h�7��+�L�1�@F�T�t<�gŝ�b89s��P�wk���+�vk����O��V��$��*1S����صL��`%����I-�����fȂT0b5�W+./��F{�O��dJ������m�����=:&"[�EG韜���ԗO����s�'�L�ˢf�m��9�D
3x��IF�'
�*R�)z���O��Fu�5�B�dӊ��O��1|n�|a�R�Iq�\�x80�
���{ͣC���Q��� �M�_��ZH����|�aHf>��&A�&�B�B~IƯ�?���h��ɸt-�-ۤ��2�b�ŒB䉰�.К3E�,�P��i�I�H�=��tK��\���8wԉ�������I����|�ɀEN�\��cI����	şL����%�
<�>��2�0hڠ��-����+�M+�e�ytȵJ��T�?�ͤ-�d���>D\�MZ�)	��2�d���7-�8G����qE�}E��'A�~�3"E��3�OϾh����$��V���RA���$�'�N�)��?��d_�ORp��WN	qφ��2�N
ƚC�		J`�X�Ǯ�-sL�)���3m]f���Od0Gz�O'bT�j$OϞ:G>|AuCQ?e�nTj�˰5�DD�PL�ӟP����L�I�?y�	��Χ��pS!޲f���Cu-�?�=�!�*{��Zu�S$c�2D��4S��"?�B�T3e�.��K�0�u��ux�vK�'<�"5p�hМ�M���� ?���h���?��'���P&�͙(�9s�+hL��S��?���hO�"<9#�@�_;P8{ժ��f@Pycf�W��`�<���V|�E@#M2i�H���}򉍖MC����dږ:p��O�R	56N40�p��P�`����;)���'c��k%�'��?���[��ŧF�����O�#)��6�D�""��`���-R���);��Y��d�9ǖ9����]���`��:r�Ux���񬔩sU���*��Wu�/��+��c�h���O��,?�& �%,#�d`���*3�AA7��v�	o�z��[	x"Mc'(���t[�,'��]���dL�O��S�l^�e8�|P��V .�:��'��	�2�b��������D�� @E���Иop$��N�8T�J �����I�'�t4��J�9|A�����o~�6�R���?q	!�TLun�#T�>3h2d���$?ɵ.��K���3��@� �4i��U9��A�5z�,h>8�c��h�v���(�nX�V�6?!�m�ß���a�O��D%q��A P5Xŀ��q�p
�'��"�%[<B���F.ӥi�)����O6�FzB��<��@�����8-�#IPy?��'�'�n��U��'���'1�n�&�˱)-I�ly�􋄬mr�X_�rԳߴv�>����۾��O��O��e�W1L)��ʳ�����[Щ�2z����t�v�\�:0$޷tN �t-6�VgH�W�V�ϻf�$!钋P㊵�w��:<����^~����?����hO��ጙ�~�=)7�&^��[��5D������Pؼ�,�R��M�F�O��$T_����'���#�8� oNFva8�i7f�q���^����̟��۟�՟��I�|�� �
#x����+l��Ht'C+=N�$Ja���;�N%�ի �rw�0���$O�LCԵ"g��i��9+�l� S4��H])r^Ū�˞(V��	�VeS�Q�
#�c�M�
�O#�A��b�`Rd��q�Hr��):��'wў�ExrcT;d�Duys�2�V�A;��=�yR	������<\�F����Ě��#i��'��I�\%(EA۴�?���6����.W�0�H��^�}FA@���?��ċ��?������Z�NX�)��Z=Jb����EE�H�p����Hm<�8ٔ.�0j	�Lb���#�R�Ey"��_<���(ҡXq��6K�=KΨE �(L�z g @�d�IZ�"��km�1Gy�F3�?�E�|�׻?��İb �>��u��k��y2L�"K�T��%�D�6^|	 �ͪ��?��'��1HVHT,�(ICn�w�X9�K>qSI{����'��W>��L�ݟ�p��|h9q6�K�y�E�ޟ��ɗN�PT����4N0�#�=��ୟ�����1O]R��0�D��\Gu�'��}�L	�f��1�Q�3cVu�h���4w:�د;\l�,�3O\�5h ,�)'_M�'���3�L�61�#�ӱA`v0㔥�5x��\�'T�0�B�O���1<O��	�Ɔ�%1X)�	5R1K���\�'��,dӼmZx�6����7��_\�k4Ć�UQ�9x�4�?I��?�x�"����?)��?��w��X��dD2<�5"խ|���5m� �'D�5��0�V)[j��S�?�|rSD�6nA���".�9�脘�F	���e�i��0L�GpH���� ܁ AGS�F�-{Aꂭ.A�}�w�'L�ʓ	���'o��O(�d�O���`�;f(ƅzF!�$�Q��<a���?q��?�ga��|j��?��ɽ9�`Y�AЇX}����J�^.�\ñi��D�>�-OX�'�?�-O���̙�2O!�+V4�����F���9'��O0�$�O|�����OB�5q�Ru	v�*#J���D^�
E���Wg�03s���L8il��hϑ��6���@���#6�b��13FǼ`��3���F0\�!U@�Ǧ}�4k�D�(�
D�Kr�G�(AzaLݯ/ƴ�˝	�Da��Dğ4�Iv�'��TMڂ*��F��J��Ӌ?|O�b��GM�/S:����20i��W'?�d�ͦ9�	xy�j^m%n�'�?��g��da�v

��Е(A0�?��}ʤ5��?��O����T�W;'��YvM0N���n�n��a恌k`����]�?��	F~r�Y�`�� `���w�P�q��i�i��K�1z�� c_&�$��J�@�X�#2�>U1OV�#B�'g�@*��2\k�MP��V[�<�21�d6�O
��s9�
(��a~�p�q�(��|¢�'�d���0�4�Д�Β)������d�	I��d�O��D�|�� ��?I6�� qt��e@1KRV�Ab��"�?a�WV���ף���Ћ� �v,{Jʟy[0��7J��(a%#�)���՛��(�m��&�� ��_zhmZ* 8XI��ʖ\J�i�'i:�u��㝁"�kT'�@�'
0D���?���z���CƘ!UJ�Ԋ�`v�A g-D�DC�J��Ҡ����
Ki�)al-ړ�?Qe�In���WKZ�P��p.�,F��IΟ$��ڟ "0Ǔ�:쨥�	����	柨λy\r�'�1.���������ć5FC\a ش,�`�������O��O � ñNN��cTb��2�I�uf8c�T'-�D�.\v�go��vg�Ӝd���cB�pޅ�g�?��	��oʹz�,��"	�OJ�j�:����DD{rF�6�@%��4A�๐2�o���in�R�
� p��%NG�P�@�	��<���4���<q�Lf�T�Pdձ2�"Q��>|q�M?�?A���?I�aɉO����^I�a�.���5�]6ۆ�p̜�FU�s��.At� ��u�f=�q�I3)8Zj`,6�Dᐡ��#�@s��X��B9�h�	
�Q����"%T�3 �J>��'VH0�@+F&
��l9�Ò>��inZ4�Ms��L*�����[T@Q/sF�(�p��q����,�I�	Q�Ԑ���BÖ ��G:mh"�OheoZϟ�'mbԂ��~B��49��#���l�f=�0�0e�d�����?�,���?����$d�3J���S�Q�]�����iʨ����lc`W
+n��7IQ�''6=-����`��l���k�4"U�t�#�[`�\ ��u��DG�1I��(6�C��'N�����?�OZQ�S�
Q�J9QJMT=���|r�'j�X��.K$c�����S�n�e�2�i>q��7�t�qM	e�\�z������FyR�(8��';�P>IxH���H��jĵ6�����J�����e�џ��ɥV?8��7팴,{��вlD6�M�'ɧ?��O$�h�VmW�HqЁ�M�#��E��OB�6�=)��VCI	M�d7�M�{���!�ѿ����\�h'����c<Z1��x�g2��$x���'P�>�͓kҾ�"�b��$v�3VH"=�$��~N`Q��Ӏ/Dށ����+�E{�'��#=���=k3\��G��92GԍB�7�v�'��ɕ1��0��d�����	���	��]�(�x����� 2�z� ��܇��ۓ!Ց@lx�Crj�F���O+���)i@ȉ�'7�↧��k?���*�'h�]J��\Hh������!B�]�-^��B�P>�s��A�R���X����y�P�E�I�.�\l����d�,z��Or���DM8W,�3� �
A�I!Sg'D�|0s�%C"�: �H��T�O0���Q�'�byrF�y���KЮFb9�[�m�"h	󥪎%�B�'�"�'����瓽V�ڽ�!e�/E�*`��K��q�@��`�	Z����֜����نAj�<�B�I[P} ��\-HO*H v�ޢ}�FJĔA?jijԃ��P�0-BH�*`��x��ؼ|=��%��`�R�d{|u�COZ0A*���ʒq�'��6M�ɦ�?�d�IO-1���a�6Oi�8���_ M�{r�ĞG�
P��g����j�C��S�'`�]y�Ξlr��(0Q( .`�x!(c��
V(��Jt�'����������r�֮if�dZ� J����A k���Ђ0	��+�脇e�l���!0R����РTj���d��,v�r���˔pa��mb,agg O�hX��'�B��$�Wh��=���#>�P���<��6�O^]"�ʌ�z���_�3�T,#��'2����Z[��H�d�:���:��H+V�"T� A��eyʟ��'�?��ː�,������
c>!�.� �?����py���2=�#�#(�v1�����4 0@��`ΎQ�1e�� f�ɖ|N����G%	L�� K^�Q>��6F�/s��!* hׯ>4�Ȃp�7?yd ����c�O��� |����N@=N%r�
0f�C�"O6�I� &��	���h�Ƚ:�����h�J1PVɝ	:@�@�K�	?=b�;��|��D�Vm�<ɶi ���I�eJh������"}۠@��5�T�Y� 
�"d*�{-��;c���8�3扨2��L� �S�/%�1�+�+�o�2��AX�EO '�t��`5�3�ɪ=\���b���pcļq�T�n������"�O��3��U�|o`l1u�κ?�ā;�K}C�I=]J� 8P�B�I���Be ˓A둞��O#Z�8C�.��#����K�b��T[�B�㦙�#\O �8"��0�|DR���I���@�e��DMx	R
K,�l]��lב�p<��
E7Q�6���X�c�>�AGʔ+(%Yn��i���L�- V�񄙸]��!E�L�s�Xݘ���~֮����'��6�o�'�܊������8��=����,D� ��� >�ġ���a��*�d�}}P���� ��M#q
|���4e.,q�̚/4���'�HJ�'(�䍂=/>��ȯ�p���hU�s�by��-/O�����#�
8s���.X;��e�UG����$�
t��e:��S;8ɸq�"g�>f:��ĉŃm!򤐠s�0{�d��t������w��B@�O$uC��_�{���2!: ꧞|r.ڙ.�6�B7Q?b+ŗ_-�)#G��)�8k�� ?y��% H�@��7�m���*�'y�� �T��LĵP�V��'f���-� \ǒ���;v��DE��M� .p��"ᫎ�F
$iH�Ⓢ��$�3�gӖ8G��<��-�6��"o��)�)x��v"OVe�w�O�~	0����Y�A`�{��	��h��Lr�'�VT�� 6�Q��j�y)5%�<@ [!����< �L�0�A[�$�طF��b�ءt�!LO�{B��N"���v'H �b�Ā
'dazb.��r����:u�Ts�Æ�	��'r�TC��͘Ϙ''&�Q�jS$9H�2�A�#n�Ԣ�'F����.=N<��c.d�X)O�	Gz��)��(i� 8Q(QZ�RA)ъM�r)��fI��?u���rt�,Q3&ߒ"��4�5)\*ם��1A �y��ͫ�'G�x�t�P�b�Ɵ�񔥝��T��՟(��N�x7�1����O�t�hٴ1��])T��)�4 F���6#>�wݢr�F�q��$c¹�4Ĵq6��u�d�A����n2�$b0j:Ac�|˄nۄ��'d�|����?y��4'ݥ�����l 3m�b����N����>�O�8)�,ofM��.J�a_04;�|�i>�:/OxybDA�0f�,гMӚ(8@1ɷS� ��kC�����Ɵ��O����'2B�PkAH$�2�����6b�z���9���l��IB�T�w)|�p,9�O�1����A���hˌ-����V�(K7<O�e(%*U>nR��Mߩt�v7-;����c�{ð�'#�l1DAtaRe�FF�.�*h̓C����ʟ$�����B�?_��k�)��R�
��c!�ά�1�RF��%�*5l�%'�O��D�b����J��u	��Yg�BD���ā17���'MR`̓c�#�' b�'r�O����P^zHE`�X}N�����L
Ck�ڐjU�2���YF5Z6�d��w2����DV�#���1�Ֆt��|{�Ef�R�2��?F����2'b�?�Ds����<��-+T	t(ڸ|�x,����\~b�P4�?����hO�扸Sn����ՆJt>�yA+G�3ӈB�IJj� 2'�Y�p~�5�E�UPX��ɝ�HO�	�O(ʓH���1��� ��%�j��Vɋ�(��e������?I���?��'�?)�����͐-gb pAP'?g��XG���U9���,
�@A���D�BC�&�
b�'�`���<8t��	�/*�`t�� "���:G�;����!�i�`(D��%n�$L��$%n�2bU�%�4AX� ��m��a"��.e���	~�'~��Əؙ)/���� y��Xcϓ�O��&�1bX�@���J�.�S%\�t�ڴ�?�.O�Řg�T�$�'��)CbrJ1�!GM��`7G�=�b�����'�*�X?N����K�k��קvӎٹZw9*y3��� h�X�4cA�,�%ӌ�$�>U�H���A����Isq��a9�͘%[�b
}��Ac
"EZ�k�N�c��s���Oj�d(�?��B���,3��@6(.	G(˓�0?�⌳)~A�HS7v�b�0b@\��x���-�<13.�, ���Т�ک_FJ���\y�ቌr���'P�Y>�FE����4}�h�d���.E
&ɧ7@,���a)���ֿS�
�PD��M��?A�|�5m߄3hY�Fkź&��ؘ��L�<���_�ZQIÕ���4;J�в���L.��ʟ�����I�����:5����7O���q�'3�����z�S�? v�``��
R��u
��jL|1""OE�	�[��̂1�Z]�,��d�O��Ez�O�R��Ԫ9&p����Q�'��Ԛ��'���'�f�� �hB�'FB�'����'�2���Ax�
	f��H�y3ꞷqZ7͗������ ��$"��jm�O�@�'����x�Q�z��+d� $�6mW�aC�k�D���'��p���Z�ᐝ�)�b1�sIU%^
 R�B�,�p�'�"x���?A���}�"b�, #�4��⛗N����=4�Cע�
e�4�2�'��楡Ǫ�˟P���4�`�$�<9������Ů�h���ѽ.�$�VF���?���?i�����?��O��ĸt��%{t���c*V#���a��`'���An4��E*aD��%O�'�&�P��#:�F�B�ߡj&�zj�-�0zPO w�<��i*��!�'Y�t},r��ę�tZ�+Q�L����!뛜"X�����T���w�'��|�n�%�� q�A�2�0�ϓ�O���$�����V�¹MU.5��Y����4�?a*O���a�^��Iş��'K��:��o�T��tl�Q0ʌ�		B8`�	ݟ|���bn0�O�I�� �'*qBp#�'�&�eMU%I|ƙyeG��E)F|��w���'����k�M�rZD�9'G^7a#�%�%��3'֪]�T%�TR�:5�(l'�O����'dJ6͇y�ӭ1��aQ�	ґ4d�X�F�t�T��ҟ��?E��eT5OA���놤e2���c����'t�#=��a��ƀvӐ\b�KæV�&h��ήN���<����?9��?A��?���D�e�xSG��~���i%���cx:�?��i�>�(��V�}��l:��ƞe�>����2���1�O�u�����M-p����*��}�t�
�C�!N�amZ�<1�O��<q�	� ��I����p!0���0Aхl��dŴ�j$�D!@*:-mZ�p��
ן� ��!����ם#[$�Di�U�f/ �#��(3�<�aǠH$o\��'ZX�yb1O���h���O�0O�hI�V"d8ɃU�pؙ�avnr�'��(���'�_V����u��~�@־r���vjESMn�H���ݟ��g�O��$�	gӈ��O��?�	�}²������۴-	����2��NɆ�����p�쟤�����$���2���:N^��#�@ ^��sF�0�$U)�4�y�Hū�?���)%���O2��?�#�Ꭽw���AnQ�,�6�X%��<2�Γ�	��ڟ��[w��7O����ӟ�F�� ��蠷�]�a�d��ؤZ��<���lӒ�	,a�Tn�<�M[5�ƴ��	�|�_\�Ҩ��\"����~	���۴X�"�'�`<ʃ�i�H6���$f��2���O"h��#�uBp�pL�-���c�����3R���@�'����o�p���~y��PF���tCOfq������ܤ�U"Op�@߁ c�s�OO�K�y�տi���'��T�IK�'L lq�`є����k��aT�i���'B�'���'�V>��i?��!'��R0�e�OM�BJ�eoZ����'�	ӟ��'�I�T%i%�N�n�
��0�I<I��Yߴ�?���Ī�,k��w� 0�ܣm����,�>�����Of�'�R��SoB"D}PV���K<A��?9O>��{,�:;"H��B�Xy��BiK���O��\��v_^���.�>����`�`�b0�ȓy���劍7���Z����\�T�ȓ�x��Bk��	8ڼ�VaF�z����P\���͓���t�c	��*A��'�R�A2�Q~*�t�"�)>��'R����p�r��`�tu��IP���O����O"�$�OB�G�u8�8`��+&�2��6o�3�^n�ӟ��	ߟ�����ß���՟P�	��B��,5��͢gh�!X��
�4�?y���?���?���?����?Y��X���:"�I8l��= Ѝ��D���*R�i"�'Q��'Gr�'�2�'���'OD����@9n���Ř"^Tnay�Go�`���OB���O����OD���O����O"��'��?M��F��	O�X�f�ئ��	ן��Iԟt��埠�	����I�����B�j�eY�Z�b⦤J��"�M+��?���?���?���?���?�Am��N��h�  ��%�P�S�>�f�'��'b�'���'"b�'c��_:���Hő2u��x��:IsZ7��O�D�O���O��d�O��O���H�UJ�%�Q�z��@$�<e$@�o����Οp��Ο|�����������	�J�Qz�
�JH�iS�&�8zߴ�?���?����?��?	��?���R�ɚ�$І3�4d$M y�p��#�ix"�'�r�'dR�'}��'��'b�XW�_�S�,�+�BK��|��}����OX���O��d�O��$�Oh���O(���[=�ib�ч<��uQ��Ѧa�'�U��E��%<H�)��E�\,���=y������';��\l��<7T����ΨoD��p�ʑ:�M���i�>Q�'�z��q>H�9ش�y�=z��(�e�ԩW����b��y��*_�Z����ʻ!(ў�S�<1F��*pL��p��ƢP�lT�0�����'��'��7�3T01OV� Z�` `���`���ļ-'4M���D@k}Ln���mZ�<y-��� d�8e}0}��Kj>`L�S�\���YFB�!(&?ͧ *�d+Xw1b��W|�xb!�΢xz� ���5,t�����Ov�}�M����SC�FC�� ʁ;x����	��M�h�T~B�u���S ;�~�X/ëW�`H�'Y7T6,m�I:�M{�i2'
@'�F���H��X)P<�u�s���`J�Kŧ~�	�р�8hq�͟�'1�$�!U��s4Љ����#�d���Q�0 ޴�F�<���E�eO�0��Ɵ�G�&���ߐ;*�W���Ar���e�O�<@C&��gEv�K�O�B���eEY�D�#�O\�	���e.�	�����Q-�a�&��:4琅���0P���$�O��d�OJ��O˓]���'�!�y"H@b�ʅI"�U�`��!�#�� >��Iz�.��*�O \o���M��'\l�I�eU�bMÔ-rZ���DU��M�'�bCN)���s�,�:��I�?��;n��0P'�M�P��dl�:W�>u�I˟����Iܟ�	`�O�6`�tEP�6�4۶�>�Ec���?�s�������Φ��<��c� H���
�Ӆp>اE]�ēk͛&�z�"�I��c��7�n��I9�8�h�횓r�N���c^3W�5�֍�%�� ��TO�uyZ�MS��?���1�m��.<�ta eM��-�����?�*OƐl�
���ԟ����?��'"C���ݜ&]�!z�	��ODN��'V������m�� $���?ɘǦضTn�H�'�33����LM�y�ԁ�w�٫{���'*���[
+���J]�ɓ=���Bٞ"�� ��f�:d�I֟��	ޟ�	D�Yy�bf�ƌT�V#&�
y�/�<���4��+5���)޴�?�N>!"_�l�޴z���Ht��MF�a�A*��oeI��iު6-ڍ&#�6�i���I�*'�� h�QrNM�'�1h�f�-`�t|�D�+n݊�ȴ�'l�Iɟ\��ܟ��	ꟼ�	q�dI�=Nl��+�NZ	����ȋ1��F����yB�'����'�l7mk�Xط�O�+�x0����1@�|e1B�[Ϧ��޴��'����Oy�T㝥ZΛ�4O��p"iĔeSȸq2o�}�$H�@k�O L��' hZ)@��3�d�<����?�Qoޑ\�,���D7^�r�Ad�ߴ�?����?�����=Zb`;?Q�Jوh�k�����:wC�@���R���R��	��M��i�jO<!挌�@<p FE4M^ �z ��O��� 
��HCV,>k�ʓ��Fϐ�u��~�@S�����:=+���+Zx������O���O����OH�}ҝ'�tĘ��׽b��E(��#~F)���43��`���dO����IC��?�yÉ��_�6`A�/T����֧����4).�6Iu�αȆiq�>�	Ɵ|R���y3��K󎞲T�1B$o��t��	�_xP�%� �'e��'b�'62�'���;P�/G0�@I�A��A�U�V� `�42p�'8r�	� =��ea�@�[]҈ �Aյ ���'��6-E¦�N<�'�2�'
$�UB�2v�P���03���+�$�%#rmJ/O� �dmE�����&����̯?6����+�l�Bx �@�J����O��d�O:�d�Ov˓-6��*�%z�3!���B!핇@*b�	�օ.��I~Ө��*�O��mZ<�M���'��[q��V���z"��16$p�x���9�M��'�r���"�/��	�?Qj��,��.ϖzxR��kT=3@�!�AaÄ)��6��2o⮉j b�(m��!h��O�I2L>�DN�"E���Bo��x%$d´��m���SҁV�(v�,�eT�7�~}�@�ۇ|j`9��'�75Mn�"nҪ`Ѝ(f��BJ
�3fS�+�����ލhB0Y@g"�!޹��܄8�I��ϼF$=�@ίt������+Ng�@ǒ�	�\
�	�$�J�
%gʶ2�]!bŅ9M�\-���ȿ
J,�N�0u�9B���2K�v(N�2io�	[�"N�?��v�р��E�c�
�����M#6�ߤ/{��X�L�#�Hmq�B�bC�V�`�i�Fz��O��і	C�8 2���2ޝR�#V��R�g�tn�3Xj`x(�8}�	JRO֞wc�x	��Ԝm���3����T(�jݱRJjp��L�"�d��Rf���nq�7�͢���剗Q0��CU#��i�FO׍	�#<)#��>-�lȻ��Ũ@5��S��\� �3�K�;6��їk�7��Qr@"�"h�)w���CJ"0J�pr��-��m����%	-�҈Bq/�- ؑZ���-mv�ٵ�ǟ}���� �Oz2�;�ԞWPYAB���j����H?t0M�0��q(C�i��� �^,�5���I�X�1U�H����$�L�����#QNn�(�&������聶u����]ƟP���0�	�`�I՟4��' ����IǼ�"�l���#�.�D�Z�]ß���x�	ß��	P����+}�bO/7���W"߳Z� PEfZ
�?����?����?����,�?����?I������V��`��J�Y|��i�ǂ����?a��(�z�� �Y�S��.)R�l���;�Ԭ�c����������B����T�	�|���?��'����C����E��
�d�E�R�'�'�RA⇎�;ј��O&r���l��t����U�ߺ/�(���'����?���?�'�?	���Iܠu5�Ի���	�Hdj5�]����S<?'�=b'�����	e�	5zHHyw��SDR�`��M����՟��I>T�|��ܟL�O��8O~����ʔ<:�2v�R�l��u��6Ø'��4I ���'�R�'�nY�T�u'^!Z1c��oi���',�n�!�'����$����/ӶWpH�W��3~n���jyrG�:J0Db�O ��OL�D�<�&l��DP�ͨf`��u �3b�X�јx��'�2�|�[��� Е�����ohd�D�K���F�*��' r�'P�V�<#�L���6F�K
a`�ĸ{�yK�Ay��'�ҝ|�Q����N����$kIc+�=R&�E&U�1ٳͪ<����?�����DN�\�i&>!��O����J�m-JQ��?��'>RQ����Ɵ"��%��
0��0�B=L� �#̋�2��Oz�$�<��x�O]29�wƔf�
 ���ǄUȫW�'��۟P��3`#|:�wV����J!��\!��1�b�Q����i5�%oD���')�tB�<�5�O9R�X&���I7���Fc���O~���E�H�S����L�ڄY�
u2"q a��5��D�6oܭlZ�(�I��������|2:T�L��MJ��� ��?�?���e~�Q��&?�埬����h�$"��;^���Q��=�Mk��?a��#!�L�P�x�O��'l*�`�K��K`8؀��Q!wێ��Q���������#�I����ԟ�zb%ȟ:��/_!Y����ag�ß���)QM<�'�?y���������a�%5��q"�_� -��D�O؍�d�$�O\���O�˓/N���e�U�v��1rfM�1z��� ��+e�'���'U�^����֟�(dK�X(nXb�.]�~� ��U>2Fb������h��ey��Q��)��B�έ�O��<@b���S�A�I���IϟT�'��'����OV�2�Ì�x.�+r��)F��1k(Ot�$�O����<�Ü�Vt�Oe`(��"1ޤ,{&��d�0<��'���'C�Iğ`�I�y��>a�Wl;d�p�R<<1Xcb�O��$�O"���O���̦��I�\���?�#��0�dD�s�̠**����!V����Ky�'�V�ȞO'�ɳP����r���!N�+����e�N�0 I�I̟���dB��aٴ�?���?����B��g�d�K4BU崑�Cƃ$G#:0�-OR��"e��$�O��|z̟.0Q���_tթƥB�+��ZP�'Mth�(w���D�Oz�$������O����O��ifg�s�B�1օ̡a��J3��O�c��O���<�'���?!��@�� HW��@�X�n
=��V�'���'"�3!�Or�'&��'�R@�{9h���4N@��W�"[��Iwy�oY���4�����Op�$�v=ԝ�el�Kf�X�	6$���d�O��3`�L}r^���	Vyb>���&��,�R��s'F�1P�$�`\��j��j�H�'8��'"2U���4�Hm���,�'o���ձҔ�ʮO��?Q-O�$�ON�ė7�̱��LB�*�[���U<�1c=O����O�d�O���<�!��;g�L՘ �C'iנ|����%M�3�?�(O0�d�<����?���/����2("s�
�,�\ʠ�)A9䉋��?���?���?9��R��+^ʦ��֟��G�;i���jۚ7�8�Um���������I\y��'�Z�8�Oy��:�f\�&I�@�'��]IT�Zd�Yݟ��Iԟ��	�����޴�?����?���#���ȝ�v/8���Θ.��M���?�(O����!F����O ��|���ծy߂M��iA�? �f��?����?�+����'�"�'A�4�Oo 3�]J�d�r�P���5Ut�ҟ�`�`���%��w�,�?CS���`EO�>$�Ѧ���?��╬kU�F�'�r�'����OeB�'^�K�2H8�)���^`��Jt]P�ǌ�3"�'��i>5$?U���Ԫī���*7h :���8��%Bٴ�?Y��?����8+�'���'a�dW+
Ě����:TON����.P�|B	�>,P�OJ��'cR��0������5�������l�B�'$��+��)�$�O���+�ƿ^ �EcsI�������G�]�����O0�$�O��.�j��-[���y�2c��0�h(�s눛]؉'f��'��'g��'�Z�2e@��TC�C�3OL�%.	 T�J>Q���?�����D»=����!�`ӂҴ5J��۠Ťv��ʓ�?����?��<D\D*��� a��ϴV���P�"&!�*OP��OR�D�<��#�O/h��S�5S���� �#dH��'T2�|��'U�؁�y��l�E
>@w8�SFN�>^�X� �O���O�ʓLΈhõ��D�'���6f���-��80"k
+�:��|2�'��%�&�yR�|�O�$����@:I�yF����t[r]���U���M+�"�d럸�'�R����3H�C4(2u�E)���?a��Rِ�[���Sܧ!o(,��q������ļ�Vt�Ʉk3^��4�?����?y�'/�'��C��
`�	G
Ma�42ԎŞ���8�yR�|R�	�O�I1+�Lx�d#�뜍1�܌�vLNԦI��ߟ���,�)��}2�'��DM���)��O2�Dk�q�B�|֢U��O4R�'��I�:��Qr H� ���F6Z&��';rĭ��ē�?�����z�
� ����LJ ፯z��(O�b�9O�˓�?����?�/O�Qɇ&B Lh���=#��U��CL�f��%�l�����'�h����\�%-�����*�GͰr%$�m�b��oy�'�b�'��Ɋ$	"	���[��� BM�l��儋�/��%�'6��'J�'7��'p`=+�4On��c&˚5��Ax��~��x��Y���՟��Igy���@�6�Ĩz���'L�"� 6�Z03�1 ���O�� ���O��$�Ǫ�$=?� B��W�#^@��N��a����'��'��ɐ[O|������"Wg��ͩ����g�@�֡I����?��(vVeDx�O��yr�&L�2$��R��y����\42f\o�a���'��T��<� ��7��xrJS�W+2�)@ٟx��˟ c��ߟ�%��>)z���(�ʄ!�/sʚ�jv��O��!�̙��a�	ӟ�I�?�O<!���P��0`x����Nea��m�<����1�*��8�D�=n�rY�p�Ƶ>E�21�A���#�׶3B8��fC�w�`K^?g�l���'Cb�'�ui��Ow����b��W<�y�c�i�7�SL��*
͟\��O��	�	̼۳�.v:X���#T�рUi�� <�#��l�8Γb��'?�\C�cͳv|�s�/��8������9D��ʖn��<��$Q�`.8I h�*o�TyAAi�=]0ݒ&�x���Vϗ�~a���� s~h�`�j� {�$�H&�]Љ�$�HO�y����5�<�, hQ�R�-�Թ��H(M��СK��@%;�F�Q��T����H��M*�*u�T��8m��(��]t*�A!h�5v����ҟ���͟�	��u��iw,�q�D	�#�=#�K� c�R`�㎁'JH,o+x�-b���]�O��b�Ȑ0珢D]Z����a�ހ�7I̟9<(:��iXb���r�,��R�?5��`� �:��wx)�Dĝ�C���1�Z�vj]�4�1?�wcD�����n����m�0;>0��HH�Sn��� ΂Z�<�󇏉d�D	�wK�	` �0��`X :A2�+��|�����D�I/�@ڰo�
��E��D%|U�s�U�'�6�D�O����O�E�;�?�����TL�U��X���y좄r�$�/L�>��☽&��-�Ԩ2p+b-��..�>����+����b'�� /�Lt��Ô75�2<��
P�F�޵ɱI
�zR���q��}���)p��"(!�-ZG�	DG�h �џ�F{��I���U{	����=@A'�#T?@B�IBhE��I�xjz4��l4�'*7�O"ʓ�d�@�i��'��V �kR�+׮��@!LC @��D�@���D�O���#1�D
���u�� �T����u����1~���p��I/�1��I�y�<� ɛ[����&A`�Qi�5��y��"^�1���@�iRr�'?��@���?�N|�kY-p��T���Р~&���	ð���'��O�>=���VJs�qsa��"�Ӄ�6�O
��3L4}Q�,�2"�xC �j���9�W��"C�M����?�,�����O�6��j�4`���-x�h�o_��M��D`����S����P�;	�t�i/���x R�K��P;p������
0�U�ģ�l�k�&L񆤝$<�MB��=ҧ X�C�,V�toV @!A�/G���'�|�C���?��O�O�	 ���ӆ�P���
d�5��C�	�`��<�Eӭޔ�XQ��?Vv��>�a�!U�q2��]�p���shT6+�$z���?��|� z� �?����?I��!�$�]�ljz�"�EE�4\�4N=-�2���3i3� ����0F�~X�!�>��L�Q�lA�-O����@�]�h�X��\im
�R�"�|��f��{��5�&�ı1A�O�X�s�	Ry�Íu�F��ꞓGd�L�P%\�@���'M�����j��'�i�|Hj�N2wS��FC��1A�'���Ӆ�0�����@&9Jʥ�'w�"=Y�'�?)*Ozt���á^B���@ĩsh�܉�i_E]��f�O�D�O���A��'
�)�:`�<+�(��e����K�@��r!�G�2���qe'TF�bL���ba��ǈB�8Ua�AH�A\D�bt�4F��\i�]�l^h�˓h���mZ�$����Z�3=�t�[�@P�D���?1����$�O���IG��I'Ł@P���h�!�ē�J1����I �68�=��*��y��!����'{�I"h��<���R�D~����'�2ez`�c�P�o<�|�M�˟�RS%Gҟ�����x�mM�;2��`�_PD#�ӺS�C��x�׭��KE���q�'H<�	7 �5Y{��q񮟔0�b��� x�(E���{�֔#��2.@
�F�a}�T�|�&��?����'8��t3B�5:����3OF�ĥO"��d�9x�i�F���n���&�YB�qỌ=�'W{�Ĝ�gO�XȱJ8Od�����R��y�'=x���o�H�$�O��'h��)��M�g�m�x�a�W�v��X���`�o*���`,�鴡�8N6]>�&>���\VJb*�g��W��a��>i��]�?�]c�O'#��rC�i$��+��*d�4�B�՟���fH2R�X�a�/�8Xi�S���BG�O||%�"}�A�_�;N<4�L<Zx�ap�<��"k�T�J2&ۦTfx�8V�\C�'�r�9��?��v�	�$� Zq�<�ui��'u����I#����1���"���n���0?9��+�����H$e;HE��.ְ�j1+��v��x*��Cr����`�J�bE�	ڄ\��(���qo�>�3�OJA)*(��@!�1:ƃ��|nX�;�ˌ3����S�?  ܘ'�Ar�ڡ`m�@<�=ó"On-SP��,�n�QU"!$x�"O.tR�ӠB$��He�!��"O
2��˥{*��ЩJ�{�Dq$"O��0A�"�d9�@ڂ=��"O��7�ڝLsZiB�iXm����"O�:���()���R1���y���"O*ʡ��*=>�V�Q"Ch��c�"O8M�AҴ[2�����&KU� ��"O�9;�c@�#����E�C8�y�2"OXՊC�Ň@F��W�
M�0�Jg"O��A�㛽r#Tؙ2�~���2�"O��D��\���F$���`٠*O^$��ٓU	����]�9'L��'G^pV���@"EZ�-�
5�Je�
�'���Ci��2��ѮK$�bp�
�'�B P��E�{�J`CQ:��|y�' \ec6�N�r�����Z�,T�P1�'�\d[%���-��L���D�1j�'�N��A¦��p�=��q��'P&ȹ��Jdp�҇��xx�'��Ee@�A��\�v�C�ZL���'��HG��j��1���y}�-�	�'��X�m_,�`�Y����a��#5��Ͳ(6�O�	�7j�D��9C�E3<I8��I(0��⦬�|�O�r�8Qk)9H`M�1�B?@t��'9Q��,3Ԑ+A�^�{N�|"�Od�����1���[���A>U�5E �;����E�q��`$!D��3�j�~��I�4 ����1����< �P�͓M z��QK޲k����'�f��4�F& �ejQ �s��4��gfE{�c�%V�DH�)N4EkA��Ј1�\%+ehŶT��TK��'18�#G(F��k���#Ø����Ƈs�x(ٱ�	�v�;�ؓ��D��/Q�y���
 ��YȑË��y�"P9b#���3�q
�z�K��yB�-<*xXyg �������∟��X`��Q�&	Cc�<U��A��"OP�����)��j-P+!�04d�;��L��-�e��z�/Y�DN��`�4�ā�X!��$��I�Kt���I%�n�ipƏ6f؈)�� S���n/*jTv-�!VQ�0a%���=�GߴF�t��ǀ7���
�I�'<��F��_��$���\�V���C�i֚܃�����d�V��A2B,�<1�C�	��HR@�OW>耢��<Q.�	 ~���B�/�F�y C
��D�$��햩�/C ]���x�D��yBER�)]�<x�Q�{��4��?+[>��b�J�����O ,����ʟz%z�ď��p�C_���Ё3a�pEa~��9!w�����P]"�*�[8b8�!�o�KG��y%�S)d7��k���0=a��ߌ!��M�����qތ h�C�]�'�飡d�8� L(�.Z��l��3�١�&�;J9n�r�(j�*���'5��B0�E&u%"�A�Ŝ֖�Fv%�S��c�	f��ӑ$V b+:��'6)�h�&_�����wv��ô#_R���KW��|�(ܓE�� ��$�>YhQڀ��H�F84̀9ARĻ�$ ܌�D���:À�`Y�%�Ā�t @�	�:qb�ZV J�vB���@�ρ�jȹs��� R��#��Q�tѥ��C,ZyÊF�q5V�ŉ�Z��@4�3�dd	ӓLZ �$
��H�[9W��P��h7����ĥҠ�P�(XB5�ύr+�xyqM](�y��B:��q�æ܇H��dI�d�(v��6-�>/tܜ� �'7p	 �iY�� �n�E�Tq�#�������Q5�Hi���48j%H��Y�� ��EC�t9�w��P�K�$J���bA"?������z7�G�f>�8VH"g��a��V�:]J���2b���!b扜s|�aA�R�a1�[��!`��)GA���$a2VcI��,1�	�d�p hw��uΆ]F|2��E�"��Sl[���j"�2O(bm�̀�dFd[����U�"��x��Z�&��CP��P�+\)��-A/������'��xFl�UT�2`�g\0�'�>��%T�ɐ	�f��fˎTK���ZJ��'ώ)�L٩P,��U����PT)3@T:t���2��Yͦ`�JU؞x���9,=��JR)���P�/Az��ca�L�4��`P��5��I&��djÀ2�֌P�mj��1�E )@�Dey ����@1R"�O��s�N�(��a�C�LOR�`��fߊa�a�w=�a�$ăt�8[^0l�U�Ys5�Y��D�v �$M�[��	� ��0�c���:%#�%N�O�8T���	��x,#c�%a)���I�m��	�����r�iCW�z�*��T��+g�7wm.����F+z� �LQ<}�U;�FB���'�h�H�1B"�����U6C�`��'�BT��HU��N�.�\���ŲD/ڐ�	��H�@�"@�~�\�)q�@���.�*|v�}�q�ԂO=~�r�(E��v���@=�ZP���3�eR�nE�Ky���ć=�Y1��]%@�X�����|�R\���Y<�M.��Mwܯ�ac�D�u!K�/l����A؟�:p�̐Ks&�CP����c�T%�TM)���8W�Y0 P
:�RU*PM}&�#𥋐������B}A@g� �dW����u%�R�:ݪc� ��J:@j�?F�KN$�j��N����j���"+N���`ŋ��u��J�+Rd�0�����;	Z�00���u�*�I"wxuj5IԊ#���˒H�b��F�����(�tz�#��M�*�b���V���l�F>���C�*S�%�qh�~����G���9���r�!���\ ��r}��jA Kv3��jU㮔 �Ǌ� �4@w�"�d�!���wt��Ja �w7�� r�V䠌(�;w��=ɶ��d` ��H3�j��ȓ6�te7IW�F(4�v ,���S�5t�~Y�l����
4�ti	בG*��� �?P�Uy�F�m�<M�p����M �O��<3�Qx	�ٛ�MS%�p1:%'ϊo��$o\0PH �0֠T}���B���lZ	E�����(O �yf�ٲ�I�j�Q$,B�'Ξ�,r���$���̫�Ǚ)+���@��#!����l�A�h����Z8��a�����D�P"��r��A���'�L(z3�Q�t�0���W�~J�D�$GՔ(��5� @�/�@�w$�*�y�`Q7��i�PG$���q&ρ*I����	s<�@r
�d�
���O��3�I-8F��A�ƜF�	e�mfl����h}�ŋr�P��՘R��@���T�r}x�GM&~�F�Q�J�gh�	��	�t�~[d�
<V��eגX�"<Q2[�{EJ�9L�����]�HiG�#e���3�!�=Y���&V \C�I�Y�x�Y�a≊a�^iw4���O�! cOՎ��d��\. `�s���9�h�9�a��_��)��Zi�K�"O�p�R�(q��]!g��,�B�O%+�>Y#�җo��R�� )}��͒w��yҊрŘ�1`:!�rd����= Ƴ<q`��;�V\��'�<$��Ħ�k�J���8y�L��®ϰ=�@�]�z�����$��6�:]�'��H��*���i�6,��kM�MQ����O0d�O? `f|h�J�G06A�b"O=�aB�%��*�F¤[.�M� �r�MH�T���ŀ!f6H�?	̻ {(	[egB�g�p�S!ZLѸL��FE���,Hˈи�.I9�Prtd��<Ȁ�'s>x��'{�����^�"AN�'w�F�!��ˉLmT��$���t��łv�n����L8W�ن�9	��h�L��1żl��\/\y2��?���/�S�)ݥn^�WgH9_{�)3�C�7+�!�� o�ȫG�M�6Q:��ѤT+/��Fy������4?�pA7��2>�.l��A$T�! k�4(rƇA��Ȁ�'� (��ɳ`~ Y�U ��<kdC�h*����J3��Y�D��GU`����H�ćȓ!�a�$_2o�؁ %L�q��?I�#�S��ӳq�D���*HY���s'b�!�\2�U*C�̼vr�sEM����Ey2��
�ʍ�h.�p����0Q�̩J�n/D��y&e�>�� �BC�h��ytcp�����uŌ����YVc���eo�z�@��/�ēU�L� ��=
�l�3�մ��p�ȓ9/��H6R@n�C�8�x Dy��|ڃ
��:��@B:X�=0�~�<Y��b���@F#P�����}�<!�Y��Vh�UGnD��;���z�<��D��zO���2F|@�õm]ryr$2�OB0Ȓ��b�u*�M*%3 x���'�Y��'�ʄc\�o9T��B8ܾ�b�'�*`97G�� �h�k�%&�KQ�'������W�T8Õ���`��� @eU,T���Jê�y�¡)�����*����$�3Nf( p�А��)�'p�b���Q�UI�h�5�ٝ�r8�ȓ��);��� 3�a0I�PźE�ȓo06y!��(U�f��H+x��p��S�? ���Q,�<Sa���1h��;�x�F�i8��Gj�Q=�{�O?7�>X$�x9P��Z(���B	:�!�6q��'���/����+�����p�l)pHV�cVT��ɻY�����%�z��)۶��\�*����z6)]-C�$��aL�Yq
UB`�L,���1Y!��F.�U@C���e��ᖱA�O0���H�7�R���f�;3 '?I Bg	*Z!$qsB������!)%D�����s��FX}ąBЧ���=#��GzԸ�ǜ�|#}�'|�gG�0v������s��$��'N�Xu��6s:�)�Ѕ��7�z���d�TB�Mc_�P�r��[��y�{�'����f@0$��|�34��	ۓN�=h�F�5�]��=F �8Dh��[� �Σ#���[�PL؟Xy�
�8n?��y��N�V��V�`�T1�m�~BŐ�j�lR�I:h4��1�N���'	A�u���Uot)y�猝#B
9��I�_M�GP}b�Y��0���[2'�V\�r@�s�����R��RO*���Y��c��BS�PR�����<�IRU�����?3dQ?����J�x s��7�����*H#�p�t�F� ��S�/j��=�f��B��#U��7(�<&�j�f�$���'{BD{L|�b�!P<���A�e`>��E�C7F�+�ҏ� ,#��_�0|���6{@�˒փx��#���H��|���E�)�~�7�'���d�4~D���lփ��	3J|��@U �x��˔���ueI[��T�ժ����O����g�,=к���u��+5뛸<w@ኳ�گJ��Ii��8R��>�rQ�<�")���I>l�<���d�?i�(���ɝ�����!�f�N)Q���~�z1oH�"�TX�ՐAE�m������>6���҆�'���a$���Ye8�KS�ͮo:���l&?���Ȑ�������Q�clr��]*d�:Ǉ+C���$E,TuV��`��=�@��U~R�Z�
2���'�X���V�;�Xh�Y��X�|ҵ��hEp��oK���;ƞO�<�Be��5�D3V)O�H�f�+V�ty�A5a���)�ʤ>E����YsF|���q��+I�ć�!"��R���d��9p��4"t�'|�,�PLO�2�l�	�<���1��rt����ƍ9n������J��En�e�n��>��]���`��!��&X�e�s �2͆�`���h¦K�@���@kě?T�Ć�m�0;�`�:�Q�@&�w8��ȓd�&<Ha���"���F4��ȓ?bd3 �FMxa@���{��хȓT}\ a�b֥.l<Pҧ�[:��ȓ2�N�xB�гD&	A ����a�ȓ.5*Eɔ��U]rp�A`�@����m���$-W n�NԀ K�!,Y)�ȓ$|����FC6�� ,�Y\X�ȓ^��qh3
Dh!$��U�ܚi�����WL�Hb脑��|��@;Ņ�q�H�a�V�Dy�C��$&X�ȓC ��
T"��]�d�R#�FV2e��f$ޠ�ټ&0I��c{�Z�ȓ}$X�r�H�6���K�?KjɄ�f�̈�De��(�n�Y���6�~8�ȓIV�<c�����RØpZ�ȓU��
r�&I��:��Lfy�؄�#۪��#LF�y~t�!�p��h�ȓ.;�$����7�`p�*	U�ZŅ�j���ai�>]D�"l�9j��D�ȓ5�2���d�(
� I;6��=8q����;�jh&�#xx��(ݴ6[�݆ȓw�L�0�l@9gBU��C�c<��Yv2|��*ټ��&
�B�����0���y�44�p�MQ�<iBGۼx�ع��ɇ����@��[�<ɑ�\�"��s@�G +�
�I2�W�<Y�`�w�aP�U/���-�"OT��⭂9_�:-Z�d�Taܡ�1"O� ���
=9�B�/}DHc�	L���;a�c�����V�N�䁷��7�<��ւWj
!�D��~����r � ]Ni!b��m"!��7=:�����D�e���Ql !�d@�rح�V�+Ka;$�+?�!�d�3j"�:�Ɖ,b8R�ÉP�!�ė(~�⠻V�N�1��խ��&�!�)FbaYe4*�H�b^i�$u�ȓ(�f���%� I�܅�W�hX6q�ȓ?ȮDs&OF+a�EE��h��HT��P�D�F4�s��DU"�ȓaĪ���.B6A�1 0�EG#����F�H}Sϝy;�h��DL����ȓ;���Ss�	S���q��8��A��h�
��O��Q�vȫ!n�+Km���u�����T΀csnE�T���m�J�;���K�
0C�	��� ��V���K���i2�Α�#I���ȓj�r��� �2O4�R%��bմ���2���
[-t�Е	q��bbP9�ȓ��e
��F�$��Ѓgk�q�����r1�p��M�8R��!C��j��ȓ-~��qhf��pq�f��?n�L��z$��Ȫ�H�0a�@���ȓHvʥ�#MZ�UPC�b�[�&`��,l�J4.xA��bT'��%�@��5��^�o�ШR�+���H�ȓKs�5ɥ��� ે�����,�ȓl����ƕ?�
y�Sj�e_V����7SLt�g�O4�֕��P9t��b����%bi/�0M�ȓ ��z�c��Q����@��"K�a��`-hh��b�E'��J�fİTJ��ϓL#�P���I��}@$�L,D�a��(�
%�!�$Φq��Q�H� ���'b�	����K��i��
�@���(S"r��">���i��e´���y�M�}�>-�"݇c�"1��N�-0$J%d�+,��|:��'��Z� �[�<�+7��L�\����U�2!<�)3����+��ӧ�ӊ^b��A�fT
=!d$�V#�"UW���ȓ�(})�-�5`���h�-T�8HP�봅·f�xCN���OE���G_;��>��- �@��V�S�#p����F�S��T9/��[�<��%�}��AgE )��IA���Q�������0ִ �6�4T���a㜍��O��(�σ>x�|�v�P��Y���@>B�	[�+J�2~<)�o�-�1O��6�ыBF��eH;!�nl�7C��Px��v�N�:��?�f-�ǣ@j�c��ԉ#��=�g�r�S�ë5�y�dˆbk��:�LA6.�i�#KS��xR��c��Xk�-@���0o qO�m�3��*G/~�B�:�l �B�|�B�4KPqQSb��$��+��0=)5,�y�_�W"��Ǎ8[2,<�!V��m���.0\(��!�ҳ�b�u�̖+	ayB-�&|�\	�rE��Kx�4R�/َո'��Ód�
*!4��B��k��]��OB7�\�5�x� �.��yi��՞��$[�Oig�	/�8|"v��[���3��Q�֝�v��"'�)�$�<Y�O�S�xs�Κ-
�XT
�K�bu�T�ʗ)0�!�d�,1���*]�NaR���
 ��I��~br� 1�73O@�H�R�P�'�tʔɴ{k��:��ψ=)rG�+<O��8��ߨN�(��<� � �'�)�H(�	G7jy��hG� �����P�*no�i~H)�ȟ���m,H}��HJ��h�) ��i��'h�+$� �)]�M�ķ;�uL�擼`�$�C#����S��YǠ�	RDBT⛦�@7?��8�����G~b��*PD�8�	OQ:�Zƀ�&�
�.�D�:�_!��XN��s�|8��<�d�7��yŉKf�y9Fc]����sw������Ǉ1�X�Zpő�2��P����{���k�f�	�{�z#}����8����g�`�p$��#U*ձ
�P[`�r ��c�*Գf�
�;+����ͳi��Ӣ. 4`�BҲ��19���65���Ӻ���ݓ)����' 3B ж��Y��h���:$p��q�,�� �M>�u�T
�!�q��x���G
��O�� ^]���"F�j��֋J�8�քB��O�1Q���Ժ�+�.�e/.|��	S�'���6ܪEyxQ�.@�&,��#_�,S��HT̀�We^��ɲ��Y����|ЋC�#[���H��<S��0�FA=8�9�m0�|ү@1RK��jV�,,�F@ ��%��FbM����=O���]�B�`ט���E��uǯAVB�)3 �6z�dI����0=�C;}�%xg��$>�z��N���jQy���O���I��Q�X�"��'��q����a��'+���q��O�aV��b�B�ZlB��4�A�,\9���Q�l�8���6��|��.��N|*%�Wx-J(��葪n�][���Bze�զ�"{J���p���e[z���`�+��3=hzq�b](�$=!��7;��1ч� ��t��F�3�?�7S>�W	�	)�������<Xt��TC�1e�nmq�:un��.H��Q���6Gy����ƾ����+�|[0�P�|�P���˙+ ����ї�W*V8t�*��p�2(��O�����'2�����N�9��$����E��	�y�%��&_x�D W�ۯ%w@�ꀤ�8�j5�f
��Zt\�n�j��V�F;�v��t%��e�@c>��p-�߼�oU�bv����ޗfW�%x6B�ɷ&ל$z2"lqV�+bXL��6�l@� �� ��Z��Y�6�.!�C�� Lrf���5Y�hG�"|��,�,�P�'N� v��GH�P)��F�P���L�("�șs���r�jE[ܴ<S�! �8��W/�2�����p�1�� !�l)�EA7sJ� 8d�']��;�x���(��AlU�F��q���w��M��?I�L�+.��]Tܧ7��nB��)Lo����e띔>��|ꆍ7��)��"�.@L�'��lnD�c�vx4��P�����V���	����'��06�4��41��T�)������ㅫx	�9Gy���q�U�!��K3���땋���� aS.!C�Q/�����C�V~~�=��N�Z��5HȴHPDEyB��*-���$�Ϸr�"5����Z$,��JN�"�})C'Boj@�)���?!��~Ph%�wLY�*����!�XI��F�<G�d�ը"�O �UfϠBj�i�܁9䌵���(�.ϻ��Dğ��~ҟw�&�!��Bݪ!���S
<������A7'�I��">fΡ9�ˀ2�������O2�͓cڰ*'$<}�����״t��i��Q�B�7�C,@��+��� p�Q��f��B�3�S#l���)�ʬ|
t��q���]44������)`���'m��� DE-|�H ��'����N�'dآL%q�@�1M��l��l۴L۔���+<������mb�'x����O��ƶŊ�hW3R�:S$m��4`miP�X�q
v4!	�)lT9i�ǃ�F���X��(3�����N��v��A_�u\��6*�ם'm�Y��ϻF��W��F8�&dע]Fp�C�'�v,��4N��4��!c7�pzЇ�D�hP���J��	�G�(YB���+Hm��O87���'M�����R�4��%B}��B��I�w��O4=��Q$hbCC�Jz����>�(�)��a�@�b'�y��Ԗ�	���*r��'q�Jl��t���9��-�IA�&��.:�Bų�cR�Y�vT`f��a�ࠧ!DK�&T���i���%"P���5z��q���G��R&
��
Ϩ]������ɴ'�upg@�o8AF�R[L�u�i�E%�Pl�ſ���A�"Y"���Y2Do(X+DL$�O� xG�J"�ˋ'=D�Q���� 䵩� �
�jx�'�M&�Γ�?!HN�Z 񫔣V�ĊP��L]�LS0a�u��N\@8�Ê��OXp´���|�a�� .��rƟ����g]�A���Y�i�,C0���L1?Y���$2نa"A����	4�Gs�'eD�x�dϫ,dSd��BD&��SN��7������Q�qŦ�+@l�X8�ԫ���LgX�ФD1A"��
!X�j���p�E(����	��дC�銠_���E��{�1[��M�9Q�ϰ4�D	w,H(a�X=c��+\O�	B�O���L�~H�-���"/��I������3�d�x��G��M��YZ�n�dM��ϋGH0!2dN�	�ɊtGEX̓I��ȈpOU8���z �3b���<ad�I48~�X��kA��Va���HJ~�Ǣ�f����ϱT�<��=�O
��!`B3oP�x�aKف��Ũ��Ш_�&5��i�l(9t����<%>5��K
���E���
�V�h;d��GQ</	X��,N�3��V���P�A�R��e�'�X6m�2O�rq���>�'g��TZG���0�P�V#�oz�ۦ�4LO�h� îw��lQ�'L��E۟@b���6����<`��Ŀ�?	 �iYƕR�O�I���æ6�A�)W�?A��L J�y�ѡ@�"��d+�b�f\�$Y�,�?���W�B�N?���	 �<�B��G�}�!����4��O��y�@�'Z"�y��b>=�F�$�c�<�ˡj���
)�!:��`9�Ńٟz��2�y�?0�O��F�g>�B���pF쀘�* v�<$ ��
4�`8	c��-�b��'�[��H�"z@��2��$P�Ё!�'<��(�DߟH �8R!+�����$���$�:C(@qcȝ�%�\��hS��'�Ȝ�!�L�V��iQ�4��*u�L�n�0x�ɇ�t?ȱs�A���5�'|�H��qw�'�(�������1Yq:Y`� g�Za(P�|� �M�T���2wP3"#^Kl�ȉ��?����ȰD W�@�glW�[]��x��t�V�n��F���I7#�!9�+s�rɟ��� ���kR50��)fD��;�ЄʕC]>@:&TW��"�t(��'����~R]����֝
W�E2�d]�V�D��� �6`ܫtMMS���jQE4\O*X�����3h����Ӹ.+��3�+�:Y��i5�ٛ�BC2*����a�y6Ļ�j3���i�G�6ŹT덝y���p��ϡ��T1��Ҳw�����'����4#�*�O�i��iɛ>�`��a�y*���m\�2�0c�a�>&j\D$�0a�i�f�\E���= _�d*wh>}�'z���SӫT�~���4�1=T2H�I�0;aiJ?"��e�K��8�z�����1O�@���˩1��TCH�;JM&�r�G$<)���\4 ļ�М>�{�d��~r)�#fG2�*B�E�jP�taR�n�8`r,C,Q "Y`�U����pI���X"͌�&x�����<� AH�aZܘ�'�~t��O�h�O��H .���kQ�@dH˯[��z��0A�%�v�]���h��!?��H�/ui�|"�K��H�+��<Q��<9�'1�����t�q��m����vAOB �a�7#VW0iX�����G$��4O�2 �S�Y1�D�
��d%*h�x�¢�|2>m�b M��?��靧+���#�öl�Е;c-J�'JnL{�M�8N�]�%�ąg6h ����jS��B!.Wz"u��<�5��?5�?��-͇פ�b��2F�j���eM4?^�}�u�'�`�y�Ŝ+C%Z��)�\�
J�
�D�ا��4Y\�&�G��\��M��}8�ѯ��B��ϓ=��է�HB�����%^�![�J�(1"�kEIY{5�p��{�$���M��	�e/�A�+B������nH-���(�*���3�+�$�;M���7㛯na�ՀՃ�*���?�S�]p�\�Č�����`I��d��4m�+���s
�v�,(s�dF���Oڀ�!%�3�l� �^��f��^��9�DFږaj�ıi_��}��s��O�Ũ') �0�����@���M�:aR/�6/d��ES9�T᳭L��� h�JA�44���]5�y���i[�	�O�8]���:\������$���
�n~���ъK2K|�q���#�)lr\�t��'���IrI���B(�Ŧ���a��F��'{�-��1�H��%QGsX��{����y,rڷga��@�<��H<���5o�&!�	Љ�%+��dO�s��,����=�t_�?,�j�,�����	�뇌����ɢ���ٴ@<~��|֧u�'�ޅ��MгewF8y��=(Q,��'��k�+Ż4Tj��$�ˈĩC!�<R�IG��m8�PP�nM��b',�#MO&�3(-LO��Ʀ	��O�]ʴ�79�n| �$X�l����U"O��X�������c�5~��p� "O$)�3ɜ�?����т=l��]0B"O�u�bi:z���Gh5t����"O �c6���XXݡ���T�bY�%"O�
T	��ZȌ�0qj��y5�T0�"O���] (�h���(Ҏ42V���"O��з`��PC|M�"��u�@�Js"O�u�H��6�^$�qFϫN�5�"Onp��́�;�>!�pk��m��X"OF�'&�N7x9��*S6���C�"O�-[�����h "IAT]�#5"O m�1�w,�ȱ��2C� %HQ"O��/�b�BVϜ"H�t͢���!!��(L��}j�CҿW������H!�d��|��n����4FH1I�!�$�,���bF��~���`���-2!��8W�R8�A�J��01�(�?x�!�ӵz������Hv��M����!�D͑Ow��ڒ!ܘ,�����'0!���r)�%�@�
ft]��ş&�!����BTYU���4��N�w�!��K]�\I!���L��S� �!�DO	f	,P鴧
 Jy��됒"�!��Z5C�f}��	��!���a䄷*�!�҈$�l�� h��zK�����\G!�dCh��}y�����]5�\��K&D�\`���D8��潅���9�"/D����&8g�@���m�,yfb�#�H+D��J���$UhiAk�b��"��=D���/Wd���!���HDi!D�4�����)2L�g3�9�j*D�� U���_-w�NQ GD�I�0Y�"O }pu(H�r�Cu�J+`�lI�"O�`���֪8�	yF��7GPx"O0����V4�M9q$�?DR�ӧ"O�l�`�V�>�0Ua�&���p"ON@�3�H��4�р*ٔ2i(1"O(a�ъ��X�kÏV68ײ|PG"O\�`�̸2,P�!\�,Ś�A"O�]B�V] ��0��A�P� �"OLuP�o�!�Œ4N�6��S "O��Wj
��)Jq�u��0"OЩ(�KX�$c0��~���"O�\����&�&�0'��$^�@H"O@���k�q�>ฐE=yNL�"O��v�V�7@����:�\Ur�"O���G�ߞ �`�.E"�*��"O(!VgU�,�����5,�NT"Ov�b&�0>��MMpi�8�"O�eZօ�9"����H1��C�"O���5 ,.>�@�!G�n\��"O(4p-��X�F�!����p�"Od���O�_�x���ǈ>z4z�"O�)�A��D���Ϭ���Y�"O�U�&'�'W@N|:rEN;:�,�E"O\��W!Q���r	��	�(��"Op�hc�Ds��؉i��n�Xc "O��T'K^@e����D d��t"O��!Ҙo�P�a1�$F
(�p"O: �vC�}x�ж�S�*	X(�"O�03u�C3[6��d�O�r �� "O��0�ܥ��Eӡ�V�X���a&"O�I�&i�>k����I�R,:}��"O��ҔA�L���b�1oH(Y6"O>�sJ�#Q�����[�ȥb�"OF@C��3S���rP X �u[!"ON�jġ"ڴ�Aǋ*|��t�"O������N��$`�e���x��"O)H���&� �Y�F,)���ӥ"O©
��B?}Lĉ��z?�yk�"OР�&d��\��)D�v9 }H�"O^��&C��[T�:��O�eT`4� "OBY҂�	�c>:`�(yP4T�*O�{�J7k����˼L����'A܈��յ	�T��LDD���'�! �EN�_d��W�_&>ܨ��'3�y;D��'�T��Qd��8�t
�'����ڇI�$�J��.�\�
�'�D�PKY5G.��i)N�R�'�@x*���pĽ��[�9
�'W�8�c��	4f�}�Q
³M8q�	�'��Qs7�$�RJ�:y�4��'7H|�-�73�� ˔A��,��'�4A2E�KGN��Gf��2� �[�'E��؃��#6��aD��>+����'�Vqۦ-�$�D*姐*#7���'W��	��$t�5Qa�O*ZfXj
�'���!���0bp�ԮB�M0RB
�'�+������FB�n���1"Ob�)���&���!�f��B�J��1"O �R�KO�'�Q+F��c
��h�"O ��rfÃ
V�A3�$O�k �-b�"O�4swd��J�(�gm�I_DD��"O����C8ĝ�%��7D8u[�"OH�Q�!gfP[E垌&�,��"O� �1c�hK��@�Zh�tX�"OL�X�m� <|Y1Q��yu�40�"O@Y��"d�H"�F@H^u�%"O�yXIZu]�&�����0�6"O��C/ Z�b �C&]�y�V|c""O�iw��'V�����-N����B"O�[e�ܪE`U�EzS(�4"O�Qd��Ll����)C.�)B "O$� 䃆	� I�qh��9�~b�"O:�jP�;GQ��9T��&��p���i�ў"~nZ�#͈�2�r��i��?%].C�ɻ��|�&'��F����o�B?N�IJ؟�(�S����F�J�:���iѥ!D��S���?���P��M.|�^�	`�$D��i�X�U�`�"#�改�
!D�Ě.�+X� �����FM� �%�:D��R���q>���(M:3|t�0�9D����'4��To��A��7D��cD��i����(�3gS����/D�`w�
�s
���A/^(��!D�L�aE��X���F�r�ذ�;D�T൨�?sh=����8u4��$9D�`C͒�]�z\��@�e��$z��5D���CƔJn��)�»a}�,C@D7D�(�!�><�,�ca�Tn^�o5D��/�24vMx�ʈ����ӧ4D���R�ɾl�z0h�� P��$ʡ>D�t�p�Q4b�B6۶	��P+��0D��3�cĕvt>e�u�D�9%&���1D��i�.Q5 �2�.�|��D$D��Ӣ�_�
Ӥ1�p���F���2� D�L�$A0_fY� �Q�At)�J?D��g�>}���F��'�6iCTO/D�P��+B �q�D�ET�0�g)D�����D�QyZe
��@)��`SC(D��2�@�g��;c�B�D+�p#�4D��FK��_���ٵbA�Dm�8a �.D�,��d6����A����Z��6D�̸��ORR�0�"!w!�( 5�6D�0b@�)H���`�f��� fj3D��@%� }�%���{��0��
2D�$s���SР�T���Oׄ a�0D��e�40�S�a��7��`1TE1D���Ec%���B�OQd��1E.D�L���G,"	�����T@��L*D��5�U�9TL��p�L�P�$��F�%D��@��ƃ~�>�r�I����W'%D�(
Q�-(�F���F Ƒj��=D���`8\��Ԃ `ϣ/_��T�=D�La��<!��Qq2 �D��uC6H=D�� fLS�m���EAPD��a;D�Ta�蔃a�A�boK�`/��QԊ4D�(q��2F�US��7sdX��%D�T�UDG;%m�(1�虜#�����#D� AL���50�+��zY�h�4�"D��!�펰.�](��I�䀃��5D��1ҪD�Nu�M���'d��#C�)D�|(�e�����@O���j$���&D����eT�Ib��YV#���T�Ұ�2D���w(H-'�L�Hǎp���V�%D���1+ډ32Bh�Wg'C,�Hj)D�X������8��ëy���c@5D��P��Ͷ9E\�{Jݟ"ގ,Q��8D��!�ѓJ3*��6�Ơ�|��E�#D�� �0,�\h����WSԉ4"O�u���R`�
t�B��j�ބ��"O��"��������D�h� �:�"O
� �Y9�Bᒠ=5t�
�"Ov�0GھO��	�P�d^Y0�"O�����]�9<( ��������v"O�aqo��l̖x�I:�\�`"O�4"�+�7�Z����_�"n��� "O܈j"��?b��qF�/@��Se"O�{��']���1lQ�\8�eks"O�� �:W��W���
.��*O�,��f�9H��䟊~�]��'us�$1L���БL��,Z����'���MBx�:�%F"����
�'�PX-�ZGTa;`�� A@��
�'qȅ��uHTy�AHͮ�2	�'�6����'PE֡J4C�k}<=��'(� 9�5$�� �՗\+
�B�'c�4��*_0A�ܰ��
E"T��'7�@�pHm�W��,�4xǡ��yo�o}v��k���hUJ)�yb�� .f٠�&	��0�aB�_#�yB*B9=媸bv��5���"�mG��y����Y<��Y��ıp��j�1�y��ڎZ0Tc��Pg�%a����y���_���:we�7 ��C7���yǕ :��Hp���W��A�E��.�y�HA$��E�q�S�ZQ�]��e��y���<| yEPj��3��y2GX�!�`L��s�DZ��yBZ;j�&LiG�C����Jˢ�y��@,q'T��IB�#��уj�y��e�Vk�(����ӁO
��y�݄!#��ZK�c��rr�Z�y�ҝ;�. ���.0�y�ŅO���g�">v(�+�y2��� ���S앨�H���k���y⥇ B�Z�aDǜ0|�Ȭ��+L�y�%��YD�r�"�����L�yW�L�R�'	���#��(�y"��/ �ĵbR��X�p`�4�yb����B�[�w`<��҂ԧ�y��̈����&!z����X�y2.ĭv�(ah��Db�(�����y.�Z�!v��k�u��h:�y"-C>���o��s��p'F�yb���uuB����ݮ�U����y�T�W�`�v. �(���y�A�����P@h�
�t���@ʌ�y�A�����K��}P�a�yRAE�"|
t!�[@��IB<�yR
�= 
���D�3[�����yR�[����ڝ3�f��aa�y��F�v�Qxpl�"�2J���y�K�}�8�2 �7o�ꇭ�(�y�.&݂��%[5n�"����>�y�Bw3��S�HU*X9Qk�<�y�M6�q��A]�F��q�L�y�BG -��9�e�.I�Ό�G�Q �y2���&D8���$̖@�FE��Z��y�oE�O.8�K�#ɽ=���Y�$�y�l�C�Ȩ3� 9��ɘ�Έ��y���h���R5l��*�1xs���y!ҤdY��'�v���r#�Ƶ�y
� :����F�&�4��Vk�F�<�"O����f�)C�Rz���-< �"O����S���#�R�)��ar�"Or��`y|S�>u��P�u"O�Pu*γu>�)g͏"'���c"O,�񴢞�����ծ�9 6�5��"O�u ���-�L�P��V"N$�"O&Y���)�
B����U̓�"O>0�3oK�E3���eAڠV��)�"O�
'ǒ�Th�����^A���c"Ov�1v��#��4(��ȨL6��"O0@h""��2ԒЏP*L&RE"O�,� ��8?��:@�
	ri�勥"O�$S�n؆M���#�(@3Tv	"�"OpL��Y#w����f_A,�A)�"O؉:3�5:4�6��1�Ur�"O�Tu�C��z�X�#	1v���"O�ɛ�L *��9��UfI+�"O�PWkK k �JP�!��1��"O����mQ5n�U�b ��o%���'hTJ�N�J���q'�۲��x��'l�� �J>V�+�$�j���'�)��.4�$t��o� (�1��'������H�!P��2�j_�a�\DH�'|	�N�d H�+C�1�
�'\��#�ڡF����'��q	Y
�'`����82�pH�䨃�7l�M
�'���V�ɱ����`b��/��	�'�.<���TB�0��\h0s�'���Ip.5���Gl\�f�+�'��0` �A�4 �!ꒉX/9��'�N����O�Ed\sF�O� 1#�'?~���	ʅGx�<*��G�Bw4@9�'�����g����e���3�\��'�������=i�)��$�P�)�'�&m@d��$WH8���s!r�k	�'�ڨr�+=8���ㅥcFLd#	�'6�����*'��01IA_��]��'���B�i�|��BΪOF$���'_V��ML#j=B�rӥ�:[ޜ��'cD-�DaįO��=��N+i_)��'s��d��4�����&Q�e����'[,yZ�Ú�W������˄Owv%I�'�"!��/�6Sǀ�G��v��H��'
NLh�nʖ4�&q�C��<z�<���'y�D ��R�B��� �H�s��]Y�'}��+c��&8gB�ȇ���rѴ	��'&R�&�ҺQm�G@��p�ZE3	�'�@����7�x�n,g�p!��'���p��ɱ:l���ƙ�Y:�[	�'At�c�޽'tj�Jׅ��z�Μ@�'q\�&#6�A�!%�z�D�0�'��P*�l�2j��݂qB	��48�'���j�eQ8CT��y����p��'��m�UI	�k�̈Pp	E�
��a#�'�.Er# =_ȸ%E��@@��'�60���L#=|�* ,Θh@�	�'����.C�?y�k�)�.`2�'n���@#Q6:�J�-Ŵ?����'�d���k�6b2-�+�bAx�Y�'��t��[]�8���˓ez�'�����90oT�6�[���q�'�d��vؕq;n����DRm� ��'+�U2щI,`�ؗe�D�t���� Le�����>��A���8�D��"O�� �W�+�pL:T �#R��(x�"O��Y��\F=(=����9ey���"O���!�l|����>T�t���b�<a�aԓi�S��/�`���`�<)%�ZKL�R%`\,t=�w�q�<q��V�<�h�6,�G�J��N�m�<9�Ѕ$ܚJ�P�6.��2�ǒD�<��c�*Q�QXp�_6~Lb��A�<�"�� l�D.K�o�\}yq�H�<�K��7W����F�RӰ��ǥXY�<�@`�qM��*����zr�X�<�@��
!�tyd���S�H�����R��d�<S蟊Z>^�Ҡ�5��G�VR�<!S�C�KU~����K�)p)З+M�<1��G��&䂵���Ci��;!�C�<���W�iIƙh�%T^�^ă�U�<��P_��`cB�.~�Ř�.U�<��Cĩ���gʉ!^�|X���T�<)��ߍ6����@Q�/;B����S�<iEi��] ��_��mð+��]E{���ix@�r0��	?yn��'b<��8�	�'D��@��!	�>��bO��		�'O�ڔ�Ԯ�ވ�
0e�@J�' dq���D8zEӠm +д��
�'w���§Z,o��pNH8/��
�'
�Qg�|��!hg.&J�U1�'�& �&G
+m�B! W�I�4�lB�'��$���/��=qQ�΄$�1�'�MzТ�S��|�@U�	��'XFD�������?�8��'a�h)&��j%d��g��:��X�	�'n���t%��w�Ȱ�C$	8�@y	�'QJ�g�G+zZ&�z��Ш4��l��'}h�C�*�b�	�4)%h7"O�!�5�͍dM*xbDK�|N�T��"O�E2gk�"|a�aꋧ~8�� "OZQ�W�µ�(S6�_,SHp��a"O�+���>d�d��gh�;G81�"O[�H�q��QG��5Cnq��"O���-Y�H�{!,��PK�e�"O���P��*�$�6�P@�נ�T�<�g�@(l��3�)�
[�`�6[�<�� B�z����<r`vx	R)�@�<A��8��[�� )���t8��'�hxe�0`Ò�BM*��!Yr�5D�Pi ��Q��ph%INb��y6�)D��L9s�ଚŨ�>6�z)�+,D��!��&AX�I�w���!)>!�� 'D�4��b����(Շ��H����2D��mO:Up����jUL�1��#D��x�N��u�Z�Z�&_��B5 ��?D�����)KZA� �/,Dc4G2D� �7$�|-��I0"ۚ
�4i!d$D�hg-�*&p |��ձO��8���"D�@9���Q4�dҍ^�̸�O D��B��R�E4�����Z/%!Ā��M<�O��O�Ȫ򴰉��Ai6EZ'EI)8�!�D"�@ij�bƀ[,��"�H�!�d��T]�D;��	Z�,�o�!�č��H���ӲNH!c�|6!�"�"���h��4�	��$��'!�d�M����`ƾN��"��'x�!�W:\!H�<�0�S`��b�!�� (�E�+1(P��/ױQ��܉�"O�(᧍�x��hq�iԶ 7"O0�8��J0!�l)�#��J� Zf"O�l�r�@3:�1�Cȵa�"O��Ǧ:O`��K�3G�q�"O2 �D�&^z�s�D�Y�tz�"Od����K���B�߳���"O�����ܤUm,!1���R�����"O��`�(��R��=R)��+��y���&u2���Q��^��C�Q �y�@�-r��Q�ê�,"&���G���y�׈"�E�fK�s�D/>�ɇ�!����EGL�Z͢Q,���ȇȓh?~��k��a)��)���/)�|���n��-&e��	,��tC��.Of
C�I�@���.]u��#��%zC�	�F��I+@�*̓�^���'��Y���
�F��1:"���'5>�ڤj �oڎ�b}:���'R�J�	N��a��%rNr���'(�0w*U5_\��ҡ�?@*�y��HO6d���ؕ_�~����]"]��9"s"OƄ+�IL!z��h��L�(B��!�"�S��y� �ni��h�B�$ǜy Ѫ�y��l�)Q�'�r��0镤+�ybB�20��D���9�%����y���$7`��I��bQ<���g�5�y2�քa�_HA�嚠�yB��)xb@�5�n����y��ה���E��������[��y��C�}X�$,ظ�6e����y��tl�hf��~z&]�&
����#�O���ŭg��T����O�L8�"Oщ��^�V5�=��#O.�����"O\��ph؆A�"%{�c]�;�6yˠ"O��{u)}F���7
��I�"O�i؀�=0"ɣs�يi��,Q�"OX1��J�TJ��+��S:����"O��˰�����u	P�R�j�#�"O�=P�c9�a11HJ�y��0D"O��j�˥feU�4�H+3[JA�"O���5���'Y,҇��U>�a��"O�u�GLI `�t��v'�n�$0yc"O�h !g��$�wf��è� "Obt
�O�fz�i�����"O�U[3���F�`��J���%"O4�Jdm̨e*^l+p�Od�l�2"O %R�Z�c,�Q��V9M]�,��"O.�;��;LP9��C�E%�T�Q"O���q�
*({T��eÕ�# �5�A"O�0+��h��@Q��c�9"O��)��̮PljL�=[����"O��bĭ�G@��" �,\o�� W"O\����T�$<�NFJ:H��"OJmy�H��'����N-h���Q"Ohp[aM1� -iP�' ��"OH\Q�#�)T$flӔM�2Y�"O�1�d�2=N$,jA��`'��"Ovlb�wB������70B�c7"O�|�D`�;���)�'�]�"O�S�aS�e ��Q��I��bd"O��0�	O!N��sƇ6i�
%�"O�@�QL�r�ΐI5_�:� �#"O�dYPoJ	%:}��	��&iyC"O� ^�9� �Pl�<ࡩR�c�z�c�"O�=�E�X�a�4ٸ�G\�B�����"O1�eJƷ
*,���x�2��"O�URc���;��Ը��O�p��"O\�I�,�.�`8HU��<��R�"On` &�o��0X�b�%s}q��"O&�C���9�|(�$�Y�X|D= �"O�X�F�Y�q��L"a�QpN)��"O�a��U%�HY��J<�"5"O2����ѳ0�ް�v�T�l+Z �"OP��th�){􊽨V.
$8��"O��E�K��2  U3�R�����[�<��a�-^7	�fn�q*8�8�K�W�<���!������	v���w"Ot��Vln����+)4��T"OXpYeQ�����(ʔ, E�"Od�Y!��0� +��\��u٢"O�5ic��2&"iȄe ZX�"OFX$f��74�͠Veةs5Ȝ1T"O�4Qf	Ëzz� Sa�صfQ؀�5"O�tIVd�k&�h�ڭjI
��"OعK� (oS��U�t��{�"O��$�oL�a�V:&���"O4]���������`�1,b���"Or`sC醏�Q�Be��y����"O����AɄ-�,P�D�]?>0�f"Of�r�ˍ�Z��i�D��)����"O�S錢swl;�B�8��� �"Oz�z�T7b0U9&�ZwӦɩd"Ox��SE@�)��-����^�By�B"ObH�d��*��t;v�	�D�u�"O��Z�h $��lX�7
L1Sp"O�PQ���.UA$���eI�� hX1"Oe(�F��O���E甦9n�)!A"OH�e�� A���Q �^c��K�"Or�)$�N �`��h�sS�	�"O�p0��P�I��Q�VHB�=>��!"O�T $�8`��L�Uh�E��9Q "Oȍb #�>[�� �7�ϓV���S"O�гm6�nq	��J5+#@���"O��1�뛬�քC�`��|�<�9�"O��`�	@H`��Q�J�����"O���MU��eȶ �)R�h��"O�L�3j�IP�U8v�EG,y "O�M�4��N���q�I	n��Ա�"OV�b�n��Se�e�3v�`ca"O�Xo��K��ٓ�aA3_X9s"O�h�g	�*�j�0�^��X��@"O ���B�@ITt�q�_�s:���D"O�{0j?_�d�q'��ք��d"O2��b� ja�̘&	J�^E�"O�t�u��k�̙k.G�k��!@"O�@:�܊,��L�ƯG�w����"O���E���@ei����X���"O|�0$�<S��dX���N�,���"O��� �E�$�$�z�$˒c����R"Opո���1o0��yA��1�XBt"O����.[ry�6��R� t�3"Op�	IJ ^�ք 7f��
�fQI�"O�-@䃕`��AHW$];S�&(�"O5�!�D�JܹA�O�z�\�`"O\�C*'+:�cl��Inj%��"O�e���  jT����(Z�����"OJ�8v��l
����� ���U"O� ࠺w I�>���@RՙE��R"O]���O-,�"��`�	����C�"O�83e&�r�������Z�d H�"O����OQ

qdst�D�����"O��Cf����4��Y,G�
�!�"O��k2��7v A7���ֽ��"O�U������#҆�.!���D"O�����nX<Y$�μ|V�h��"O��`�& 3/8L��G�@#KCt03�"Ol�Y�g�:b�tI�,�q�\��"Ot��
G"z\�)rP.?xb���*Op��AH'%�l���~��3�'�"���I�R�",�++t��Q�'p}X�Ƴ/��6o��)?ީ��'���	&��EM��'�/$��5q�'6(�5�̼/�^h���=F�����'�La ��!]H�ć�h�
�)�'k\��0M�)H�2��%�B$g_`�	�'� ux���$69R�Ѕa$S~t{�'��H��%�3���j�/K b��q�'�TӲ��6�~��BY�%���8�'s����ט)�ѱ �#�I"�'O�9�wAM�	ݤ�2Ǭ�oL��
�'�Z|#���W)܀K�CG~x��
�'�h-��m�M|6�h�)��i.��
�'��;6*�N����d �;
�')�Q��'|�>����$QdQ*
�'(�q0��"��HK�k؄��Qq�'����.P�ipZ�2�����>d[�',X= ����P�taB��U|r<!
�'��t��;�d�`2+	�\%�Ȣ	�'} ���%% ��aQ�ѩT"�B	�'`��w��!̾p#����:�;	�'�2���� H
!�� �Tp�'׮8!�C������9s)�(�'B�EC6K�5_\}��R	\Uz�k
�'�(T�@ ��E2n�
���8� ��	�'N���eج&�6�8���
�h�'ΐl�A��!Tp�ly���!1��Q��'%�DjӪ�+v�43�#��U�2�'g��H�jvCЅi�^K���'E��H��$n�E; $��n� T�'�\�r(�=G͈
��2�B�!�'g��j��ێKz�A�G�Ҁ[�IB	�'�J��Aϖ�(��,�VB�R�c�'@�X�J�2�TL�Q镂Nl�Ԉ�'�YRc��\�|��UJ�?5����'���9¢X�D_��% �@����'����a�FԀu�%����'^�l��o\�oQ�(�l�*la�''l�С��G�T� �3v�h�'�N2��ɾ�TLr��[�l�;�'f� fGV�n�A���;.>0b	�'CZ�	�IE�����M%{����	�'�F��i�|\�����^rι�	�'܎4z`�C*i-*LSe�U:Sef�	�'���
�$ի.��q#�Q����'�A�@��B���2IH @҈��'�4ٹ3gǾ9S����	�Q��'�B��C]���uc�l�
�R�'�IK���lڷ'�9f����'<�Y�(��!�&�0��� �'��I�� [�4ɉ6h��t��'~&8�!Ը<��0�R�uwB���� pA���S���ɴ�ε
�Xh#"OZ<�5!S�~x\5 �45�ڬ:�"O��RH��|,%0�&@��U"O�x�e�ߩ4��y��ֶn���f"O�)�� �JD ˳ŹXV��r"O��²,��}J��s�A 2愢�"O U�S�,�\�2�o�X�\4��"Op���E�.*hJ�.�w�z��"OҬ�v�Z�r�M�8#B��7"O|A�7�߮)�j����٫U5Ȩ9�"O>�3a��!fV���C�jFىS"O�[W蛕A6�3�n�*tXEPG"Ox��������ٵj�Z��Тv�<���0�|����Ej8@xrFu�<��ϊ.��0X��ı����s�<�aᖎu�4s��X):��5���o�<���K�ih��po�"\}^�۵@�m�<�"GҪz`�(b��	� #�	�<�G�2xyլ�V���;ՇXa�<��D7Ƹ��vDк+�D����y�<&
�m� ѨA�̯6�~����r�<ᐂL�|�����(���b#�NX�<� ��)	Z�%:��E'Qˆ�:���V�<�&��%��D�q�ۋ]�`Z�)UQ�<9�B��`p����E(�u�<�֧�}*�� %HlJp�H�<)@G7�F��ZOfΌCEo�<�墂�{���8D%�>vE�p�S�i�<i�⃳q�֤�,�0xi��S��b�<��E� X�n4�cMRj�\h�&��U�<	)��DjXq#cΚ��1�U�<Q��_�V����F�
�
,���OZ�<�(��&���ic�!A��y� L[�<�7�вH������M'zc<���|�<���^(z�RȊ@JԠ6� ,jd�o�<�ʎ�*�z-Q���� Kő7G�n�<�u������PS�eg�<�Gۛ�Dy��TA�V+cEzX��f�Ȭ@�FA�5:Di�g�BN�ȓ{נz����{����Λ�s�j��ȓO�8�v.�>xt)�g� +4M^a��ς[! ��qY���?>����LO~PF�.,����wIZ$ ����ȓ ` �a�R�R�"����e|T��ȓw_
o����B*�X�ZI��2F�	G,�� x!��b��@5�$��h��E
U�W
R���4�U
�8�ȓ)�X�tΎ8g��E�z�܆ȓ0�����v����c�eֲ͆�k��1B����l
w�ЂX0Nh�ȓ�h�� �=�~qÁ�O3+ZL��Ck��YW�J�)=z-KС_�bP��`͆���-=FIԔ��*�i�H]��Iz��E#�.m�af�j�Z��ȓA�yB��2$�B������� �ȓQ��zP ��my�	�3��!
䨅ȓ,.����2Z:�9ԃśH�P���r��0�vU��Qa��Ӛ1�B\�ȓq6�,c�O�%O���T�L�AO&��ȓ@WZ���̃+��R���_�\���Y��1q)�>�Bw��E�����	R�̠$D6!���B�Fj⡆�4�VU+�n	38�L�8��ȓ`|�2T�>t`c�]�m"L��	{y
� �Z0�9LI!qB6f����"OFۧl���L�aE���j�"O�C���2�N�AQ�J�W!�}��"O:�#ϙ�W�
�r��9U���"On��C�Ç_z���-�:\�a��"O����*N']&���*��Sw��sU"Oڱ��n�"l��c$��!$|�r�'��������M, 	�3'U!	�(�.?D�hhwB�D�AɳS��FAÁ
=D�Lk���(��$���K�X	;��7D����ǜSL4���Dc��T�d/0D�@��T!>�4�?Bl���.D�h��Fė@\T����Bg���P�(.D��)���< �3�/�RZv����k�PE{����Ol)**�,�����MW��0�"O��j��� �j��׋@�m`�"O��D�ͣ8(d +sɚ�K�Z�"Oj���!/u4|�`��~@P�"O��"���15�^���nz$Xb"O^J�!�� ��Lr]]p�a"O�0IF���2���oO�&[R�jb"O��#b�I��\Ђ-
YX:(�!"O�� ��P�Zg�{T��#4�5J�"O�-J!�P$����!Ҧ;Ih�k�"Ov�I��.y�hŀ��Vr?��	6"O�p˛� ��쳡���t�`E"O,�J��	 \4�ar�E� �"��E"O攠��Zg6 ��FM�"���+�"O��y��$'t,XYD�ɫg�4��"O�0c!ʃ�T�!�%O&}J�A��"O`tc�n�>�D�+�5DE��B�"O��愐"<�#��<0HD�5"O@MW�ƙv�P#U�^��*Q"O" ���ػ&.���5�5�"O�����úS,��P��m�@"OQS�G�%�\y;&τ����15"Oj(:VCʢ �yJ.��.�j�:�"O���nW�4��@#��+Ȗ RS"O�4�w���T�N�pPH�8Q6�X�'������@ =|�Sl�,8lh�'$xl���,cK�HxgQ���h�'۸�[Wj�hi�g/���
�'���b�3UKxy3g�]1pq6�+�'�J!����/Eۀ'�χg�ΰC�'�Ę�2���&�p��JҴa�^�q�'%���ⅰN��T�,��
���'�l��e1A L�g���.�3�'~0h�AC@�=tЃ�&E@<d�'ձ�AƼ8�h�vI�B����'ޘ�)p�\�I0����g4)�
�'(F��ਉ0=�ش�f9\x*P�	�'�Z����3x�tY��&O7Z�1	�'�&թcG�v�PPpG4M����''�����^�x�7��8
1��'�&�o�.���WR�E�,��'ب�(� 4�٣-
��
�'(��)1�i�.%S���p�S
�'?����k�5|���	�'۪q���k	�'P0�{c��.Q�^�ubG�=�BH��'�VD�#��8#��u�T)48X� ��'p��� ��:�m�@!3�lЙ�'\,�8g�G"`����$A��{�'��}ˁ3�
(h$G��-� I�'�,� ��D�RԊ� ��y��� f�s�u��p;��i܂��"O��!�G�2D���ã�I��pj�"O��da֝h%:̓��]�t6X���"O���Qi�{ ��H�`�)H:�)�"O�xg�DxM�0/]�w1��"O���%�(J|���KA 2D�t"O�Ȃ�"������l����"O�� ݱV-@�[�`��5�^d�"OJ<;B4U[�\a��8O��1"O ���G�L�ѐgaL�7�8<@�"O6 �� 4p <�Qf���\@(B"O�`�DĂ~2���L�	�M1B"O�eƇ�o���c��.�h!Yf"O~�1�j�gol�Pv�#�4�"O���7 �0z�6��!NŊ*�>� �"O�D�a�.s�*�1t"�"_�J�ss"O|ġD��+�^�5#	6����"On� wB]�!X��-�h�����0�!��(1���-��f`I6)F�!�Z!K��!�r�B?}��4򪔔�!��P=V�LȜ^Tzt�u��8~�!�W�;�����O��F�p+ N�c!�DI GL���,<�����7E!��w�(�i��Y�e�z���@/L!�W�P���#��.l�r�xZ1��U�ȓXXhP-�o�4l#�k��w�-��B��c��;p@Fذ�Bz�r݅�/`PQ�n�1��x�����P��8#Xs�*$B�Y a�"�ެ��p�PXsk͇4��9��!Jmt��!��P��%�$ G00��в4~���j�JĘ��=Ln �A��Ʃ�ȓ,�lݠ��R��$�!#�6�: �ȓ]��T����43�Vc� <�`Іȓ!�LJ�뒆Hs����Z��\��;�j�`S-�;pJ2U����2Dm$4��<uP�e�-*�X�V�[�}�t�ȓ^��rF'؉x��1;��B#-�zA��GPf�TnDe쎑BF��8(ʴd��~��3�[�˶��E���>0����.u�F����C�0 �ʃQ�<���S�	I��^�d�sR�S�<�'�[�w�4�B��_�/���O�T�<!����UT����,X�tU���Z�<��5zrEz��OF�5�@{�<�(��rѦX���E��ra�t�<	��gV�\ʵ�2P�2�n�<фj[�\��#cK�x*�B���l�<��JҠ�����a6nD\��]d�<��CY5)�JԸl��<��p ��I�<Y�f8,J�!Q��Q��yVI��<)5���j!���&W�w/8�֣Zz�<���Â]�T�k�`��[�i�R�K�<	���� Z�̘'p��D��`�F�<a�EX�zU��G�e���`�C�<�R�{��z��\�,�@сJ�<�&�,��c���-�\x6�Zj�<#�_7��bR�՞��KӇGd�<�U$�:ݨY���כ}��"h\�<���b}HЪ��X�e�
�����T�F{�j̆+W�QuF�a��a����yRC�<���i�mՓO���+��y�H�0)��d�Sc��x��f���ybNN�(��1��C�X΁/	<&Y��S�? ��@�R�q�v��.+Ha��"O�	Ѓ�����:T��z���"O�Q����>B�(�`���oi�H*'�	cy��P��9���H�ʁx�E]Te�B�Iao"�YF+��Dh�	� W��B��g�n]z�F�5V(�gF��jV�B䉘gBp�;�b��W"�"��,e�B�I�u�zl�.�<Y�ZE��I*	�B䉌J�|���ܴX
��cF��=��B�I�� +�)]b�.��d����TB�61�8�q�B2j$���#���p�RB��L ����F�+���hfޥc66B�9L8 ]qBWkh�	�	�4}�C�	�sW��2�m�0|:C�JG?9�C�I�_V����A�5�`�g�C�I4B��=9���A��8�ҡ��V'rC�	X��x�d�+v_����뇁�"C�	B�� 0JE��b؁�!�I%^B�I2{�6�+�Ut���)��c&B��^�i�&�ݩp�bt��_^B�-qhq�#Ȁ�vt^���_�B�	�*L��f'��g�F ��aH�U�C�I�0v�c#M�tTx�u,C�}��C�	�mR�ې�W%w��l:���2�C��D�~�HB���h�9 "L'.��B�I/u�I�$ٚ.�I�J��M=�B�IZ��PҊNp��p�M'��C�	�w��!)��_z̡�-�A��C䉯����0B��aRp��5�Oe�tC�	�-w�d{'�`�n�:Ę�\
C�ɢ[uH��W��F"�����l	�B�I� Sv��cO��%��
��KX5|B�I�G�D`�RW</F)Q���#�pB�ɜ2�paR�"�+@9���]B�	!`Q���t�Z;�$a��S "�DB�I>)*6D�c,�910F	c'm׾�@B��+t$I��G�W�0E)�ϊ.{�B�	�	Qh�[EYNMÄO��&,]i�'��cĞ�u�Xr�&� 14��'z�	� D�*����sF�#F8�1��'':���5������
t���'�F4�P!�1��9�R`Y�n�P@k�'��i:�jˌ[j���H�j�]�
�'r��a�&�2ݸ��Z9&Ld��'��L�����';,`��]�ِ
�',������a>n���cG�ct<��
�'^�<� �A�Cf�d�C�� jg��	�'���j�$I�rc�q����'�}i�V/X�����+��d-� �'��0�UK6ہ��\da�'��2Ŋ�o�Phx�D�W�N!y�'G���t�,��(&@�=��� �'e���/�$I���5oK${6��
�'-ޤJЄ�?���M�(�a
�'}��
u�^&a�,���&W�Q;�'?�E��XeiG�I?\l��'��V�ݯ3R�i90oݹ3�~y9�'b1���|ȫ ��+����'ю����ݝL0\2�Ls?�h�
�'�b�����bW)�B1&a�'��lAd�Z�[�^!�Ql��@q��'�$$�⏆(��� �$u����'6�Ձ�jR���M�@�8��'.��p㚈y�IJ�MǊ5zR�Q��� �pA�S�K�,��I�8�-�2"O�A{'N�2jΘIJ�R�{d"Od��р�¥�T
�!����"O�;S�ƿ8Ԑ�[����D�8U�"O|0Z�bZ) �����Oŀ�X�S"OMYĊR5g���S�.A�~Q>lK"O�41�Ιbl� ���x�Ԥ�'"O�A�$���A����s�"��S"On�5o�Фpbe�1�DQ�"OL8��nI8
����6��V���f"O$��&�nT�1�BH�Q㈄��"ORx�cJ	a��11 �X����"OҍB�d��*��)�e ��7h7"O�XQ�Gq܊�3B/j�j�R�"O>�耤�8=��%�'��!�Nܺ"On�SF%��B	��.��e�Ni��"O��(rCϝQ�PЃ%f6x =��"O�4�W�������<Y��À"O�P[��@'O�j�A�ԣC�-b�"O49�dW>�*�3�H̘@*��a"O��g�'9�f��)6�s"O����
�"�>q
4�U�lxh�"O.�C�9LQ6���1�FyIR"O�X�-(Y�|m��iܣwy852�"O���B�	�¬�5��'yd��&"O�`A�[&/�qY
3#P���"O�!F�T?JIJ�(^�-��e!"Oni� N9¸R�e� �R��5"ORm���W�U�X�cV�	l4��"O�hj�)�� #�[���^��թU"O䴪4�Y�cC*9�0nҗ(b4��$"O�{��S9�J�%H�c1й"O��ϒ \����M��.�v8�%"O��o�7��c�+8q�<��"O�tQgV����c�J�P���0"O��QCu5n�A!��$Vm�\X�"O"��R�C�:�H�bW�6d@���"O���0[�h!yq�~J}�a"O�	p�A��@<�;�o�
>_h���"O�ER��BI��x���[B:��t"O2�)Wǁ�Bk����&��SW"O\D;t��j�"<�0Ă3�>�#�"O頲mM�x'���"%��K�:A3"O���򆓨�ddK`d��V��"ON 3Ў����K�L��|*"O�-�񠔰p��q�`ft�:�Cq"O�%�܂	��ܛ'�C�]�d�g"O� 
w�䜨!&ߔ`T�m�a"O��i��R
N�H!�'�x,,���"Of4*G��n�9c��[�n:Љ��"O>�� L,7x�H�j��j�9�"O�A��E�F����UǛ,/)t�:�"O&�nɂ`��	4DԹM�l��"O��HQKO�_�n �#Y�2(�*"O�ً1V�=x̱��D�3
MH��"O�	��FO�Uq�w�S�c;> Z�"O�`1KM�2�)�L	&*��R"O9Y�����@p,��8W�!�"O�5��b4v��8p�K��B;�Q��"O�˄�_%T\��%��Jf"O�yc��I���1�
"�ika"Od�z򬑄x�鲑��_ �"O|-2i� ]F��HR>.��P��"OܩÅ����^hWÏ~B�z"O� ������v�b��d�H�k�"Ov��^�|�̠xa+V;;zB�ò"O~ȹv�U#y�^���C\�Os�\!"OR�C�HF� rh�2eE�Q�"O�h$�����%g[�
lB,"O&�	@�G�qC"Ls��՗\~!�g"O�YK�B1u�� ��.�v�! "O���%�bhq
ԁՋd̂�k�"OhyEP	t���ţ�7�|��#"Opy�d%�l�� ��GXy�"OR)Z�� 9�J� �^ZeD�"O��H�"�58sn�E^Q�!z�"OuJN�ZT���T�ǵҌ�3�"OZP�Ԍ��|v�a���5��
�"O�#i�1p�eJ���>u�^@�"OZ��Q�K�)f�iz��g��ȩ�"O,���E�.�l��&)��X�����"O|��$lS�C%Zq3���VJ��"O8e����2��c��k�z�26"O�Lka��[���1ƛ�L��{a"O*|���-"�,�6��al 8�"O����x����.Sf*��%"O�P�ը�=x��pA�]�'����"O��S杬R�赫�O˃M�"O U��H��F�b��ρRJl��"O�pI�J'a��Вaכz�"�B�"O8p���3���"�G/��!"O���S�\E�J�T�A"O:A�G��8�N���iZz��9�d"O"Ɖ��k̜(â�μV��Y��"O2�Ѣ�O �� F)����U�"O�d���S�O8@A��-!W��T�6"O2H�ӧ�
++��,S7Dޤc�"O�B��!:�}����}:t$¤*O�V�6'��˥��)�&}R�e5D��+�B_}S�0�+K'��j3�2D����r�ޱ���h���1�0D��x����>�X�$��B��P�-D��aA�M�̹C��N/!�ʱ��-D��`7��W"z���L�=�i�/,D���hܓTG�h�%J�hY"�H&D��3&�[/R��c�j�T j5h��0D���u.�#F$�L S�Y YgB�2�b#D��a�C�>��E J<z��a��%D��y1��*�� �0��/iخ�X.&D��#tK6
�F�!a)�	nPT��2D���3f�2!���+P̉0:8��(.D�4ô��a�E���=�Ȱ�n8D��z3�F�9�F���c�H
 �+�8D���`��?B���@�R�Fs($��0D�����&,��$hOS��I�3�3D�|��47����Ł%+��q��o'D��	"nA�Ln�F"�%	�:�Xc�2D����_,s�e	�C�[Plё�.D���Gn@� ����E\}���#�*D�H��&�c�%��ƫ?ں�	�%+D���p!W�o�L�w� !"��sv$D��B�,8n��!�Ԩ�P�`�+�7D��1���-�#_�T�I�]6<C�I�I�KT&��%�
�0H�%w�\C�I;�$tIf�L�Pg��DT�W�C�,4��Ȣ�,�6��ġ���:UqHB�I
��c��:B��p���6!��C䉚b�T�*!悾;�A���Ԯ8��C�)� ���f��7z�sQ���'A:u�"O��YgaL�>�����I���5"OtC)U5f | 0�0&�<���"O~L�ߗ8��i�S�[T�t
�"O>ؘfg��0^4P��M�^<�k�"O6�ʠ�(~b[V�46����1"O
m!֭��Q$� �μm��"OVabG�u���Vn�8�}ib"O܅�ê[&$��ZwL0d/=i�"O�|�A��}#V�*���w��$�Q"O\��m�/�X�R�U���"OH���K��:�>iZĄM8#�<HH�"Oy@�HN&3��)!��ߓB�4��6"O��P	�W� 00�G�c��l�"O��BG��a�X*�U>!��"OB9ۡJ�:"�b��8�X�"O0��
:},%�Q�ˍQ$�4��"O�`*�$	�D��|� ��=Z��B"O>��@΁>Z�����ϵ!����"O��6@��t:iRUL��v��sf"O�TA6$ �~)��%�Rm�9�"OV�
%�§Z;1�vČ�/Nƽ:7"O.���/
I��l�G(/�HaQ"O���	Z�Z-��@�MX�6�̸�S"O��p#,�^b�)"�,��C��M;�"O�� B�N�N,x���&�:��"O*YVJ�Bl��X�+|�B�"O�-�j�g̪1����i��1q"O��#��8�z��F)�TGF�`"O\H:ˇ
l�6-	�)�R(����"O�8��ޢS� ����ޯ^
F�p"O$�i�+����!�%���"O Q���^�[��yZǈMA���	�"O(5�O<�f���)�|�����"O�Ip�Θ	f���A�&�¡�c"O Hc��	%T4�E�#�]�Lx���"O88i��Y�`E��RL<�Qr"O��Zg /ﴹJ@m�;Wj��4"O��h��7)���t��1a�dA{w"O��2@�8*D�0�6B��'x��)�"OX�BBF�Ѹa:���*�$�3"O$�k�i�'kz$(1J�fM�0"OT�:��D�_��Q�䌱Z�t�SW"O��P�k��yxQ(V�;����&"OZEH3��k�"�A6�/-1�*O�irVg3^읳v��)�z
�'%��u Ώ$ ��E��nH�<!�ퟷlrF/HM�nP��h�<���I������H�c&p���j�<�pȀ�p�tI1i	+|���h�<�K�2	ߴ��iWWq���$��g�<i���A!N�q×�)�64x���k�<1��\^��Lb�F\�ڽK$�r�<�v�!��zVd	J��`D��m�<� �;T�
4 ��BT9���g�<�a/H1[���L>P�� ����e�<Y�G�,!�*��uf8	���ZX�<a�θ8uNTXcg�0j�Q�,S�<	2i@�B�nӃ��mR����R�<��%
�{�ѣ�jK9Ո�炞J�<1VOC�j6H��*L�2�i��OR�<�e&��[�����&� ]��|�e�R�<�d�Q/|J.�:~8hiu��U�<��Cʁ7�n�S"�Q���)4z�<� �� �ۗvȮ5ʷI3M�<�x�"O�,�v�W��@T��Ѓ;�tya�"O�x���Y�m��(�	0$}lm��"O��v&
<��I�;FвXq�"Oε�c�/�~틤�A1+��1��"Ol�ӌ #tو �*��p�W"O>�aw�14DF��gG��}D8�"O<aR�쑥L<�dфƋ$3p����"O�����)_�p���Y�	M����"O��@�Q�4q8�1�5H��i�"O~��*O�0DꈘE�[A���"O^a���#]�>�1A�+#��8B"O�0@ߔp5��s�[�:b�3u"O�
� P�4r��b��5R�8{�"Orb"�&FP�+aO��;<�-��"OШ��ĶA���ROˬ� ��"O�Ы�cAu�ͣS���b^�`��"O~H��P;X5&`���/R�-�c"O*i���%��ʅ-J�E6�=��"Oޠ��B�L�L����0B�"O>5�Po�?_fͰBIn�z٢"O�m ���Q1�c�[�^�K�"O°�/hRx�caT�?\��"OxA��hɞ]��1�FϛV�Mt"O~��%͋�C�����%�k�"O��i�MJ�}g�=3�*�z��8�U"O�!��i_@h�Pa�)�t��̊4"O��ö��m�� �
�" ��KF"O�U ��^�6�~Q8wdA�P�8�	�"O�B}�v8Iĉ�>5��h�"O���#H�n��(���[���"O���kH���8Y�j�J�d��"O�%�	| �剘�vj��4"Olh�4T"nU��� �G�n� �"O�۵o]5+B��H�I��yd"O�M	��߳ǂh@�Oy���A"Oh���Z�q7�K�"��x�Z���"O�yӥO\��p��-{iZ�Z�"O>(�'�0����FN A�#"O@	:@��#D�'!��)j����"O�s7`/�6�����@Zhl��"O�$��(��Ul̄� \6d^��*"O8��W)��z9*��ýet�qCB"O�!�dɘ�@bY+%ꂤ|q�DI"O�m�wOS�'5Ф��?s���#�"O|=a��B#�T}1V	5�н� "O9@����\ŨQ�a��3+�4x�r"O���h�?V��KH+`���2"O���U�T\^a��P�*-@�"O�E�cmi��]ul �1"O����B9inl�Q*=B�a�"O�y��"���FbP0�"O��(�a/T���4mL�-$�Y!b"O^�[�g����kPˋ�Uu0�`"O)d��6j�����)Ɏ_�P��d"O���W�_�<�Zx1����(�H���"O4�����X���	��iPP���"O�}����貰盁$���'"O<�2�],k"�Q��i
�a W"Oh��f52ݦy���'� �7"OD��BH�%ZD��җj�Ѕ�D"O�]�s�<#�"�)����7�=:�"O�)�PN��	�
pq���Q�ƥ:�"O(�(�� J}��� ݟau0m��"O� �{ǈʚ�Ȑ-Z�CY����"Op��';"sh�:'MF�iG��2G"Of�Y�GW6fI✹WNL�^��l
�"O�@E�T(\�"iq��I�5��A "O���	լ5�P�!��&��"O�]�C* ;h^5� �Ư>G~��%"O���M\7?��(�e�"e���"Ob�{a	Ѧ?�|(�UD�Ga���U"O����j�"jz��R1��(D�u�"OT��JWP��d���W*;��U�p"O ���pB�;�B
/ m�"O�@��]U��BAƷ\��س"O��6,��A�A[e�b���
�{�<���3; ub���:�@DeDu�<Y3䝹�t�B�H�86h1���p�<s/	?QP�$��Άt��i� G�d�<y�	��!�l� �����K�<���%I��t�b$��v%0MZ��n�<i��Fc1I�!r����f+�o�<!�fA8'�tc��]�)hl�`�F�g�<��BI6S����R�&kc��"oN`�<�$a�R��TX������8�r�ZZ�<9t Si��QX�%��8��Kp�<ɳ��M� CR+��0��9�w�<9c��7�tD�U`I@TƘyu(j�<��- �A�Lï=suЌ���\Q�<�&����� �R0	N �֥XL�<�c�F$Ne<G�L]�l�B6��F�<�B.#}��d6瑇~P����y�<h7Q����f�j�R�r�<�D�
q��`Iq��uڒ,�q�<��&�66�8��#���{^�[tD�F�<�Ī +!�Lx��S�j��pd�E�<����f��|�g�(h谪�A�<q񍙋Dt�	�˝�[��=��|�<!`D_ :c�5[��86��0$�t�<ٱ-�]N�zӨ��}���ht�<i3���OH��ɡWt��!p�<ɑ��
s�RQa'L!0��@��i�<��g��d�f��:��#�)]n�<�$��y#Ωbj (Z���Do�<�$@V�u�8�ʖc@(�'i�<�Q@��4L���Td�_�l9��^�<�T�{��a�U��_p����W�<IV�ם�%Z���80��V�<��&�� ����I��=���#A�O�<�wMO*Wp $`�5�(9tdCL�<YC�?X�@)�6�,��@�H�<��	E�/���%ȴYJ�H�+�J�<�rj?d� ��k;,L�ؐ�*�D�<مK�1pxy��'��' �0�uv�<��^�fްI �Mטr��8�-�o�<��$)�`%���Ԁ��	��S�<ЇH�Xz�ŀ�%����@K�<���$�P<8S�۹K�|���F�<Y�`i�Uʶ�\50(N����^K�<It�����hRgD�Oz�a��@�<yh�"2d���:����r�<�BN
!;`�q�E�W�e;��@d�<y�m��w�\��g� �q8�&h�i�<Y��@�(�����=��Bl�<)���/4H!I��	/�qӶ`X^�<��X7�@q�#)��y�d���e�V�<y�!1�|Q��p=��aw�<� ��0gW=L�zL�E xUyb"O6���(��Ua�ή=��� �"OJ-�O���m�"�H�`�`j�"O��%�WP�����n���ش"O�@Q�L�9M� 	T̚�"OD� �=>?(��!�f'V�"O~`"ҏ��T�Eiq��7ch�3�"OT�y3k�W�����oŚ"^J��Q"O�b��_"w� i{@$��4H�A"Op1PT�]P0l�ە%ũt32d��"O����CA	]�����Li7���"O<(Z'#۹�p��&U�`z�bU"O��`�`&���6rmL�cA"Ojp�WK�tZ�Qţ����5k�"Oba��b�K�T��\�K4'"O�I5�_HԠ�Õ�,��"Oz%
"�T �:p�?��s�"OV�s�$!*��y��rچ��3"O���򠅈8<��d��;J�jl�S"O�D�Eм2�]��Ŕ[�F�"O�#���&AŎ%҄C�:E�=�%"O�P��+��&^�<c�=��"O0�K�l��MIz��SE�.`b��i�"O��`Ĥ�D�)ЕdQ%20���"O|�adǅ>��(wC�b"�-U"O�IӅ�<@Qc�Cǜ-!���"O@�p'L
�*�AȞl�6d��"OnLh\rWz�	U'�1LNH�#2"O u��aD.(����88�!�1"Ouj�)�`��ɘS�@�$DAR�"O�����#[�M�A�#4�j�b@"O����)�#$/����@K�n6N���"Oz��6�?'�p��`�HCn�Y�"O�B"K�Nd�5)�?��E�"O��b��*'֔b�ʀ�����"ON�x�@R��VQ��NOO�h�"O�,����Q�`|���"< p�x�"O
�+4B�#sx���%�K�F,����"O���B�
}z5R�E|���3"O� ��	�[����Q^�mz��'"Od8Ggj���I0��4'XDCd"O�}2 �X(�p�_��>@`�"O@=St!�;k�,bZ�4�4}�d"O�E���<7=6��Ö$Tt�"O���2��k�H�RA�]�5VtX"O�����T��Tx����"O���bHE���Z��8�"O��`u,H�p!�B����*ڂre"Ox)ɒϑ*K��݃D�Yd�j�"O��"n֡_��2��U�=8,
"O�$8�
XGeD��fo�GN�,#7"O�����dޘ��D_�Q=-h"O<�#��%�*4Q��TE�1"O>�+֋�/4\F q�@=V	�"O*� G�E���[uSP$T��"O��Փ@���y��3zP^Փ�"O�pQp�íO����5`H,+5쬒�"O�sGΙ%�z"*���*O&!���0Ϝ��gR��tY�'`��IE��XF½�E��*8	�'�P�R�U�n{$h�Jq9�'��Q�� ��JYc"j!�Ba��'��aG�F�A:�쑱B�X$��'�� �r�\u6TbB- i�!��� �e3�*��jD�Y�un@�ޘYB�"O���J�Z�,���/h´�c�"O"��B@�,St08E݌B��0�"O�(���D* ď�H��"u"O,X�S���H|����N�b�4d�"Ox��U�&H����ǝ5g�$��"O�E�F�B�;��E�a�|S ��"O�ѱm�f2�Q�ae�?2�8�"O~=�M�!Ȝ̡ƤW�R��""O\����ת5Ә|qc�	G�|��"Op�
9���j@CW+*p8��v��yrcG�B��TS��@$8u
��yR���U��@b��8b.M��B<�y�-�0&�­jC��2����Ξ��y���2B�T���1'3�-1�a�3�y.K�6��B�㺡���D/�y�F_2z!^������t._��y�ǜE���b��y!$1�B��y���lW�$�dC��k�8��A^8�y��@�hӨ@�t�U�\�"Xi��[��yB�"L{@�A�G.X{02�&�0�yB��$-���{��ΟPr��A#��y��ɠ5R�����IJ��3���y�����
Ǝ�.t����S���y��T���hs�ךk,Z��۝�y�lB�"δ�I���.
+T��y��Z47X<����!��u㣄Å�yRIV�xo�d��ز.�#e���y2��l�,M�1&\�9���҄	�y&AG���Y-dJ4� �H_�y����� J7��.L(2��K8�y�JїoL�9PpkҀ�ʕ`cD��y���*��	��b�c/�y�t��D���	��fa��&��yrC�*�쑖&��e��@����y�b
n�x�Cɕ�c�r٠�g���y�@�+{_jub��qAh��V"��y�D�J6l]XGN�x�fΘ�y��K<,�lHE���&��uQ��y�"��iF�"��#Z�����c1�y�,�,��\E�]�i���1�昴�y�f�lhvi�6� s�t��7G$�y��-7x�Y���n�\���^��y£T$�X��0k��A�U	�#�y"��v�������=I�LI"�y�O�:��yT.�?'ND����y'O+CX���O 0�Q���y�iS#~2��0�.
����s��)�yr�I~��UW�;��g���y�dͩf8��˷���h ɇO���yrҔF =b�&&!�I���yR���mz�탛	�i����y�I�	m�}#��t4*4A����y�a�Oq�V�Yj��;��C��yR&�\�e�F�P�c�y�/�=~-�D�0*�rO(�5l]��yr�L�X\|!D��.�a�:�y�㑾p�=�䄳T��q�σ�y�-��Y� � �F8	ϒ��q����y&_8�l����V�2���y���0$t���7~%��U*���y�(] ��a��+S�v���q�o��y���0d�K�fI�lx�P8�˅��y�o� ���%�aV�"�՞�y
� 88*$�6A2~PT��A�0�i6"O�,5*�2�4�t`�TԤ���	P�O�6|'D� ob��G�8(2�DI�'�Ĉ��/܄D(�$U�!����3O� HGDX�F��]P+,C��"O��+S�PS�$ɉ�m(8 �s?O���D  V&xj��ϴP,p����{�\��A�*`X`,L.��)�0?<�����������^$rpY�5,�Dy��|����c���i��nȁBf�U~�<9u*��cd(U�FHnF���4�A_�<�٨0�Vݪ��=
����\�<Am ��tŒ4�06�iP���U�<9�*�k&��Dk�Gb�JF�P�<Y#�	ayt8��@�xU(j`��a�<�a��"8�yY��A��MiqLXW�<A�L���]��@Y�&���R�<YF��Xj��3�M�	�	�W 	Hy��'W8�z!b��Dڜ�CV)ʻDX�k���Y(������l�)h���R�´�ȓA��<�DĆ�8Ǝd��fʃ5�~��ȓ2v�;�
�*A��$���!����\o��h�##����L6=Mb���?�.QI�+[8�X���Ā�_����ȓ��#1'td0*���)x7�'��&��E{Zw�<�(�q��y"�įP;>I��'���l��qPr$_�3�ʔ3�cҳ�yB�\,��4�� _�+�*p(d˖�y���6�dA���� ɯ�yB/Œ`ײ��G�K�ZLK3��-�y����PJH��v�	��ĴX�AI�y�����̩����xa��R=�M+�On�ť�,w�N� �B�h�!Jf"O2���+�4��u�V�(�r��1"O�dG�~FD�p��}��`q�I�F��B�dE����/�|�B�A��y�	7/�<4!���y�l���	���'�ў�?�����X����� [p`(��Wz�8oZe��`��aA+C9��+�Kw~$�Sr%8�O�O�aq��#.p������d\죶"O0�� �'����|��S��	L�<!��W�m,�IYj�4n�;���K�<����?��{aeB�#wz��Ւ.ў"~�	j�>��!j%x�F�ZPCO�7�rB��o'8�!c"F�ae|���ˑ�0C�I
5И�g�0<6z���λ�h���"��.D)��K�	�`�"���_z|B�	-nYH`��V�V6Nʅ0����ȓB�FY(ed>2��)���_:�2����ޙI�e;G�@�c�˝65Z��%A����iP1�ҧ��.E�"8��Vt�*�}-\�aF��<#vȄ�p�����m��0	ԧ@��"L��fZ�A&�N�1�x)q -�5��������"j���p�������i1��V D�<]�Ť�?98�ɇ�@)ҵ�ǭ�:%��s� �?�h�ȓ\�d�R(��Y�Ļ����H2h�����д&C�O�2y����4P��ȓW
h �玈�PNǲ}n��ȓ?��ٰ��8/v�ai��X�#J蠆�	˼$�g�D�� ��d�*�5�ȓu���@�i�9�H���ǖ�t��6htt��   v��@��@����S�? �%� aT��,�1g�	9J�A;�޺�䓢��s���jQe[�Ҡ���2hK�0��8D��s!L��)�~H⇊E
HԘ�� 2��0<YG@X��2��ÒR0���b��f�<	&J��w�~	�u���A��KW}��'6R�{3�ʴ4��10VkR jd�!
�'q���V�¦	F剶"+?�(�	�'�4AE�x��!�����d�����I�����2X 8�43D��1� �D�U�!�d�>u�U�'��Jn�	@L�K�a|B�|J݇q.PZ3KK3tK�<�eS��yB�_$�z$�[�g2����*F���{?���%a��4Z�RG�_'h�N$���w̓R>6x3��@�]H�Bqh�VL�<QP�'����	tƠJ��^�J�
-��r�)���*�	�듃b�a�4����y�ᒁF�B%{�����r�ƍ?�p<����,��ٱ��%Y���船co!���.��R�iL�@M9���k�Y���?*�%Ϝ,���&aҭ
���� �/D���ōt�U�v�\UΉ�  !�	2�p=!G�ʝ�,%�C�C2N��,�w�E�<91I�%�dX�%.�,̊҂C�<�FIЮ�A�P�^�`�0������9�b 3��y�0��#F�z`��=�lJ%�A�a�D)�t��, ��҃O�j�)V��!# �ԩ^�ބ��'G�b�{w*F�q�E1����KFy R)���<�v`�-��#g�'�Z x��O�<��΢/J�qj��S�(�ęChF�<Q���O�(�z���yb*��`��jyxґx����s!0�)3�Ж)c��;wOW�Mma}R�>y�/ҬNTN���N�͓�C����'����)�ӽ,��x*�I�6����D�Rt��?1����%E��=I�@�. "��0ԥ�8I6�|�'2�h���.,�Y�����YI��r�n"<��a� �*�EY��t�Hy���F�<���ж-�0{7-߂N�<!Ҋ�@̓��=ٴ��&�IP!4(Z޼H��S�<����J��d�a��{�.L���z�<�����-.$ 0��.9&������P�' a�$�Ag���������R��%�Py�
�q$�x�!6kO�Td	F�<AE ������fc15e�8:�B�<.Z�1t�fJ�0X�q@ SA�'���$ql d���)ORZ ���HC䉢G�����
�I5&�c�Ώ>
)j۴�O?��~&Ľ  �*' �蓡��g!���zT���zX���c!�$�*|�NU��-��n4Y�ӏ�N�ў���	 #
�a�R)��K�����<-�8B�	�B���!"غpR�5����DTB��7@�Q@aMޤ	�������G*B��[Qr4���ݷE5fY��U6C�1L<~@`�JZ�v@�bg S�B�4 �z=��N�p�oQ�N]�B��5Ш�R� [u�\r�DE� ԴB�I�4�Q��5p;F�[�C�q28C�I�T����/ъ9��u�Sc�G5C�I�'��|�G�V/�Z좦��4�B�	4zȎ|��h�O0��A#�5g�B�	�ќ@����5
� T��7[1�B�'a� 0w��Y�N��t�Έ<��C�:d��BV��=�"]	��R�t�B�)� ҹ����U�_�0��x�Q"O"��sFQ�gFZ��7��7=TR��"O m��&X4�L`�OÙ)Ln�V"O6�#�fų(��a�bn�(���!"O����J�6�����$=��Uz�"O�%[f��1s�����t~����"OT��6�T
"�� A3v��"OL��BɌ�M��\S'�(�(�"O9k��,P��kc̨m��|��"O �R$��lx2��#��2.W�$��"O(��.Y���G�J8W���"O	�V�	�\����ʋ�m�3"Oz<;2ϓS���"�"ƺ�Ja"Oz���/�./1�ݚT�X�B�p"O^��E�j���(��V5j�8�{7"OR�0Ԍ
u�,�y�a��Ln��p�"OZ�ВcǍ<�Ȼe`@ 6�\�"O�ђ�+�[cd5PO��JNA��"O��4'�.lPZ�&Mɴz�tE�"O���S*]-��!O�]�J���"Op���b��N��0XvmX
6��C�"ODB� �|9z���a��/����"O!�avH.q����Eu\|2"OĠ���7z�\�tJ���.��G"O�e� ��seZ��F��zpXݹ�"O\� �l�5�~UҮ� -f��R�"O�8��\�%;���"�q-�9�b"O\�ۆ�G���H�A	�t"D`�"OȬB	��T��
�˅y6�I�"O�����.ET���g�h�p��"O0l�&-@rI���tg��H�h�CB"OHY���� X�`Q\%8��Mb�"O��%�[?�K�'( �c"O��R���n�nmi���%$Z��"O�pBфR2""���Γx0��q"O��`�[�8��@�*q�Ժ�"O|�*G!Q>P�3_�D��""O��J�͞�P�ruH��@9	�ڽh�"OH��#�?#ɄUG�/m�"u"O����0F��;Fӆ��A��"O6��Î�T��eX.T+~��!"O�mb6Gվv
�reʀ?3�H)�"O����%Bf��H����!:�"O^ݩT���Y[�ѹt��?|�l�e"O\D��޹����"�6�Z��t"O�p�!_��P9�&�.�
�t"O��ӧ�H�)��iI��v�6 �"O�$#pbߩ8AС�&CE�Y��a�"OR��P �)���9�Ι�g"O�����H�hS�B:Y���ؑ"O@��a�M�bFX��R��D��}@w"O��(�3�&�
WkP&*��:"Ob]��(H��Hi���/���ؑ"O��Zd�7�4�a�"W�s��"O���i��+������zj�-3w"O�1�`F��]��h&�E���[G"O�%�`�^�=���	A�ٿs�*�Yq"O��y1D��!>=���:����"O.�Y'��m�J�B�>s����"OT�����CiH�#DB�KS�1!u"ObY�CB�0�f���Ό�K��kR"O4X�G%��8Ȟ�����B%t�#c"O�-����Uu�!��+Rc�6��"O"�!R	���B�\�4���W"O� �@�`H_�l5�D)q��#%"O��{0Ø�v��uJ��'Ig³"O\<�0P������M�H!K�"Op�Q�-$ n]Ҧ��*74����"OVݻ@�E
��J��`����,D�)4��
�d�����-�E�$'D�X�T��xt��`���I`V$D������LL��C2_Ģ�BW�/O�=I�MM/E�)�@<
��1C'(�\�<Ap�I�zh����>B�N�Q(Xc�<)�!��S��|Q�Hι/�ly�r�`�<9t�ɫ��#��DJ����f�'H�y"�\�<%��mR�gF�iy�)�y��)X��Z$+\�\��J�ο�yb�����ԆS,"�|����y�ÎM4�@��g�.t��#���?�'lB��UHC$[�(���B�6&�(�'�96*��E:�9A!��&͆!
	�'���Gl�]2p	"��l��'P�(q�NK>�`�`�H$��u1��$&O�ɠ$ܰ8�.����ίHx����"OҐa�%T�@9��mM�/Y����"O��a��R5t���BP9b�+"O|�G�1 0��<���W"O�2��K��>Qi"A+�d�f"O��Q��P�9�8Y5o!�
H۵"OtI��Bi�I��$F�%w80�'��DF�&8�p�aY$����Q�W�ab!�0B �d��@�G�ZИVʆI!�L'?�\��B ؟t8�@�+!G!��u�`�4��LAJH�@	O�u(!�S(f|�䒲���h�ٓB�.!!�D�A4L{F�O�b��m�V�
k
!�d;�F@�Ge�ep�`�働.T�򤐲'T0mq�C薂�`�(�?y	�'0���c�;!3�4�1���-3�'/�p�3N�|aN̲GaT)\	"���'-Tu�ra��e���h$�A�X@>U�L<i���)�)hfh���O�zjYZ�H��0�!�$��1�Q�6" �]d�Ъ�ҬY��	P��CWOG.r��� ��v��Y��<D���G�Ա!J�	+Go= ��x�Ѭ.D��hf��0JXN��#�J����XB�,D����V�G��i2��2a�L�0dI D�,��]7K��5��cR>vH�!@>ʓ�hO�#R;&��r*��a(��0�?j��C�I�6�9�� �9 4Xvo��?�lC䉾VI� 楛6?̼8�!�\}$C�	���ubcnڽ/ɪ�A����D��:(qa�<l %��,KM!��J)�%��(B�;������~2!��O�a��	"|��d�Ug���yw/N�������dx�'��w���n�yb�9&W^��Q�s�%(�Q��Oh��$�;0���k� ⮙�#�Z�%�!�$�t܌�L�-}����̕J!�DB=H�Tj�\"Zg}�̎*.��'��|�\c���b��-�,$b�#Ʃ�y�D�0 �H��A�{��U[�.����OR�zЏ�F�������Zqi�Y�<i� e��R�)^�tV�Ű%T~�<��C�Ѫ�����S�FX��b)qƱOУ=%>=��Ě74	I �9l���X'�5D��(�������[@ Q0s���! 6D�� A0�"Չ`�$;T�̶h����"O����Ӫa��9�"�(%�y�C"OlM"�*��\�PY�A �
E�r8�"O`��� J�
$�m�ύh��F"O�����ʿrF���M�Qh�D���'���OxB��
Qa��e��.�d�e"O��*��W�}>�C@-�0z���R�xR5O�b���}�IǬT}���_HH��F � �d�ȓqB((p�q��0	��Uc�'�ax��]�$h&i��2;��8£R
��Op���O��Q�%����a����2h3���'j�!���Udd��ׄ5��A��'��Ja�?~It@��+�:.)|:�'��ja��:GA`��&��)��I�'����č�.>*��Q�
����'UJqf�s�p*�Zn�8��'Y�]�����d�z�M-fʎ4��';���{�0 $���0���0
�'D�G�Ҷ1h�@Hc�{L���'��.��h�z({��S�a7 D��yr��<V:`(җ6L�)7�ְ>�H�l�G�U;�(�6�� h�����3T���`Û�%�|蠤�N<R�rQ�u"O�Y�Q�S.`�p�¡�lA��"O�}	�"�&7#NX����5��]��"OZ�&,�i�����Fc�*y��"O�p�Ձ�?3y쁡���Q�AH�"O�Ab����}{�N�0+���'e�]PD�=9_���Y�~��'�x1����E��U@�D�T��	�'Ϊ���D��1< ���	� ��	�'�� �s���Mڊ]��f���5p	�'a
b/F�5P��c%!{���z�'M���EQ!Fn��䁎;3��+�'W�  ��Z��hYG�Ͻ0H�3�' X�3ר��t$H��Ed��(@��i	�'�� ���0N�f�M�x I>�����
(cur�р�
]<U�
]��y�	f}�0&�?.]��� -*L�C�4
�|QZ�ˣ|��D�r�@w�B�I�D!4�IQ�QRg�@]%(<��'Ad�B��g!�5�f�8"�zE��'�F�9���`U������B��(��'#n��#j�"dO��ID,����'#�kGe�,b��D�ƹ.�I
�b��	���pZ���Vʎ$�pxŃ�P!��"\�1�g����0!�$�%E!�^f\}�Ր�<�:bK�k�!�D�0W��h$&!{F�UfQ�ak�O��ė-��	��ڕxYb��Ş;U�~�O A��F�+�i���E��d���M}h<Q �_�~���O�B��pUNL���'�񟚨ȒhL8!&�A�CXRd��yr��!LO��Go�}V.����H�v��6`�(O?�� D�p����7QD�+*N>C�ɢkH�t�CH(Q���pG�ڙb\�dB:1r"?ю{�U?9�(�uHD=�c�ˏ��=�����Ԉ5I� H"�"(4L#q�N�!�d��h�hM"WI
�H�S�|�!��! L�KfƊ���c�B�!��0Cr�% ʻ/�^Y�W1q!��R�rE�
0s{LA��i>c�!�$��6����,p���'P�!�ߪ%jL��g`��4^��1ׅ�)�!�� �|P��I?x�t���)��E�"OV�adF��ti"�+\����"O�ER$�<t�SS�Eeݎ��"O8�Ҋ�(��Ѡ��X:4`�p�c"OP|:2,�(>.�QZ⭝'i7>0��"Op@�5J�7���^�I�찚�"O0e#���\N`C��7��{�"ODL9�m&C�x�y��7lU��:�"O<���+Ɗβ�+�(ސ5u��Q "O��)�����5��J <l^!sr"O���b�[�D�e����(R�Y�"OTq�v�G�b��e�V�PKH&�A�"OF���(X�6���DU�Y��"O��(î�FD��S�튕6�� �t"Op�j�ȅ�K-T�I�� R�&�9"O����-�/ �8�)��sr�� �"O�ذs H�3a�e�ɇ�c>�L(�"O��b�π$M!*� ;U�@D%"O��KA���`��43�O�"��q�"O�la ��|g��8���:�bx{"O���F	�3v�NL�dƱ,�<� "O��F�ۛ)EF`�C��
�X́ "OP1B�.<�
4`e���)�"O\t���
�xp�N����"O���W� ҈�q#�o�Lb�"O�8��Hp����P�F�$)��"O���� qh��+��6�ձ�"O���#M�#R���3/B�X��@��"O�Q���='������ �ĉ3w"Od��ߒ;��D�C7*��(`"O�,�m�6/F2x���Y�5�#"Ol�$@���)Q�+¨v�\"p"O�h"6l��l6,��,��`B�q�"O�I�d�<�� qf�y,�T��"O&��ԖJ�☋d��.�I��"O�@(u�>z@���(�)PXu"O:@虧
��@B(�0i+>8��HR"��EҠ J�#�,���4�l!��
Je� x@`Ѓe�!�d@"Rb��F�Ԝ5�4|9w���!�?^�bFT�r��=顆�'9�!�d	9�@� Ɓ��\Fp�롤A+e�!�d%��rG�> vT�Э˦m�!�Y3����p��?'�9��CK)�!�r���S��E��=+e�(�!�DB�B\��,M@��ŉ--��4��'�>�(�$�1v�޼�`"�7m�д��'�����2_�n4��f?�~���'Ki���f4DׄѴ�q
�'�z�A&�;����A��Uk.}�'�0�j�`�Y��=���#Lmڰ@�'��8���ʺ.m�4o�6�0;	�'L@�.i�F,��
~9(���'՘�X���4HP��	�ho�)�
�'��H��t�	"!gQ�fٮH��'-5k�	nPF � �H�XZ�S�'�d(*��5�,����H� @)
�'� (�WhK%u����ˍ�T ���']f��Q���^����s�'0d���'��X*q@�q4��p�-��4F9��',>][ʆ(mF؄��'�'� �'��y�7��8{��Uy!�ˀ�4�+�'����-,�0�Ǥ��r��S
�'��VK���8�FN
�s
p�;�'����A�Fx��ޚc=�CIY�^ĵ �K$�O� $��W�CH�m#*�]X!��_�1���)!Hp�On�5�[�_����OǯJ�,�#�'�8(��C��t�}��@�9:Y��O�St(������e>ͣq P�&h�v�ߌ\��Dr�#0D� �VC�S��"�]6pNI�F�#n1�����}�q�hZ���'��ˆ�Y%!o���#�Oߪ�I	�o�̼�7�4C`��qS�ڌt�̢��BZ+v�z�f�3��P��'R��n��A��P;��*�(�э��*^D�%냈�o�*4�"��%���� Q�~�V�=L8x�����y��?�:���ǧ\9��ҥe�y�+S�KufL�E��.[Q�0��\������;x���A���*�rpJ�"O<uU��46qX�q#�=Kx8�U��%T]$Y{#�E4U\�ۄ`F _���K��l�z�AU�ͤ0�N�:�MK�
�6���ɅA�@k+�<Y��`��+�V�@�^�����cE�
PjJ�����.��=9��"Av�U�EAU)J�tp0�Ï�'%*�b��O2M�6�R�)Z�
�|��7BR�E]n,�u��p��ETE���'/Z9���أI2Bqf�����#�']�%�4AҢhx�ӱI	�v&H�E#�����5�D
Rn�R�P�GṆ"OJ�e��!� �o�;z�)�vG#X=><I��@0,���QG^�lx�S b[�c��c��R��HC!ڣ���a��-�O� ���(��ˇ���<ڵL2=��pc�:{7��N� X�:83��'W�Q�I�R�v��FE޽x�b����:iU2Ea���Tڶ����>S%����&(jd� �J.K7h�hv�G!��[��F� E��&y�"(��n�	>��]�AM�P��D�W��/⬬�c/�H� e9� ,��.	?��nC�@�H�"������'�;F��"��D���̓��YrgQ+t������*���$w�
�!ʊNe���L����UR�� �_"�YT��6-b@�K�/]9	���
�hM�yj�q!c�3���x  ��&���vH�g1��4jÐx]h%p���*m�
,��Y?E�:�ӓf\A1��2'��U����45�"a��`D�!�O�-$㪵�g�C1���H��u�����[z�"� �Jڙu���J��� �(%RtB�*��7m��\k�R�'༜��b*��J��V`T��Y��ʻ*���1��+qt`0&�[�f聆���+��b�g�f^ˌ�gf��5��k�O��M$H�Nm����h�>6�Zh��K�.����K�Y"���bT�Dt���Z���%`��&R=�։N�>ݐ�a
\<��0��Cj�
�gB�jI!i��ʆL��p���2�[��P��ȣ"��i�P	��J��xꥌ}:�a��t9q@��q��U�P�B�|Aa�+֑¦d	�
ݴr$�{�'є��'z@|���ڥ4f���O�'��ta�'*�EB��/������3qVP�7&;x��'e������+y䠵�&h6/I���� U=v�HMSD�ۖ&�r���N
Mrn�v��;zi��x(\����GW2nzT���	���$�Xª��N�%9P� '!�;(k,��8�$�xP�ш2h��jАSa~�H	*x��%��=�"���\aN�P���(0^����)�ά���Ռ7;�L�R��z6�Z.�+[nP�(�/?@���&�o�$�Z�RR(̈�����O�R��&%6�mä��� L��$�# �
l�t,�7�P���SdͫV��J��9��Ԛ+H�%�a�־oNPɄ��0�F��>��͊BM6���6U�y�����<)���p�� �۔
��]�3m˛D@,�xQ��	1Z�M� �_>ڪ�-6h-�^�$B�쀨kI:��5�Ekb�cРp����Ff��#��D��S�*)��N�Cm����e�B��S铀Y��;���>Q�U�O�V�>����>Ddkl�%��k����k6O��W�a�
ݧI(�Y������=I� }q�\J�l'���!K�a����I�D�Xa�@	�,��F Z�yx�x�T���!��劀 ���s�[; �(yBq?��*�b��m������:d��d��RݸdÂ��.�vqJi��)J��;��ʴ(`���b.�'5��$�2$Z?WЦX�2&?���t�xei�~��ȓ�D<0T���1���~l���N��� UAA�����a��87XHZ����h��a+��5@�ף~<dA٠쏴
x�rH�S��<ّk	�=��ԋ��]d) dԒ�� �(H�zܜ�AeדIT��	�<��ث�͙�[lP�����[���	)����7%�(3�TH$�2D�����Q<C��y@ȑ�Zޔ��U��o���c������-	<Z6�����=A��i�4��5���'1�1�P�עJyrE
COے�8Ŧ�e���r�4�rW L�F ���T
\o�Z����HL �􏅑-0Z����!�M�3�B�E���8��.$o�p�ᑤz渴��ύ�Q��x�CD����"F�1YRY��k��N)����EELK���8t�݁�K�IYD�'�`�)�kD� �1�OL+0Ɇ�0�O�=Rv�^Po�1K���.1"r������DS�0���é$���e��C}!�$�%
daR'��2(M0��%�i3\(R���q�@<��DӰmX����ӟ2�g�ٔ=x��	6U���H�)�U� ��	:���C7fX܂uL�<C
Le*�� C2�C���^Ț�KT`�$6��
דQF�ig8�V�{���)��Exa�>y'�ˊ<�N��$դ"��)%�^Z�? :��3����a��+��X�'"O��W��.�ؽ�� ��7,8���{}Ҏ�X���ѡ��%��Փ�	BW�'�y'ʖ4qVV쳂�K6�H��-�yrNp[ެy$��)!��P�R�G���0@��D���l�.�n`���pY��g�>`j�I������Uڐ1�e��	�QV�[f,7�y� )�ZKh�Y�F$�B��!�xp�ۓ��4X�����8��S�ԎѸd�?�a�:?9�h�+M$��c 5,���|��BB��iɴ��W��Vv!�D#!�XQ6d� �r���2{�!�O��s�a��{D2�S޼����J]A1�S.B�P`����p�<��kߩNf,�0n�m�D�9���/j���4�"}b*���*�I,�Dk�/� 2�l��ŉ�z�����7|O,}�O<)7k�'8������@��)oIO�<���\�(���4��%,1�U��K��+�^�<���r��	"�!�L�D���C"O�D�S
��>�X�@RG% D�h� ME�'�>��>PU�1��/Q������^�0��C��#8��p�Wc����l֖G�`�D���?����~Z��c/ʑDb�5c d��Y�x���DYԄ��$Լ�:� bS�y2hR�\�8,����N]p1O�)��'/��GyJ?AR'M�(�ن�qfa�@,D� ��9m���ʕ$�(�"�A� �(O��}���<�eM� ^C�����&QF`�ȓS�Y��*��$d6 �������]�a�Ȁ5�`yr�Բz�82�B��0>��x�oI&=O��lˮn����dΛ�y�X�Ny����fP2qW������(O��=�O��=�"I� :��q �W�?ɂT��' ��pc�>���r���31�D{�'�P���i@��d���bZ	!�|2
�'8U�'F��(uT�z6������)O�܅�	*MR�{@m΢C��8�b�(U ��d�+�Ğ�(�"�
A-�$K9j!���"p!�W�|���j7���R)��AB+�;n�Q���w�-w ��2���]�S��$ ��h�5iT�i 4AC�C�ɑ�h�E��e��I�D�0]�ʓ{��Ŋp�ҧ(�|�����D7~�i0��Lۈ���"Ol����K0C֪����y�v :�"ON0j��@�m;��Ü<�P��"O�L`���r��vM��,�b��V�i�8(r� � ۪��O?7M��(d,  F���2���&�"}�!���%�6�T�V(�c��q�W�O��1 'J�@�L�5�|8���%eE�
��0 ��(Ey(%�g�6�O@%��=`����҂Y	s,~��#h��6��Kq�_w���(�OXr'צzP��hкM�ȀP����,�:@�/N�42�Q`�ӏbN��$ˠ/���@AC.4��B䉘o%(pD�%2>�y�*)!�R��&�C�D=ujs#��*�M5�g}b���}9����9�J�Ȉ��y�*�_ݤ�Ig)���X�
�pH腭Z�q�좑�0~��X��O�y��3?���Ƣ�C_2� ��'�P̡�J����a"�B\��d�֬U�l"�q@�<G��9��oK'�?��N�^�Z�K�� ��t���Y˦�1��P�{K��K�{���U�O[�L�R��OC�#6'�: +*�Ka<a��I�D�rw��˃ Ǆ�(�`/�]��i
�iz� @����ͪA�'��x���>�5 Ý;[:���jUK1��S�p�J4����
2[6�~���9n�nT9����l��3WjX�im<�Ӗ͇UwDԳA��v����{�'
�=y��*?���+�+Zd:R`&��O��Ĕ��+�-+C�$(�iH�w@DT���Fln� r�]�
$XRц�'`���R7^��䒍w#��9'��v7l	
��;UA8� G��O8�Q�W�V=R�;�$R�w-����d�]yN�󃆃^o���z���6"�"3G� ��	�iO<q��ę%mS��c��*Q�d�v��:A�u��E>˔d�E,�g}��Ջxp.�*D䝇nN�1������'M��a!�9�R�D��J�.����&J,a4��XQ*��3�VD��(��k���Z���l[��O� ����!Rǩh��k�`��'�؛_,ѠN��!�8���+�(����u�K\�U� ɓ���L��� &���B�'*hAZ� X$	
.�H2d\�#�P�ɧ�֤7�I����>9�b?�*�i@�`,�|R��8�R��!F�W�����@�y�<�	�1<\p-+V�[D7�`�7�(@�fヅ׳`���XD��>E����
���#�-���`�lZ�J�Z���e{��D�J�y��A��>b��}�'WHŻ�`�E�[˓]Z!��G�|0D%?nX�ȓ&J��i�:O�ޙ��� �����pD�PeSS�$DV��un.}��F��9�Տ �:�ꔫ��;�n���
�����B=)=�m�I�XoR���*���(3�����Q�. �ȓ2,8��A	4��U��A�:-��݅ȓvZ��%G�9�p;�'�6�Z��!�r�2���	�T���7� ����a&e��#Y$�Xb+��#]��ȓ�Y�gV9c�{��-A��a��v����"fP����lN�;��ه���@e��=
�%����M�4i�ȓ:�4y�)X�lᮥ*gH\>D��ȓ�D���G0�tr1ƒ\���{�ܭ�KF1��05E�3����`��b�S�^�� ��ʆB*Z��ȓ��� 2�:�� w��k�.܆�iڲu��g
�Ix�+�#��?W�8�ȓ)T�%�b퐮*<�h�b� �6�x�ȓI��lؓ)�Zɪ�,ʐ|���b�<�t%�` 8�%��0�'��IC�*ņX�n�Y���4��e��'��8"VN]�+��T*�%�3���Z�'�ޙ`�녽l���ha��:_L��'[��r��W�=C�1u���b�'G�;�'�h�Jdht��i�P��'�2��0���8/xM�c)�k@� 	�'���ȇ�H3��ip�1�����'3�arJ��l ��pG��={����' l!���͌u�����V�4H�Q�'��M��f��c_Ԕx���.d���
�'	���G�Ի� �:b&[.k���
�'�6<�bc�&T`�\ö�l�-��'a,1�Ps�8��֏f*d]y�'���q#�\�R���whU"U�� �'. �QA�m=h��.C�ε��'�4�"J�M�}�e Y�?�ʤ#�'E��BHF�n��<2����d�BL2�'�P�ك�;�hܱT V�wC�]�	�'�I��(6��p{�D�
:��p`	�'21���I�St���ˊ(DV���'�Z``�e��੩��� YP=�'��4L�1�.hu��A@��R�'�j�1�C�90�d8Ƌ��<8�'�f��o�7�*�����}��'-kd��7�6��W,��ft���'m�@Ⱞ�
E��Ж�N0gF*Q
�'�B;����p&������RϺ���'���*ݿy��H����X��
�'��{��D5/t�Ye)ݞj3�'hк7���F�
�"��^�Z=<A�')��b#_��:�&lQ@��'�� RƋ����֣�7UR���'P��	��V�R���,j����ש�[�<�`�z��L�a��)������K�<Q�F*R+XH�BjV�@H����F�<� $!���Q:I�]��)�҉�"O^�:d'ةt����a�<ȸ�"O���4U����n�2(��1��O���Nc9� icN,�%`3�+$� �(��LR؟0{��E69 2D��	�2���7��"���0H "̧�N���/�0����I.1�����"OԠAG$�;�D����s�X-"�P�(�f
��`􀣕�љ�0|:���?XFl�c���t���VG�~�<��oM�1��S��.���IV@O3k���'W��bg�(���O����NS�O��� ���7�r�)2�'8�� ��s����ϊ>�^��W��%m�]B��Ow��ȃ�5�O�${�@���Tu�6��G�h��	�m	�#�U(��ݓ���l���@�'�����O8̆�(@���b&!��	�j1��l��(K.ɼg�����,�fK�12��;�����?�k�c
"8D\x
5�۶}����>D����(��C(�%�áĦc��l��̞;j�%��_=DHbfm�o����'�ly�,ܓo��䚐�XU�b�G]��`�CN�^Ӟ��T���!~�:��\6|����,P�Iʰx��V�p��i�ۓ
�����#4���[���E|ra @��@u=Y��93�8��7V(Q%�[��|�i���ye�e�*MȀ! �H8�v��-�yB)R��%z�jE nx����Ef�"A���I��r��"�	�$>7�)��B�0�!��W�XR,��Yi����v�d9��及 �xL2�� ��g�?�T�+���l��E��|�"2��R��D��G��l��@�����O՗%�|�pɋ�}=���N�=�NM���\�ӓ5�l�y`#�w{���E
0�x�D|�F,5zt:2��eӠ�9��l@�z�a^�p��%p�H�$X;p�`BM��y���9r��@O��	� �9x��eR�C������ �:��J�$>~��O� HR9�y��X��I ��Q 0� ��?�'��Z��Q20���bYȤ�Rq�(�gj٧�8lA���N�:�I7i���Ap)��dI��y�@��D���UTMn������O�z��d�>�Zc�4ޔ���"*������K�
Қ@jSE�G Ȍ�2�-h�����H&5�X܄��55��]��� �T�P�8L��I')#$�WE!A�%X2m��n��T��"�~]4AP��݀#ܠ���\�UȎUB�h�^��Ђ���Z�!�$Hd�N�Cb
�(Myz�h�GD���� �-�8'�਒$熏eyH\�q�	�a�@�cB*O(Ot� fg6�~�^k�A�� ��d����0?�򣛭4B��#JQ�]����_1aq@���g�?�5�ɞ/A�[��Jr�,��*� X���*��p�p�����ףv�{��nۦ�G|"N�35Dɮ=O�	�2�F5iZܥ+@LŪ$��!"F�{�<����0p𐒰�]=-|���	;\����U6<��-Q9V!2�i3�fd�$�9� ���R1|�8��� ^ �͐�����*G1��;BStr� "T�@%<4t��)D�XHt��\��٣���<E��Y��JB*壵�X�~0:�s4]��`4d�����/�sK�w��(0���*�Q'I��b(�+�ꀉy�$�L��7��8�����'k�T�pȐq��)/��dB�]J��i��M��&��<��'�Dy6�Cǌ_ I����R�'��P:h�s��sԉ!%V��8򫎧'c�i�u��2s&��B������&_�\�.@�S�,�*t�	ӓZu\���ã*�F�S��6���ϓ^�6$�2I�95�DY{A�8\xFъuI� ,�\�c�+���Щ���\r�s���->�s�"�q�vP�ȓ�`���� �H �H�P��4r�a��jhElҔbM7�h�ysG��n��֤`݉ cm��h��)71� Ҳ� 6C������Ϣ=`�� ��'�Piĥ_�K�MH�ʞ2>س�L� \��OQ�D�ء��¿R�P�Ъ��O�i t!���'cN�!q��+Wn�@��*q X��	rGV�B�h���;" "�͈;s�!h!�/*yNp`u��L���� 0���T�a{bI�C��h:V$�R���+�"�����2����7��a� 1pȗN���p󪞸zHF@vLºK��5vt���8!B�ȣ-w�<yҠM�'W:}�u�S4M�x� %E�%	҄[2%�\#2]�4�\D�"B@͸%U�=���w������?-촢�hԛYQv���'0�*wa�`(�cH�#\YJ��4��+u�݁a��0��)��UJ2�:W!b,c�	�ă�dI�EY�r���'	3� )�$�:�J	���08&���gڧkp~��7
U7a� �♽^x�z�M�BmhUQ�L�h̠�[�d���0<ykJ�`y�y�埱"�����,L����M
�*�J�∫"��@�ȓW"��pQ��~�:4�A>+�v=�';� 
� {Y��4*E("�E�T(�-L��#�Pa�S�N����� �a
��:E��'�L�h,jD��%7� �d���|����� @�1�1O�Ń�k�}L��I��r���(�O�ճ�k;��0���T4k������܀l���؃�k�Vi��ߞ�p=I��ÉY��A"6�çbҼ�A"%�`�Ě��R3$!�6E�,�����j���+'��qi���GFǠ/WC�7Dl���f�e����&��` ��+�ds'-�o�Vd�&��"^ޢ|��-2����G���K�м�D�u�<)s�m;���d�����F?6�<��6�
+N�ق�.�g���|�<YЀ�&F؂�q��Ki�Ĺq�(<yp��z��9S@N��Tv�x��HٻC��)���]����q�H���=��h�Q��"�.	�J���a��|X��y���h�	c x���#P��ɕlܟX>X��#O��y"(�6u}.���M\!}�=�#�����|�-�c.���TeC���ɥ2CH0�]!zx�)a0$�" !�D�*2Dś�L�! z����Z�5lI�<��5Hi�"|�'@~t�g���h�xX*��4ba�x�'���4%�ǰ�5C�g�P�I�'�������mh�Z��U�Rj>aB�'!�6��;������L�i�'��*榆�0�(}�ӄ��2|P��'(�P@��'�l8T@���l1
�'��P!7�r��؊ E�"	S& �	�'`­#����=|�Y0�
�Zl`
�'���Z��;"�6�GHێH�B�
�'�:0p*�j�#��Q��j	�',�ڄ���m�hԘ#��MG����'Wr1B��r!�U@�&DF���
�'ҘX��K:o��<���,FC�i
�'�$}'�&P٦ux�i��2���'<Z�G̕�W��Ő �/\D\��'�Z4s���g�}#�LP*����'�>�؃aU�T����ЊP�2�z�'�ᴉ!v�0[�ۥ�r=��'���� nB6������]�p�����'�(���
0=/� �4� ,m!���'ʪ���O��r$rd+Cd4Zz	�'�T���98i�S�X7��q�'��D�R��~^��㇝�S���B�'���l�O�T��Ѥ�II`\!	�'��	�d�*!d�j��U�74z�:�']�e����c�踒Ä>*o,0�'ovE:P��.�~Q  Z2/���y�'D��)��P4D��P$�ԝ)�D��
�'Hp,3+E\��@��ǘ-�2��
�'ژ�i��ʒ��%K�	�P�TMf��0SA%�/��l����"~n��D'�|p��%jT��p���R
vB�	*&�US���O�|<�SMJ2(��	�$5vh��cٞhV�M��S�YK�d�[�>u�����Ȇ�I,yr�8W��à��W���ot�9�
�*�,����}�C�	�;�者"S�����b��$ �ɽǐX��^x��	��'Lh����$�'H�R��˓;Z��ȓ9�6�j�ϔ� ����m7pE �ӊ�(r�^͠�b
�(�ZaG$�A����@!�> "Q�ͬfL i�[�M�!��� n��C�&�q�l�7��I�J�	Ҧzq1��A:d
 ��`aE��u��$�7A��7��=���+G��7�a{�G��{��a����i���Q��� a܀�ք�-ֆ<�ѵ!0ĭ0�'v&�� �_�t��t+%�����ٴ[l��.����L_�{8Ẑk��s��hGe2�)�2�n0{ҥ@?h�����H5J"�z��; ��hr]�|�E Ĕ�{3��4R�^l�BKB�S�J0Z���90��dk+ŗ/�,"}�'"�drq��'TP+�
Ū�Y3�y����ucWB�f�O��@Q�3Kb��!J� 嶅1A�Z�#
!ac���
�i�N��u���@�f���EN#F��}0��6?���ߟ���
nh�����8�*�H NX1I��h�J�%g�A�w.�#��uJDޏt�aR��>0��:��H�g�f��c�׽C��4��Y.4��4�ɨ;�r�c�H�?6��"�j��d�b�� 8$����!yѢ}0���4��}���'�04�Ea�g�0��F@!���65e��R�b���	�0Z&�EA��ts$q1V��X���G��z٫ਜ਼b�8�u�P1O> �ũ�[d�Q��)1�L4c̦p� !����*N'��S�HB;�HB�)QL�:��4��p�eY�i(�
T�U'�e����EY�	A��>�dF�+O �=��O��.� uXy��h�Kw��9a'�$<(`�5�O�����؍f�b���I�$B~�R�Ϗ�
K��p�Nj}�K��x@Mhl2u�XuP���J�u.ԃ J_5D����1���Pyr�b�n����ߙoa��D�:�fE fo�j����&��>E��Wf,�G��>6qnY��>	�:	�ȓr��ౠ'F���,i�BC8*1y�'0x<0'�3�U�	�7Ŗ�w�ҘzZĄ��@�8�蕄�UQ`u2 B)�M���;"�܄ȓd�|�I�X�&��UW���'X�"���$\H&0ڀmA�q�r�
�'��E2�g�#d`���h�%�4���'��a�#�<}f��B�@B
�'�xS�i�+��P��-ڸ
�6�H
�'���H�/�����'�=�T�+	�'�~t��㑿*��S.�. t(}��'�l�d���`K\*cLͮ캈��'H^pċ	<B1�d��HYEd� �'���1(&Vo�9�g��+y����'���3$��	 �r�It�?q�fy��'���re�H\�3.��y��!�'MP�[f��&g���r���$#�Aq�'�����'D��@XGG>L����
�'-b �$EW�bb8�����;t�L���'j$����}g���'BX��qk�'q~�;p�B,=�*� �^�z���'d�P!��}
�98p�;I <�q�'O�X@K w��8�F��E�ȡ��'�T�{5O�N`�u+B&�2	�'d<�A(ߨP�`�@�VhA
�'8x��o�1+��'A/���'�j�a-	��踻"钩
�Rɚ�'��U#í��=��������p��'B����Տ q&�9fǘ�&Ji��'ne��%J�U�`ҥ�קvV(���'�"8�GnG���Re�خ3g��'xq�R��eT���+)EL�8
�'����-�)��#��_%4���0
�'`
�h@g90<p��� �$>�U�	�'��b 	�1�"a�p,��]�lܨ�'��!�	8%���!�ͻJخ�aP�"m��+�I�axbELJ\����X�G�ʥ��ۋE&xK�e�<��pT�*�Ms�Ȁ�oH��q��?�~:��JG熕�k�ZFv����E���ytN);��<�uD�.�\0��S�*0l��VcƸ +$d�Ŭ;(Z6-�{�h�@�l��q*p'K�OT�.\]�.I����Z a�Ȟ&#������40������E�&��}i"���'��HЪFC��(��$�5-��J�� �h08�kȲyLɧ��$��s` l��-Ϊ����n�=?�p	�,�����$	�|�:"O]�-96�Zp ��7��/��+5����4�� �b
�z|2hU)�}���&�`��'���~B۴{6�9ɴc\?e�$��%�G+0����'�bI�k�VapW-�i�'R�
x�։@�G�L�ې	UJ�`�͓j�
6�թp0���O?aq₇T9��[q�/G�z�ғM�'!�#J<��S>��f�Ũ$M�a�>2��B��o�X�"Q�x��V>��'	�F��C��[x� �C��z�'���	&��j�'��sӸ��u��?j=2�S� ��i^���И>�dA�ҾL�<��pk�)$w 0f$�gy�=q���^?����#*8�<E���L�9��]����8�G�J���q�#k1O��iݭq�} +Dby+G#��}�:`;+�7"ȱR�7�䓙H����.=*� I��֭	]��C�57P�ҳ�)�$�4jl�Ѝ{*��6�7,����팯S� �nB�'��9	 F�����π n!��Y�j����E˦\� �q[�PS��bY�2ٞ�E����3I�:��eLU_�VѸV�
S]n8���i���C)Nםs�O�N�q��ɍ=��$�r^�i� x���I<\��)�d->���ءf�<yC
�Y�Tx��X�6��b޴bJc�4S��s�r�S��۟K�hm�'�Y�z�.�iv"OP@���'d�H�p�Ɵ�J�إ�t"O�T(�nY�B� ��DK�0d��X�"O����$@8|���׼:l�X��"O��b  <fU@P�'ѸB����"OB�E��(&�V]�w`M=�J���"O�Y:��s��Qj���	�zh��"O`�0�I�%!��Mr��%+�V�hw"O>E��t�
2sx�I�W�G�8�!��62�l9���ܠ'ˮt�dɗ{�!�%tC�L����	�|m	�HjS!�d�{F/rq�����$@!�Ė(b ީI����Ma�񂐔~#!�YL�zuڲd�>5�]Qb=]!��b.�r���^�����r�!�D�4%�ĵ����E�>��7�p�!�$��y�L� k�6�f��c�Y?sz!��	#����H���P��W�tm!�ӕ0�F�S���5�8��h�7vT!�D�`� �!Jɸ�f,�c(�!�^���B��T�b�1�D:Qe!�� ��̘ B��V�҅{TGǳJA!򤙪t��%��	�x�&`i���V
!�O8bq�@ �z��-H�E�M\!�ͧt�	q�N�5Xz@��f�8	;!��%��x��#ʉbW�-yt��*!!�$��Gvĸ��T�������;!�:(����>{�Z��%�]�$!�d�K���ٴ���T�玈�!�̫>5v$X�L�0/}L�2��V!�$R�*ЪM�f�42�;�	�G!�$ܘ5���kۙ�����"nL�ȓ;7���#b�	t�XP��`B�c�n���4�����ʈ�� �4!Q�`�j���g8��YDȁ�'�\��@�[-f��1��9ޝ0�KQ�,:��B%�F�$�4��ȓy=4����3v�\�R��U2x�V!��8��̧g�^�f��*A��h��ch@��$��17�Ѱ����h��I�ȓ[��p$$X�,hdOG��  �ȓW�p<��Æ^>���k�eJ��ȓx��P���+"���`n�4Na�q�ȓl�rPU�Q2x��L����
�D���R�aG����^�b�/I�����ȓ3��Q�ل+4�)im1��ȓuFv�A#jE>+O%�d�C0��ȓco�@�7���4�j���ˋ���(��5�Ԙ�6p���@U휽���ȓb�I��A�:1���8㢋�	�^����BՉgi�<�mpT�PIJ|i�ȓpt�M�b��1o��1�
�r�6A�� 1��I�9�ѓC) m%V����Kp��dvL�9�ĉCT���ȓU�܃�	р�%�C��r���`�(Yu#�'n3 ��V�^�^0���ȓ:>�A{�"V�@x6-Y���V�9�ȓ�����
�5��@�Ξ;����2`༳�ML.e��L�'U7F�2�ȓ2���c��<b� 8p�
<'hd]�ȓ~�)��H/!�p}
U� �QP��S�? ڼ�d G�K�pk!h^�=��"Odp�B�'e�)df^2]�0�j�"O��QE ��&�I��4v<*�"O���䊭J���	�cVc�쪒"O��8���y�:\𒉑(%�ݛg"O-�p��oe��q���W"�E�"O@��FE��#cıbu��V"x�c"O,���)�#P���U���u"OA��S)�W
{�r8Y�"OH��!��`�r��;}�p�PF"O}h�F�'Z/���N��g��ˇ"O
5���ǚ\����K�^c��r�"O�a��R�ZV���K[$ݱ^�������8y��#N�`���ZT�C�ɘF����e��c\l�����C䉭;�h�P�HW�X���ϴM@NC�I#�츊�ONh��8�W�r3:C�I,9/�٫�@]�v�l����9�C�I�k�F���l�D�&Y8�'�jD4B�I WO��8��C_�z7���B��,;��\���%la��1�L�
װB�ɸ�6ܚNY	50�4�t&^4S�NB䉗�x�R�+x�\rƫ��f!2B��:@�ΡA�ɋ���4�3D�( yB��46+�!�Q��N���eO���C���ɠ�^�z��X2*�K��B�	�:w��Ci�0A�l,�ЦJ�`�C��0�@��a`����ĸ	G�B�	�Bc89�v���"bH�$ �08B�	�C�B�$��9%h#���\3<C�IN�� �O�S�<3� ��
�dC�	&}��:R�M�~6��+�(�$(0C�IiJ��ьn����J�q��B�	��
�*�n��EA��*r�)�B�	8��9i�N�P�p	�l�
w�B�;���b��]}f��O��6>�B��N�I�����2e:�ϛ�u�bB��7��*P�؆��eJR(�CH�B�ɀ)~�Tr���0r��G�5<��B�ɑh<�h�⅁ +h�:��B7,� B�	)ʘc���O�8�آ��8�C䉯'۬@q���;_�`��AJ��3��C�I?[��1q��64�@�kS�-Y��C�?�l�E��dR�+����C�ɬTd��l6�~�
�J�33DB�m��8"D!�lŒ�e�-.�4B�	*3�rq3��G  
^��ă&�,B�Ɋo��Y��ä;�f�0��
�B��	u�l�
M
U9�C�3
�B��:M�̴���O_,�z�^�6*B�Ʌ@�*�V ݵ[#:�QC�ν<<�C�I�n2y�瞙~+$�dψ�d�C�I�I�����U# H�s�E�mhjB�Ɂ?���aqƅ`g�aL�Zw*B�ɝ�DP��Pby��r�i�x�BB�	�T�ҽs-�B���R�eO/�B�6@��X˂�]4�V�+'��)g��B�I� w��(�Ý+H�>�yfo�1+�B�I�E���Jf}�%����ȤB䉿|�B}���̈́F$y ��\B�Iyt�-_sJ�Q2I�c�LB�ɤ'� � 6��J=��~kRC�I�H������~*��C�?l�TC�	�7�Ib�K'������d�6C�)� 
�3LH�/^�����I=4��݃�"O�5d�"�"�;��� 㠹A�"Oks
0n��5ECH�`���"Ol%{����$(�7#����v"O��Ȗ��/f���A�p���T"O<X���iy A�cX���$"O�p��U2}��E,���j6"O�0�%�:iE�� �ņC�ґ�E"O@=�Uጀ	R�,��L� |0��"Ox��6�A6(Z�vn�	gh(
�"O�H���7��h��m+L,˂"O�<iս:���,E=2�z�V"O�Y�*k��c��*aK�514"OH��
�`�xP
D�nD�m��"OB�	B�O:9բtq�	G"�Z�X0"O�	S�&B�� ����U���S"O�q�@�	qH��c� �vI�V"O�t�#��nu�%:�c��]\�a[W"OT9 B��Jy���K��{\�P"O|�"�N�ZX�A1 J�#�^X�"O�H���AvFU��H�d��D�'"Oֹ��"��)��苦�0�X9+V"O��Q�hA��H���T:]�H� P"O�ݳ����jĻ���j����E"Oz��B��#S�p��� <b-��C"O:t���X2.h���'�0;�Ɣ�p"O��"�̘.O��es��
��D�"OȝC���) ب�cf�Z.*4ӂ"O���dk�2���bR�V�
`�)T"O aYWI�m;�Dkp�D	<��YZQ"O�m�$�9H���¤��C��,�r"O�i���X�g��
��nr��'"O:� �%�!�r�P'#�K@���"OX�q��Y[L���D��T���0"O��@g	�2�ܓ�#;M�B��"O~�K%�Kt���i� �dp2u�b"O:�9��U�ep���! `B|� �"O�1���"N�!�OP63BX��"Oju��AV\��d$� Q�,J�"O4=Ql�1E��HDd̤[� �(D"O��6�ߝVz��c��=�J5kB"ON<��B�O��tJ�델T����r"O�A#k�9���jػ}��d�D"Oj!�W�Z'n�R����Z0O��`+B"O���6�G�|�@+3��w�d|��"O���p0g��)zǜ�M�EK@"O�8��N� H�l��e�+G��`�"Oh��B�v.��ve X�8 7"O� )��c�j�
R.d�"�"O��B��I�6��{��$dQP�"OL��Ub�#z^D�υ=6��Q�"O��1 	'\�2�II� 9D�0z"O��$�D<g���$'��QD~iYW"O2X��m�'@������V4lbƽ��"OX��(Ţo2�hP�#��tCP\�&"O���5S7��Hk�[�J�<e�e"Oެ��)�ah��[�᎕P�<�"OJ�jWa۠KUd�Ʃ��$�H%�V"O���u�/#��\1F���ZDY�"O^	�un�9t��C`X9����b"O`u��hף(�*D�a��]
��x�"O|,J�j&R8T���X'#�<�[�"O��ڕ#Ĵ c�)��+!>P�1'"O�Xs�n��l�~�9��Y	4�@"O� \�#u�Ȥ/V���U�]��]k"O�0�#B 	n�˔�J�\9�D"OX��
цc�.C:>��Y�b"O�u8��	L7�C��K�w�DH#"OB��.E
7|�Madmܦ&���+B"O����f�@z��*I�N5��"O��1� S�!�l�:C �
Y�̸��"Op� b���a,l���P�Y�ĩ�&"O6��f\96/��PE��W�ڵ:�"O�����В	*��c�E�=� �����U��4����O>�H{
�P�IV�iZ��>�T]�� L�����c��5n���R�H�x!ȟ��ɚ��y']�lt�%1s�!sb i�`H�\�8ɷ�S	?6�R���^gT����|6*��H|JT=�1�p��3iJ����ތ>���cb,���޴2���b��#|���ص
$�^8aNP�ZN!<��օ������	��	8l6�cV��*t^��N�u�➠�ߴC�6�|��O)���i��Ԣ��>4֊bʎN~���i�O�Xվ��a�O����O2�d㺓���?��4ou\�i�B�۵U\
��7Uc�H9��U"���[���FG\*�VM�BB�= f���%&d�����ՀlA���-��	�jHe�m@캣�"�c$�6�ծ��,&�\��EP���(�wʏ��dB��-B�i�nio�����'X��x���nY�#�>�� F�F��~��'eb�'<ў�'��Tz��S�9�JQ��K:[�ubq
��A&�|1�ן�9�@c���6�4Z-*d�T�m^����I��x��'�&���V3�L+VIk�`<�G�N�#���3���!��!��K�}�0\9r��'�(O��k���;`4H6�Ed�� j�C�o��sd�	&�L�i�i:D�x�j%�0(.I�>�`(�՟ 9ٴi�uʆ,_ :�Xu�$�K��x�р!}��'|2�)٣@@I���RY��"�&!�d��l[��̼LdbZ��s��x��4	�F\��y��MS���?Y-��X�@F�09g6YA��/W>�3#�=iF�d�O��� V:H��É(� �R"� ���-D��"SZ��ZR勨_c�ȉ�hJ�u�b�x��铟2��9�EּE!G�>�0mPQ�T]��50��3��Aw�Z�A��0�2���Ʀ�B�~����	�aˏU�
x##�J(*�#��T���?Y���?�.Ot��w*J�:�(9�l$�bO�}R>I��'ў�S2�M�w�i��	:^z ��fR�'`Z�2w��.J�����6%f���'�����+?n^"�'��i��4hsoT�=n<��`_j����� �&��!�eʃa>��U��*��I�|��'a��}��"�Q>8���h� �PE�ÅA���]����+�^�p�
Q�/[����j]>(��:)�n�̻#P�p3��/�8�!B����;�'��<q3�A��?��}�`��$��jf���V��q�����?�����$1��g�v���U�
h�"�b�S'��Ɵh��4o���'l6��Or����7��91��H%H��V���8�"N�K51��HY,�B6�HΟ ��៼�	���	�O�7�I�5����#qǘu[F*F�9Wv8cBa�4f$��kTU�S�"l���	�zd�*��"���6����ȋ$μ5b�$�0Ks�\h��
=A�L��Mؿ'jl��u�a�a�)������%�$U�0V%HU�F�cq�����T�SR� #a͟�*�4ϛ�'9�	ҟT��쟄l�8i3R�ְ�|�"G&z�\{��'����,�9�L��a����Em�<��H�i���y�v��@Ʀ5��g�ǟ�Nʘ� �  ��     �  !  �  �+  �6  �>  �J  T  IZ  �`  �f  1m  ss  �y  �  P�  ��  �  %�  h�  ��  �  0�  t�  �  ��  ��  c�  6�  ��  |�  ��  � N � � �  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d�OJ�=���!B�Z����lm�%i�DRw�<��&ޢ+�6x�cJV%�%y��M}��'�&88$lݽEO2��!�M� Z਄��v~r �>0���#E����� ��y�F-�`ݩ�kR:A��a����HO���(� D�3�V�6�T��	E�����"Ox�cd�*l|-H%B܌|)�I�>O��=E��/<���C|�����y�EǴE4ά�G�1?e��ѩξ�y�"g���q��,o���!m;�y�Nɯ6��\`GȖ: D�`c��y��׊#3@���@�B$ಞB�	8k������+)����qN��Ib�C�ɒ��=K&�7F�*���n����C�	/V�����͆\��;�M3{���$����w&�!�(��âۆ^yh�8#�6D���׃˺{���r�$�����3�,��?���iK�I	!�GD�k�����0D�@�?0���i�n��M` �<D�l��H�:|t@�/B4B��Yc<D�0�bJ7�v�Qe'��#��)�`�8D��D�)3^հb�'f@��y�G!��n�RV.,��tP!%@dh��K��>������ߢ�ӳ��lWJ�x'��y��	V���)�B�4bE���U�I5#�C�	&=�z��@D�S��,��!Ļ��B�)� �`ZO����֎34�"O��:*ɫkk Q�FH�v��"O2,y��ǝ?/jy�,�0t4���'���'�����تF�⒈L� j�a�	�'i�ɡ��B��tXуڸ�>�h	�'�r�H��FI�J<�$��WV�z�'���i�-��3�ܡ�#
ЗQ6ݑ�'\�F�)�4�����K鴠�d�"c�:��ȓG�J�	R.�9y��L1wb�7*j��Fxr�I��=�EʀBvBH�W�=)�
�2$�"��~��R���Vx ��`�M�l_~�F|��S�~"�ic�D!%3R��m�>]B�Ƀ6P*��c}|��T�Ҽbd�B�I6(A�9�w�T�-.�8Dk�r��C�
P�r9(q�݅,�.��ã
�]���>Q���p��Ih��O��������r�<�pW�Ni�(�I�*q�eX"�Io�<��)?��2�]R�u	��g�'�ўʧ`�0(R��P��H�([�IS�ɇȓ��#-��J��AP.ݿn����1�]�t���i=�\��`H2z@8̅�	4�ȡ�E�D������L�ȓB}P��g.Ɉ �,@�I�G2��ȓ#t, �`RS��a�A�'[_� �ȓ3��� h�.1�n��a��+liV@�ȓdz��j���83J��T.@(���ȓP��1��.�"}���p��N�T��L(��qp�� p,� P	���@�ȓ 3����)v��8 b�']D4��i���s�^�K�`h���[i�a��I���%�в$e���/D:8���/ �7)�Kc�Q�.�>T����'��AX�� 0��uوE��(��'�hrB�' ܩC�j��.J� �'��0/���|Չӵ�F�X�'���[�H�2�|�!db�<'�][�'$�J�$Ή���H�h��U�01�c!�>�1�|*����M�E�(�S���7s-N��(Z�!��k�<�G܎(#�=��%�{��	u��p��
��n=��*�A��d(���EA9�O��, �R�֧G� ��.2vv:0�ȓ��h�� $bږa§�$��T��\XLL0ӬW�(�p��� (�t�� �@��g�Gx:؉��Ȃ����;T��"~�u���+F��a\cul4� �[�<�ѥ�'�><�VKlS�d����W�'|a����	qW��;`�%;��T�ba
��0>�x�H0DpH��n��9aB��"�M �yb	��ƌ���-��	�"a,�HO��=�'��1;bĎ;?Vp�w Ò1���O�3���k�`�XO�7/���u�i�ў"~nڡ=(�l���"_��ׅ�4D�:B�I6;xp �c�܀^H�M�D�@?m*b��F{��TC�?N�.�hf�1[T��'���yr �H��|��@Ե`�������
�OZ<��I>ܤ���: �H����C�Mä�y�!�&y��h�C��4�N���'T� \�T5��!�Y�����'��s�ΝO��|A���p����HjH�P�����xHV	Y�ć�r���`�^tJ�`�0�ą�	m�I�5-�"p�	O��Q!c�7`hC䉓fޮp����"���jg�K�ng@�<�D�|�
\�+O<D�eJ�_>8�cG��<��S�? R-h��";8�h�^?<b���"OZ	0�c�h��1���^;�E�D�'���p3��#��b y�c�s���8�D2�S�4a�z�@��]�2�`z�mR3ԨO�Ox���0E�>(`d����nz8�s��H�O�ӧ�g}2�Ư��:�Z�n��.���ē�hO����ȣ�F0j�t
� �?$b6d
2�'Hh���I��P9�֪��{y�J����|�N"<!�4�0<�5��6+gz���@G9'V�"���Oh<���̰klL�%^>y$hc��Ȟ�y"D�/9������}"u�ӝ�yB�� d0�	b��,�d�yb�J��"0z퍻t�.m�F�����=�S�Ox1x�̙<;e%2+�_��x:�'��q��+;$��:!.v�1wbC�I�/��)r��(�hh(Dl!1z�C�I�Xb��Rh2��dr����@��d�O��"~���LLv͚�(�}�V9��S��y��H	���3B۲�ڄ�ŋĐ��$xӖ��$݀c�X%�&��6��\�Ꮣ��!�Vxl���h�����2/�6Y�!�Q �>,B�o��[�����W��j����ҡE�k���cU�s�jh�*D�  $ȶ+%��i�CV92��@�5i;D��q�!��P`v	T"B
�H�8D��3��ʫ()�ɸT��!h q�q�1D��"#,�?Ebl;��0���l4D�DʴIT�q�b�+�RZ��3D�H�W#,l&���#ň�� ��,D��v� >a�qUK�ư�ҁ,D�8S�	 ~��e�~����)D���B�xWV���I�Kp�ԛ��:D�,���	z�Ӂ'U
 �n�J��.D����e�Bq�$� �w�H j��-D�@"� !)����g�0��� +D��2�G�>k�NE���[-;{̍���%D��s�ݵ`JJ���c��Ɲ���0D��`7吰�<��O0���K�K/D��X�$�i�F�Ӯ(�҅'&.D����H3��"�#f��<s�6D�� +S�d8P �kåeE0�#4�5D�@�	�H�	2ҁ��t�1��C&D���v�
�IP�x"����ɉ��$D�����.�c�]�';Ĝ�g0D���#Ȃ�EM�P�\�6ޠ�c-0D��x��6��e�7��7R��L��/D�T�ǣMN�y�éֹH�|t&/D�ܚ 	�� �ȇ��T)	�(+D�<*��1I�����,��X��$,D�[g*Q� �8j!��M�P��=D���cE�&��"r녳N�
P I.T�dSF��8_^ZeAa]4p��L �"O�	RL����5��N�pl��"O��r`��.,h9R�����ɇ"Ov�7gԨy���;am�S�5��"O��
��׾���8 -��~T�"O���`c�$?���l���B"O���k��.pKթ���T�ޭ�yb"�����ӈڢg�Vy��/H��y�<v �؃醳N�0`�Y	�ybϓ8�M���>t��RE��5�y�%��d�\��a \6 $�斩�y"c]�<p�v�P0?9�D{�B
	�yb�8��Q�O:hL<)���T��y
� Dy�)I�i&l����џ@RM`�"O0��&S2-��1l�:gD42�"O�}*�!�0 ��, *"L'tpq�"O�53�*;�Zƨ�O�ڸ�u"O�]�7ؼ>7j��ׇ�8Y�́8V�'���'d��'���'	��'�b�'˨-�taӌ5�}���&��c��'vB�' ��'���'���'���'���[������bD�|¤��A�'���'r�'���'��'�B�'�p��p��63� �Hm�=��'���'R�'���'	B�'YB�'�����pj�0� @Q<���'�B�'��'z��'0��'fr�'�ti�	�<ޘ���k@@���'���'T���m�I柘�I֟����Hb��׀c���#�)�*
s��PS-����I�@��ϟ��IΟ(�I���	��0�r�脍#d�ܨ����,��Ɵ\��̟|��ӟ@��������)���;&4P�o̠*\0�&b�ɟ��	�������I���Iݟ �I˟��%����Ś���;�b����ß��	럄��� �	ȟ��	۟0�I���pl �����g[�M�bU�|�����՟H��֟p�Iҟd���D�SI�+��a�iPj�"�a�k��l��؟x�Iݟ�������ԟ����T�ҦY�R���C�0<��t�����X������	����ԟ �I��M����?�a��fMy�e]�d��xc�h�֟�������������';8qk�,V�SVx=���E3<��I����4���̦��6�3E�a��ᕖ,<�K��2�M��lQ��
۴�yr�'�t��N��k\�X��O�@���3�`�y�I�wdF}���d�OD˓�h����F�F�*$HZ-!T�<�G-���htF(�	q�'x��w(,� EԽ!�dL�%ܖ)��!��b�"�n�<�O1�~Pr��fӲ�	�v�Ъ��5�~��b�3Y��I�dXc�X�S�8G{�O	R�\2,�x��([�t:�@Җ�y�P��'����4hP���<a��I�wtH�"Q&,A8���a	���'kP�u�FeӚ�J}B$?1����?^�{SA����d[;Hq�����1��鱖e�q*��7��+B���B0<���]ﰈp+O˓�?E��'�}Z�N�����:���'��I�'��7-�?uc���M���OMBMXd̀�;<���AԽϓ%כv�g�@��2y��7�!?Q��=I�]¶�.����G5+$zPhƮ�7�2��J>y.O�	�O����O����Ol�S6���=����-_GQ�p�<)��iu�`
�'-��'���yBș��H5�Ӏ�n�<H���ϸe���f���eӒ�%��S�?���u��ظ4H�+)��a��,�y2�(חH���'N��7L1Y���R�ILy"#j�+��g�Lঁ�8�r�'6��'6�O�ɺ�M�FA��<A�A�?�����.7F���T�<!��i?�O�8�'�@6�����4M��0� F"��
s'Ix�Ӄ�M��' ��75h�"���D��I�?a�]�y��M���
�&AFY�c�V[������Iϟ���Ɵ���l��<.�a���8��:䔵o��Γ�?���?k��W����D����Ny�+H%ft��w�P�S�z��v�ԱS��O�Xnڪ�MS�'yLPh[�4�yr�'��Y�aƹE�Vl3Pa2Q�|,��,S�I�*��P�*��'��I柤�I����ɮO�Њ�-�T:��dPD��I���'6-��Z��O\���@�	K"��ꈥQ��@,�w��	���$ڦaP�4	������O�xT)[�v!��jQ�R�Pt��ӞH<
))��� ���I)OD�	�3���sY(,�Σs�ĭ��
V�Bq��b��?i��?��Ş��D�ܦ]*5'��CN&�P&�	06��!H�RU��M[����[}��q���lO�AEA�P� �#CQ˦��ٴ$�l���4�y��'[nx��Ėe.H+�]�ܑ�D�|���+	�L-����b�Е'�R�'[��'�R^�據d4Z���^u<ԣ��j��i��M3&h|~b�'f�t����j���g紵��n��|	FA�'��.�^�l�&�MC��x�O��$�OT���i���B:�'��)gΉ�� �b�ة��U~�ȝQ@�|�S�T�����A�FL�!��CB� v"����۟(�	ܟ$��xy�mӠ�@?O��d�O:8@BW��z��M:UƲL���Or�O��'��7�¦�YO<�!	입��X�}j؃�	T�<�� �2#�
S����-O�i�H�@���? rx�R�Ʒlw~T�#֖�?A��?���?y��9�Ի�:�<|��� �l� ����O�5n��O���6�4���2��\�E�xZ���~����5ON)n���Ma�i�0�� �i��$�O|�k��%H��Ū�
ZFX��2�GX�[��};2F��bL��O���?9���?a���?���wKP�q4�2S���iБ
m�-�/O\�mZ;H��X�io���#���Of�c`��L��xI�G\����Ls}�KlӴl��?qN|��'��t�U'{�ش�ӯ�f��x�눜u�-�D�,���^�'H������
�,����2�0MAR�v�J@�/s�4i�D�C�#˔��'�J�5`�y;�g���0��QF��z
H��o��"��,�P`D�O��30/�0�M�3DJ65�2�P�7׸��3�;;�܍�mo&�x	Ⱦ.� ��O߽Zʮ�㍒:%X\�a -�-Jfk[N�ȐǠb8��QI2� "G�&J�� Ô�UL3�U�B��+d��9$�5B=p�(��Ҏ$�ukG�>{����ؖC��Ըv�i�Ƚi�APx�4����z��C7f�>���?9O>����?���<'hA���SR�~|8�d 'N���'��'U��'
.� ."�'J��@�!嬑�'�W5�`��6P
�6��O��O���OP�2%K���'�h�E����$�A��j��4�?���?��=t��R���?i���?��'�B���S�:�� ,RҸ;՝x�'+�"�
@���q�y����h��1D1��K[%-��	��i,��'F2����'m�R�(�SWyZc� ���Cb%��۱QjVxr޴�?���"�~����u�S�'4�j����� �8As�� X�l�3cn]�	�H�����S�$��E�4F�p�2Q+
��x\�ݰ�O�y�d6-G���������|˄�9Q�� R�D�nʄq7�Q��M����򤕲����O��?9�'V���j�������M3� �I��'�ɹ-5�8�I|����?���x�DH#qܱp"-և'iX\��a�i!��@�"�2�';l�'�?	N>)q�ܜ1�T�VmN��F%yÄ��!�ɽ�*����6?A��?�����܃B5,4�Ò�zlf`�!DR�5ll�ßc�	���I�IdyR
����)h�m��tшc1,_0S�,��y��'���'��ɑs&PQ��O֑ �S�Q�4� ڵ$��O����O��O���ܜ�'it0���4C΍Y�#�
j�0�O8���O��$�<�v�T�E��OB�C�˛DUh�
0�O!a�����fn����O���?y��u�
��~
p�J�| ���C�UC�:�yA��Ԧ}��П��'�����K1���O���Ʈ�  -����O�m��$3��i����h�	���#|"��k��X�{���$�� p�uB�}Ӟʓ^�&=醽i����?�����I�L<"��ŎYk��i�E	ۘ~�7��O���׷<�*�S�4��ēn��XB�G�&�|\R�cVfМHmZ��T�3�4�?���?)�����T��Ld�h2�A��l>b�c�d/K�x6��h�	Ryr���'�r"��*��y�g�<�*"��B4`�t6m�O��D�O�)��,HN�i>=��П�bbD��.r�Dr�O�H��f`�����Od�$��1O���O���K�������Y���9U���8���l�џ(�SEժ���|Z���?�(O���BΓ%
�hl�c/��� ��Fʦ}��&w��c�P�I����I`y�ѩ>/&��%�9c�,pFM�sF �s2���O����O���?��Pqf�I�.�q�4�X�î�T8�a�E��?a���?/Of���	�|Z"��3����A�!.2��q��K}"�'��'���؟�I�z.��Z0���a��_Bp���ʲA��i�'���'b_�8��%N���'u0���Ο0 y���F�J���C�i�"�'q�	ߟ���"l�0c?��DOYH�y��抰ӊ-:��y���d�O��D�O����KTަ%��ٟh�I�?i�3+�6z�T�@�㗙0\���"���M�����On���<���I �y�禱��	݆bDQ"�H8w����t�4��O~言 U��i���@���?E��Ɵ�A��M��HB��K���"W�Q���d�O��S� �O��ģ<�'���&�t"5k�"B��`�☺-I~6�ׅ4��`m�ޟ��IП`�S�?����� �I�4�^�������E��B��h=|ejٴ!~�|��?+O�i �	�O��(B&��B��"p*�#P@�L
��������؟$�ɡv5�Q��4�?���?1��?�;#�Ld��W��P��3O:����'��	r)���|���?���پ�P�hӁd13a��1�qսi�҂Maު����O�˓�?�1@�.ԉ��g���H+Cp�8�'�Ȩ�'G�I˟(�I��'��e�$M/[{,� ��2U�l ��C:6��ꓼ��OL��?���?���
H݉����t�^�kq�J^��M��?Y��?���?�,OR%��J�|Bԍ��[�@9�E J8|��Ó#�Q�'1�\�T�I���	dM�I$c����֤�,.��Ԩ�H�2g�ʙ�ܴ�?A���?����?1�'���f�i���'���q�%�M��aj4# '�uk�p�v�$�Od��<���R�D�'��#by�ȳr*� `Z�3P���\9�@�a��OF���O(�$�7e�J�oܟ����4�Sy&��������&eM)B2�9۴�?�-OH��$g��Op��|nZ�<���eh��z ra��$Љi��7-�O��܍t�	nZ��H�	�����?�ɹ`��B�J>#�PL�u��*:�J]��O��D��F7T�d2�4�T�Oޤ���H�2�J�+T��6�ڬ�޴O"��/�M[��?�����'�?1��?���ŞDZ���F��&uu���?����</���'��i>i'?����⑎�w[lI���"�rX A�Q��͟@�I�
�<(ZL<���?��'E(	�TjɴWf�R�@]��l��4��d��-�S�$�'���'�&1��!�*TK*����ƣV���DMq�6���j���$�x��ş�'��؀[���`��> ��@�i�=��u�4y����d�O����O2˓iI�YK�h�9m��xv$S��%R��8��'���'a�'���'@)�"�C�6�θ�q��'F:-�3�' ��'&2]�`@��������
�c��y`%�ѻ%�@���@��$�O�4��O�$e�
���1�<�٦��z^-L�7��\�'�'�2V� 9c`��ħ}�LC%�/b�V��L�]����w�i)B�|��'(� 7�y��>� b�p"�C�2�|<a0j�#}��`��iZ�'�I�~Cn�
I|�����"B	�誱�R�M���!�O,��'�R�'\!��'0ɧ��)2pF�U�ٰg��86 ��/ݛVV�X��o��M+�]?����?)�O0-�$�#q�@	���c��i�2�'�D�h��'mɧ�O3��{��(�QR�Z<fn���4X��a�5�ij�'���OL�O|��ݣ}��i�R��f�Y��-*��o����I�Ix���?��)�$�(	tN׍~�m�1��+�6�'�B�'	�y%�<�	ڟ��u]�6EK8o�I9�a�2|+Io�`�t_�8�N|b���?��C�Ūѭ��H�17�E�z���i3�H��6�Oh�$�O�Ok�B�ҴsC��?-T�h�n�B��	T����fy��'m��'��	�G;�@3���f`�&��e�$�Q������?����?�(��I��׽K��i������K����<�,Or�d�O����<��	B� 	��Jg���5;D�apAOI1 ��ݟ\��O��ݟX�	����1Z�d��C��ն�!ʵ̒h�'B�'�T���rm�,��'/��dqQaX���u�K!�µ��iOR�|�'NB,���>�R�þ{�t�I�P=P�:���������'e��ZU?�i�O����>]W�%�Ӭ��mz���c͙��4u'�������-�S���.=�`����� +�W+ƒ�M�-O���vOY������|���d��'C�={s��]�RH�!��;	̴��4�?��d�f�����S�K� 8�e�K��Lq��$��<S�n�X@PԳ�4�?A���?1��u�'|rđ1s�D�,8dd�#�
�6�S8	��ħ<Q��S�Z���)4�~"��C� �q��� B
�yj����'n�!8��RIJD	�t�.ᾀr
������� ��-�J��լ��oO"ɚ�*�*Z:xzB)��J�b�Z������Y� ��1�:8
T���{gri�1(� vb���,��Ҙː��4�"��3�֒x9�Q������Sѫķ$O�)�c��
)�X[��9�r벥�l�Le(�e%A`��@M�r�D�KTG9!��	�������'[�`���|ʦ�K"v��c���rzu�֩��A�"zfjĴ&1^mz2�׬�M�n4�Oɮ����3�iZuB�ք`��!ᦁ�ad�bFt���4"�z�;�-)Y^ُyre���?I�]	�Mj&���'Yf�)s�[,��p��1ON�ж@T���#�F�,'�VвÓ�hO`��6�±N���JƄ�B�ig>O��l�����'U��s&�~Z���ID�
�.8Q�?i���?ǜ�	���O���O�9�0넀�А9X�� 0�A�
R1 ����()媌jdZؘQ�����<�bo��6�֔�śZ�`�RC#1��i�pi�Q�I!x+����/��L�Q��Ӵi�O��(��kVn����
sn�ab�=���k����`ぼi�ZE2Q�S8O��ш�A-�O<�%��a�Η�a������m��k�m��R����M����?*����$��O��$�O ����-���G�U/ *"��T�_�Tl���G�x,�qc1����'���?�N�v��X��ԩw�VdX�G�~h60tM�5ț���8����O.\�`�5_�p�	^�m�E���4b�$�O���?�G�������v��w�^Z1K߿߄���?��X: ɻ"��B�r!��7�T]#��I�HO�	�O�8�rGϟ dB&��q-SfB�OX��K/��m9���O��D�O��$��c���?p�Z3��3[pt��u�6.J�2&L`�fASj��g�'���F5���!���chV��^�RD�r�Jr��P�������dR/O���'P�B�N�)ҭ�55��ĝ=y���'Yў|�'o��)S$��[�^������.�(�'QD�8}�؄�����v�v�#����HO�	�Op�ROP"2�i���w�I P@�lAR�ˋF�n��%�'�r�'Er��\��'g��v�<���֚{�p�St"��:eVؐ�\1}|�TǤuQ�ࠠ��)5����[����F+ʿu��A��#@��`��$��v1q���-Jи�sO�;� ���d� 9�Ҡ}ӜM�Q��,V����B�5pb�,��A�f�ϟd��C�S�D��?͜`�!�{�lY�����y2m�*��2�l�0���I��ybAmӄ���<�&����	៰�Oc�r�%�n�}�Q��8�j5�pn�4%U��'�r)�?���RR�\�By�J�̦�'��3��"Wj��4��[�JDyb�Ș5���;��C;#w�	�_��'w�*�$������a!L�[k��<��f_��d������I@���_�o� c��#^�x��tB���s�xYF �8�䅨у���4d��;�O0'��XƧ�;DY.mc���3~�cHe�8r��ݵ�M���?�+�n �k�O�������o�Py��A̸P��s�%E9_�*�Z���otK���3��T>m�|�	q~���1�G`(Y�5�A��>ѐ!G(��}A��oO��#�F
|ЀR�ܕs�a.�Gk�&��ܔMJ��&AH�/���E���?���������|h�,kڬ�S�S��`���R4�y
� Ȁ�r�Xl9t� �%ga�}"���O^�Ez�Oe"��]�|�U�8\\�1�T�$=��'膕
aG͛�'=��'J^�]Ɵh�I�dM�	$`9��*���*;��ٕ�i��⟈} r9�ËKF{R�ۍ6�����F/`��Q�1*Xmڽ?`1��="(�3џ2-����}�� ϔ2y�	�9�H(�,_/U�}ؤ�;C;��� e���d�f؞,`R� L�vahg��6�9i�?�4���MԊ��fA)kd�պ1���.m�$ ��4�V�=EKP2`��S5�H)j �0��N�<Î�(ѮD1��6fb~�Ja�<��H*e����d�s����čQ�<Ii�U�V(�c撕_����G��X�<��$O; ~���R+�Y��DbD�P�<�2���y=����ፒ"4 ��+AM�<q��]SX)��k;�Z���O)!�[1�貢��|b�#���Sr!��\,l��E�!C�v��,cA@�47�!���wjƥB�D�$bK��q
��!�	7+9@t�q�M�G3�PI`w!�$F�$V:�y��:et����*d!��[���I��`
Q��w�!����Ip���_<@CGaȗ"�!���2�$�S�HQ�$[�Es�&��!�d��A*��2��H�C����Ŋ9�!�_�0��Bɍ9@4EzD��'(!򤈅�r��sݮ^/�m��E�9!�ɖf^�T ��܈>�ف���4J!�d�=%d,�̳G#�����^G!�dI�Tk�c���(m�,X�K�!�+-ᚥ��n¬|h>8��́)l!�
�>����K��{�P��ԣmP!�d��%��4�X6C̶@E!�֝7"�����_16��)���>�!���%b��i7�T�2����t�_6e�!�	`Il\3��a璤����.�!��s=y�F`�>[������X%!򄍱1�~A�n�}C�<!�Ē,kA�a���p[`����=G�!�$�2]8��	P\�1(&� WC�%Pz!��0i7xT8')�qHAC�Mv!�$�}5����"�	�>� %�!o�#�?9%a~�\�ZJpR�D�!`�x�cAEܗ��=A��;��DY��r����
'���$��Y!��H?xY��q�g�'��S�`ȗc�7-�zN�M��<O
-��d��>p����6����ζ>}�Ug
L%J"OlP��.�4;k8E���p!i3�'h���
6��ںò&�{�:A�*����R�P�#�,U��D��-*O�y�+�lզ�@��j�H��4ę�y�@;B@�'UL�rS�3F���/�g��} U�w����R��)��
�?:3��㶧�2�'�fY��e_92�dA�f(CE�^���}i�8�ł�C�x-xV-I��y�G)�� ȷ�E�P `�͔?X�4�p�"�<� �?�'KPb�ń�yG��X��s�&ԡ+z���UH����?1���T����m
�8����#O^4La�3�>��O��d�h���oF�3ޠLCO��D̄�"�4`�"F��i3<�F~",� ����4q�|L���M[��9v��0���>��P�˕%�~�a�.cz����	�/\�"ce�� ��@��!٦ʓY�:]���9��e��j�+W0�Y�>�S)K���6�A����7#��^JB�	"l��qІA�;8a(��c_�]m!�� 
'-�Լ��1?A�O�IQ%^{b�h�0��&�:��ܸ$`�0l̼rO�"��=fL�a&�QC���o��d�[��& />�m"Gƚ�M�e.�q� ����Ԡa8����"l��E��B4����Oر�	�^����U��lHť�u���39O8�QU��Y�'���ƙ~�O<�0�n�,b~�3JƝh<��V�`�����=B�'�L��r���禹��Ob-��ZP�)Z�T{�Ό+�MKD�U��J9A�'|��� �q��@��Ú/E�ة�
q�`8s�>}"ܟ�t�g�? �ŠuT+��4�Ů;���3�(�OF�E㒕6C�Q�Ͷr���2�œZ�<�IP���Y���~��'�jT�d�ݰCh�I�� �:���f	�5���Y��$�3C����B�W� �o�p��A�WH&��Y��G(;��l��<��nGy�֐Z�|��`:�~��'#ۦ��֫|�NM8#��w�j��0N�";���9u\�PK^�1��;�E '&��|�'8����1sc<����W�P�1�4T"��2bf��2X �����s�pYG~2��$A�����)�;F�\�G�[�
�L�A�;L���܅:���\��S�"騉��/�"G"X ���1R�,�"�����0>i`1�$e��HV%[�֐��!�=)e�,`�IB�Z
dT$�,b��Ɏ�r��ӑX�j��&#�$A��mF81�0#?qQ��t��k!J$/�Ӂ�X̦���F���`Z�	wjh�g�(ik bP;�yr�i`�I?�RkҝZZ�ɉ�NY��Y�`��kg�P�(dlʓ'Q���w��)y���u�U����l:�i-�v,��,�ԁ�ӊq�d�RW�D�i��h��E�:��DV5�J5�r 8�<�89a�¤h�T���(�.(L�����3&,M�Au���)���ڔPԡ�|JC��\Q�
D�Þ�tm��\�4��x��'dB��=~l�7��;uo=jA�O3,Nz�A�Oц<H�u�ٳ6�x4��'�	~M�3�xᗨ�$� ����s/,�>�4�7>	��C�E�[Y�`:��b�7͒[~��3��M��6�I���:�����o���5Y5a��@�.l�՗��b�Y�\ڬO��"c膃Eܴ�#�I�QvՓET�,ࢅ�?�:�����bzt����D�VF8�w��'���"�y��/�a\j�8v�3=Z�Ĥɨ
~��­&�Q:(`��ߒ/	*TP"a_;k�(a���!����R%e����R���������>%�R�	8o�tE㠳�jǑ�/9T��0�M�
��yWNI�U�� %G��kAh9��d��4e��X�(	+z4I����=��H��D�ɮ���]�s6�XV��020��K� fazRY8Y���J��] sn���E�'Y�!��-	�R�([�)� (s�YX����u�"��t��A
�t�'���2��4h��*����P(�y���\]Q*s�Q*��M��c����9ORPR��C�)��Q�Q�O���;P��/5�	�[%�����CUZ�P��IM�v��1B��L��QXP���a��Ӑ`9X#	����Erhx���(e��9�'���Z��89���B���)wF�D���ȴ�q؟��WjJi���b(�O�	�3�;%��b�'�x�0�'%��(2o�?�۶������K�V|��4LOBY���3�>�QTΖ��K���b0���m݅��iK�(��?�'��$�O6𵯱�:�6���z�kиBzX��~����<Y��%>;��kGa
�8�)@��`��'��Ԡ�_�<��AC6��Y��'���˷#�0t�@`񔠌�/6�#?d��Y��9G#@18��Z2��:�H�Q�N�3���e�e�l��gyR<O��9d��ݙ�!ާ3V��೨ 5a��A"�νɰ?�"ۨz7l$b#��*�s� �+°��s�V6r�I`�������RW���9}����
q�4y‌JV�����x���zӤ8�4�ߓ@�hP��=������>��%(K `�5��厾z���� %>������dω=���Q�ε�6�D��	l��'�l�۴�����G~h�w��6�S�$t	"E%&���jw������A�O�7�ʾmn�:d��:�<��L�\�'�08�S -֤@u	B7^��:Ũ�#�0жh]* ӧu�Oq���c�B"��Q�w�� o�>��Ta��~�(u#�֧5椒,B��	���oS�)B�ɬ�O�=��dx�8� ����"�K0!ݣ~��H��疲�l��dR�}L����%���00�K���:���-��{ Ȗp��ڴ�!��f�9���2��F��1� �V��	��:*@�sjԠ)�4i�2c1�dĀiU4h�6k� ����
W!qO(x�uOٛ= J5� ��_^J��7�i4�P�&�����[	?u�P��d�4f\�L!�@�I��D��2��Ma���P^)�E���p=ѓ���\���ȧMnuPf�}�|�:%�5�Ok,ȑ|�:�����#:�s@�J;1a~R���X������V#\�t2���	�5���)�p<����?"h%R� ��&��� .V������p��m��KF(E�">��ɚ�_1Аyf��<~�
�`��<�ES/Fr��!�טQ���+Rn~RKB�q�����G�=�a���Q��O$uk��FlAR�O6]Τ�"�'yh��� %O�ea��\�k�$ti���-fp�����P��<�Oݗm�`�YI�
�ד�?��!��hcc��{���q�ԟ�"�S�B0|ON��;'Y��Jw@�Y~@�1`M7z���'�f��`���� �!g��ܸ��Ո*j�`���#HX�'_D�',FUS��m~@��'�n�m��0`2T/�'C@��W���iI��:9�ɂ�M�u�#�a RЩc���ϓ!b�K��@ .+T�I�Mv�,D�'���R/��v�ؠ̓|q+���oz>��a����ő�ڷE�آbM%��
�mI<I��|IU��jV4P@u&��P^�N"�!ov����ۚe6�9�E+�6uv&i��'���[b�k�h�ۢ���u�+������ܴ.�J�#F�_�%pa���37"��V��"D�tZד��� ������l��]� F�I|�\9u'��]�7��K��)�5�i�N��'KYL"|Z���1>ؔ�Ͷ��=�%]V�'���Į��추�ɰni����4'�8 #Tˋ(ufxl韒�n�q6�ijx�F�,�-�Q�J��0|R�#��D^q �)vA��ƕ`}�)V�8I�' 
��MS�+������	�)�D�1@�y`���Â�"��eB�OPm�Na�,�)N?㟈��'��:A�T�!W��n�(�k�(����]��M�T��͟�ٴlz�i�6�T��D�l�z��Ȱ<�b��Cb��N��Ī��,ހ�'"6LObԬ񦅪g錱+vԉ��BS|jAC $?�'�j@A4�����s�l2p�*W(�a���V�':� ��d��;�T�@5�<67*<�5g1֧͛ǃM��;Dg��r~tљd�Lu�z=ڈ���O$	�s��e��7�H������#^WVy�F�U�ȍP��M����K ����Af�:7���`��k+���I5.иs�����P�ު���7O\�o�\��ZU^D�W��+������K�$� ��ťLʀ:f"ڲ!b���EB(b�Z]�O��=�����Y}V�+%2�l��S�ML�M��o�0!=�Rד�yg"�&r܂��Z��5�� �>�8�	���!��)���Bh �mSrdj�&�l����0<��(��3�[�h��H�h5򲅟	DZ�TKeDE�z��X�֊���C�]��iI�譻oURS���Y��8[�"�s�,ԑ��F#t��4�� �8{�2��U���k�Q�5~6D����z2��j��f�dc�O3��ɴK7*Pi�ȗER��A�CF�f�&L��'ž-�V�]��4I1i*�WB\��iO�E�����ȳ-=|�3���99��X a�<�R�Vݺs�^�l�'�\o=��<i��?��L �o�95?б�����C�-b���\�H�1�l�s(ԛ�&ܢY��Y0�ia"t4� �9�RͣTg��K] A ��\�Y��$�:K>�G� �3�� `-��t��-���B7� ����2y<�aw��,tbĔ�x"��t�`��e�3 �=0�DW~�L<&�
n*0��APÎ��bx}R�	O��r����F�r�t�'����+q�S�G]��$���C����+�R7<Dx�-����X:�?LO������@IHQ�LU!-oHDQ&e[߮p
����<����O�3?%>�`�'��\=<$ѣ�%L�=i�+%�Ov�Z�_�?xZ,2��F�\3�`���L���ߴ����cv��o3zp�s��b��������Kw$mYC鄣#��ɀ�	�XN1E~"a�:
�t_&ψ��v����uG��"�T��K;p��d�W`$�,���[�;:����4!,���xb'�S�p���C ;��$���9���/A��`�@��cf�K�����.�3�K;;��ɶ����l�o���E��=7����#\O�<CADS�'n6��ß��XQ���<y�n�ڦ�1�h�!\���g}����S"z �9��(�-"�A� +I5�R�C:�J3½`{6F�$�D|iTC�)BJ1Ƶ`'�� �y"C4�);ހ�N�*��E)��џ0z��A�`�����ƨH���s DH�;s���y"/��m$F��u"��qx��#��H���Dǩ8^��o9��S�Ol5�&�
8�~��n^�"��,q�'ź�z2�\�b�u��&G(I�aK�'	���i�?Wb����ɉ@�X���'���`�� 0�� ߤ<z�J�'��i�,��&"0�f�P�L�
�'*
�"F�z�r��
�JB91
�'���#r�\%4��K�d�0C��T�
�'|��h"I<~ڱ�7-�5�d	�	�'�"� ��̝�d�H��3в@�	�'�<r�IN%W����1Q��l�	�'d*�c�-�$m>�HBQ鄃�=2	�'��q����U�z)p�#�����'��h���@̰���	:e��ѻ�'Ժ�eۈ#z�P`��4*f,��'�l���͊Xz�H�L8$M�Y��'4H`�Vn_`�ށ�W�K���,K�'L>��%�g�F!�'�D
�� z�'#Zi %3�"�A���x����'6b�I���.B�t���G�l9#�'� <�'(��.-��g���m��%B�'��8� 	 늴�"cǆ0����'��$����並�!� �Y�'M؝sU��^�&բ��Q6���p
�'�4�U��E�<����g�H �'0J	 ��T���a�U2u�!@��� fQ�4�V6G�T�C�2Z54̑�"O���w��Y&ݪB��!d2�"O��2�AY*#�&���d�P��"O~M��DT>^��*��M��mi�"O̴�q�Wj����/�(y C"O���OՆ;�^(8W.�QTaQ�"O��zB�[|�F[�M��5�S"O&�Ku��,8��AS7B��3�"O�|AD�K'HFd�isa�&e�i�T"O�٣D�D�.�q�`J��\��"O����O�Kp|!��ѭD�@J�"O޼����s�y�g��+:'d(� "O@�+C�L�`��ѓ勠/!�أ1"O �eK�#����%�����j7"O�T2b�9m\5yP��  =J�"OP �q �acF@$C��;�"Oz,�WhY�w�!��Y%��D��"O��!ǪM�sx�k���T}j��"OJ��PQ�g��I{��,R��"OdS�`�N7ޜ�pg�.0�)��"O
�A.����s%�!��"O�iB��  )�٣D̍'dq2e"O2q@D�{pH�a��6c�a��"O!��L,��]�T��=R�]�"O�ؑ��G�RBi���̗=�&1"�*Oxܨ#�۾M,f���T8����'�ԅ�v�j�%:ǩ�S$��x�'�@]�AK�tL�W*JN�j�'n�e�sł�Xr��a��C��X��'�j����Q7c:U��J�*c�!I	�'���3� ^7j6�)��Ɏ�^%��'"�lcN�4~���Q������'M���2۱�4��1��'R�E�	�'vҽ�U�#ifm*���x
�'�z��
&6j�)� �#	��p�
�'�(�$U?@��Y�#^��\�
�'l(*��";����͠y�bp�	�'�b����7�n��s���m(΄��'�d�3�㏥G�f���.�:0�aP�'Y Ȳ'+�6�ɈQ��2�z�;�'j��xcI�-P���E��ht��'ڀ��	�,tg�( HC�\���'' ��@Q�R��0W�CUT��'�.* Ā�hѸ�P!H��e�
�'(vX9c�X�,>4�X�f��l�2�P
�'�\L��	��d����^tb4��'��c���3vgj1PJl�tu�'�A�JX
(`��k�e��)��'@4h���
�pȆyת٨ho>�
�'��m��V m@V�G���3
�'�&_,!�V�6$�+�ȡ��'�ГUP0<z&i@��ϡ4��Y�'LVT1Q��>PN�R�$[�,mf���'�X���
=�4 �� ��Y�'�x�;1-	�#~̴5 �3��P�'�|Q���ժ<.a��D��.ͣ�'����� P�B�H�#�#/����'d����#bӘP�wj�4sȦ��'�<=���~#�塷�%���
�'x����hS�[��廇�N	dBV}�
�'N@�5
�1+�`�g�6eۜ[�'f�H��g�y��{�-\a沍�	�'�`푕�*!V�p�*UTx�
�'1$�y�����(���2DG�];��� ��[q ֘8�R`*1%�(r��r�"O.��v�� <2 ��E>~�vd`�"O(�z�m_�Ao��7 L 
:�"O��У�`�Y�����6�8M��"O��s��ٛ3c�a���!ٚ)�"O"]��'D�*@
�٢9�6���"OHtq蚇q��L�I�8H�"O�ڂ�!O� 8�êڥ8���q"O*}�u�ά�����k�a�$8��"O�U�r��g��q�)֋
i��"O�0i2�D�m�e�T���xM��
"O�8�@�=M��M����8i谂�"O�3`�?a�cd/[�	�p:W"OB������XpIq!0#�L��"Of�PHÒ��l�����R�Qa"O�[W�	b��CJ��F޺ij��x��)�S�5��Б�/W�E���&�V�t۲B�	2"%Z�ْ��_v���U-7��C�I�t��pT<LQ:�1��;��C��=#�8��$�?8� �E�99|C�I(L��nB�F�� �%��+>C� 
������q��;$�
3�$C�I�86U�`"��H,��R3�J�4o�C�	�b��{$�D�H G)��e7�� �'n�< ���|��Ȃn�%	�Du��'����c w�\T�Al�?W+����'u��ZFi�L@ ��D	�x��'Mb�錂w�
!�4��,>j�h�'�FLåK].'��Dӂ�%J	�'��劢��.�m"Eew}�-��'u���ħ2o����t�n����'J��b���>�8�'�({��)"�'t��a��7?C�H��I�\�h�'��Vd�L�D���Iy
�'>~x�V,M(D���L�Y�����'� ի�3H���9#�ޜ��yI�';&$�g�7��=(���{��Ļ�'N���&c8ndc���%�zY��'1�6E#��	@a�[���	��'�����ż�n�e�a�`h�'�(����#e�ȡ�3c_Gz��*�'�J8 B䏥,dֈ �oL8�|0�
�'�ބ:�ϗ !`��T�݅,�Ơ
�'�Tt	&GD�u�P)����v��ա	�'�~�Ac��4?�ŚP�?
�a��'ܲ���:���S�F�=0���
�'�@��b�"p�L��C�%�ءX
�'�Ҡq�ϑ�F�2H�BK�-fT�y�)擵#~���
��4	~��d ׋D
VB�ɽ!udY�n�x(X��I�hC�I0�<0I�"�G���)Tc�T.C��<+.����]�T
$ͲqC�	�~�"��b��'h�U�.�.�C��<X��K!O���$Q��»
7B�b�~� ���	r�x�X��ܞA��B��.T]N�`O��T�XA��[���B��*� ��C1F�Ryj�!�3ʐB䉭*��z5A�8&[F��N�B�	��\�{S,�P��<07��-�B�ɯ4�Pq@遇C��\#PLs��O0�=�}��ᎁ+��h��J�RUq�`�z�<���B5���Sԫ[
j�^%�b��x�<	�Ő.��(B�� 
=����l�<)�kJ�[u�y�D�E�%+�Lk�<� ,�Z,4NISQ���� ��"OtI����X��`̼�����"O�D�5�;뮅p6`�,`%��)�"Oz@����6�� �Z)A^�ٔ"OH��EH�Q%���uNC�7��Y��"O�Ѐ��ϻP�HgM�v|Ҝ�P"O*ى֡��y삠�'˒>�*HPt"OP�ƣQ�
�`���՘a���*�"O�Axף_7(�< �v�\�E �0"O8l�����i��&�x`�"OP�k�J?��!j�A��Lǰ�p�"O:����=�� ��*E�; ��9�"Oؤt%_�a0����=�ة��"O��V� f�qc�� i�T�"O6����	5t	$���.��
|� "Ox�{�l��Az�,��"L�`�q"O"p���]�8v���N��*����Y�8D{������d�Z��6`�!�$�X�Du��i�"B�L�@^=Q(!�$"`���TN�tt.(�_� ��'BLph!j�O�А�Lv,(��'N��(�#��e���^s}ؽ��'c�1"t��#x�\�1㡚?i�=x�'�H�vg�9k��%��ĢtrP,�'ў"~��#A�z�*�ǃ��F�a�aZrh<y�)�T�KCn׊ ��2󤜹�y�,ވs��t����J��)���yҭ�7p�|ي��TW��wl���y�˰#谩�"Mƺ<��M��j��y��P+н��'�'�nX���� �yr�AVO�a���+0h�9v�;�yb B�5��x��%U�ije���S��y&H��`	J�n�l�%S��y�"�
<�a�oPb��Q#g����=y�y�c ����rR��?� �re̴�yb*B"|*���p��;Ih�8n��y�2Hq���6J�*�s�`V��y�@�h�~�yS�x
��c�N8�yƗ�E�IHs��n@Yc��&�y��N�,��Ƀa�D;�2$zTMX��y�dZ�_h�*�J�j���Yu�]��y��ҝ3101�&\i��ȣ3KD��y�Ξ�7���!!%��r��d	3G���y"�U"��_��)�b��y"`W���5��&&�+�'Z�y"a�&.�� 7#H��H�����y"`^6f{X� �FQ}�>���D��y����D��C��e�D,��#ߠ�yR�F�HHP��0��q�Z�y2��P:���k 5+���5l�>�y��:������jx��̰�yҪ@�~��ā�+W-�B�%؇�y���=x"2�cdHL� ���Q	��y��L6]�X�[�C���������y�#GpGf�Sr*�)k��Ţ���y���A��Y�`�ǅ��`�l��y�7VX��1Kԫ0Ez���y�Om��ऎG����gL��yRLхqP `��׸e�����I�y���w�b��S@�
m�,u�ƠK��yBAvDR`���X'5=��Ҕ
���y�F�0C��Je��0�nI�Ӂ	��yB��Ќ8��#/o������y�JD�b�Y``��7��Xx�&܈�y
� 慊"�)=��,ʴF�:UH�}p1"Or,17L"+[(��%B�U^�j�"O<I� H�4дe{񮘘(�^0�"O��!��R$u| `8�M��'��`�t"O��S'�<���k�����  �"Or�bD�>�(�𑭑Z'��X�"O����L1]f���,�1C� �"OXa1�HWSu��T	ըC���x1"OЩ�Fd$\�́E(@&	�
`R�"O��KQ�4*Q�W�,dF����"O¹�����f¹�p"�
�`(Q"O%�'��3��Yx�Fƻ6��i��"O���Od3u�Ě����"Od�AE��"c��[�Y2D
�0�yB�E�IL��(�^�x����yҨ�' ��Li�N�S��D�R��ybJUtA�P"V`ӄ?�P�4闗�y��?Z��I��BӠ>m��	4'?�yrK��0���
��ڸJd B����y2.B3k&����ӿ3�t�cVn���y��C2/<<�u-�to�����y2��0R̬���D�[��H�ʉ��yRb�=v�*�L�`E`D��yҩ��z*���y(���0LU��y�KL-kTѶ� j�|�w��y2�ּ]�( `�`U9hϠ$����	�y2��bT�9��Щc�>Q�R���PyBG0a!:���ån��$i"�Kh�<��xh��N�el`�5`a�<��V���q�O�� D���_�<�W���?�Ѐၟ�x�^1�C[B�<��@ɭH�Pq���Y��] 6͋@�<�3�T�W'��7M �+\Ɣ�']H�<�t���l���/���SfC�<�chԛW&\���4ªE�T�Ae�<��Y�R��� H�"��)����v�<YP�0^t�c���L��y���H�<��ٖ'��0U$�.r�t�Wa�O�<�@�
�iQx�2Q�F#�P�@��s�<�������դ�>VY`�ǔl�<�/$U,f	�C`�:&�d�YmPg�<!e��x��4"�mU�e�"$1��Be�<���#��q+ `���Q]�<9­
,w�L�pć���	1� N�<����T�D�U*^#p$\����t�<��^��Ĺ�Qu�B��aECl�<!wȗ�M�v��ʿA��)ȳ���<�e��llr�MD;}eR�C��{�<I7��yft � �0�l,�E/�x�<R��2PQT�)V
��9�N�_�<I�LU5VI�A�5�D� ��[�<),]�*&���l,L���$�X�<�v$S�>�q�oԃZ��c���Q�<y�ș��2N�(yJ�ʄ�QN�<!�K	�zA��M9�:��0�FM�<AbaY�/�¹�� �4rҰ-��S�<Q�Ã�sM��#��^�&˼}2�^L�<��e�7ST ��NB}r�h2�m�s�<ك&j#bxp`�_)W'^}�Ä��y�
pШ�Z�b�9GHX8pC-�/�y�e��{@x ���]<D���`�@2�yR�M�S{�1��&Ұ��|ꠏ�4�yR�����+t����&�i�K��y"���ET�+uK�Q{v<s3�A��y
� <cP��]Y�H�8KkXP�"O�	��˛�\"$�1�.�tT�9y�"O�Ɂ��8R�6u����>.����"O��A7�D-i���G��9�"ODp�t��Q�,��˅�(�Nu�"O����=ir�Vd�I� �"Ov����ʃ4D�vLzj$�2"O@��$CFB��ѣU�wY<,Z1"OF]K)�1�챧d�Lb���"O|lxT�[O�0���?E=6H�"O.�H�g}���E��b)> ��"O0�x7� ���٠m��~F�e��"O$�g�X�>]du(�
�>->d!�a"O�u�EhR9z�fY� ���A��Zq"O�0���ax*��%h50��S0"O��U�ҝ_[^����V�W�(T1*O� �Ñ,�r�ӊؠj�<  �'5��H5�Ȩ�:���q)�LH
�'�>|Y�	C�b����E�f!��h	�'.9�Iׅv\Z��g��0[��<)�'�.e!�< �QP�GG�'���{�'6� 4�N9����a����H��'�:�E�L�4i��ǈ(	�0�'x���.�kTM���Z�q[�'z�8rF�8-1�f�8��q�'�,qba�M���I�fɫ�4}��'
d��w-�G��y�	�~��d�	�'��9�s�Z�O�jXㅉ�� �	�'"\i���H�T�hT����sF>%��'_�� ׄ�O�dt�Ǫ	7�d؂�'80���I*R�R:"o�(ij��	�' �%�·@�� ���i��t`�'������G���bL��V]ڑ��'��Sq&�8m��Y"H�6e�ؼ��'���s�X�z��)�0�b�+
�'��\��-^�ΰ����/C	�';�y��\+L�`�	3�ʲ �6R�'Ơ����6�@�
ŉ<*t���'��y��(��o��uK%J@x�f�c	�'ކ��OT?y;��
���sN��'#�̒ׄ��T����eF��
�'q�Փ��^���	f$_���(
�'�P�j���;���`�ĴM���:�'P�<��N�y��9��
F����'z�@�����K�*}[�=^P��'�f})�$�~���[02���'˪�)���k�&H*CIǰr�"��
�'�nY
�,�o&�b�K�cY�
�'}D�!2 �>O�A"#ȸb��\��'���}�alO8J�`�:�'�x,طoٚ44�D1�*;�Fp����-!6ɂ
TY  �*_���i�'��"��B<{;��#aUX԰��'VT(��� ���iBi2D�.\��'W�+�CN[-8`I�g�:j��Ԃ�'{���1�'w����٩I����'<r���lݜE5��Z�Ƅ!�P��'�TKTȜ�]����gd߀R��m�'���J���? 0�p��懨KI����'�x 2ą�7/>�8�g��G	����'QfyV���8���ȏ:�*�'T��B`�*�𡙀�ظO���'�H�`Ȥ|(a�eɩ�E��'��y�A��`n�p�,϶�\�	��� R����,#���Q��=4�Ȉ@�"Oj,``g��!2�H2dLEC����"O�q��ҙ�nA)kZ��"O�Yc�_�(�!@*�{��h�w"O�hz���V�r��Y��!�λT�!�.'*�����W7j�ī@�	��!�D/<P�PLT�uM�5��9*[!�@(hJ8�c�i��S�4�Qu+�Y[!�$�hG\���0ؘt
�i>O!�d�OVt�f&�"S[DiY��ԐI(!�}а#��۸aG�=z	��2!�$-*�������-Aג�!5nտZ!�с��m+�H��@� \@��x�!��B0�ѹ�`� ?A�!R2��Dq!�䑈<��ذ��4Yڀ�Q@T�!�D�=V�bD��)�����pR!�$�m�4x�	D�S,�uM!��!����$�.k���[AE�(!�$�7v�����U�<چC�}^!��0�<hHܰ^�iԨ�G=dB�	�J0�
w������ h��"O�����V=/K������Z�Ĩ��"O֐�%�Dܜ��)�0݈A��"O�X������!� %�d��"OPI�W�Ģ	~2��)h5��"O���qJ^�DT*��J`�����"O�U���_	x*�1`ʯ��if"O��1���R��<���F��<���"O`��3L�&�:e��C�9� ]�%"O�𻵯֑k�v,6)����"O<Ÿe��W�*m�cG�A�,�)�"O�=���ϴHyx���Œ�f���Ӄ"O�HAEF==�"�j�M]�K��=�D"OD}a��C�Kxv���Ʒ" �"O������w�l�1k�$6Z�Jg"O<p��a��f�y ��&e4Ԅf"OEڇ!�"�����,d�S"O)	vHR�P&^Ic���mBLK�"O���-���܍���N0eMĬb"OTd�AC�7`g�u��ǩI:��;�"O�����\�4{�!���8����"O����5y�V�X� �J
ƕ(�"Ot���N`6�Xr��L�P�7"O����"3�݈�(Ɗy�V���"O��p#�NGT!�	W�[��@�$"O��PÏ�Y���Q�
n�@3"O����e^�O��X3��Di����"O��2R�Q�����S?>.x�"OX�R�JX5B��];s��}}ȼc�"O�H����jՂ�b�'
`H�b"Otd����o��zYaj:��ީ�y"�3`@֑3EC�j��pfM��y�A����b¢]�e�P���c���y�"�HǒJ��Ǧ`�ly�GT��y2L�#�"�j�͇�N��}Q�j��y&K�g�V�17��=�`|B���y�+�	��C�ɡ������y�d��:]�%5��6>�z����y���m��Ųc� 
�jԺc����y��L�H)rA�{C��%�L��y��l���ąk l0B� S��y�銾l*�q����^ê���%���y��§Z�Z�����UK�$�ąD��y��G1o$<� s���R����H��y
� �ڲ�
��h��ʊ�e|��"O��@���F�td�cJ�+PJIq�"OL��u�ݜaI��%C �!���.�S��8	K,�B�E
 Pf�{��Ŵ_!�D�)9��Y��)�����ʅG\!�d�0���� \�g0`<;`�W{!�dD�R�VM�WO,.~4�c�Z�a�!�D].�ҍ�U��$a:Ib���]�!�D�>Sps�G%KP 5J��q�!�D��!K&�� m5�$pd�L�nW�'�IX>��pL�0L���a���Ra��'>D���$�D�0+ʑZ�M_:[���P��:D��p�,�#r K^��v�Y�M;D���R-;7���26��W��K��7D���D�ʿf��p+�E�-��s�a D�(;!�۶��d��(_�aW"D�X2�A��]���3�ֺ%���#
�OX��D{�O��A$ႦO����mʄpu<���'���1�4T��s��i��߲�yB��$�p�2�˛(`��d�㮄�y�/̆$�~x��oD�[��-�C��y"��Y��e�u���J�HM�,���y����:�����!��S��I�+��y�ML<c�T)�K�5Q��	�bK7�y�
.!|�ȊЧ��S�c����y�%��n7��z��R�A�8x���M��yB��vS��ҧ��Gs\i�D�H6�y�O�"1�0���;9f�"�y��"���CK�h1�)%#̀�yb�x�ƭ��i f (Ӥœ7�y�DC	��٢G�ڥU���p� @9�y2��88��LcuC�*J�ZH2Wg��y�('v�ٙ"M�Y. ���2�yr��&x�h���o�K�J9IC@K�y�8*��!r�M"A��IWK0�y��D	��4����?w���Fe�#�y2	E�&`V��eH5/L�=�c���y/��*:��YNQ�Q,�L�aɛ�y2aYU�SHǟN�J����y"%�a㦽�`�O.2X�Y�B�'�yE޾{s~�SV�^�8�B�Qⅆ�y�nJ,�6�I`���-����K���yr�8C1juP2%]$˲ ���#�yR �">������AC��yb���V`�Q ��A�2�e0w㓮�y��� O���sd�d8Hv/�y���4B!8tI5�ɒ"m�E��
�y�A� p7��Y�ûh�LI�2h[��yb����^�QF��]^<#ŧޢ�y' "��頦�[�N|<�R�bݽ�y"�ҏ_�`�1�+��2ub��G��y	T�e��k�!ѝØ�������y¾X�@�r���K�l̈́�y�Ȅ�?�^����*
�,c�\��yB)�05LFɘ#�0���[��yB�ϐwJ.��'���"�:�iR�ɱ�y2$^	�4�)���r `�`6�y��Hx�<��L�k�64�R�P�yR)߹b��E��Y�n�v4�"�+�yR!ǾZbx����f��,��ʂ��y�KI�Rаy�p���_��e�n���yZ�U!1�2
�1��С~��d�
�'�:���l�8V���:v`�o��ѣ�'[�a��Q�T�8afN��Y�.���� $8�"�
@���yA�͊o���0F"O8�z���?CW>�@KG�2F���"O�٠2,�7
.�p��G�
�� "O�QƭT�%�`����A>�:h��"O�	ҧ[�M� �!��5�����"OM�E����F]�E�zMS`"O�����^1|
f��@eɣB۾a8�"OX�H��6�
�cעB�Ĩ#�"O���b�.�R��"��5\�nP�s"O.�P�F�+�0� ���<��H#6"O�2��GG��)3�Z�M�:tjQ"O|9�w��� (<�����
�1�"OI	Gȃ�\�Ĳ�/Z<X��M��"ODq�W�G�4��e�����"O�u&B� '����$�1��H�w"O��!0.Ef�p� �W��&"O�ܙ�Y;�6�j�K[�1�4��"O�ԫ�f�?��i��+E$@��e�p"O��[G��$7������d����"O�0�'۽r�`@{���%B6��a"O���09 \��H^�/;�D"O^�1!ݼn^@��'2���"O��ʐ��(*�����'x�6�*�"OL-�C��Ҟ�Z'�Ҥ5�(�1�"O���#�6rH�řcZ�dߎ|J"O���Ʀr+~ؓPB +����!"O<���U�T�=��FЌ0���b"O�衔+�/�rP�m��B�"O�웵aÈ�JUQ�1��p"O�i�%��R�1s#� H�|�"O��a��YnP���� &�:��"OF�z��WǪ�$m�Z<���� Pj�<QƋ9����Yr�T��P i�<I�aI+lF�p�#�ۧux���^�<�#@��W�Ll�7��!�$A�c�<�s�܎�VLԘa�T!�@'�v�<�0�&Z�( @��<7C�Y� Kz�<q���y���Ek
�q����Or�<Yrd˛.�p�#Ř%A
��j�f�<ar��$u�^�[��
��8�Pb�<ɑ/��p	��y �
�7��P�a*T������n �\
�=�(���.D�p��eO?����	�n��ؓ�1D�0`�a��P�Nɉ�*�f�|��!D��`pj۵1��݃�Ș#l����$D��Ȣ"W�<�R(���$d,2�C"D��je����I�	�%if.���C4D�t�씕~����ĀD�~�H�
�3D��zѥƏ=4��3�Ƹa�|-PB6D����ۼ|y��Ə[�`���3D�D2ƫ�o�	��kE�LuRү3D�\ᥭ�;�x��e���P�4��>D�ĸӅ�)3��7��[����J(D���t*��མ���6�<=)Ê#D�4��I��x�
}�h֟H��	C�O<D�xѲ_&=�H���T5x%���-D�채H��^�MR"SW��J E,D����T�V"���p.�$j���(D����!���ab�1~f��c�(D�`�rC)1B&�֡W��BYk�I)D� ��G�\^�ɣ��(}qH�!��%D�,�è6#�1��S�OK��Vi"D��Au�K�n�M2/�;'ܙ�C�O8�=E���%+��b&�@+;4�:�Ҡ6V!�� �I�#�29�Y��&�&,,X�"O:����M��t��7���d�'"O%r�枘Y A��W&~����"O�}j�M�Q�x���H��W�>�#�"O��3�L�s��ʡ���{:X�w"O ��B	�,%q	�f�.[%��1�Z�D%���Iv��<�ŀx�����O��{LB������y���u$-c�c�r�~t@dh�$�y"�>J�6]CG�֕WN��1�×�y���N�!p#B��y� i���y� ]�P\��JCDxL44������y��T�4FXi�Sj9s����P����y"��%��K�FØai܁��N�y"��79���*�(��t8� ���y��"\H�X����Q���pX��yr�X�uq̨���YPH��� ��y�Ǉf��a��EM�J*d���&���y� 7�niI҄ȧU�b=1P�O8�yҀY�v�L�� ^�I��:B���yB�و�& �6f�_�4�����y�J�o�!s`�;`����yR	�6�� ��R�- Ì�G�<q�NR�AI��W�U"j���cZ�<ɰj�Z�"`k�O�T��
�U�<	� �B�0�T�Z�_TTPr��@}�<�$Œ9��]�w��3���b�D�<�Q�Ɏ+y ղW�<N�	'O��<)�.�bjӠ�..Pp��Q�
�<����.�x�! W4}���TR�<A'�ʦ2{�AZ�,��xe��P�<q�$ůG�xxG���+��HV�L�<6��8H��C��C6I~�[�HF�<�"oз94!�p�K
zp�T ��m�<���+D:,J6�U
+89�!SN�<�FϨb+����*I����	��F�<9㇅�F�Pk���!kX�0vmJW�<�Q������LN8�RX�+ R�<A�ޜ7�|\S����T$�T�i�<��+׹D�0��ɂ�i6�=��ɟ\�<q��kWuY.�\��d����]�<�dk'U��I���݁]�4D��ǈZ�<����I�0*R��;9X�ӗjLW�<�ũ�'
�ʔ"5�O51�.�cKT�<���ע~���*�
c�b�(�Fu�<��d\:Ͳ1���XP�-p�<��ݼ{��pX���$h��D���k�<qĬݙz=S*!o:��GhEQ�<��֮5�^EK1k� EY�S`�g�<i�$Q%#'���Wc��g8��mf�<aeg�<`=J�.�d���WN�d�<�d��8ꝳ1g��F�:G�v�<�#�!/�)�6`ߐo:D��r�Tk�<��,r
m;�]`�X���}�<�SŇ'�* 
p�܋yd����B�{�<dF�y�\���F
hJ���v��B�<ytL[�1�� �P_���q6č|�<��F½=InȰG*<,K)y��u�<��o֘A�:�с�߸3h���7#�p�<Y�C]�*XrBk<b�:= ���m�<a"(^�,���f��`�$�cg��N�<�� ]��T�Z�Ə t8����H�<q�FJ�p Hɂ0#Ѣ
bD��$#CA�<Y ̎&(#�(��
!��\��JBS�<�$�O�+ ����F�d�1���X�<� x�����%�"�� e��q@RD0"O�T��A�(4�T��D�t%��A"O��1��ۊ;v|y�㖟��*F"O���ХL�6@� ��U�x�7"O4 0��0# }#���jd�<	�"O���,M �����&H�HA�}(�"O��ը�G��� ˗�R]�<z"O����<S�����j\�wH
���"O��f�<�إK��ӜE�
��"Ovl8��UQ7D}ؤ)C��X�b"O�P@ȱ"܎�RP�ĝ!Z h��"O�� D�s&��#0kܺH0~���"ObQ� nC�@ǔ��Q�1)ʨ{�"O�G�( �%���x
���"O�Az��^ǸH��NN+Rg6]��"O��B	��J�\b5�ɷn��(��"Oj���2PU��
cLɉx���y�"O�#*�	z5@����j���"O`�P���& �C� +tf�{�"O48��B6����e)��"[v�p!"O��TKY�'��04�n9��"OJ0�N�;1�j�$*?R�0ܱ@"O��{WG��F�����#p�΍1r"Ol�FƒY�F��,����qD"OȭkE�+E���tMU�3��p"O�APnj���`n�{�TF"O��4^���-"|� J�"O@E�4'�,�E��FP%v�d"c"OZ�2F�^(�ЊVE�Nu<)
�"OH�9Ce�'%Ǧ���d]�a4���"O�q����>p̅B��D5>f��b�"O���Ǫګ"�8ѻw�ˀT�@1�"ObM�̰d4���k�!d5|`��"O�)5@��sHnJ�K�)����"O0��2�i$�D��IȘH�"O<I��N�"� E◪����y9"Orh�bmO	�����G'�p�"O���A�. 5$e��H	�-��� "O�=�I�S�j�aq���4��"O���w+_��(��V��f��Z "O�0�
ا2b��I!͇�|0`P"O0\iRh�׬�bt�! �b���"O�h3��T#��3`]3�����"O��9����'�t�9u˨FvL���"O|�@��?o�r԰���01v�x��"O["�:���� .�5�A`"O�)�D\�*�u��Ο���Ib"O��c璦|�Ij�(W�h���f"OX�S�ez�#0�]� P�"OX}qE��&;J��!D�
 �P"O�tc���]AF���Ɔ�:��!1"O�V(��>���X��=9��m1�"O�`��A���Xe �5 �X<Q&"O�����?+!�e�����A"O�UXa��0RL̐�3`ǯ0� "O�L�5�8�]c5��!7��:�"O=�dg_�C���R7S8��*`"O>�j��/�J�R��@$�d��"O��rWf�z �������	�$�t"O�hR�e��'�L�37k�p�@�"ONA��՛q��yrPʞ���}{�"O8Y1%e�z=a�i�zYҕ�!"O�e���-�l�p	�Vf�j"Ox��%�F/V)Q�I��S�l���"O� ���g��6q��I�	��.��]�W"O~ ��J?NH�#*ŠV��@�"O��CՎ�h(p �T�V�@�x`&"ODeM{�4a0Ѥ�e��"OF}�R.��H�!�ĲX���a"O�=#R�<x��Z�A@$m2h!�#"O`�p��?Km`u��	�N�z�B1"O��S��D1|� �;Q����$"Op���	s�f�-u����"O:��e <��	A1���A��:�"Ob|��퀲wJ�d�F��?]$�@�"O�u����c �X�'��S �8�"O0���Z6Hx�HC���j$<�J�"O���EHB�G�H��fK�
P���"O�(�I���y�$���Px�"O��S��EߒV-H�1)���'@��y�Ch����Ž���3oD��y�� �
GƐ�r��-`@�-N�y"HN5yc0�0Ǆ�-<dB ݶ�y�[cw^,۶��8�:YV�B.�yB�L> �Ա���ϖ _�Dx��$�y2'L�
�R`"Abر.H���j�y2���R}94ʄ�,�D$�ye�'�-:��� ��dDK��y¤�WB�=��h)��l��-��y���T��)*%C��5�2d	�yrE��@ؠƇ�:uuʀ���9�y�F\��!3h�nP~%��F �yrf��i6�!��mj0���A��yB�֬X�tL��G�f�� K��1�yR�^�@L�$�ď1��p0�e���yb��?	" �$.B���m���(�y2���|��Ąv�������yBj�"َ�
�k�+pnfe�*٣�yba��VLR�@a�ɀVk�y��۷sC� �L�%>d�|�E�U�y�!G^`��L�+�
a��yrl�8Q�fIs� \�u���y�T�t� p�S��T�%�K��y"�;B����ׅȺ.+J��m���yҦ�����S���!#&dȠ�ݓ�y��ŏ;�L��эOI��K��Ҭ�y�Ñ3.�]*sB�q�i�Ԯ.�y�O�l' ����o	�%A�>���F� <pq�9����҅�
�����N'>��BHՀZ��ey���;�����FEp�	C+bO������%<ʞ��,I�0!��M�om>�Zi�/F܇�A-��Ç x��(��K��+�TՇȓB��}�Fm_<�R��-�����c�� ��פ ���rJ̧9�Ԅ�?Q�<�e6�V H�R  ��ȓ7%ȃ��)@Jj��n��o�RL��-�Pꂭ�.INB�C�A[:3S�܇ȓRVf� �۱g� ���5�j=�ȓ>���(\�~��� iřQ ഄ�D��F
]$cD��cw*��"���ȓvE|�k��-<�D+#���5�x��c� ��@΀�'��Jbi�^�����V$���݈X�X I��	(s �\��k�ɺq�3dR���W�k�Ԡ�ȓ�nM��P�t�����Θ}P.��ȓ�f�AgG�t�M���9Mmh�ȓb_�<P㤀�;� ��B�?����S�? �p�O��4~��%.'����"O��r���%��� �E�X�	�0"O�X�C�T3ظ���+��,��ن"Ot���1>u��Ȅjֽ$�����"O�P�����b�&|Ч��4��"O�"3�@{�����N���J�"O$�i��QpJ��r�[�z�b�"OJ�B1���
��2+�!�0Es�"OP۷&Z�K�I��(	�2�����"O����L�d�๛��ۨ�
��"ODPH�lP�H�F�3ŀC\�Y��"Ov%ر(��~� �kuFN�>Yd
0"O��3WJͧ8�<98䄁�dW�*�"O���ei��@��|H�ɄIA�DE"O��*��[8�0!��O[�c�\DI�"O�IJS��;��9A�N�?�T��"O���siٛz:�(cN�6 �dj$"OX�Q��+`+p���,83>�E�f"O���3��]�J%[��:|8.� "O�Y���*��l�SJN)m3�8R"Oyq#��'q����1����"OH2`�$� T�w�7# ���"O�|9�G08�n	�wʄ�>!�E�0"O�� ���I�^�C��]� Q "O��̸(�g���T��
�"OH���&u��x���k����w"O�����K�*5�DǙ�e��#"O"!��֐Z�jEb''�#lN�Q��"O�u�!烤E�BD��U?@6x�"O�;� 
8è8ے/��!�T�"O*tc�Q�Al�b$�_O3�x��"O���E�e��r!τ5dX��"O�s�#M�!޲��[31�P��"O�<e\�:W�˥+Ըu��a� "Od��@&�h��o#"s�1��"O�l�6˜� ��:��91T"���"O���"I����huGΨ]d5+B"OHy�œ^��ܪ��qQ�4�"O��bB������E�m>Ya"O楱Uj�� b�	�&B� � �"Oj�9$+A/�IR#��p@P"O.�z+G��(�+d��52�d�"O�P���,pDp����["�,��"OF������m���,�j��"O�E0��C,+�LaA�.�\��P3�"O~j�oQ�Z��`Iw��"b=v�2�"O���S�_6o�B���R/	;b��"O6`���G`=0�C)�|��"O�����)
��CNQN�'"O��� M�, KB�&gX n	�mF"O��$!�"6S�ʂƍ�!��C"ORYJ��[<?�`8��*G�d�^�b�"O\Ex&D̷���3f
ҬK|d��"Oލ��'�62[�4�%��:I�)`C"O���0�:-!hqaH�6WA`�C�"Ob��*�6.� �w�ΐ 6���@"O��E[!0�LICcT<.X���"O@�  ��-����qha2 "O�4J�f�V���цgѣH�%�"OJ ѷ�m*�Vщ�m�W� t�ȓ������Gn٠g^
k|XX��.|�� a#��A ʅAf4���KB����ح\`�#���$�PP��'%��Tg۹?��-�$$I�jǮ��S�? $89�`�</e��0��NP���"O��UJԕ.��D3��=U�x��"O����[9#�
A���MC��3"O�X��ƅ!Ar�5"����b"O|t؂h�T��D;�M1��E06"O��CC�_�Db�+�`��o�h��!"O6ԃh]�:y�!� �Z�-Nz4�6"O�\�f�BԘ��E�P<Nؑ "O�=`f�X�U]V@�a��$;.���"OaC4�/�؃�EP!E��h 1"OH���F�f�q��"Y�f���"O�w�@�
b0��g��-s<8$�E"O��0c��L)�m���1�;""O�IB�ᛖ30��{�@�P+n�"O�IA���'��8c��8Q�!*�"O��+ +<N�ɨԎP�P�F1��"O��� Ȁ?R��4�_�3�� �"O>���� a�p�Ȣ&Ւ̴��"O�Q�[0o���)WFR��T�A�"O8p�E�H�kȌ�a�C�)kJ�ݒ�"O&�;� Ӆd���0���$i �#�"O����m�> �"��M�����"O�D�VE:�<���e
B�h�"O��wOߔ75����τ	4k"O��kd�K�*�R��:�����"O�x2` ��JT�p� �|���"Oh`dd��t��5�WE��]�v"O�H����r�PPRbٟR��9["Or<�F��?���ؒ�_#�$�2"Ol@���N=oPLX�6ANYҝ� "OB�2�坲_�Q��ͅ�
m��y�Ϟ�.���+K.HXU��fA'�y�Z��:H{C�,u��@bA����y��TP����KK+R�0SD�y�΂�/Z�Ҳ����p���y�+������4.ȹ9�]��y�`2��Y��M�����DK-�yb��*o�V)säa����e͔�y�ܸE�8(�A��'pH��m_��yba
D�,h��\�x�d�Qe�"�yr��=��<�w�*l���h�'���y�jK�SH���F`=UQ��� P��yN-5T�E0��_�T��̲P���y�S�Z�Q�(�P�.�j���'`��`ˇ�5�X�
�˟ �d��'����CƊ��P9�3��(����'<���@��M�ڱ�B �t�~P{�'mژS�C� R+�`s��R*lI���'��|�D�X�g�q�D��]p���'a��!�Ɔ�Ap^�����-L�I�'>�� � .�q����nzBز�'� ��a&���W��:a�>AY�'X��3��^��1�f�ˊ*{�X��'ظŉ�`��1�\�8a��!�0)��'?�MX�ő�
�~��q�Ԗ^4�-P�'ޖ��0�ݍ	�hZp�����y�nƅ&�0���h�#�5���D�yMVԠգƌ�� �<D���*�y�.LA�c�� T�hGo@�yB'U.!�ds��K��Dm��,�y��s�tH��E��kZN�ۡi��y� ��u�cӃ�aVÖ��ybBΌ�|9HRm]�ub](�I��y"*۹l.4��'� �b���L�y
� p| �*�r3�RRO #
x(r"O��`�;\ި�]5g���!B"OF�3��Q��P�3p�S�`����"O�� j��RI�����.P;��v"OȄ��RB�2�br��6x�����"O� ���I�*�H���8J���1"O��jP��&(�m >3;;�"O��x�F�j� �Fe(l\w"O�(��-Dg�*�a!���l #"O�R�CO�Z�l=A��;=�
�1C"O�i��F�~�� ����<m�"O�q��O$��hxf��E{v1��"O́r�T�N� �Q�K�']�@��"O|�)�/q���V�T�NR �yf"O�+蜺.�J��� H02C6i�a"O�����J$f��m���c@0{�"Ot|x�o\����1��� @�ա�"Ot����5"D� R��,z��`H"O ���_B�B�D;nɞ�2�"OzTQ2��80�^"A�ߪ�`�"O~	ؗ&��l���.Υd��ʖ"O�|��n�4+��!gH%r��Aї"OR�����m)��B�%/�n]�A"O�B��	(d2XhR.Ͼ{vDTK�"OZ�{SN��Q���8���XW5��"OX��3��PX��푯"@Hy�"Ox����(���ڥM@�b��"OڴJ"G�Tk�AP�K��h��"O�8�g�Ԑ`ь��Y-B�h�I�,�y�'@�vטּA�n6b8 ��2���y��1&�i#	�4_d�-�D�ܢ�y�OR�:.D���S�V�xG��y��%~P��!aQ��m(�.���y��1�*�H5j_�HIرj�勃�y�i��=7���4�'Gc��FC���y���+�����n�X|p�O̲�y���*x�� �&�Nh5���Wn��yR/� �#�,�^<󆣋[�<�e��$N�v�Z�Ł
9#�1�`�r�<9��Pzҵ,!qZ��BЏLn�<��F� �:�!ąy�乒)S�?V!��6��ܛ�B�~�X`��PX!�D�?֠2���5�(�(@*JB!�O/["��B/̰U�"0@u0!��A!�P��4��n��遶%�2,!�T�q��ŊG*� E��.CC!��<Hh�	��� �d���d�+�Py�֦C��$)�
�R��Ы��yRFԀZ�Rls�	"U�><"Ѡ�,�ybw��Dp�휂K�F��0M �y2(ӛ+e��B`k9E$��HEM�;�yb�߃��Ű3�ݻp�֨���^��yBj30���*s��2cr�`#Q/�%�yR�Z�0xRA |[�H1�yB��4&3 �s���L���H�yb�()��� *B�v�("c�Ә�y��6P)�1���:КZ��Ŧ�yBmK�Nu�
vmP� �� �c߂�y��ts���#)�i!�����yR�E�Y��Q"�%?�j�+U��y�لy/���$7CJl�7� �y�@�n5@���`45��!&B��y���~H��+�H��� G�L��y�δ�<)��M�)K�n͋���4�y
� D��$Ԟ��<�cI�\^��3W"O4�`��*4E�a���<g$n��"O����֔Bx���fh�T	`9�d"O��B�K�z#6��Vb�Ν��"O^��3�?�`��W+��O�����"OP�jK��:�VKA�_g�1�"O�<�q�_i�Bq�Ȧ:bx�d"O��"��X@Q(C�64�8l��"O,Z�`�)-��ɳ'X��^Q g"O}�V&D�7�l�J��u�l��"Ofx��/�"6�X���/dn�@@2"O�!
䪎��TѲ3NV k`� �"Of%)�a��D8<I"=F$M��"Od���.+z�`�b�FҺk@����"On����f�6�[��aٴ�R�"Ob���_�~�ٚB�P�y�xy&"O<@�6��)(���jƄ^� C7"O8��q>y����ɅV�@!��"O���b�%*�"��ӎ%�\�"O�iW፱Vt��E�X7*��m�"O�Uⴂ��\���!�2��`"OԽ�CNJ�(�v]�+Sj*�0P"O�̻4�U�.X����MNv�b�"O�2�$��*�)�l��`1L�%"OfM+� ��+�\���L�u>6��r"O\yKR@��$U1���#�V�j�"O��a����!�Ə�.��)s"O��S�I�s�!ys��p�"��d"O����� y:L�pß�*�J	��"OV����W ��l�!�{�`u��"O2 ��N��8C�"+��xU"O����IU����F͠}��d�'"O�0P��^<cx�Y��g�1'*�9�"OfI9RAQ�&����U��Hi4"O�h@6fB3=��i�$H�g�!��"O���+�p�H�ĨW7+Uh���"O�H�$,آdV���GӔw_
�B�"O<�J`�
�V:�㒧��HE��@�"O�*��i��ͪs��V�dq�"O���PlQ��Y*r�P�M�|R�"Orh�/ѣ-������Ǌ@�,Z�"O�9� gN !� P��"X�g�T��w"O��(�h%�Qq�9|��`��"O���B
!��5�8��u�s"O���N 7�xʤ�G��x*f"O�(�ц�"���B�ǩ9p�My "O��;DL�EiX�u��9!D�uЃ"OD�8B�:@�@�恘=��pJ�"O�� ĭ(���с
Y>K���6"OF*�ɓ1g\+���7l۔�"OT�5��l�xT��:~����#"O�U2�%�:MQj՛壕�/�FȰ�"O�̘F��:�� �t��D���)A"O��)#nR <YB�#�܌+�"O���޿"hr��"%
��Hс"O\�	W%s<�T&b��$��"O��!1&_�%�
�a �^���x��"O�H��\ WMvD�	O!��M!a"O����}��k����DH��"On��͆8h�ܤ�B�}t��"O��aS���)f!K�
��w�UR"O� �d�.=�D|h��*h�L���"O��{�LJ�6�^�JBҰi��D�"O4tK��T�qED��Rᆵ{\d�P"O� L�QC����D*�"ίM�Ȕ� "O��ڱGG�S5��C��w�x��"OD�S�k�!s��41� ��"O�3�ĸ\F�e���wuTi	A"O|�GA�P�,��1���2}L�"O �qD��=�Cw��s��"O,����:H���r��J�Y�*]"O�i;`IU����2*͆/}�i�"O@H �k�=	�x0Ôh�,vd�l��"O�@�FT
a׎��g��7\���"O̒����^�HMZ'a81j�"O`A�c	�]�=��kIDB@�q�"O^�#T,ێb�p�P�+�' �(��"OX�r7��RĂ`k�=>�:t �"O�����)jP>�0I͈��@	�"O^`aKH3mp��(�� ��m�"O�z�ぅ�:�#��ecF�� "O�m�7�F�/��D��-�7c�(ç"O�m����p:T|S�BӴ!K��aA"Ox�:4�[�
 Ԡ�ִl9dћ3"O
�Z�L؝i&fȺ��O���!"O�|�'Pz>5Ђ��/�y3�"Or�A�=��@�GF�}�<��R"Oʁ��J,^�܈I�B*����s"O�[�&C�mHX��%F�8�"���"O�Tr��6��0�"$ ��8�C"O|�:d�ʖL?(p[�aΟY���8�"Ol�H�aҦeY���.���y0"Ob����)5��q:MD*>3>�I�"O6q�o ��X���^�<͑�"O��P��<��<���$�
@�"O\a[%�ͷ:0�]8���v:x�G"O�h�#���i[�hޱ6&�"O������PݱD�Y�R�Y�"O�mju�O���LW���y5���"O�Rc�M�q�0��r'E�
��"O�m���$K��)��ە��7"O�Ń ��WG������lh�"O�0a�J@<�<�	��=���`�"O��s�I�>i�l�$����Mʅ"O t{p%>t�r��� �U���RC"O�p���Ќ2GF82 �$�v	��"O�l����Z
@h�R��t�,�z�"O��#B��7�b��v��%����"O�M1`��'�mr�Bd�z��S"O4�Hp���x��t*�#T�B�(�"O�͑��?�@��c[)��y@7"OZ��F�ϕ,�� ��������"O(ɻ"�V1'\�<(�B�c���"O�]JD ��]z�*OF�h@)��"O4�a4'ڷO �uJ�@�t���"O���tJ =����'KP7��8`g"O� [� R�Z7 �0P+^�y���q�"O��kf�l@ek��Ә3'�\�u"O4�)�q��A���[���"O<�`A�"Z�����u�Z��&"O`-�4FֳoC�h�/�,}��YC�"Opj7���)zYh���&s�9��"Ot%�āݯ`�؍��/R*)���1�"O���>a�0jb�[/\���c�"O��"�hϭ���0�	�npƼ(�"O\�C"^�G��pQQ��n9K0"O �2EG�5TiR�i�dIH F"O�%@L�ݲGW�_/,I:�"O� l�94g
�?��u� �@�s���g"O`�&!];JC��� cˆF�*��b"O����N�c���!R�=_���U"Oޡ�4o�	<D�AЂ�P\���u"Oppф�ΐ5Bpo�N;�`�"O�,Zeb�.],��.Ś:���7"O���.ӊx��̨r.e0B��p�'�ў"~
��ۣ1�v�ж(
�j�ab��yR��!uyDIBb�V��u4��y"n!|p�s�!I�?������?a�' �
&b\h�r�Kߎ/nL���':�Y㳋��!�B4�)�,���'}�Js�G�1��0��
"}y.�q�'_�M����AYz!��)V)	�8��ʓ>L�ЙӁ����YDO�<@0�uEz��~ڂ$݆�^��cEJ�l�����i�<�A�s��Tk�
���!�e�<�l��n7F��ʁu��L��H�bH<!#C�Z(��)�JU�d��edT�Dx!��[RG����āj1`^
:g!�^�K�܉S���b@K�;�!�$A�5�,���ȋI��A`1�J#H�!��O�i�N�Q��^���T�I�I�!���.ke�@���([fA3AO;8�!��Z�`Ze*3F</U�̣*�!�$��� ��Y3\�A���u����F{��P����#)ҁ��葩0R4��"OT�2�A�=7̦�h�F��+P�!@�"O҅"����,4ԁ��K̑;A����"ON�:���#*�$�Д[���G"O~����q���(�ɀy��m*"O�TJ*�#@_ H3�+X-�$и&"Oxf�˒�$Q�� Ra�%�c�'[Q����A��0E�|,%����ET2!������2�֭YΔx��G� e!�dT�S�x�� o�=�&�8v.�)ua!�$m�T8�1�)8�̵ P�ϋBj���>�Ec [�pM�#��MdKD��S؞X�=A��'L��d�E��!k9�JJy�<��G�;1�E�"��r��`����r�<	u�������C�u���
��q�<��VM��G�����R�&p�<A4C۹o�L����W�@����Ɗ[n�<)^:D4�%�D�;)�mT��i�'��y ���ꘚLӊm?8m����y�ˍ�Z����[�`Ĝ�f.,�y�`R1JK��8d�JJ����%���yjW<n��c��H]\uۑ�ع�yb�� ��}臣�>=F��1fЅ�y��ćc�94`^=<\�Q�� ��hOT��	�2��lP�e�:��&�)��C㉋^�H)��H~Tru�7n�89����{�X��AɮX�J@H���y�^L�-D��ʳG֫c7<��Ї�mPt*ҭ0D�|8@H�]��c݅��@I�j0�O�Ox���C�pJ�z���.o(��Q"O ���N0]Nd�z$�L�}T�(��"O����$[J��g��!O.H�t�IM���fM@;O�`��H����V�"D��U�3a���ʑ)=3�}��)!D�����H�Jf����l#��r1�4�`؞D ��XR谚��̲OYD��2*3D��Jc��NPCqB߉d�n�h�(=D�Pa���9VCF�җ"��P��RDF:D�� >�����4h�Ή�[�&�:�"OD!���!��ѻ���[I~]��"O����Ǆ	"Kg��l�q!�"O�M�$�����St�}l���xb�%�S�j������"H��]�T�N�8f�]��	Z�	6hK��ϟ;T��1 I1|��'���-�	j�Q��q��	�"!�"JN*� ��}V��r�g-�30��r�i"O6��5�U1b����W
B&
�X	W]�X'�F��'7 e�e�,QmY9���9~��M:�'U�˔��>��"bł�� �'�&��q�/;��́��6��'`�S"K�7�u3�ٰm�^l��'>� ��"bn	�Q)�e��qi�''�h�刚&�Z�;�CR5Z�"���'���Z�g�:/X.�A��R�&�
�'R|U+��c>JP�(Z-R3�m	�'�b�1�'�D?�T��-��L8�pb���3��Y,��/[#��H���<��ȓ8�$�K�PM�\��Ͽq@�=������A�8�R�cw�K4m5��Qg �y�S"�谊W��^���k�#��y¥�-.^��WN[W�9�Cс�y�J���U)0��-^��kšǐ�y�ȏ0^�t;&VL�F��q��y2"+3g�9��,�F
�H�6CR��y��;��BaV�:���k�y2b��F)�A��0���V��yB*�P�j�q�jӽUl��[6#�?�yb��(�|�凃*"I�m���y��
c�XI���*j�4D"0�[,�y򀆾z����u�ɧ.]X!*��V�yB��P<�*"&�6&A�`�O�y�&ͪz&��Î�tkd���y"�Ѣ'��酏���R8�aE��y�"my.�!� �q.)!ա��ē�p>IwoS.yR�{�Ǌ�[N��2��p}�)ҧoP"`����n�z�)�.[-{����ȓ�δ�TM�"u�
Y1�j� �X ��D��Q���#QJ%����:�D��r^���J{+�x�э��ņȓ�ب���� �����1�x���o@�L@�.S:7E�c�F�՚p�ȓ,�4 	p��+�P!�G�-���>1E�)�D,S�THÃ�S�`T�pz����y"�N��1y��O�#�ڑ��MK2�y��iF�[P��Y�� 	�ذ?1�'D�U�kL'2���M=0:�E+�'kp<rR�ǰ}�nА�V�[U�	K��D���[���؛&PJx���&���; �!�D�l�.�yPe��B����w�٘=��I�<y�}R�x�O�y���X���V��ba�H@�OJ]���Y\@�q��@�Z�vL���O��~�u���3�8-2rH	�x��郒c�gX��[t�PL� ��	*�"ă�A�>,�V`�O΢=��!�f�,5�׺`|R"$��G�I�L�?�~b@?3	��%C��l��P['M�F�<�Gh _�:����R�AX�|�*�B�<���o��ĉ��J-!�� ��nRC�<���O=���"X(~I�i���B�<a 'Q�0��|��h@!F�raP�Gs�<���?m@�)H�dP=�}�@v�<�7���R��t�T�MK�u��Vu�<� �5�8�A��	v~Tz��z�<� vm��m��y��t��OH5���W"O�E��ߖ�:��( w ��"O^�����u���$-P�Vc�-�a"Oh����6
5�����<� �`6"O�=xg�}��щ�IC�
ÞX�"Ox���ϪZ��Q+���"�~@i�"O��xW���m���Q�^�.x��X�"O��	�n�\�*3Cn�A�"O�cc���O(0p���t{
H�0"O<��j��QY��+�^�4��"O���R%c�(X�H�"ŠMC�"O� �fi�%ў����J����"Ov��'O>O^�}*tb�/_9`U&"O��IU�D&~���Ӡ��NM(�"O�@�%�J$|���P	Z�B�L��!��@�L	��f��W���P��qh!�dͅT��=P��#�|���&E!�D�ܰlA� t��a�6� P!�X'v�|��7K��"�29:OM& p!��[�tZ@�X-A�u�7(��gS!�$�,XM�f�M'H�\s�M��<Q!�߳.OX�������~bl� ;!��M����%lC�_�^�A�ԤEX!�[����x*��YT䆖O�̉�ȓ5;�yE$�7�0�8M��&�e�ȓI��=+q/Jx��pO1J�B ��:�F�ˑ*K�Z|�V@աE��\�ȓ+�����%����V�S#2��<��ՁٹwBUss#��cH���" �RT�
�'SH���#v~���ȓ]��@�2,E-��%��dH�-"0�ȓ%_&�Q >��`C�#_()�ȓF�f�a c^a�nHʵ��;@RVy��|��9H��J6,�D��Q�\��ȓ8@�q͇�@7�L����M�d|��	�p= �yr�T�VM�I����O�
��3�V�$�RC�ɫ��Α ܔy`*�n@]��5D�����R:gf��A�T����j/D�����ӯ�"��qʬ����!D������F^���'�"�V�"+D����'=Тe�#)� O��4��m-D��(p�!@p��ABn��t�/D�a�� `]~�1�"C
2�tz�;D���f<s��y��+�P|��;D�t�t����w�Q�B]:��9D��["@L:^��Q�F�ұE��X��0D��0�뎧=8��*I��~��8ؖ�(D��Y���H
0F��81�d�B2D��"��?l"��F�� ���*K"D��k��RY�Z@sÚ���6D�ȡP�Cb�ΌJ�$۹O��@%,2D�a�GP�:�#4�V+B�>��C�3D��񥈍.a"�4U�S5*IX'�3D��!d�A�,=@��t�΢<�zU��G$D�(96�ر|���`gV�1X�KW�1D�T�Q�Վ?Ht�� �&jn:�"�a,D��D�M'f�d��D2y���d�8D�,c��4YG�P�$���, �s:D�@I�A9��4N������;D��`�,��0��@'%�kx��xQ*D�Pf��6�	�F��p���%D�,���Ǽ$)�i����3`$�J�ih�+C�/���|����p!�������*:f�4"O�aY�!
�0�X�v�[�c/���i�8H�PF
\��}��O?7� @@��BNl��N�$Q�͉s"Oj5�d�*8�6�QH �@.�Ȱ�OP��)L�ADZ�`�F8�p�#�w&`а�ѼPK`D���4�O�zb�Z�-�6�����B�X�K�jH��R��P���3dO�ԓ)&i�����$z]��������u�y��H�8�uf�a�S:}ȡ�	��'��i��~~NC�	�Bhp� ��iêD����.S-�Q��%9
�Ȇ�K�z@��2E0�g?a�D�2 ��X)�e^V錭A��`�<a�a�#@�� Q� F�7If�둯JT�0"dKO� xpC�<�|�3�2ز�H�b]ST48���+�|t��Ƀq	�(��)�45ר��㋘l%,�#F�gvjQ��J;:�KL7�����'\�zIT@��@\ ��c��[��Ov<"+�H�(�rB����(FAGb��KT:-���d
*,YX��^��yrfZ/T��L0w#ͺQ��-¤\�gc��
E*�t8̐cu���#KčJF&:ʧ�y��"q��t@���U�n41B¨�yB��|���Zi߲�>��P �5��`�ǯ/�����&d�'}���Fy���2v�\x!G�1uؤ;�ܔ��=�G�;��q�bBT�+��Q�Թ7�}ʷO����P�b��@\�� #�g8�0�����_d�9���"b����&�I�7��8�c��`2����ڲ=O� k3O�?�`+�3L��}��T$\�����0D�|���!fs,�Rf��#�\�H&�Ŗ]w�5�g��(j�C�/T
akVd�%�˼;��&-����P�����g�Dx���'�B�d*2�L�+F�h��ЁZV�� %���Z��ж&�T�^S���qexQ�ɘ:�ȬPRb��}��IrM��"=i�L�O`^8	�M
?^�4�֏�Q�衴ƕ�;XX�$�]�-�X7Ce[B�s%D%�5k	�c|����V�k�Z�$�D�iLd�:�珑\(b��k� I�D耆�֪gu�<��l�D)Ȕ酏jH`�λZ\ؠ؃/ҫk|Hʇ&���XY�ȓv�Zx�$$�- G2h� ��.Y�QK'L�NJ��B�$��(���u�޵u�^x���@<t�pb�Z�A�;f��	s�\^�ࠛ+F���ɝ 
��񄋲b��8�D�;��Q[s!	3(�^��DGK����JY70���*)EjxY���8���<Q䨓�r�(��-���L��VP�IZ��J������Z�c<�$��.'�Ij ���|�p�M�	���x��ԡ!=0�b��F��|5��IW.����ˉwÏ%�ٻ+٤E@E��=]&��Gd��U{���-��Q0��E"

pFҼm��tS�I��J�7/f�p�֜`�(�Z��E/��8��(x����^�C�"��w���ڂ�V����ԛ�ċe�¯9t�3�h�'9X�[2n>ۿ�qb���Fe*���!��Qa�����=	Bk{!�BA(��c`�A���M�U�S%�H�.�--F��p�ߖX�(�x���	�,䪲d 
��y��,��*��O���a��3sJ�����x �!�D�4G߂\�WcA�a�D	���^`;t��4z7� �$��fF!{V�( x.|�V�ƊGB��2���3eC��:�G�6hwj��d@5<�r� �;s��ɤ�H�'� @�Sh����g�K�X���;�l�j�Nр=x����A��#�t��h�gi��@$It����E,��aa�O�)f	̥8-NP��$D��X��
�g��x�sB�yHJ�� �����	P�)M&?"P`�WdE
�l�@�w�H���N�F�*٨2�!���Jg�'^���,�;O.N�ї$�9��I��B>�3� �OKJ��C��n����:U~š$DT�<��e��X�I$�K5P��hBf�yȊ�!�_��a,�`��X"�ّ}��<�J�[��)X�A�� i����ٺV�J ����S ���,+p��S�H�>�P�`#JԺ�F���-�q#P��a���`���M���E8l$a��L�z�Ш�DE�;�N���@�|,�4�w,@OFD��S��UjJ�S�B�4'4�9��O�j	��q��4�OZ��bI�$#f%� �Z����Ed�-�8qRB��
T��eJ[^EJ��ғ!(t1���TY����%4��)�a����ЅN���j��a�'?�,$C4A��HԀ,Hy�M�ϕF'�q�L�	Bf��Tg�V��d�b[5C��h� -J�mPE�Vy�ǴbΉ�6�O&o�ʽ����O�)Z�?��};�"��!D����)k�ʈ+".�,!wV�*��K����F��:!��R�'��g��d��j�'sh�J�g�$|��lh�/�����)��#w�ݑ��?���3b��=w�r�:s���\��Q㕨mNLA��e�G,-kXTذ�O���3�W�<�pά<`��/C��$ޮ1~�� � ;h9�Bd
�t����p\���yb�@@���@���4��k)D����hQ=_xm�U
q���v.���U�e� "F����/i��'_��8�'�_���(��4q�� ��xaz�Z�$c�^�5	"(H1�ɕѦ�!Ʀ�<��XZSAH��hQ��
`n,5كN�4ay�g�,\ |�����	3��D0������?E�D�� p���F��g$�y��O�j����\���0��
�l ���75��[���H�� �$_v���ɾ'����@˳��u��GO	57q�"��O���*��9� ��a�">��-�O�� ��U/� "���(q�șw&A5AX�X�$	"�	�����ӖT��g�'�=�Ѐ�<�px��F��=��h�	˓r{$�=��p���1<z��7�S�3�G�3�PQ�|��h1�OYR��b�8qhѫ_�=V���a�x��y����f��c�i�
]�����V>R�ټRn��U�ҵGр4� �9D�x��l-[���D̐�m�d�#�,�����/�!a��t�u#����+y����Bh�*��C�E�,�c�n���x����4�I��ٚ]�Z	(�
��"��X��s �*~n|�@�~�>���G5s>P�gM
 =܀�Jm�]X��0e�xrG;�:`���àP�ʹ#�� �H�\ѣ��6�<��InF:�*S�·_8�x�Z�CO�Ot�ь��I�)5��A��nw����Ƙu�!�	<Ⲭ!½mC� ��kR2dͱO����,a�� ���w�̓<-�lņē5<X��kן�Q�CC0�$m�U%4���M�
�b�2VI!<pС���>,O�ɢ��,��.��s��Ǳ	���c��yR�ĥ3K���Y�	md4��5��,ܢ<�~b�I3~f
I�C��t����g�<q��Ȓ&�:Q��CI<	uk X�Cߜ��D�xt���q�Q�j/<���>eg!��n�L���"��E8��60c�`��'�F�3��:%�p�9�h̛ �1ϓ%��OfLx7��Q#�aP���nz%R"OB��eH�=vH�{1P<~|Ya�|"M0�S�'$�RM��� z)Μ���.T�&��CP�rMO7&�:�Jt%E ��Ex��'r��1��Dbd�ԁ�:"�}�
�' �æ�ňkג
�M�G� T�'n��*5�w#<o~}K�f�1O���Ќ͏ ����5Ί�
3 q"O����X����0��&d.X�3��{`��OT�s�Z���0i/͡X@��'� y!!I�3O8Ҥ��.XF�+�/�4�C��al�)��<������0#�kͲ_�eRT�<�d���n���:��h��XU}�Ė1e�l� �fx��Ju���w����-��p7o2D�\����U�yA��X�
��ȓS�2D��	բV)[�T�gdه[.R�f�/D��I�&Ԃo�Ĩ���T�;W4P���L$kF%��=�L���	����PT��1EoR1*!:�p��X"6���P�_;�=lZ���U@C�M4\��[(6nC�I�J��"�T���pa��.�P�O�|ABO��-�\�$ ̿+ Q>I����(,�c���T*��)D�yS�_oJЀaϊ@jVP�cC4����F���6
wb��~&�[""W�~�4��q�z��K1�(	ѫ	!g˒�;�đ�c�
�Qz�2&;gF�YР�9$����ć"]x	�ǖ�K���)��EX�x2��X�:��s�ɞKMI�&��+1�<jVE��c'���C��
~䥳
�'�|E@P���"�k��C�.Y��N�< ��WQ��	eMج8�cd:��?9O.hj���Ww�HH��˻p*���䝮aT�A�y��1	�Xa`�N�.SC���b��j�d!�lT�3�z�d[�.�x Ɏ�L>���?��ĹQ�ǃ;�<�0f�x~Rp�eA�|���O��I5J[�È�"��ݻ��N0���E2b4��R"�?_��!	ϓ6K��qc��9���+�/��}��!B��>��ߴ"��{�O4�x���H�7�)�!2L�ŉDgT$v�|�(��G�)+&��� _�ɰ?q@�*O�$�zqb�V����iЈOG@Lb �ӫ ����m�������$�r�⋼T�������h�J�z��Q.=t�E*5�IXh�%z�
�(D��ODx�a#��70\��bEL
�<�*@��$V�0�L[SL,TƠ��c�Ö����X�"b��, d��Ն�R����'��,����}oD�O��6�	�ą�xP>�h�È.g�h�y㫞�wOL�ӷ��S1��"vh�6��y���,����ad��Y��T�5]��'��3��+ua���=@��@�;*�L�K�E-๤K��q�Čb�/�$T��i�"�'W.��K)K|�ch��"��TN�7F����`�<)�L⊍C��z�C�3� BH�F�"c�T�R�]
p��S3�'2��Ɗ+��'���Y�H��#��ZRc�1E8|�uHX�V������<	c�����ɅU3qI�~��dà��P�B�ɰ:�0]�C�1q��bW��!���Ӵ:@�P1S�(��=	A�9�Jĸp�P̺@���m��X��A��/�nt`�O�!�ׅ�&U��+3E��ڄ!�"O�g�H"�t�!��-=���	"Ot4��h�tX����#��"Oʅ�BbY�X8�mavg��.���2"O~���c=r����GsZ�p �"Ofq�۫?/��
��"@�x�d"O@�
gERjlTK�%X �<��"Ol<�`�1%S�x�!!�bs| ��'�fQ�� ŇCSNĀ���4Sʄ�'�r��ZU��y�G�?-#�3�'!��	���R�0I�q�a��I�'�!�4/[O�L��!ʖP�T	�'�ʕU�A�JP��2㖧!s<�I	�'�e��a��B�򐘄N�&>Fl��'h�!x�j>X`��D�0�@!
�'�rı�ǿe!);�$�=r̔H
�''� 7=��1�������'�rLd�7z���N�%?V�	�'K�uL�l�8�@}!V���'X�4������z�Ƞ+��n#*���'����o��J8��a�
)~Z	p�''���v�[��:��Gɢ,�����'�3�N�u+,A��蚫$�K�'�8�4h@�D U*DVo��Q
�'��m�cݞB�r�DD�r�t]��'U�Y��/�{b2!B1��auV���'�:t�tL ��g�ț��2�'����),!�`���O�73��� �'0�`@��0b�@�./΄"�'�TB"�F4_�Ī�`�$ ���	�'�. J���50M1j+"k�(��'_�V�8I�� ����U"^M��-D��F�!Op@��&[���J�?D��s�mI_��zEE�U��azB�?D��v�S'T�MP/�(���y6�=D��IqLZ0-fe%���V=�1�;D���fMP�`�dM��)�#-��r�4D���C �-�P�I��n��z�/D��s�
M3�"�q���&���-+D�Dp��1t����@��ح�
4D�d�qj�r�x����T� Ӑ��+0D�Hy@�K%�'�AV�1գ=D���#��f�V��� L�5^�@�*%D�<S&�N1Nf��!gV�u#|2v /D�d`�E��Z��v�S����4�8D��
'L��&���e��I��:D�P`giB����j�Ǎ�;.�T�/8D�4�$oA�LB�3����f+D�h�#��>C�>�A�iF�o���Z�(*D��AӋ�8X�R/=-�bѫl&D��5'��yJ�!�(��X��$D��{@E�D����A)ya(-`�.D�$x�^>��vhB��¤N��y�j��9��!�D�V�
�S�M�yj�`?�)�Â%y^��*U�Ü�y�]������82H��
��G5!��1����4	
;���W/p!�$W�(�$%��i	J�֠:�K١$�!�d�[��EQ�[�i&��G��!�� ,x2��L6�VJ¡�)6Q���"O���Ӆ�)U�8�y$��?�6!��	�'/�|�E
ա��OΎ@��٤e����f�Q	f����'hT�ˣ�.HP��d��Yz�cڴszRm#��	4��秈������i&F !�ߘO z\�Z��y"���8������݊;k�j���<�~���Z�iC��_���$��-�2$����FK
A��-��Ga|rhʅm��� �)Y��h�ĤDx�Ҁ`�N� 8��qkH��x���P�CMǄ����F��'����-?)�,X�g�><��>��#(O�$p���+M�,�"O��H��QT,�2��A�V���CJwX$�B���� |�!�	E??�>�	�bd5�ȥd�T��HL7gBB䉻2 �D-V��k���?9�� a�Z�R6i�~`5���G�?�>���"*��"��λ^�d���n���ۀ��%���c�^ ;�񚦅N�;����� �I00P��K�.kY�<��I261����#��tB�ᡪ-$�r�<���aa|�1/-���Õ3��I�5cr��aү �u��
9!�^�G?����U�Q�J�`���6*:�mBd�X�@�`UՌrOq��c�g�O8���2$�8�F�׏��dz�˸):!�K! F:<��S/����P��� �4: ���,a��J���U���OD2$����U�1�@{�/�=:�f��G�P'N��{���]A���+6��bB�$m�xS��2x3P���A�#��h�FO�
�p>���� f*�{6��z&pT����m��K2���eM��8h@'̉>'�ZĐ#O}��$M()7��n�`�i�eq�<a�$�� �ig�߅s�x� mdN�}�q��qi�a@��@��D�Q�d:�'�y��TϢ,���_C�t�fL���>�v��!�J���+��J�aj�d@�)X�
T�V����Ԁ��D(��[b��9����@Dy2�h!�2���]"�$�5ž�HO���O	6�H�e�T�H��Z�)w'��7v�v$�pM��orL�)���!}��A7H��Ӱ��'!��ӧΜv�$��&��<�x
R`��;{��Y���[jx�C@�$���#Gq���恷=����%p���O�k
���&�7}!���2G&n���f��e�Y`2䜬'l�8K��	Lbv	���"K����3F&j���Vf �EXB\�$h�Y *��zb�ڧ(R�R��.o�{"@U!(�н�b&�.y��1�, ���v�	���G#�T=!
����!�G]3}D` h��U Q�xQ�� ���2�˩t�Ȕ��G!�I33�,#�~�YP
�(F���r7���q
D)plG�{�L��Ӫ
]��(����7<�x�W*�:>�d����'5��A%���pP�.��"�n�˙P�6E� �F&G�t�@�	��s>��9��4�nlb�i&"U(�>�ʄ�jW=���V�֟�l�"O��8$"Y���	@�dB,3DF+���e(�o~�ɵ�@��Q+�X.=pa�@i��ļ[�|b,{K�,9��p����Γp�B�c 
?\��q"'W�T�S"CҺd�dЋW�t$�\:��T�#=:�3��>*D�ׂI�Q�Q�����	6]�
P�{H�{$� ���p�J0�7���=�P����#o�<�P��x��i��޴!(xc����zW�<qf�y{B�C&3"����L!Rt��Ɗ"�^�9	U%�� ��֢Ux�P
�$�N�(RN��]j=z% 	$�H�yr���%��.
<t�u�� M�u���E�Lp!�dJ�Ub��#��R������ 0U�$lfl �M*e|Pmx��U
)Ƈ�'�
�:v'���a��?G�mIp�<G��`���Oma|�' "<�Pd*�&�re䡕�XqlAۅb�4�*�ª�FHХ��6X#|�3cL��-�dIJT�4ғL��[�b�46��(1�Q�Qi��Gy��J;N��4Bֶ2��y��U`����O8�Jd(�NƑJC�,ɒ%ٗN�
1�&�h�� 0�;��յ��� sJT�]��o� tX������g@�r�K��`n�`)m�Z���v����T�`����>�v�җb��ϲ�qA"Ob]S�do�}kd�إnX�)��V46JX� �B��y�6a�2�f��9�',�6�ތ��wd�ԁ
�s��A׊�Q?�X�� h�l�CIȹ�4e
� ��jPi��ID`^���p�S�BX)�� Ԕ�Z�hV�ȸ�<�=���f��l�̌�'BvJ�FXP�'U���)32� �qH��bI$T��%��+7�;%˩G>��b6����CݰU�����l�|��HC%\�x7;g ў�`C�[��Z�Q�`��8���^?QZD�#"� ��>d� ����6D����N.)��HdĦ�X�Х�O���bOO�NXP���Y�
�����Πi8����v�Py�&ès�C�	m�J|��ɕ"j�������p,��lĶo�X9�V��g����G�|Fy���6��xa� �U3��8⃃��>)�CC� ��CmK�A�t��d#P!K/��\�40)piV�J2��� ����Q18.�穏#j��E�s�I,�NM*D��L�M�sh�#cS��V�V%��L
#'�����G
>_pB䉘>%�t����|� ��J=|��Ln*������-���� �������bg�	;2�T�� "��@�f��ah1D��C#D[�x)��!�.�x{���80E�ف��@�"���@5r"��g�'fH|����w	D��`gʢ*����	�*����ᦅ%o$\��B��Hʩb`�F�����)̖š�<�Oꍉ��Z�iݤ0Ё`�)C�ȩ���=0�~M3EM[�=�%�R�T%L>{���C�o������g+�&�yj>(O��1Ǣ������
�2�~ǎ���}dF�U����� *bް:UB�+^�:tr���8z-B�I�"������^�.�ä�%� �0R]���4 ��P#H|�>����
_�`��uo�"�N��e�Z�������WJx�D�J\T��p�����E�P��j@a�!�Z��E_^�y���y�ͩ2/�m2W,��J��3b憞�yB�y�2M��N�@��KWb �S !�D Y���K� !�$I�aQ�,!�]�'�$"�����.�
!2!�dE�T V��	�/�`�A��=/!�d��&����s�	:/�Z��!兏k!������Ge�/1���"��R�!���K���J 
X�UMl���L��!�ݵ��6v8��e�+R��l�d"Obx�烱k"�����!	���"O֬PB@(6`AI�"*+��<�2"O�"T˝@�"П.tҹ��"Ol����?i��� �5A�M�B"OH�V*ף2"Fq��C�W28(J"O���B1/sK�'�����Ş>�y��X%zj2�s��%�.t��O�y��'N�����D�r��D)���y2�ϋi<��uD۝i<l��
�y�/VxČ�yv�XOj� T�Ҋ�y����!N0�
1��R�����N�y�hX�	�$q�Lң}ͨ�8�.�2�yBc�*���j7��a���"�y����TU@����\_%�����y�e��J!oαrshղnG�CC�C�I)W+n��IɍA6���ŗS�^C䉹G�|�r�"߶Z��(Z����f�6C�IZ��Ib���J��
�kF��D�%=@��Ќ�4a�8Tإ�	&x�!�d��i3���b�)yR�W�ܒ�L.b��� %|O��C��;DD�`q�G%|�L�A�'b����#?q�ʰv���A����p�Р�G�"Y����C"O�qd��#�2�;d����ē��|B�%��ܣ�ʙBs 5��� ������ضy$��!KQ�Y�!�� T�q�E���m$�as�*B�e��xU�іZ���f�ilVU��l6�3��ԓik��XQ�C�t'$�ʤǆ�)^���	�7�"�:T
۬	#vq��E]�6�\3��*G���ҠBV�8Y؅r#�'j2�
V*_���%���9���	�|�H�k7��&W�ZL�O��r[�Ru�ݨ�H�xbAFN@`h<Q��@"��Ly���g� �BW�j�$�2A�2-0U�t�:C ��&��\i���VC���&O�8�LE0X�p<A��H�>��b��(ҡ�v6d<��k�:��Z�	�%� �#��
�*�+���>�O�y�uLL ��u�L 	h��c ��p��C�`%��>q��&��a#PJ�)h�*����9@}@EZaص�J�궍�hk����-c[�U�nζL�
d(��Y�ekDѦOr��B^13������H�D�A���av�U,`_���G�̰�V�ы&q�q �/;�O�y�uo�?9�ȳ�MF@�0��O��:g����J��?����m��Ѓ�>9�����O��\�j��Ԩ�Ytx����%N� �E¯�!UAp��ψs�.Wȵ	Q�#<ҍ� ��<3,��%�����]��ի�C3�3�d
�%l�y��L����Ǩ��I�s@.��r�!Y �S�8H�� �)�$e�3����`$f��T��A��NY@�ic��4f]J�h+<OD���K���J���;� \���_���1|]�@E�?�)!�����3��.J��K�R\$nD,��9���:8����	-vÇ�1m��)�Q�Vk���4��PÞ'w�Q�&.M���1n��#|
� �MEv�z�
�{h�C���A�d2�CTT��'��r����c��x`���x1�p�f�+$��@K4<'|�T���>i���+�$��C�	|��&��j�<�Sf�v,����(��H�"-%<f`!I���k$�E�"�'�x��&� CŚ� ��X�~���&?D9*�AF�0����::�9�̅s"]Cň��B�*A�Ҵ�U ���|�G E�|�C�	�D��Aæf,\LŐ��Ί*�C�	��&]Is�M*:;�y�J�>�
B�I6�����U�n㚅�"�J�u�C�	���f�dQ\����ޚs����f3J�x4��%X$e�% O�Q�ظ��9V\��Ua�Aѐq��Y�Dԕ��U<xI��Ȟ��p��L9�a�ȓ�ޔRe�'�|E)�h�)��u�ȓi��@��� ���n�, ���ȓ�)����8��Y8����:5V���d���d�.}�
u�&cQ�t���ȓk�
�2�GQ�w���aM�:�$��ȓd�
�@�2Lɾ��ӎ�h����ȓO�L�e��?��s���&#��T��������e �\��*M:t(�ȓ$O �1᎜)}߀�1cΙ91����ȓwsp��e^0h ���n�;����a��z��1p�Th��JM<$�����kQʽ@c��-|�[yD�q|
��ȓ�,�S�$���:��0��eD@k@�
=	~T���IM�1:}�ȓ`�@�Ԣ�a�d(pi�4i�������5�K�3?l�$�
 "�ȓ}�P�X��V�jm��23iTu䕆�&���:'#� �1�U�8*Ĭ��Fp���1��/�H��56�VA�ȓ�ĉs�FE�v1HI�6�˲�0Ԅ�~���k�.	6xHi�o�)	��ȓP���c����!���[�A�3o�H���Y�n�`�-ģVx4݉�i�7��Ʌ�>�$H�e_�8*x��h��{;�}�ȓZ�z؉�K�}{�MS�@? ������gFJ�j&#�%c����Cߓ"��tB1(�	O�"<1�	؂dJĀ�>'D���|�!L«#�e���AD����b�?�&�2��k�I�ʋa.4��O�:b?� �#K!
-.�I�JY��\���� 9�����t��ѡ���OY�	a�O�(�ڰ�ٛ�i��]��:x�ஂ*ʚ���IЦa��Q1���>m�'H��m�m�Ҙ��?���`�!��U��mӘ���O?ejvgA��0�KDCT�I��m����O�(S;D5F�OQ?�0�m�W�����tZ��\�<qa�>��<��d�#��Dr�	{CQ�_c�]0&.	�N1�'b��)��z���*��Z���d�.�؝&�$�'�ڙ�O<e��9\/哽%G@Ir�GՎ�a�5� >k�˓U:@6-[,q�]�OQ>鸁oM�N�Z$��BqB���,�O�p9ٴX�Fy2P.?����O���{1��P*21�t�"W�m3�i�Ou�3}r�S:��� �c6x�b��Z-j��eh� �OX����O�$Y 6F�fy(���QphP�h2}r�_)� �ذ 1��IF�r��e�(�+���I@+	<w��	�DVpu	��6�)�'%y�4J����c�@�怉�^|��4�=3oJD��?=G����-D 9ij��q[$X�c�_,�$Г&���|ʣeߒ	'�43��M� �8�� g�L��)�`���ē`�l�]�Oj��{��ӕ��Qm�a4���{"�����Y����@;����G5��W
���h�D�Td�S��O�e�p��c&FPFl�:g��E��e����8vbDa��S�T����π ���Oƹ-���X^�������0<���� ?�v'�R��~�N�=&]lI����
&�$�E�	�M��T�4�6�&?���MKAHEŞ>��	�`�#fv����P�z
i�i�P
t����P�*�����cҸ��V�T-!�D��>�*�*���6nJ�p��	)*!�$F1Q�zP��G�δ4��*�S!��Q�_T�j���䜊a��-K�!�d�/:�4x���I�p�	!����!��6ffuaR��(l#�bу^�?!���
�
��F� ftNi{"�=!��V���:��N2Q\�����!���@4��8CB�!� o�V!��aN������8R�+u�؍O@!�r�p-��LX�^ts��A^�!��1A��K�
Q�>5P��
G�!򤈢f/"4��f�{�L�� �	i�!���*�x�ŌF�k��`�/Q �!򤜘m�<L��lF8'� ��� !�$��]b��7CF4��aN�9�Py���& ��Z'���{�����%)�y"�ɪmzt�b�אs��$��*�y"�����!�V�Ϯ5Z���� ���y���3�y�1`�< �a�#�S�y""=Vf� �u�*�q�f��y�G�>y�9qh�jj��"����y��3�(`Y�n�iȒ	1Ƨ���yr����Ц"h��e�5�]��y"�Qf�,b�B��^��a���W��y2����1Q���3 �|�KO���y"�#_nR���N7,����%���y"���f7ά����vl����y2�F_�ڐi��"UP�a�y�lO�5=z��0��*| i+��O��y2��1l[�E���ޗu)���Uǌ��ybD�>\x��&��V�l9j���yb	əH�)�K֞��T)�����y"��
it	{Ǧ��K�Tz�\��yB�\JH]c&�؁(젶璌�y���!�]"�T5"r��&HK��y��L�|QiP�-	"<`�$��yR�8!�p:�OyPhPHT�J,�y� F	e|��cL*wC�p)g�H��y2C�6xTM0�f�wk�УLM��y�W1oYF	
��̚%�c�J:�y�h��+� 8p�m+��@ f���y�ݐD���
ߔ
s8�	����y�g�Fzmc�,�&{mT��a�ų�y�F̾H�T�#�eU T�Qǂ �y�!�� i<ā�Z f��� �Ð�y��T�_�q�Pk�R�\�)�(�yR�,0�zt�(�I�=
�����y�S�nɢ��@�+?fr�����y���;@�ȨZCf��?C ��l#!��`���0d"!�G��vP!򤀔���!��]� )D����w3!�d�a�������n�refP'0!�ӫ��@�Z�EU����8gC䉑1�\|�0D��nFd��㔿NB�	�^�D�rl͖~/ZX���H��B�	7w�ؙ��L[�A�,,i��M�w��B�I~"��6��;c��-[F�@�B�Iy(����Rk�z��sH�,5-jB䉽Z��!��M$F��R�PB�	�W�lr�	��]��d��T8/>B�)� ����i��i# �!����z�"O�I� R�\���bޡ/�J}l*D����j�H�Vi D��?�,l�#�*D�����ҿ"���;�A�&�4���`&D�(�qk�8���+��%�d!f%D��� lt�h`�C�[��0����+�!�B_r���� RCi���!��P��ѐ�D�Y�l1�b̔S�!�!R?�H �lڿ0(bWa�y�!��֮[$,0�"�OT'L�r�ފq�!�Θ7����q�xaC%/�+L&!�$��6hK�nB KE*Ѡ���[��ޙ

���t,˿�����,Z*�y��O�@֜pR����z����y�F	>���g�UQ~|�����y�I4B��I�rI�Q-�a��M2�y�p��q[�-ͅD�8����y���k�e�C�D�>3���	B��yB��Ҥi��eo��I��P��y���~�a����
��$[G����y�)2����o�*nbM��V�y©�K���!j_��p]��h��yb'2�XI���zFu ��yR�W�R�v��D(�ƐaX�y��ܗ|��p3Ј�/��x�!�
�yBaR!	e�an�m0I�%��0�y��
j��P��O�&wjlH�튠�y��ݼm�r�zu朤�\�a� ��y�
�Bhq�0���JR.1 �F���y����4
�R/؎D�8�CJI��yңʭ�e��(@*P��@8���yR�T?wђ��E"N�N����$��yr$ԕWsR��'d���"�+N�y�/� n��Avi�s�$��T��y������ɺ{�2��R-ӕ�y��Q2HJF"P�'���R�޺�y2��&}����%��Z�h���y��\�x+A�M�8�0�5�yb��j����ǃ4���˄�y��6t����n$�ξ�y�7`�d��:�.���'�y©S�/�h:AN�`J@�ZF	צ�yr��?����Q�><��-Y��y�,X=j ���,Hk���[�y^�.X�!뒽@,�d�f��y��(G'`t���.4��yRf���yB�$'td�ff�-{�Fm"&nG��y�H�l�@H��ʧnp�xf�_��yC��'ڦU��*ޗcO��95�©�y"��zMTtbr�G	a�4pd�B�y�M�:pd��O��N& q������y�錃h *��D@O�}�~ �	��yr�ڝ{gV�a��\�x��e����y/��5�ݳք2q�h�"s���y"�A	Le1gED�{%&)+EW��yR��.R�, 
��Y�t�<J/�q��'��p�恫E�pG�Da��	�'M�9���F2L$CUI��?L�3	�'�������!���^�;����'�1zD�˯�D�+%��85@�)�'A��a 䂈5��YJÐ*d�x��'>��h�oOv�aBF�V��]��'�*e��Ǟ9�`��aL�Q.x1r�'�LU�JҢ8i�ZA!
�I�P� ��� <}�P�ϐhc���[�"�Y9U"O�b'�I�]���@Ms�"OP)xV�H�A�"y���ïc!L�AT"O�A��#�*����X9'hq0"O�d iX�h�d��8�\�4"O��8¢Q�S��0�W@��-�>��"Ox�2�IR�)"nP˦eP/D��b�"O�MqG� 6��	�۬F���"Oz�Ҳ"̄b
"B��.(t�B"O"�y�ꄂvR0��Ê�Z���"O�b-ڢX`�5A�U�(S���"O�`c�%_�顗KI*�#�"O����'Y�%Q���'.����"Op�9CH ���$��&g��T@B"O.0�&�o�8�j���]��MQ"O�X �F�L�UaC�ݖ*Ԧ�B2"OFD�˛;kDZ�s&��28%<��"O@3@��p�h|�BA֕ke"O���F'�(I��2c;>؁1"O�0y��Q2��<�"O	��0;�"O
M��%�Q~�F,�=�(�2&"O���ǉ-@�� ��� �p�"O:�DC��B�rwi�Z����"O@03B D&8���G��D��J�"OF��g�ܼh�~�&�/(��(:�"Ol��GD)�U)@ƍ�W�r, 6"OfD@h�7Sp݈a�sZFL)`"O*�&�f8YR,Ώ3HLy('"O�1�,m,d�K�
��.#��Y'"O�]�5$I!�>�"�Ci)A����yC�V��(����+
@�r�E�+�yf?V9b�q��˗&w�,
�"X�y�Fٷ���{Vm�o�D�VF��y"�TF�`�%��ltx��l]'�ymN�?Y�q�z �	K�,U��y"���¢� �zf�Y�����'!ڬ�sɞ�J��qZ5���N�,�S�'^XpH3eA�oh8��iڟL����	�'���׍�5Aꅚ�I3$����'x�}z�j�.}����nM0��y��'��(������!�'/٫#�v��
�'ﲀ�!BP�PHъR�HhH�'�RA�6ϓ9
z���L�)�';V	8P�_,Ԑ�v�$9"��'��C�LY�k�D�:Vm��BmK�Z�<A�Cօtp.8��ԭL�(M�%�Y�<��n�*J��P **������|�<��Q�xc�1T�Q&NX�1Cs#]�<�v��S�d��B��Z�@�¡�BU�<Y�"��u�j;�K�A$�)�#�\F�<���Wi�F��(2k��Xąx�<I )�:�l�� 
%D���ԧ�N�<!�@Þ��)7'��7��i�K�<�h$U���m��6�X(Pi�<�p��T��,R��(���mD`�<Aam�84�~�yr$D�^	�tI�Ƀ\�<��̃IF���פT��beQ�`�q�<�J�[	f��  �F���c�B�<	�Ɂ�5�<�Y�D���!�6.�j�<�H�/U�t���ec���&_k�<ф�#?N
UX��Yjc|���DP�<�4D���$0t+�G-�ؒ��F�<نdP�)�V��6>����A��B�<i7���^�cU�8BѡcG�@�<� �l"�#�jc�92�Od�&��B"O*���ԐKV\Ah����`���b"O0����Y?�6��D�*dbPC"OJ%��B�]9��6R����"O�X��I�;�x�A�b�%P|�Р4"O�Z��C��~�� M%?h�<q�"O^���mA�2} �z'�	�V@��"O����n�	3�\|S�↴��ဲ"O]	�   �P   �  �  X"  5-  �7  �A  H  SN  �T  I_  �j  �s  <z  ~�  ��  ��  ?�  �  ��   `� u�	����Zv)C�'ll\�0BFz+��D:}"a�ئ�pgm�|"��f��Aj�
6a UQ6�Q�a��!�d"&� �c��V�EaA@�t$Tpa�N�ٺ�Ħʹ�jԢ<�����><>�k���J$��Vg�h+T�.:6.CF ��4o��h$��c`�N����	�OaZT"ϧB�$s�,�$�df��״h���Y⟠9w=>���ᆢT�M����?����?���?�c��-q�|����|��JI��?��H��F(*Y�I埨kR�L�?y������U��UH�LZ���k�UQ��U����`yB�'�"�'|���4qӖ�[%j�*��@Cg��$̰;p+�	_B�yD �4pF��ɺ ���ɢ�P���>�I	+4 ��WGU�Nժ�#�����"�l}5O���#�?�䱫Ղ��<���G�$�4U�śm�	s�A��	Ο���4�?���?Y���	q�	zd#ٛ%KXyLŤ2M�t9���O�tl��M;Ӽi��7-�O�m��S-�9�ݴDT-���X�Lt>���y'L��7�܊%{�q��鉟}��Ђi�<�H�cN�Ҧu����D��<I����cOD�8�� �pdI6A-M��%#?/^H���	��M� �ik 7��D�Ӳ%	�J4�F�b~�d"�
_�U�@0���:*^l6͛fI8�%�������f��0Ǽ}ae�E>`-j�m��M�Q�i����J+WP�3�M-[qzM�d�L�m�d$;�$���7-惡0�42����bQ�'�v�
֋&Cf�m3��@�eM��y��9pm�|�� �8>��Ĥ]��֝�Ķi��6mGΦa�IϥD��ak3��>��m��Ĳ�2��E��
���"R�s�Xp�4n��AӄbP�a�Dq�`�//>P����'���L�?W���g̾y�&)��M�X�8q�'��NrӖ�	��H�I��M�r��O �b��S�%����C7�����O�$_��$���O����3�*��2m� s�n��l@�qq�̵qUx,[Q冿b�8�-Jt�ԂQ��Q�!�bU̦�2�(�5J�eɴ��.��	8��ϕZ.0Ɇ�I�L�vʓ7L�	,N��H��K��_V��[E��AGB�d�O��d:���O���<q��$�\�)A�Ԕ#UB�j�O� �P�y���?Y��ېf��I>���f��O���$|�������,e��P��{��Z��[��A��M�����O��n����!�A� ��,rѥ0���'�\dqm9$}|�)��l�j�"�8�7{f&<hU ��\��L9�G��#�*�'����A��)��@�ș3�J z��^�T�OΒ!rh܀4��{�٨����Ob4I7�'�6��_�Oc�ɝ![�$���ܧNBA�$�ˊ<q�'��'~BU���|a�],PZ��
��Py���=� ?��x������]�'E�8QF��	Ahj�ԃS�v�V�[ܴ�?�-O:|��D������O0���<y"CY�J��q���~w���GT�ы�C�l��W�D�	�p/����d��}�P����
��$JD� �_�nh����Z��e9�%J3����KŴJٶ˧���81��y��ڐ�@�`��ht�}� ����6d�<�S��ğ���L�L>YQm	�l�x�K��X�^h\3 
��?����d�O��?�'_n4���=
R��Q�A9w�hu{��?Y��i�6M?�4�V�ɮ<iS�T^
���N�>���C�_�i��DI5��<���?��R���Oh���O�ՓA"٘(����j�-Au�ͣ5O,c�&(��,�Ysǡex�$9�&�����2���AG�ʖk�2tu�	R��$n�(27��_�ʌz�A1�"AJ��dI��T"��/i��2U��៤lփOÑ�Fx2E�sF(�8U( =����e��*�?.O����O>��qO��ss,$yN�,��LѦX�d�a�'Gj6-�O�Mn�,�MC,��i������	ɟ�S�+�&f^��0*�\.�r�!�ٟ(�	��X@�I��ɦO.V<s���/)�Zr��6�klM�(�f�x���W$W��b�axFH�_i�8Z�/�Z�ܕ;��im �2�.�?�l�cA�'=�F ���0;�xlR!gC=e�'�zlb���?�ĸigU��D��V }���a���<_�I[	�i��M�i�%�~�DY �(�"��#g6FY���D��hO�I�������F�D�Hď���lR�D���M�� ��ve��6��O�˓�J�'�?�G��^V��P,0KT$�sF3�?��������CL:ﲠb�i��I���[�n~X0+�邃��a#��]`��&_��s0�ݫ��H���RL��Q�߻	��O9�l��L�ZX� ����3Z&%;�O����'��6�HF�\�'q���X��H�V	Q��4Z�|-%����{�ID�'hL,I0@��~�Q3��( �����D�O�o���MK>�r��_����ӌA-"k��6��:v�v�'2�'����/��N���'$R�'6�NE.%��)�gL� ED��rJ�pS��([pT+A�	��U��J��ϸ'��Iq���$L}�6mr������}��t�C �-\�F��J����Y>R�E��睙\�F0qD͛-1�a�����m�+/��ɦx0���<��Ot���O�h��燴F�x+�؅�:t@�/��O��d�]f�2wg=A�8�ƅ�+B`��'q�7-�ǦE�	:�M����"�'���ˊL����d�=#�`-8Q��%i��а	M_D��d�O\�$�O� ���?����4'?�z�(qK��j�p�
.
=&�8�:�'��U	��[}�����*)wP�p �U'�x��X��"gԯJ�H�a�,l��ka��bJ�\y���˙I�)�L��ybE��g��!9)�6F���O���9@�ƕ|b�ݕcm���?�
[�5J��Ck��6�ݣ׃T�?��8T&����?��O_�}���߰n���EY�h�B7� Z���H�:_�zt�GŒ�B��4�'�1�%N���qD,�;e�$�zC[u<��b/�6��WHD�VQD�f�I�+��D�O�{:�0�I�z}Hlst/C�}�z'�8�	j��x�6� 'D�ބ�m�A�U�ea7�I~���D$�O�0�Q�&NtU��J�'��ͫ&�'��I�_0(��t�'_M0a���B6��#�Y:n$DI��6��4Q��?��O	p_��`�Xn#�T�(�D�E�|�	��R:���k��	��ihw�M3#f�ɠ:g�i��A�v�8V�� bҮ�3��:��l���?��r�͹#��EX��צu���P�-?���Q����V�On�dK��0�mWf���c��ե)g!�d[.tu$a��O�.�6d`��[m�ў�����HO�,k���gF�պFڏ8��x����)�������#=�H��3$���0�	�x�����t/V�J��"޲Ƞ0�7�5b��q۴H�TRF$ՌT�.�/�����>(�l�G刁2�a#b_���D��Nؐq2ΐ� J�3&j5Q��ɉ�G��x�'�&h�d�T*W(ث�b+Px$���2W���'�T�b��'�1��I��2tJ�>%B�9��\�R����#g�s���0=�D�A�b�8��(	 YO�S n���I,�M�i��'^��OG�IX�h���Y��9�+�	���pġ�R�F%�	ڟ$��˟ [w�"�'��)ٜ8`
	"��j�v���ReЈB턄��ָ�MK�L�V8�䢘�j2��y��-w��p��A�%d�8�fTT)�HsF�G�jw���%I�]�'q�)�a9]�t������m�4)s)^ �?�a�'}��I�,}1�Av#�-+�fP+	��'���p�FP�rج�Ҩ�$zf��K>�%�i9�'\��Pjn�f�D�Oj�K2�67) ���e&�R���Oh��U�U�f���O��ӧ E�5�6���uO�D{u���Mۤ��"@�6��3E�+7��!$j�Z�K7�>�W�2�B00D�w��E��&&9:�=�'H�AN�� �H�����30�Rh�'T"����]�'�T���fةss�}�π�V
��1	�'v@�z�Jh��r�ԶLH,�	�n�R�98��a�����c�d��h�\���i"�'#������
���bWJ�0P��`�5Քq����L;���П��<���	��l����Q��QmD���D��Gx��ɄBl��K�I��07��f�ɗz�
���`�)§={�q`$G�7����guL,}�ȓ������ "ɌEa�#[��dG,!�'j���i��Nbޠ��-��UѨ޴�?����?1��R��>�����?A��?ٝw��Lh7��"�|��ԋ�]z&iJL/ �r�:�J�hPU6ИO��[w��IR���]�xP���2܁(�XP�#��P�<!�4"͎�!�SoE <;>$�O ���y�gΦIrU�%�S�	���`JZzk�'���P���Ϙ'�t�:p%�&��t�����`����
�'�(	�d� �/�X� �IK?Rt�U����?e�i>�'��� �?<��B�@?�~<��M�Gf�TY ����0�I��h�I��u�'��8��%���ȯ5�Z�L��u�6T��O��>\@+j	�H�L	X��ϟg����< �D�x���S��C:03�0pÚ�~d�4�L�v�0�
#̨8Zr�a�@A�x�$*��N�U�'�P-x$	J6f��iQC�I���ؓ/Q�?!��'Q��XoL#N}�Ya�̹0X�Lz�٘'&m9�>+�)�mκZ�b��K>D�i��'#6E��d�|���OJ}����$U�,X)5��%E0��;��O<�D��e����O��S�b՜�X��=U�Z����y{�\��S84��@"�ː82xe�e���M��!
���36|�@�(ǘ @���V�J�z� Ѥ�+L푒iˁPN���L��y�����:m@�dE�& *�aÉԡrqތp"cQ�qaNB��-7]��
6�� y�|:0 �>(�&���ҟ�f�4
�0�v*����֠+���f�&�o�՟���v�D#Q/ V��	5�!���2�Ӄ�Q�a�"�'��� ce)h��'�E/Ir$��[>%�O�ҝ�iȇv�vUA��y����O Q��
��1�X�@`�^2D�z���(�3��D�Q�R����)�{L�)��b�@���A3<R�I8.ł���F�)§St�}	gGV�[r�8�d$D��#΀�G�xY�b�(���;E�/ړ�?�鉁Eba�&ȁY��e��`0K��O|���O�e����>���D�Or���O��]�$��a�"�׮Fr<Z%��8��������y;�	�[,�y���|��'Ͳ5yu�t?�i��}d�!C-�B����@��)ٶ�:.�h��P�V;#��$nWR�G�4OFp (�w�qj�hK�̖��g�haS±id�7m�O�����OHc>˓�?�4	�Z`𕃒��pCD�p�ڕ�?9��0?I�
Q�0J�rs@��l�<�j㉓���I��M��i��im�������i�|��C�B�r-��!P�)��jݣV��pŚ��?1��?��M����Ol��>1�Ug�.Ͼ����&������&>:.U3�V�J�ؓ"�ȶ8��xR(Ŧ� <�l>�r ��i�y0���1q�š��D0'򠙅Jz&����Ön(��2B�ՙ*^�`6���< ���Oz�=щ𤑁8��E��]�4{ܬU
���{��`�6�Q�nJ \��]���P4N��'vZ6��O��:�j3�R?���2
�X��̐o���0�N�8������+����P���|B��!5o�`�3IG���ٺ�'D.c��@���{�p%`@�,u<�� �q�H����5�"�A!��jJ��!�B8*ڕϢpؗeF�2��,)���T�#���'k��	m�(@���afU���ʃ,�ҒOj���K�^C\Z��z��Qg�^�`^�*�O�]Yb��Z,���Z^�����'��	:^�q��4�?����IA���'֔��$��U~��PP���B1�'�������d�C!7fL4��ȉe �Sj���D9L�2�AfG�'7�|	�d�=���Du�A�XE�()V֝�0xh�6Q����D��F�rNO�1����qh^"Lhh������'�r��<Ѣ��*y�'iڅgZ�� V�<�d"���t�K�a�-/^��k�N�'<RH9�=A<]��*�C3 ��2m�E��M��iu�'�V�F���R�'�R�'�=���͉;s�m6�=%��� �d�,��cRQS�a�!��r&1�1OV�Z�m7k�6M+�CF�=��ix�����.���J_/b<��ȝ���]+�
�|c��@t^��;t�*U�*R����@1�B�`�
��@~���P��d�'��Uh�%6z"�X��b_�h۶U�`"O��/��=r`
��ǃ�x��'�"�8��|����$�1p� �*���US�Eɂ*B-S�R<��ҜuU����Ob�$�O���O��'(8-��C�7�|�G���I�m7� �(Z=�p>)pc�<	?��"VMCr,�#�0er!���4r�~��w"�BT��R��hO�xp1	I�W��sV��.L��z�JĘ�����l�����'����$,?V6�r�.��vk��C�I��R��� �Hf�@�Ŗ>D,�O�\lZ�Mc/O��{��O��d�O$|��V�GYt�0�c�17�P I�OH���6���O��S
p-��1b!F!zb�	I�H��ZJ&n�ӧ*�.XI8��0W�e�Q�V�/�()���>V���D)��>�B}8ŢM53���s��ʵ~���T(^�'+�T��?y�Of���ٚ6�m15C\��JBE�|R�')y`@�gN����b`:H�� ���ߎ~V��4�T�h��f-@7�?!/O�!2#�O���Op˧6��@��x1�XB��B0!uX|��(
�^t�U���?�Rb�:}�~��&a�i_HXB���X��'��霝.0�P���(@�����S���	�f���R!���`b�%���F�%��u�iٻ@�b	�N�7+�T`C��%L'�I�nV~�$�O*�}
�'yH͊�Es��zu
�;h���'�bّ�I.:���*t�׌8�����o�O3�"5mE.�-k@J�琉����?1��?���7H9B��?i���?�w����aD�Ӟ��V��d�R7H�,(�6KR�&Rzh3���G�1��hN��Z5�*T��:��
�w8@��a�E�RK��H�j$t�"I�(.c>�Ĕ>��ܙq���`F��.n���%�ПT�'Z�����?	��� M�Ƭ���-E�@
G�ݜ8M�B�	�p�D(ہ!��LT8x��٩#@�ё��SǟD�'�J���ݢ'rxu�E"�h�%4*`Y�4 Z9!��'���'��4�'�:���sg��x��L�b���bA�'��%�k�7N�5��m y��I��D�R�Z��d]�/�ڡHVN�(* �24O؄[/�� mP�d�FA�AFܯ�O�A����5%���ůU#e�� R�ʽf�r�'�ў8Gx�`Y}���R�8a�H8Z���*�y����̡XG#�)e�B7�D���V����'��?����L~�3�,6{aH��O�eP�[U������	��`�	�,�'�uY�JʽVpH�*F�Ļ?7��� (SG��L���i���w�%?��e9GL'ʓ[�����WZ!*�d�<?�e� ��2�ơ�q��3n��P��ם>�H���1�/�=�	���')�P1�)N�
�lДAV(b�1K>��L�H��B��\���)��7qR	��I�?��ǂ2P�DM���11�գ���ݟL�'%�̠��v�����Oʧdq­��`=�葢F"3]����ܖr������?���L�;y� �dU�NQ�F�I�vv�y�tcL�o����� ���������)w��)i��$���vk�8@Z�:�0��Nw8|�J�'����#x��I�M4��Dm�)§ �89��H�#�l�3ЪO�E�>`�ȓƪT��刪u
��T�)�|�E{�'*#=�MVm�c؇4����f���?�L>����T=�u���?I��?)�OP��f�15E|�	�J�(�j��`�D]TsPD��@���c2�+��O�Q¡m�p?�@OK4���ʝ-��8��R+n��W�
.�.��bY�@_fq�|�"DUt0��)� bhf�<=��O^1�!���'d�I=
,��O��=��,أ��P�F�7^qV)�qkD��y�C�0S�b�J�d��g-��ֆ�)��Ćm�����'���nޮ�iR�5��$�OK��]z����`^�)�I������aZwF��'Z�	Q|.pS��.F|��b��[�\� 9���O0�a���P6q�V�nZ=0��]p��	�`&�h�7��BY��Z:6`C1�,p���(��O�#odu"�4RFD���h:ʓn��U�!� �X�"J&Y���Zo�۟|r	��(H+ n̨U��"&G29l���R���M�
�X�A�.%8&�$��ߴ��o+���d�i�R�'�j�͙'�8�ie�L�Z��'��,Y5���'�)Q<3��	`0�W��7�u'��ʖA��<:���֙b!�3Op�y��ё�T�AD{���sFDd�*i��/u@<�3̀�,��i5�<ړp�������L3P2�	J*^D��dY�v�D��
- A��oT<[�FA��'�4��-�?��4���I�,I�Pd虝tI�tB��m�N�O���OL�?�3��Ꟙ[�I�{��x��D�PR4�Jaϟ��	�_3� s�C�g1\u)�O�{ql�P$�H5d=��O z�Pg��B*Z�e�RX�c�O�q�-C�$m|�k����@�ɐ�>�;H?͛l�0nr�1����jp�	��i"?YR�ȟd�IH�O�$Ȼ;m"Lz2�D���,�� �!��:�~���c�>N�U'���?�џ,��i�$^��1C M��%?��pr�Zs�B�'��	�G06�s�/V����ןp���|"rn��C�B�#2���44ǜ�H')� "W�`H��S�J�<��|b"�_*~���	�Ǫ<f��q��e�W��)_"�i���F�PV������x0k�ژO	>E9��@?���G�	� ,0�J��$��ᢠ&�͟��'Nb%���?9��$��X�v���
L9�Rd�*� XHB�	�k��,���A9DЀe�S&<ʓxґ���ȟ�'�"M�ҧ��*�ʽP�&��Ջ���;+ax����'�"�'Ҧ=�ip>Q��@:J.H��.��^�@9�7�A� ���F@�~-�t��F���a��^�}~Q�,��K�x��H8��
^4N�!�*�+A�x��7iI�Cߐ��wG��k̢ c׮[�M2/V�'��'
:M���͐CZ.9QS��"\��5U�?�?9C�i�76�����O�Lh�o�!e�R�a�IX������'N�������ԭ)S��
?ۂK>����?y(On�HpB�F�t�'��p��G	��:���
�.�@]Ҵ�'k��!	�R�'[�Ië'�F���̗�������;��w�C�l�8i�k�9@^F�Pt�6�&�� �ٵVǚ�h&E�[�čR0��/.ra�R��h��M��<s����ڏ���e�x�4�?Y����d��(��M5 �j� $�1��'�a|f 4N�H��>Ш�P���'�ў��?r�L�ے(��-V���GF���'t����Kk����O�'E�*���kv$e7F�*�>5p�CڣK��I���?)�^5?|���G�	&��hG@V����c�W8�����<\�F����W>02�Nn~B�L������G��7[֢�����(e+��{>����� ��ZE��W��L٥�9?1������J>E����8�qcU䘉X5�L��g���yr�_�S����M`D:�C�C���hO^�Dk��ug���hX8��g�2B�4��3�] �M��?A�l]�e�C �?I��?����yw��1� ��^j܊�ŗ� Q��3 ��4g�N]�B˶
^�ip��T�|����M��� b��Kv& ��I�h��-L�9G���W�������|�k�Kjp�v,�q�촋q��=��'�䴻���Ϙ'�T�ɴo��h�I�G�����Xr�'L����l�&?���fH� �|Q�.O�Gz�O��'���s���	z3ܠ2��X'���:7Ô/K�4ɗ�'�B�'#r�1��8iS��ĕ�	�j��]�RĎgB�UZ㘁��ĠV���
]+`�Gy↛���kt��h���
� :��[7��,q!�}Ȗ̍�`�@6�C�T����8�N%$�����o��#DV��^-!b� /:�D���p��D'�t	,d+��:(��x�b*�w�j���;�2��i2+�	H'�ɹ>r��'����4�?9-OM����Ŧ��	�+�� ~���@��I�N�S$F�ܟL�	lo�����Ļ]�0��@�z��w����(�kP��9+�ݹ��=_#:Cq�1{8 �@D4ʓ.+�M��\&l��")@ЄX�F�'�25�C�x&��� N6R�m91�~�j�q�y�н�?1c�|"�:�����?'n�Mb�"Z�C�Ɉm��	�n�V��� Y�NG���G{�O��D��q�ލ�vI@�$2��H�"`��'�ȕ��ih����O��'X��5��e�.y8L�]��`��C'>8�8����?Y���d:�����ΐ��yX�K�.��/�S��:{���G]�q!�t��U~RN���ȑ��Y��8������ĉ�F6 ,��s�K������D�'�O�%�"|� �X�u��%x�$l�E������"O�U���-K�T�҆�� �r�h��	)�h�t�#%J�4]��2vGVu�f��"KӦ�OX=��"�Dn����O.���Oz�n
�c��X��H�0A���#(�|�8Q���`۴3#��$�ZŢD�X2'B�������p@<��.B)S=��$1��3ľ�M��E�� FT�g�Xz�:虉�$tޝ٢����t 3,�N��� $ݦ�.O2|��'��D�?�O��"&Ŏ�@h�nL8)�`p��)$D�y׎�5ϤT����L�<X��/�<i��i>���RyJ�@ ����f`pYz£�*����4�Є���'�'/��蟀�	�|�uߕ�V��u'сИ\X��A�9z�Ē�l�lW��q���Wo������Qb���Wj�(=�mXq��2n|4�C���B���RK!t*��aΤ��O�*䮄?B"ȡ3I�J�-16���L`�`mEz��	�5�ZM� �ڹo�yǠ~��B�I�O(�`�ƍ��:\�$BŶ���O�m�ʟ�'"%�h�B�d�O.̚Ό^�a��B�#�2l"�`�O���^7n#R�d�Ov�)2&u�5�3��ċ��kk%2pD�)GkX���u�2R!�ÜvTF<W�	"Gi��(5G�ܸ[��F ��0���3b`yG�\�6���B$���Z�`�	C�c��z��O'�Ę�)�9`\���/o�ֹ��! D�"��:Z�Ypo�L^��Rl)�Id���D��OjI���'+Hx��&œlA� ���|��PNT6���V�>��'|���أ��F�`��R�0e�~4�'�0e���8V���AȚ�$��D��AZ�J���X�L�[7��������$Nϼl���W;����p��(�U�uL߰@9R���O��TTL�:3������O��nڲ�H���"X����-K�j���k0��r�lB�OW��ЕEX�ad�I�ԍE,~WZ�?�D��,7s�	��&ބ P5�u�8�nZ�~�$��'���)�Q>�< �F�� LY�-�*�^,b�DY̓%Ն���� ?G$xZ�h��4�Ӡ�(p�b���cD?LO0+C�͛���]�6���Uk1�d]�6�����)(�FEH!�S�()����ǯ]!���>CD�+��-Er��g�I1�HO>Aq0��0r�X��Si��@�H	��F%pJ��`�O�`�̌k<$=0c+��M�d�#P�����~��F"AS˨p����C�Z�b���OJ�@f�O����Oڔ���S�l�Gg�s�ڜ�@G�nCJe���F�oB��4 #`��=�d>�yqk��e�\�#b��XZ��;��Q9�`^�_J�u�Q��,D|G���?�����OiTy�uI^�%m�yc�)i��M(O���䍨=P��i��Es�X�E�҅d��}�d�<�Ā�6b����Q4u�X0��Vpy�B�[���'�X>��F+��T���A���2���cS�q�an�^�"t�	�<НB�㜌*�<u�&)B/a�,�Y1e>u�|����4Za�&��-dx�y#��U�<��'[[�|as�%�/U�Z���fP��|z%`C@3���FE�M�X8cA�\�<9ÞƟ��	~J~B�O��ӥGǸt�&��0k��V��"Oa��ȯPL���g�����@��>�ȟbQ��%ӽa{�RÊ}��E��Oj�D�O�墢hK����O����O����O �xE�QzO|XD�Na�!�cfgTXq1$"
�vG<�`�i��*+��'�@�D�&W�
Y�$� A\�!����[� e��N}Al�aǇ�	E��'#�L➰��iS�9[D���ی5��Đ��1?)������In�'����/|��p*
5%�r�� !�
!�ě12��Y#9�|�	TO��"�#��|�������sL����3g���I�
[26�t�r�޾~���D�O�D�O����O��d|>�j1&�~�\P`�G|u��,�,Tj�A��G�y�g$��C���S۪x �"�aR�� �E� /�=�U��*i��e�� �2Y$��!dS�[bQ���fK�Oǹ���3���#+R'&�d��Ot�=��P\`����<Ub�����!�dҨx���'D�#O\Y�f����	 �Ms����$�?0� y�Os�8�
���"5e�b��J��jUBT�"�'���:��'�R�'��b�N�s��4z4�ϔj����/���Y$��$=��m����>�԰{�$����E���< �d��
O�>�*�N�",1Xh�]�M٘+�DX:j�n">a�%Fʟx��_�'h�n��lZ6::n�6�ɀB��'�a~Rg,��m�����X�K��X2��>�@V��;K;}*>"4�D\P�c�<Au@��?I���?	+�%�f��O.�DǝW��p���o@�H����f��ĝ� ��e�ƃ�tF� ae���':!q�>��b>��".�,��`�X��*P�x�`���*o/���NR:2uȕ��>.�Q>Y�E�?0�h�wkL1�]x�Mw��3i�O��$<?%?U秀 X,� �р��J�����
�x0"OĀ� (�7cf�cb@����E�ɲ�ȟʕ�΄aM<%ڶ Е0YL�yD�O����O:���GC�pM��$�O����Ol�i�O�����0�����7'����i+����EV8��,p���1��I�㞠���^����P�G�
`�=�J�1x;p��E8ƪ(��S:k���pB�@����~2�5��f��~-���:?QE՟4��x�'��E�]��a�Wl!nA݋�f��G!���r'�@%H�/`�-��+V�n���'��|����䈲�nTX$K?U�h��4
��/|�!WdK�L����Ov�D�O��	�O�dk>�XÓ�al��c�ΩL��s쇣f��-���!-�,$��`\� ���k��ɶ�\���/�4��ŘG/��Z6R�Iւ!Zr�2�o�I��\8��H�dJQ�z���O"�q��
u@|��Z���A�
�Or�=���D�� Kƅ��N��&I�f!�G�s��$��Eő �r�����3�剩�Mc�����ԗ.�lU�O�>��=i&�C"R�:�iW��]��;��'.F�KU�'���'�*��u�I�D�� ��aR��U.�Ԡpj߭䀍;�EG�u20�v�	-`�Qʖa��a�zP�N?����1�T�b��<�@�I�l��DNs@">�e�\џ �	X�':���^�(����G�4 ��'_a~"ևo@}Y�h�1EȾxI�A��>��R�ģG�Y�z���d�Y�3Xc���<Q���?a�����|j��y"N� �2`Bqm�,a�
������~�I�HO �8��[*E�|E�х��zt�;%���xD�O�|q������ބ顤���*��y�fNn���lZ��B���<9�-��x�	�?���?)���=� �
R�Կ+�H5��#[�J�����4�?�u��?�D�'��P��M�;M"�����b�T�BuFIʁCչv8JQk��ϰ.6���OJ�K�&t�4���?���r��y���L̒ï/p�����, �j�0i ���?y�^9�?��'�@�j��M����I-B<mi�/�m���TG�9�����
���OZ�[�h���']"�O��iK_�H���.ޑ.�6��ǆ�)�(�D�[��'#�A5�'�F����.@��i�(�"mT�.Jp����ǹ ��UPw�Y�!�6�i��h`�Op��Ş���I�?����=A���J�'�|T��Ph�5�l�ϓrvD��	ޟ�Z[w����O�a��ҟ�6oP,[��  ��J2(���ON�0���A�x�牅�\�lZ4�M�2���������1���V$��h:\�ar�^�r�nZ<�T�Γ7BH(��45����O��2O�����T�0��	 wB��s��_Ezh��~��)y��������M[P�O�����맅Z�$�$\�T���Z@�)�-�m�!��ϸD�����	�/!N�`!+|���'��T����p��o�H���!�%H�@dE����J���'K��'��'�r�'��Sg:���v�)3���&��)����妩��dy2Y����uy�X���q�H+�,��l�u&���N�MK���?qJ>����O��`���{��L��Nd�H�"W���W�'��-n��sOC>؁�Vԉ���%������D%���'P�� 1�>��0�ڕS���(R�չ6��6��O$ʓ�?1��?�*O
���?iJa�'v :����#g�&�u�*D���h!(*���� ��
o�q���4D�t�֋B;<����ě����Б1D���&��v)��� Y�h��5Ђ�)D���$'ax�Y���Õ�.%�k,D�d��@'b��4�t)�$�:�T�/��|�Dp1��w�}�&o�yn�9!WLF��􌁑+ұ,&4JE��7V�$aI��hu�CF4U=���1���؈q�,�~�D{��⟃W����Ђ~R�y���ݟ��'jpqc��H
|L1C�=H�Y��2|g�� 'A��H��4F�'��Q!$��3M�% ݵG�A�bH~�YY���`{,u�,�<U0v��,��I�f�G(��� ���@"��7|��чm���[#Tѓ#�po��AEE�.xNYlZ�zs�I�XR�,�1���R� �ȗ'�'-ޮ��hO�)0�	�{�0II��<��,;e�,�C�ɢI��$�F�[b��{V��CTB�ɜWp��M����� ��/p$B�I>c�m(+�god E&�4EXB䉹?����ïD=�,�$��&�@B�	�^����,M"���dM:#�^l�ȓX6H�P�\�NH�e;v�W2n��X����&!	�ۨՓuE +}�h��y��Ӫ��S����@�]�~=�Ņ�H�� 	× R����d��z��Ȇȓ0"��Y��i�&8�3�(F�̆�J��)�u'*_�� ڤ"��00��S�? >(r5I�i:��!T�ġ3����"O�qF���K�b��K�?*f!�w"Or�3"hӊl5޸P�'�+~(�"O��H7oO��E`��Pu(�"O��cE-��Q�׌БX�H`��"Oҽ�tmS�C�h�"�Ю>��ȑ�"O��g'΀I�R�,N��t2"O�Eb��$���ǟ"��)�"O��W)���y6�ɷ.�>`�a"O�<� ��'������t�$�1"O�A��U~��*4&�4`Zl!�"O�@�u'T8,�~�q�$b`�ѫP"O�����+�|01���QV��` "O��#T)C$)vQ�T)�8$V�\��"OfI��I��sY�M����EP�"O,-؀C�U�:0��hM�0?6��"O�10eg��7�p�U(^6$U��x�"O��rƐ%x4�jť�Z���"O��8E���r�:����	�Qad�cG"O��i� +"���;ӨցkL���"Ob5�sH�A�8��I�>YD��z�"O���.GnݼQ� �
�0,* � "O��r�� j�&r��W�f?�1��"O=��	R�]�y����e��Q"OH@�&��p�� ��0Tm<I"OT�Y2�[� d@E)7I#
�$Y��"Of���Ü¡Z�@5d�zآ�"O~$ђ���'i<a����fYKp"O�=����Pz�0�۝<��="OX8�!H�)�V���n�?�~,�c"O����)6o�j�i�M<S�$ŀ�"OxT��BE6-����b�J�7�h�3�"O�(�H� !~D8P'lJ�,�)�"O2(�+Q;{�!���ښL�܈b"O��9U@�\�
y��o��5�"O�H��$M�B�, e�_71w"ܱ�"O6q��A��=�!�(je ��"O�y�$ ]�Z̑�ΙU@u҄"O½��K��� �6�H��l �"O�=B��ד�����������BV"O������E��{�
O�fE�"O�"e���8��q�`��?i�n��B"O4���*>,�����[n\�$"O��J�lŏcBBՐ`��mC��Bs"OJ�b���~��4�S$P�iB�Dj�"O�hs���Z�61�uL�/.�9a"O ��E������9i�̀�"O���납u���rC�,sq"O��a�Ҽ��i�'�M�8�pو$"Ot�d���:L)@+M	0�*u�2"Oҹ�F�ңe��%*=K�� kV"O�(�C臌��a0ţ4Uh���"O�ZK��c���w%��$	k"O�0�@J�2�Q�aE�b�qE"Of	����c{��� �W�-�@l��"O�����4+X��`�^
�n���"O�ղ"�ğm_��ڷkC0o���q�"O�,󧄑g& �g��<Ũ,�"O�T��@�t�U�u�;J�6q#"OV��!ʚ.M>�l
��.]��].x!�" �@@�
�
��)|�!�D�~@��p�!b6!�`	�[�!�d�_c� Y&����T�w��1�!��	;t�\4�Q�d
 ��GD�XE!�� �Ȳ��P�sxL$(q�ʟ|���z4"O���ӄ%Q̥� ��r��C"OԜ����w�0!J�{�a "O�U �7UR`"��\�7�x91U"O8��DDL�3�:1k��F\z��F"OP�ϟ>��sRQ�dv���"O��pBԞ����ܶj�^�x�"O���ٛՔɰq�Gv�9"O�ᨣL9Ѩ�k�U&@�� 
�"O��{cL;ob�E�Ć��{D�`�"O�r�GV6*�d@��$͊?zv]�A"Oؐ��I�d� ,�SFͶ~���"OĹ�B�Ѱz�E��%[�P���!"OI�2���F�"�A�f�f�r��A"ONY:�LC�L�6a�"œ�!﬌�`"O̵�6@E�&[`�i%��
u��T"O���lr��Cɔ,Ϊe�""O,���R CU>y1��f��eR�"OҴ ˴.��� �ѻU�r���"O�@����L:<��!F�+�0� "OFI���\56^|;B�٦%֌�"Ovɚ$���7�x�q�(�~��"O^��E�B��بLC[醜��"O<�jWNO�O���)R�6�ިy�"O �Q(ؽG�`��I����I�"O}��a�/-x	�a���.T�$"O:��b^~�
dq�O�9q�X��"O�h��+�-Q�e��N	4�BHI�"O�݀�`�w��P;��U;`�4�:r"O� ;r- ;�i*D�w)��G"O����A�$^R����U:�ٸd"O��#�J�!ʥ!Ѐ��u��8�"O(|�ƀ�i���B�)�;uڝ�D"O~��6c?��4g�=f:�js"O�9��I�iYMHM�nUVi��"O��G�ԟtL9���̡d�@8��"O0�@�톯\�|:F�ό&|�9�"O�y�bჵH]2��d@��.`r���"O��Qe	ϣ4	���/�$cR�L;�"O֍����1/ҭK�N�&��UKe"Ot�q, �2�!�-Jp{@0��"Oq���[�VܤDR���pd�yÕ"O�j7 ��H<�$��67��.�!��?,�]$([3l��lۧ!:?�!��ok�4���m�@(��o��,!�ϱo���k�l�����9�!�$�Dm���Z�S�~�#2,�1M�!�ܤoϦ��e��(f�dH��<�!�䟦^4�A�&Pm/�<�`�ϕb�!�䓿
���W�Ɖ/N��uN܄)�!�$F�]��"3

��0��o�!�DBE�(Q��e�i�U��
X&z�!���
<�����c<$ �u*%$�!���96�@a.&H+���vI�e�!��*Ҹ�G�=4&�%:q)�?h|!���2F���𗆅�*$��0��_!��(�(ZS�Z� CVQ��� C�!�d�=lk�U(p��7t+~<C�bR~�!�d��+f5ⶠNV�}��� �S�!�D�Nf̰���T�ʀ���-^!�DV�:�@ Q��Qf7�(x��E8GR!�$N�y�L��"GN��	����!��=wH�����ֲ�pH:T*�&,�!�D� ]���a��e"�x��e�!�� Е[7��4��&#Q�mn1�"O���6b�l�h@�ˏY ��#�"O�ᇃ�
�NJ�)ˬ)��;r"O�����qL��CNLF�"< "O`�i#���&^�z�7"���"O<XZ%OƟ٘��d&p�'"O��h����{���cV��Y �"O�P��+�V
���bדD����r"O�%"�mt��S"��z�H�4"O��P��<hhL�@�Ӿ��Tx"O�չD(�5
�: +���.Y����B"O��I���gق�rS��$8�"Ofl E;^q$�N�6�@R"O$�6H�;�diCƧ��?丰�"O�IV�+��F�X�h��S"Ox:���D|����п9�`�� "O����"鞬��!xz�1�"O��J �zZ��z�LR0 hE�"O�����
�-0�y�L�6~6I�A"O\M���Ə1֞��&��Yx�x˄"O���W��Dr�ճ�(Q��_!�D�"�XI[��P�
)&����0eG!�dY8>y���@�-
a��& 0=!�\8g*x��HL�.�4}
��@":<!�JԽ����x� (�o��O!�߰K�E�F��Ayh��r.�O!���J�]3w��Se6���͐R!�䁸9>zT�B��?�H9*ׂ�0!�$F��^L(�*�"g��\��(m!�d�w����kГ{d
���̗fd!�ĄwT�Q�6(�1L�q;�"O����(�lp��]�,��XA"O4)�:s�p��
�/"�"O�$1p$3+t\ۧJ��_�N�8R"Ol�җn	)Q�زG�σ0� ��"OnyT� ���D ����j>Q"Op�ѣ�H�($��(���" �B"O�|j�A�7{	D @4퇒N�*� "O�=Ɇ@C�E��u!(�H�3"OLP�3��Y��j��Rmty�"O���1�C"6���3f�їD�F8p"Ol�G�I�l&�8BȚ�c�.��"Od�!�V%0�RH(�$J�}���Y�"O"��8n�qS�[��@+�"OF�C�&�h��I�ɍ�|X�"O�쉁 �N�n����ܶ,Ն,�"O�us�jO�h~�%��@J�`9r"O�l��ŗ��(��!z�ڈ{�"O6���:K68�䝕d��"O�aZ"O��"wtm�1c��Ta�"O
�s��83�H-!���Vxj���"Ob����Z�ܣ��'Y��c�"OT�fN�:���ۢ�:)$�r""O��s5Α-|���K�O�4K#"O�Щ1Ǖ�>��|���&L���V"O���قJ.�� �Eҫ/-D9�"O��`���8n�0ʧ�B�BZU�U��I1+�*�+$��O/Fq�6�Y.U�'{�ʓ�C�֭0���*��P��'��ɚ��]I������'l8�A��i�J����u����'ut�g�ҒK�z����=h< 
�']a������� ���'Q���qk�iT�L�BBJ.H�Hi�'X��lѥ���ME^������ �@�i��W����Ҷ5��@�"O��)�'E�v�&-p���=iʈ�� "O`���Z	�B�Jt&�&e-^I�F"O�ň�IF�c�.�;�f�.'�%ڤ"O~t:�P!�^���oV���H8�"O��v�.XX���4��I:�"O4����wO��˲g�"�\;�"O�HR��4E�>�1��.����"O0R��Θ[mZy�qo�~��;�"O�Ei�)�"�x36)ܝ�$��"O�����?1{N�R�Dd��cV"O8B�ͱ0x�d͂���K�K0T�Xn�^�,Y��E��V)��9p��������jfA�qNj��;�O~�֤�'�~���ʨ ����G�G���녺A���8��94A��ɍh5V��P�R��U�� 0Q�"=��N�:�Hx�Q%Ͳ�Ly�	�����d{��Ҧn�L7x�:�cC�MW�B䉳�dqD�#~<L� (�6m��ȼ`Ƌ��I�  "��&Go�����y��hY *��Ӓ>���"O��K$�,b�b9�@C8���p�H�$<�oZ<G^�he�PN\�'B���Qe��gц(j�,��<)2hH�+7�O�dђ�_��52�`��.M:�jc�Y~�	��@�v��֬S�V�ހ��ICn�	�F�:CL�Ӫۺl��#=I6)�1�D��
��E���k�eEƦ�ӝK.�'*Pl�tF�X������'9J���29N(1c0oUN��̻À�-ϛ&�5FLf���M��9��a�	�"}�1}~�0���M�<	QL�s�̅F{Bϧ�,�E��"���˴i�J��bD�
o��.�$�ɴm�j���c@�>���Vv�'�8��4AD�1�I�6i�)�0�Í��D�wd����)�92������*dθ���4Zm�S�Z�B���1C���&�0>�OC11��������*ԝ�t
T�<�I�:�(8�6Iͩ
��U�GK!��O'�Tͧ�:l�u��:Bw����"CN�E��ITpF%B'$�6$���H;|�̑aAԘi9����_2J���i�<Y�D���K���$���0��;��ό�r��#GşP��c�+�x��0rdslE�Y�v�x#O>�ӿ9�D�`��=e �ay��U�����G9A&��P(�Ю�S!@�~2G�Qj�!bHߦ"�P��`�N�S�X(���a�l(ŞO�5���Z�N�M�0���N��Z�P�o׍I��tڐÈ/i4qxu�]|�T)GG�*"XԀ�$^�Bm�7@g��`4HU$KQ���K�~��T�����Tc��T)eD^�b�� ��b��D)�	�.H��,PUk�_�f�1�ߋzyT���W�M�x4�a/�p���O+].z��ЀW\���0��N-��1&�Z.s7.�@Q���`����>q� H~�8�J�Έ�*9�ܺ��/F�F4$��E#M�Y���0�^
ŉ�=ipd�IUd�rqͬ���	�|�'':�a%C�=��t�@�A$�r$Ks��![�2�ڗ�]'N�C޴$i��z �/Q��biR3
�Z�	',�"&��Q f&4�$�Ũ,���%}ԝACoݔ\-�v���#^,��94t�L�q)�")G�+5��=T�@-�$*$�l��]�l��aI�M
&��P��ٜ9M��Ĕ*lN��k�(_�ylY`�Ɣ~�����a�Ajr��%V��M��?ݎ�2A	�F��YE����4v�ipЀP�7�LAF!ˈ8�"<�M�)l
����F�nI�N~r�MY!x�ܴ�c)�Cg
�pb&>w^����U�\V�9v��/g���O.�導}�fH�T2�R����>
�+�f��d�5��l���U�N1�?��'jx(���
�X�&��?���鍙|�H�W S�K@�8[p&ǉkޙ�s���>�0����4��	s*O���3]�-�p
�b�B-����I�P4������|B��i�B���o� JӦ8U�����yҮg����%Dh�3�dغ�(]@ƬX4f�����~��%$L
Eb�% A�i���Q�@�""@斡_kf-��f�E8��@�
4gfX�('����iR�k�+��,��pԠ81��vݑ�$?O����Q�:
�Uٔ*&
h�j��>������dBU8HROњ��'�jI#)(b�4��p?Dֶ�1��d�	,>�l�kv݅��{*��t"c�
��8�S#�9t]��Z6�Zr��ٕ�����'3h�!�dF՟L��BS"ت��¿8����B��4�4T"���s�=a��N _��Јt�R�7���e,}ᐅJ�na9���g����,O��c�"P�B�#6��+;�&EB]��	��(�I �dT���L��$J1��m���HGH}ipkS�H�݋p��&�s����2ߴ]ȼ܉t�h������ي��[Z��|��c�/r �h�]�|@���� ��.�qzx�E��O�{�@�e�8���747� b�ќ���/�n%��O��%Y��]��܁ @d�UC��?��Ʌ
��"<ͧC�2��ң�6�ݡشt:e:�Zgdpy�K�3%T�5�D�C�S`��rB�T>��eԞ4�{�? �QJG&Q/~�x�n�'�0�� �>1@�4q�@`��I�
i�%���O�i� /�8�l�"�%+����S�<�����,�h��
�8Z*�I&�6ʓ4y���iK3�\����ϱB���K��
?1��3�'���%o��+.zL�M|R��1t�/.qD��bH8"]�(�r��N΂W8��D]�aDz�:��@:J>����[�a���B�׉h���K�Aڼ4�H]\��C�ӛxP�!3ë)��l���3�&��	L�m���,sj&��5ժU#���v�FNX�)R4�PQ�J%b����f��+d��D�}��<Ӥi�;�JU3�b�Lv49{��������(�����������U�<��[q�Ή�.x�A�Oޕ����5�l�y�������-�b����É�X��x��l�syP4)B"X���'���'&�bP�΢YOL�@ר� m����!�0�����koVq��߿�(��I�R�؋�D�k!j5@K� ��䚝Xˤ7m-�ijs��l�\�o�$cVJ~�C,�q��@Ŋ�A)�<�/\�<�G��PTRL���8:F\�0ř>�ΌG!�K���a��8cН��OV<�Ba%n�p���J��0��`"O˒��5w�l48�.J-C(p	A����LIzXqc�V�3�"�3�� t�axrbU96��³� J�"��B_�0>	�ĸTz��	�(dR�*¤V�<�����W�C�	-qԲ�[�� _D��;s�כG�`�C%;�ɻQ��	f�u�ve� ;�f|�	�.N� E�`�$D���G����$I����(~�)õ�?��$9���(� �Gv�'1��Bw��"{�遒��j�9�ӓ}}�A�ŃP�Mq�I��q�+���8{�C�.��I19r<2�@�S���9PIR%=4)Q �>�ܐ��$~ݒ���C$TR����uK�0l�C�5xnE�cD;�y�I�5��)�3Rbt�v�׸-$\��M��M�eNZl�S�i�1c��ݒ3�r9Q�OB�6�� ����C�C�ɖ�h,P�@�����"��Z���\K<�AB�>ׅ�"U���ɤ�?��;��`��/I
���BA�&#N��$֟�$(�Wk +E9��:��~�V(#� o��`h o�P|Fdx2h�"2�� �p��f2�q�clӆ�	o x�CS#9���)�C?y��,'7l�ΙPm��f)�b�D]�s!�	`g�B��@���6�Ӻ���/�|o������XgM8�M���ȏOv�����57�,)eXw�'��񲎇j��uoS�\`�d�)=okx٣��`��b��1c�nmi���$��l�����!K+][�,aW�K�[�V���'7��Q�
&���zu.s��AᲥ�n~��L\f�`��i3��O�L6
�mv�*�U�'�.��r�@?̨]1c�,3�>��$�C��1�r͜P2�e�왩8�L�'�.��}yb<Vz󂏷>�·iv��c�ip��_6D����s�C�O��aÍ�&iؑ�劒R	2k�x��[$e�,�\�l��	�?��t��OźL�X�jRE\��>����R�u|���ͪ��i1}xXh����ըOZ���O�D�~�;R��(�#ìU�	���H�U��nZ�M�O��"B5��Fֽ=�vy�4��@�F����	�d���e�w���2�.j��zR"L�n�����*#^�r)��g��U���1Q\��|��w>��'tMhqR� ��J�����îqD���� e��}��igӞ�ɕix\�j_��PXF�0X|]�r�ו@+��Bu��U�Dq��'�'7����@i�SA�<6[����N�40/�O>�1<�)�˘F%�!k��\?N�(���)k���jT�
�6̄���ԯψ���ˈ��O쐘���C�F̰��/2280A���I����v����Å�6�L����1Dc��h��9Y��!��J�ܱ�UFA�$tfy�F�2F�����+���$�h��r'X&�>�IBB,�d)���`��D���1�-��~$�0��%"#���y7i>d�8@�O�1N�����ܐx��w eC��$P7��z����wH&d�@�sD@U��a�A��>7�eE�$z�%S1�
�Z�DƀC�`MCg�кk��;�+�z�ay��ԱU�F�u�O.Z5F�vD�;=^�H��CįbX����h��D+����%��?�D�(���/f�K���+�Q�ĸA��J��U��w� txeI%�$$�6��Ί�x���qU凅j��@��f�N/,��u�?E��)��џt:����ӳ9�R�W,��"_���D�'�.�Ǯ�4	�<���]�u8pf�B>:l�H�Dc�k�^�YAM�3G6�����it�=���U�UT�8q`�R2��&U�D��	��J  ~��I�Y��y� �?��6".,�@��j�%+����Êĉ ' !�����X�Ы�Ȝ
v
 l^@��f�K=J��ņܹ�~�ύ�9*y�1d�?A�Ƹ����Ÿ'#\��PȲ\.���S�Ý�K�����Tؒ���;�l�18[�$Y h܃#茹p2`��cO���Z�E�<:�ƈ+g�֨8�`%�΍k&'��JF9z��5�p���ԨF2�i9�`��go0!X�W�|�N�h +��c�F8x�
�u�����V�c�n�L��WN\#��%`�' v�����)7�`��W"<n�n�Rt� �t���p���?�B����%w�AHфW
���Q.��t��T��s��ۖ  2T�� ������O��z2Dȸ^��d��ᛠN�� $�SF�@�Z�Hi��%[43뮔�K�$���ǋ��K2E1��Z�x1��RD�X�:<�h��)CS+.���'�ŀ��̩2�nM���ی����(Oʱ�1��OsָS �J�Zq�01q��{Ӡil�:7��QV#4A�.,���X�:�aR)��)��X�D�s�Gg�1�Gx��-��O��9����x�F�y�O���qb����zX)��o��g9T��D'F�*�:����ƹ�;u��čY�j���z��3}��aHE�LA��S��X���+�mܳ%�be��%Ɉ��/�_����T�x]���!|Y��I� �bc��{	��+��7Թ l��!B��	HY:����\�S���p�'C���v
B�N��a�A'_+ �ԭ 2� 
g�f��3�
%8p�'h浣q,�V�<��X�c�
q��mFZ���ڿG���?��N 4�X�F	�-n��� ޟ@w�U�/ ���ꆿkA0���F0���D��?��M�ji�6_13�!ƭ_�\c過��l�	sb݄�I1Hd�ApC�$$tLb�ɕkPz�Fb� $��IAD�A�]�(�&BvG�44�f�ٵ���(V�&D���D_�le@�e����ݷ!�xU '�ŇIW��)w�� oe|����5��]�w�Ox)��T�u�6�ԅ� �*q��0O%��	������J���IrԤs�JL{!a�+/"Q���&�Z�Mx�KvĔ[�Mx#e�;b,�ۂ�D��8 HE��?�@�jL�']�$����4���;�OY;4oF�z��'0��2P�W"r�v �@@)qV�Rc�	Cu~$ b j���k]95p�3R�_2R�� ��Oʨ�7��1-Xf1���͟jιɵhU�D�}ЀaS<�"aۙ{=,eKȏ;q����KǴM�6����J�@|���R:	��L�&i˹;=�e�1���G�ļ��-�>,�T�dL��0�`&��y8�h���� GgnxI7��=�fY�#dФʺ!�f�L�y��6��<���ON$�U��4]D�X�!`ش'�:!�d����Ks�
�o�1W�
��2ғHL	�����ywT�����dEn��r͌��Xx��(�:�d�rbL�|��q񑅍�i��|�1�QM�Fd�uM?ax�s�4�ZNˡd�@��Q�R5�?9�@��`�HĻ���ӹ�����f����
���49]!�SXJ�]���ڠ�`��'�`(#rA�+6i�U�'�����g��1־��J��:��< ������X0���.��V#���Sd���T5��9�0� ���O�@mZa���.Ȝ�%(�A��| b#��4���D4.�\�*tE��9D��'��!PQ���J�9�Fܰ���<уK���(�`d�5gM�{.��h�"V:�h]�"O�� Lܖ�(�iA�/� `r"O������)F�z����$�� "Ott�unSX�v��A�6 6"O��p���8�I� � ��"O}I׮�Xz���#�3܊P��"Ol�)�kB?L*Z�i"�z^��#"O�h�&����(T:# �(*YD�j"O��YE@؆���PP��?b\bm�%"O�tE_%i��%H6�'
Zf4��"O�,�3�Z>'�`+c������Y�"O�b!���R>�Y�D\k� h�"O.,�����P���`��@�"O.���C_�_ƍ{	Ei0"OD`��Dƕ������Mm��H�"O��A�@�A��I��o��(R��it"O���L0H�m�5N�r�2"O.eJe(U2(�sW�Ee�^���"O �u&Yt_zM�&*M#l�����"O��	�+�8���J��4���"OKE$D�RDє ͱqH~4��Ý��yRi�c�`5�,5��<:%	���y2`��%��4�S�@C (<�Q+\��y������8@�ZY`�H��y�3����Ȁ~�B�IA��yB,O�}��-��!I�H��u���>�y�hVsb��� y�HHq0�ς�y26�D�{��U<t��T���y�GR�m��d�g��z�0���&�y⤜�p#�̛LNJr����)�yOU�*���h�z�ޱHs�A��'�ؤ��� .X�U0�Ĝ�`�ЪO>	 .�X=��rCH�(Yh�[�c\l�<I��C+8�d�+@ Ơ^Mڽ��c�^�<!�&܎7�������E�X��C�W�<� ���-G7���3p�&z"��*�"O���$�)B������,+���`!"O��󃝀)�@]هi�9[�&���"O(<0`b

G���"r~�xR"Oh`k�G�4��0y� �3s�8�R"O����)��,��PY�ڬ~j�1Pw"O��pS*Y8 �T��q���U{$xh�"O��j��[*N"B�J/jh!�"O�h�Ɗ@�`�lm
TJO�|�BTp"On�i	�I�4����3v��;a"O|bY9Y�E�1S�7�Dt��"O�����̘0��M:A  j0TpXb"O>���o�Ơ�rM�0���f"O2̳���I^�5p�KͲu��1S�"O|��F�4���:
�yڠ���"Oh� �G��L2���
�4,��Y�"O�5�֋�#�C�)�%���#"O24�ט$�D	 ���B�"O�$`��Q,�1�چ¼�ʓ"O��
pOORgd���!�R�I5"O���D&��k�S�~�ѷ"O�}�d������
K�g� ���"O��F!^ݠpJ�W�>�2�q�"O`h�� n8�P���=��`�1"Ò֣�����X�$�zp.��c"O����9J&�:�Bؓ"�T��"O<�)d*Yz]F��6�B�"O6���dB!��g�� W�*�F"O��R��k��pcG��D1�4Yb"O�`��B�)��A�œ�0$� &"O��P�K�-�>a�`CɑH��`p�"O�y9 왠i�0	�6�H�p���"O�x��Βu�L�0D�"�.�2V"O���ہ_*��b��p����"OLsf�}ڐ�Do>m�DѪ0�$?�S��~�l!;��X*��!*�dOd)�B�	t<�hk����4f�պ�H�2;�B�	�.�	�t�Q�r��a �E���B�IB��%�{<�) r��C䉏Lo�M���
�#F��2��C�IQ�pM���G�x�gΊ�lC�I�P]*P:$��(l�Q���F&C�XC�I(X�l�B����,@v�C#r�C䉓d�\�6e�~��yI�N��z  C�	:Qʲ��1���;X��1f����B䉦 O��I�m�1o�� e.�(r��C䉮�9�ٖ,FX����*��C�I:	�J\����U|BܘV�ˀD��C�ɡ:�LQ�!.E��C��Q,B�	"6���I�0���J��T)&�0B�ɚ�Y��a-�<eJw*�g�8B�I+mQ�<�d�/S�+�Z��*B�	 %�B��T�,β=2��3!}>B�I4#��,Q�╤b���	GFCE�C�i68�B�͗�|��U��p9�C�	8 }�u��L�H8�Be@ $"7<B�	3".4�fIf(�x�ȸ�B�I�^��X%�@?f�ҩ���YB�	*p�,�!�Z0'��	v(2{6B��8��� ��~��i�Dd� �bB��5L9�	�Jε ���2!F�SGC�ɋWI�D3G)ԡI1R-�V0YC�I'�KB�P�Q"=�f C<jQ�B�%j�FIbG���	H=;m߅.�C�)� Z]�Dkީ`��h�M)M&��"O�q��),��U�m��e��"O��t�-����L%��a"O��q`̟�J���J&a�/}y�	�"O��+4C��A�2�u��4:4"O�����a�DH�%_�4&L�1�"O���h	!Q	8acN�P0��"O�Щvk�h֊�� �ޅB���3"OV�Ť�&��XaHʓo�T�Å"OƱ�5IZz{�z�a�>�-�e"O��Ⴇ�.c༤��/@�t���S"OD�� �+V���W���#�"O� �JߧP�P���j�v����"O���w ߫I<�@@�ju�!��"O���ɒ�'��`ڷ"?�>5��"O����6D�y`�Ļ� PS�"O��Pnقh�z��.�&zv�ҥ"O`���L,'�(t#&��Q=��"OR��F�خ�<HG�U�AM��7"O��뢇�+8v0���N�dKLћV"O�}Ӥ�ݝ��C��h2 �"O���3J�;��+"x>�ؤ"OTH�.0v�^��U X#dʬY�"O�E8��_5L��Х�6G��hk"O��Wː`�`�b�D�W��p*O�	ا�\.3/�|i��$5���'�xQ�B��#��s ,�1M� ��'�~�h�a�$0�j�%J7z�X��'G
�BD�@�Y{�����>3���
�'�b\;�+�� t��G_��FN*D������eB�x���sD�3�)D�|(Bd#���V3�����'D�ث%lĄ��JqG֋��M+r'D�Bv%9ap�K��ǄP��*a�&D�ٔβ.H>�`p�9s�hY�#&D�Xy���`x�l!#��X�t.#D���'/͏���c�Z^aP�K� D���%��aΘ�`R��0'��B��=D�l�Co"`��tr�ԙ}R�q�8D����7;�Ej���x�Ja���!D��ʦG.�iǥ�<9A�P9��"D����ȇ�3*�9�K��ON�t��M"D�ԙ�̖~Ӽ�3���J��(C+5D�8"�B�F����r�D�B��1`2D��%m�{��	z4b��\p��A�0D�0K��PP(�3.��k�pAӲH+D�|S�� �>9dph��Ѽecj	��"'D����E�)R�R�ksZ��3"D�44��de�p"�5���2n>D��I���G���i^.|B��S2D����$��۳ �,*��%���5D�\R$a�!`�
�ȶ(��s��� 6D�Ę@ B-:���M.� yy�1D�����=Ul�*��I��N��f<D��CE˒E*���m�>�&�5D�8�  E{'�TRD� :�)T�>D���$ңI�*����:Ґ.��C�ɶ:aн�ǃ5
�@�Xv��2L\C�I;_��B��'�P`���*]i<C䉱#�h��&H=M�
�QA�0��C�	:%�b���"߃������
�QE�C�ɪ*�d�9����+!/�}+�B�3��i�ŝ`��i� �6g�C�	�)�&(�w��B�j�VF�.Nr�C�)� Lx�2��>w�(�[Ŋ)����"O�X;���+M𨓹��\r�ɇ�p��Y�̯?4��6Eއ>����ȓ.(d2�!b���qχ�q<����z��" LI,�v}��$�8M�M�ȓe(��uk�j�����Q0E�Ը�ȓ�b�A,W�Xə�$ܓY�$��nX�)�X�g�A��,T�&����ȓ[Ny�r$؄>�f��G�4.�P؄ȓdG8dY���>�t����� ����V�J���刵���``�M��	��|�����)U ��pW
˴dd���m��Dq���O�M8w��8%{,!��"�&���p���8z�DX��L��c-��W�2�3�,��n0�H��Gy�P��B��E�rH2A�_�1��I�W�N:�B�����9�g"O1	s�J�$|XyW�P�2�J$��"O	s+V���tJ���K�,���"O��I��a�8][� ��:D��U"O��cB��>$mK��2YLT�"Ob��A�9<�6�j�o��B�b$"O��r��	k	B��W!F��nh�#"Op�P����6�����������"O��B��Y�~|Ĉ'@��j�֥��"Opy��n�EAՒoy���"O�DiT�Ӓ4�%)�,7h�<�"O�1��
�,������`�]��"O�]QkP(+��a�!}>��ؖ"O�i*D��i��2�o�E����"Oz��ĤŕI9�U�o)V��Q0"O��CT��:���t�Tz��p!"OP�ZU
��(��Ms�.�/>h%C�"O�
"�$eJVxG�ǢB7�ex"Ot}J�-Ȑ�$0׭��� ��"OKێyK�x)a
�}�#ʕ+�PyBEE�bp� CDΖ¤�h�cVt�<y�H�7Kt�H#�+ڒ&J�]�hC�qM��AT�Z�`�pw��h�6C�Ɋn��Ty0��;Y�>���ɍo�(C�	S��4He����� �A�C�I�~�z����^ODK3�8�C��9`M�'��9��#��J���C�	>}�HD9���]��y
'AI".JB䉙C���8�/ǥK�Q�G�4� B�	��&I)@M^��9�/�j�B�	�Ԧ�-/f�\	��C7:
U�'���K���W�H�3]����'`pH��>�N�i�/�9r�'�̴���ԟU9�e�`NU)2cp��'!T��	�������#XF�6"O��t�]/m�����̝�Y�X�"O�*�!l�!iUi� :1*���"O�����&r�6����^+_�����"O��1t�F>k1Ru:��JT("Oz5�qÉ W�b<
6�/K,)`"O�D�k�u<FmQΞ"��ɛ�"OIPD�20�1O��V��(�"O���qQ ��)%/�|ު�K'"Opua��nJ�'.N:X�`��*O^��*,�^0��F`��1�'��MS�c[0�}E%+d���Y	�'�p�H�#�!r�0б�݆\#�E��'u4m��%6Vh��4��+!i �3��� ����`5R�Qs��+ƾ��"O��r�חS�*�����
��hk"O޼��ÐUH�k�&��W"T�H�"OB�A�M*{��12�L�!��@"O}
�R�Pሶ'A�fU�1"O�Y�,��1���*h�,\ݦ1G"O�(y�`]�u�%;4F��=��qj"OrQ��e�> K�۞Qɬ���"Oxt�`g����ij�cT�J���Bg"O�Tk�C��%F.���� Ͱ�"OhP�釹=�(� b���%q����"O�)He&��_0�R���yj����"O��ЭS:Y�^%Rw�W^��w"O"T��"ަ-��
��A��"O-�w�ʏ`s\�(��J$6F���"OԴ(��9��1s`�`+�1��"O"Ҕ�]�e>H�˕U��ӣ"O�=Cn�.AX�ZsgI�b��T"O��9��Q��(	1G�)z��%9e"Oı˕gɸr9h-���l�Ltx�"O���$�&�xY�� �8��""O�P�ˎ	+#p��E�G�C����"Od�a��B���f�w�t���"OԴ�riI�.��A�E�#�B��yB�,���'H�(����&��ybM�xk��ơ�b�TA�9�y��ٮ�����փn���r����y⢅>ʥ `�d�4� ���2�y��|�T���H5x�(�4�D�y���v$��Ѣ�@/ OT)�D^��y���''bt1���p����i��y�K�$vn���@1=Hx����"�y���Ji��B��/��-��Y��y"�m�d��5�E�&����C�E��yh�1�)�߬o9z-���:,�!��ȅ������'b5���-�&|�!�ě=[F4�,�-(xtC��4v!��W,$H�zG�� g�4� K��MT!��E��B�LJ�;��ap��$"!�DY05`�9#�/�~ ���M��!򤋀��z8v�qW�ہB�!�P��dܫR!�-:n��uh��_�!�$Āv���z86�;f��!�!�ƅ2���Ӧ�^�K��b�Ѕ<�!�J�|�Xث�I5n<����e�!��1�TR����\ ��˩D;!�Ă�Q�2ђ���, ĥI6��^�!���3�l��aO9�P�3���.9�!��܅�Ѻ��	}���$|�!�d�k?�8�(��{$`6�C)6�!򤜯z�@t��CZ�\�e��/>$!��<|���C,P�R�.}0�! )!���Z�<X�B7q���D@%"A!�M�~�<uy�L�7ٰm)�A+f>!�ٱH��ب�bJ�8��'�A�!���4>܌d+V����e\&FF!�D��W�12�E�VȀ����nJ!�Ԕ48bԺ4�ߨs�u{p�`�!�dâp���0eX���ve��m6!�%�����I�/L<\yq��#!��Z�s^P·��)y�Θ[��]�!�E�M@4��D�~��3U�A�4d!�$�6[�|�sf^�2�Hы�-�!98!�F�k����(�;A~��⋛!!�� ��0)�	Q�
 9s�/.��tY�"O0	�]�Jd���D��-��"Of��#U�z��0��/.�p9y"OnE��J�;|ܼ|�d	D�Tv��G"Ot��@���T_dղD.��1i���"O��P���-�t�
"'�i�؂`"OF�q��X�;����u.
ET�t"O�у�B�'��!��fW�3&���"O09f�%�^)�u���OB��"O�t�Ư��g���o��D�g"O@��«ц2H�xy7��9Q�̰ha"O��p �/?ԙ�hλY�Ȅ�e"O�JT��)�e��	1Vt	��"O�����	�So|M3�,8z���"OJ���AE N쒕	�a�%��("O�bf��Z{�����A��"O,�0�W�B�pu����.NZ�( "O��˂oJ�>mJ9*�̟�z+N�Ae"O޴15#T�x�����l�
>(���"O�Iz�$G^�x���7J��Se"OhA��b޴A������
�"O���RI��sG���Р��-ȘP��"OP�:�.�8L׶�ْcB�)B"O�Вr�͏?���D���%�ڕ�y�J�<��uxBc.h
���s���yR�UYZy�1&L�\�h5���^��yR�'bƌٻ�f�!M�聪3����yrI7>^�Є�_L@��qT����yR��V�j��.	�z<~,�Sh��y�N˨��M��Fѷs�"�K���#�y2��I���7B�m]�����A��y"iʥz��\2��fx��8��,�y��YQ���p���R�3�yr+��Bز*vCU	H���I̗�yBgų
b��� ��K�1J�"��y2�ޯy&(Y4��7�E�����y���V��P����2���`���yrݔ?�VPV��(^~���E�y2K�.Z����:�p�p$��ybiIʚ���i#��M5�C䉸I��B��'2 ;���=b[�B�I���Ҥ;aP$�%��'Bb�IV�)D��&�,y	L�`7�ݺ2� `h'D�HiGn�U��i@�%Q �}[p�$D��R�'�F�D��=Z �)?D��Pwi1Yʽ4e�+p"�:��2D�p�� �E*P	;�*!i�m�׮.D�0Bqoȑ]����q��e(t�Y`�2D��I!n�2'�� 7C0�`���2D��R疍Fb��E�Kg�1�//D�����H79,���
l6���f�,D��8��"�C�/ף'ڲ�Cg�,D�s�*O�K��1+%V�^3����b+D������1=��13N�)fn-[��=D�tb @�j�#j�$Y����o/�B�	0y`]9pLDA@6���{ھB�1m�HZUd�]Z>��DӑY�B䉀~���	"�(w%&��P���Tr�B�I�'��|�W-�� 	�A	e�B�I�|��t���޵ �*x�5��+�xB�I�|�F���Q�.u8�@��+�zB�	ʦX⡀'_�p����C�	!A������)�6h�o��4��B䉿`�bv��&=��Lõ�IL�xB�)� �1!��a*Z����܍Kb�2�"O� q%�>;9FRƞ�;��9"OD-�E��)�~���Ɗ��~�8V"Oƙ+��ùJr*Ts`%��X�P(�"O�yY&�XK=�ٸ�A�5Ȃ��"Orq��I��HJ�I�"��Y�!���]&�=1�%̶)��l��*ݩE�!�$����P�$�ds� 	�>�!�d�-I+�(8�e��P�y�D]� a!�� ��;�N� X�^��#\!��9�2� E�
#��*�<�!�Z,B��U��/_m'R0����F~!�$E�0tQ���"y��r7G%9b!�D���rPC�!D ���%�rB!�ɘ`2uKe*�#��k E�%4!�d�9LBpu�Ek���f
 (!�R j�[�b�(t<���$�!�.���qJ�Yo�]3��J�!�d��)��5�`�E�U��\@�m�#�!�$O�S|x�� "d������\�R	!�dԾ/e� �%♓ń����L�!� ������>j�B	���]=L�!�Ď �Ya��&�@��w�9V�!�D�'Myb����Ðw�*�!EAB22!��_4�vy�񀙵��=`�^U!��E�,_>�HF	�4����΄�B!�D�s��hA�pX-#g�k+�!�$L�*74�`�D\�2>�`JsM'.�!���a�R �I��0/�2�+ �!�XY����_0Z)fJ@)��N�!�D�O���j��8I�rL��?�!򤌍P��8 #�߈n�
t2���l5!�$݌D{j���o��]� 朔>0!���!Z7g�zؐ	�5��=�zC�	���h铤Q[���?bC䉂�P�pqͅ!̄A)�ǢL;B�I	R8p�Y�%�4Ό\*Y��n+D�D(�d]?>�D(�aE t��:��'D�X�&��w(d����O/���� D���
45C��r
 �-���P��!D�\�լ�>�Dq��	\��*�*D��3P��.��5�c�؉I��ez�)D�hh���7}[H$�!��>���KC�*D��ٶC�,9B��(��h(`(�D)D��°��.��iH��T*&ھ-��:D�HyD��h�d#
E�%�B-3D�p�b-��/���)��ұ1��}�6�4D�(ӗ���< ��9��%I$N�(FE D��y�Jű*D�r`޳>���s�8D�ԘŃY!f���b���Po�E��/:D���Ͳ+�"px�#���DBe*;D��cI�!Z\!���Vv��Ca9D� ��&V��Nhy�E�N7^�R��1D��UΖҠ�[�Þ=��h��4D�PR61�`���}ߠ���0D��z���l�2�P��@�g�8�Z��,D��#��;������=���*Oν�mI��
��ŧ�x��w"O��Z�+O����O�?�NA��"O:QA�/�g<����2� �"O� �3�.BD���B9d�t,	6"O%���rD@Z��	8� �r�"O��Q�ьC�:]��#w�JY*�"OX�UFC^P�����s�zy	�"O� D "],<�48w 7�\Pr�"OfI����2�)�π@�d�a"OҘ�!rv��"��h��	�"O"����C�_� a�ASzQ��"O�����>�a��ԇL[��IU�I�DÜ9+u���'_�tS?��ׄѢQ^L�r�
R1�h�a�b��=B���?)��rCf��6dmD���VEfh!��6Ty0�?E��|*%#
�5�K�ɊWl�)�@Ѹiڕ��C֒k�L��O��y�'�)B$M@-�L�jH���ʥ?tҥ`�4�mZ���O�,�*��:`�
�iI�{�pA��)�O^�b>e%�t��b�^?�0�1dάҵ�2k �O�il��M�޴Y�2LѰH�":I���F��/�N���sq�-�S��6�?A�����@������O,7m\�n(D����8XNX��L��_^�ኔ��S�u��c���d��F��3\F�E[u^M�t�O�klѹ0|�TYh���8a�W�'X�&��'�m�1���� c��G�s*T��P%*M�8!�~�1d�����C	!=�T��ɔTE��l�Q�\���O@�����i���I/�G��5I��W�r�'QB�'M\��`$�D��1��9A�zY��d���M�аi��'�����!��� ��ځhQ=hss$�۟���3f�ݑf����ן|���u��'9�fS.L�Dm��ȝ=5D��%&��O4�YS�J����Jb`XhH�f$�FM��O�5h�'n <�A��t�A$�Η���( ϣH8Z|�"�֜b�8s����)�U��j�ϙD����BL�a@�YY
�e#J�;���Z����b�L<a�/7��>�ƤG)7(PH�鎾M�ekW,Io(<�۴N�8pSk�'���E�0	�D�4�d���nZs�i>��S~y��ݬX�(p��E0d�����+:G���P���[Pr�'���'��x���'�r�'�H)6}%> ����B�vI�C�`p�ɳN:�l�GN�8>�� F�ͅ�(O\�����#ˮ} �����H����:X�xE�W+��,�����l�>ՠ����(O�t	��'Z�,0"hڠB-h1ؔ�N>}���kpk@$#�7��O�ʓ�?��*�d)�^9qd,�Ѕ�J�P
��"O�D0�4 �9�B��'�NܨRkJ��t�شwV�fY��aЀZ��M;��?A��n	�D�8�J�{RN^Q�V%���Ɗ@$���	��@�	�n�	Eg�$-�
�r��S�c����7��tKҬ&ں\����5L@�<��D� �d��|"%�W�L�fE��*�6�< S�� Y�rݠe�c�0PP)�Q��ZZR�4C�x�g�5�?I��i����6-<?������Qu��joM�OUR���v�S�t�dR@�4���A<�>}Kt�ϰa9��hO�	����4�MC��M�A*�-R�D ��d�M?�� �2M����'�Z>�h5�Ɵ��	������
�K9B� ҋU�	~ ��d�/ �z�����X5�c��'�pJ�qP�	*���)`���Q�R �B�2�nƸ{T�<���pӐ�C�$��dF4i!��SQl�o��}�� r����U�4ř�)"�	n�1�b�i��8C��cF�fO�<��X��MK��'���U�tހ$B�d?����D.�S�Ĩ@|"�HDOV6ƬD�֣+�(O��nZ�M�H>��'�uwC�z��$�N�
H����J��07��O���čo� 8  �   3   Ĵ���	��Z��t)	�y�����@}"�ײK*<ac�ʄ��	ڤ´�xbjR�7퉧H�8*fe�_R�l*e�	[�R����&cQ����Ŧ%����u�.R����g�6w>t�r��O`a(3�C�r@<�f���c;	����!Vvyr��(��؀f>}j
/#(�QR�aͼ芝�[3.���%^c�\9�'\��a���;�)�-OX���BA�a^�|�d_�й��6E�N�ː���Q�_vX�dY����L�j 
u��s�	C�~��b�"w_b�
�,�	�	�i
c�F r�'F�y��`����'�t�4Y��pzTT��h��/s�2���J�6�!/��?�6�ō��=���d�(8Ԣ�OT�K��x��XB�P�����ƒ�Y���{%�,|
كG�'�
�Ĝ�
�8�PP>�I/����
�`��1.Y�Z�@�0�4	�O� ��,AB�'���[��0iA��_E@�hҬ]?m袔��%� I)�I�>iJ�S)�DK -�F����|��VY6z�C�>|�hqN̚:̄˓D�g�I"f�n�C�d��L�'�%��cܟ�q$�X�'��}+6���F���ր|�:]ϓB@�3�>	30�l�����w���P�@@,AI�k��hqI�֋,S/j8y��2�>*x��(+��.S¤0ۓ  ]�e�͊�K��UXs}�D�ҟ�y�Fƥ.��	��?�����:�T��p�,�7+�Pa��؟Y��$A��O�d�E앃���şy�L,p��O0���M$a�![�!j�ݲ��]#i����O�@�O>�N<Y"�r���סU�
sT�������s����g�)L`����nX�}Q�QR��'��t³U>p2픊dL���A�'J�=���E~r$� ���N>���*��i'�\���%9����R�@�d`v��>FBl�"�d��X�,,ڃ���5g�T��d	".�8�IO�p����5�7D�,��   �PyR�-W$���M�	����S*�?�y2���E���1: �TÐ�ܒ�yrN��O��a��%x���3@I��y2�@?`���x3eG\���;��5�~B�'O��)ǡ�}Bq@�fי=�̌�'�,��!�T�5Wh����+ ��L�'�@�RE��/Hsh��C�%�1��'�V�����t���Q��'9H���'1���	�єa�W$�P   �  �  U"  6-  �7  �A  	H  MN  �T  C_  �j  �s  4z  z�  ��  ��  @�  ��  ��   `� u�	����Zv)C�'ll\�0"Kz+��D:}"a�ئ�pgm�|"��f��Aj�
��EE`	�l<�b���^�Ma�Α�61z`��V�p�*�i����s�� �:@�S����a��rձ�/ԻE�����96@|�`k��7�4X�nJ^�b��W�(/��.�'"���O��
�+#��t(�����,d)0)�)�D\�y�$zS��)}l�dm�<}�tq��ߟ(�	ٟ �I3�8Cc���,���%l��������.]R�,E�'�ҏ�Z��'��s
��4���P��D�4�r�����L�' R�'�����M���{7�]�E��ȥ*Z�t0)��X�*F��Q��Qɟ�A�h��DI�l��Nb���p�� Z&�tȑ��hb
�(wn��]@D�'���%�I�hj
�!���Urt���$.�J�й25+�).�nI�e�O����O�nZӟ��	՟X��V��7���3qNΨ.g\9��`�s�9�1�'j 6�DϦ)ߴy}���'��6-�`YT@n�B�ṯa��-G�\ط�Y� ��5�ӄ��l��P���*#S,�S��
 N��aR�j��lz�y07������P� ��:�8!��ď��z"j�I&�a��H¦��ش"��v�Oc�i�Wfy�2LZ���Á�.p����MvH�%f�5�@�E#� �1aعU����+Q+
|^6�N��޴O��\�G��w�n���j1�`Є���V��t�i�\7M�����ꏖa�`���cD�W��H�� ��y�6���L*b)��̨Gg*�WnMZ�0�G���M[�i��7���k"@�H�xh�=�ta��Ph9�-�B,��0��'�)S���֦%p����P�|�8�e%DЂ�Z���?� .I�>V���`iZo��亶l�(�hb��,�?���[ʛF�O����h9�j��
�ҋF&���)gp�:v	��\���'��P��'���'��\��'�V]BP��y��Eɂ�Q�����dNG7e ���P������GV��r� ��6��;����ϐl;�)�n�Ulm��B-O�h�1Y��-Op�J�1;kK�'ub�Ұc�9�?����?iN>q��?�/O����vhicQ��1zt4��ߴFf����O��XpN�SQ��Oz�IW��瓯�?a��EML�{�j�<Pb (��ɟh�'���AA�h�T��"��ʼ���ST�=	d)�4(�y��̈ß����i��Ԃ�甏�F���4���������F��}�tB�
n�n]�E���a���%���Ů۞L����/��?��㒋q�ӃUM�H�f�+GvX�q�շ+Y��U���	�M���|*%�C*lz���g�@�8*�)�^����	ݟ��'�1�������sr&��"
�z��E�V��ğ�ش���'�p7�`>��VG��#���y0����� �릝�IyyRG��0��d�'���'d��:O��1{N�KB@#PfP�x�&M�m*%� ��CA4+�y�WlO��ϸ'���aa�+G(�M脅	2,����@�F.�5��$�Nd�T�n�/�|x�RS>)(a�ǣRp�]�=0di�m_�E�A��B��s-بn��򤚬�B�O�3�d�
ƌi*��[�:s�/C�I���d�O���?9��L��9i�v�,A�풖b(8�fC�O*�$Ԧ}�4���|��'����D�p2F��U�ʕA��A�qA2]�$J[9�$�O��$�O��	���'��B�1֬A6�M�Q�(��	���Ї��d�X�	�)z����$H�]厁;qf��A���0�A��>���hT"#	F��B�ж3s��)�Ȟ�?���Rd��v�Y�� ��q��A;�INb}�d�䦩ȍ�&�\�u$��x�r�������	nyB�'WҐ��{B
�P�=1��U���rj�8�?	�i��~Ӧ�l�f���8#��7��Ol�dӏb�ă�(N�#x�Yq���,> ���O�-�Q��O��$�O��`ΐ�)UN��RɠJ2e�]cX��:f@.>�%�'+@��j��Ób���+�/ot�t�6-� ����g�K�RaGoa�B�8���z_�l�����B�z�M>���	����ɷ�M{��ӂ�3բщL����*ў$.>ٹ/O�z+�Od�O��9���9����D4�lٲFdG:]?���D{�O�7m�O���D�8z��Hk�"b
�l�����4H�Y�1�iU�P�S�?%�	�Tl�A���u�#�a�o����I쟨i���F}$�����M�Fj����O�V�ʖe�.G֩z�Y�j
x������f(�.K�`X���˱c����c�#U�Z���~��F݈z��)@�ұ|����N~����?�ǹi;4��c>Us�MX" }A;��E���1�'!�D�O�OP#<�0
�dE^��ǯ��H��@�F�'B�f���oC�	5�&�Bp���1���O)N1�iX۴�?i���?�F��#d� y���?!���?!�w@h����T%!��uKֽ����S�l��Q:�� ¼m���Td�D�ϸ'����N�cn��B�ɫ�K�R�R���3 �����LP&wu:�(�_>]sa�O(r��]�,�U�Ǝ) \�#���G� mZ�#��	<s�f��-��O����Ov�cpk�>@$
tp@�@:�K*E�
�O��)LO<�Hs�WÌ�p�o�3I��w�'qR�zӒnџ�i�4�?��'�z(�lȣ�#�4f�e���Q)lx�mY�m �\8�I�O����O�������?!�O�h�A�V�(����yT�=�C*�x2,[:��'tG��{t�պH�\h��i<1E�ش~Uji���,+�Kfφm�u�I2��?ٶ,	^@	�m�j&�ԉa�Tc�<!�·�C��Kb.��j����	�F�I$�M�I>�U�G+��ӟd�%�A1�5Y�O�m���ȠH�ߟX�I��n���Ο|̧hR�8�R^�^y�CΛj��� ��I�D���J%.��K�'!�����86j�Q2S�L :$I!�yX툰o)/�t<2�j��r#�u���I�W; �D�O��02�8�KƾFy�@��&��'��IP��D���D�d�H|��<y���1�=�	V�����O�`�H�7r�)��BD ߮M��'Y��d$�<�	`��}a��i��hP��D��[�t��>`�K���?1e�J�l��a{U�#T�� D���gɨ� 6*�e�I �=��c��PoH\�a@�Όz��I5+�B��b�	�������B솨���bH	��I[�?q�t-��v�^̋���8$����p�2?�'O�ğ$�	i�O���[�?��P!k� [&�Q�ւd!��ݢb�<вBJ P%��@D�S�-aў|�	��HO֥`3�C�����s����5lRP6M�On���O<�zrW&�&��O����O��"t��Ӡ�H�J������*��e��4���M�pP]�K�q����?���#FÔ	E�@��]7��	�#Ӧ
� S��
�+��V?rc>AJ#*�gZ��a�b���j?�:��'=P�rd�X���V���� �<)��w�4�gj�9��� �[�Qzh}��2�'�B!��bR�v��s�Δ'er����?��in�7�9������)�<�A���v�	�kj�Jp��[�W�\	����?���?�����n�O���j>u
��I�T<28A�a�ƥ��m�58e3�%G�l�"pr���S*]@�r@JN V7h\H3+`��TsnJ".�8�c�EʍK�0B�l�(�@�=9ш�2z�J
���w�bQ�O�6x
��	��?�T�#?�� ���	2�2�´��O����<I��O-�q��%P:^�L���eN򉅡MsM>)E�0B�F�'��
!�R]��
�@���{�k��BF��'�zEi��'�b2���� �׈V�4� ,ڦuA� m��:�� ���6�00 �3O��J_�u�Q�H �/�<9�t1��}��ܚ۴r���3k��4ܢAp�-޿!b�< �&��
ܚ�<�����`�M>9'䆶|��1�0o˧e������]z�<�4��-k!�E�����:V�$3���u����,�t���$W:p)p�$���#�f�$���Q�7�M��?1-��̸�+�O�9�D�J��AU�AL~Q;n�O����*����7�|�O�}xCВ_��V���E�@��$`�+*�S�OD��� )E$8�lE	1"��p�2#�O�ɊB�'�D�O>���)(X;�q	ì�<!����5D�TcWB�_�B(0�$.~��i��"1��n��>�+�	N�@��D8U靫X���	W������	ߟ�����p�i��?i���?���yG���=\� c��: �Ш�-��r �����!�3�4������+�uw�O�*t,��}� ���˅bj��x��S3w�Aضn����,H��A32a[��PD��O*�8���w.�����k��!y�E�����|���?ɉ��y�c�+T�TE���:oz���	��yBM��j�c��2]�.�r-+�?q��)�����n��3{�0C�@�?��!0��2g�L��0!ʿd���	џ��	̟IZw���'��i�'ތ��H2���gӷ`D�B�� 3wtBD�r�F�9)�բ��H���0���A�W��*u�x����ͪ(��QHJ�k�+W���SRă�,V\Y�W���Bɮ��x�/%`Y�5��l3P�U��t[�i{���R�-9���ڣ��@����L���=��yfS}���Ю�1~�|0#�K���W�v�|b��G�6��O��W�(�<5�����me*ȳ���A]����OF8����O^�du>)�u戣J8�LP畅w}�Q�]2^L�y �L�8��i� �O�ް�� 0�Q�y +@�(�$�q#��	{���"Ӵ:�B����r�����$�hƀ�0��MQ� ��G�O��%�<�� Т%�&hC,E>>��&*D�xS�lT�^"~$(�.�62-��4�O���	
n <i���F�Vd�瀐�V�O:= ��ߦ��Iʟ��O8�	�'�$c��Ճ4Ȭ�AwdX�|0���'��-RB#��QKI
jaX��(٘��St��� �c+�9yqϋ3E�����H,����!���	�
hb�j�NR0�rF�)b���&f�bh�iU�4Q�JM�(��Đ�t"���OT\&�"|ZcGj�ĉS�#|E�b*��<17.;o��]H$#F!�8�A�'�2!$�vHh�,�}�tHs�C
=�%+�Q�x��՟�1եݙcJ����ʟ$��ݟ�λ;܊ؒ��Ͱ%�f�	3��!k�0���*�-Oc�@r�ψ#tIڶ�p�$�OxFD�fN��~��k4V�H��%_��@P��E��(�E�ȖD>��
ɁNw��������I�1��=��fF��BP"�� Y��Z �q�޴l՟4HFm����|�'8�)�/"#FU҈6NlH8F�%/��'�a~�l�TY�`ƀ1"*���4�?1��C�Lgӂ��]����?�Sk����p�LY�!�r���&~}
-��	��'���'��Ɵ����|�Fnx��HB�g70!�rnÎM.�)I�n���ص���h��.Fn�� J��7��Z/Ryy�$\�B�ǧ��};����G����3@|� ��E�yZ��O�,n��ci�1�6�H 1o̡p��˵,-��O��=�����(m8|���Xi��%��)i�{���.6g؅(�M
/Mƍ��1SK�'�86-�O6�!�`��Q?��	�Z�2�GӞS,�F��&/lX��I�\۴gӟ\�	�|���/zv��E�=X��M�:'HN��K�'Z��x���Q�6X�(�9�T�ACY�tʴ(`6h��>:ZHS�#��2G�] v��1��,��EP)|:\�>C$̟��I^~2�D(|�֌-7]�� �1K)���0>����4��uW�o��`�
�X��tb��BHh,
�����ĕ�7��*k����dy(��7M�Of���|�a�?�?ل �f�� S���+rx���e���?i�8��X��A�}?�q�B�>p~>D�+�(�D�p�4��E���C#ڜE�'Fh�ñ��qV�!"sE�(�������({\�P�e�2x�DE-����3��Thh������F?����h���ɱ1�pJ�ƶ]��y�FO3(�C��
,�8��ӏҡ	�Xq��FQ(f' �=���1ܑ�p����\���	�*({��Dj�-�M3���?	�G�^�(g�D�?���?����ywn��Zwҽ�b�Bz:�� {� ��Г7�(D�<7��pɌ��yB�*X��[&�E&I���C��vr*�+�n9CC���D��{=�+ׇ���:4��I��Lp�	:�NY�@z� ��g�ez��c�O��
����O��=Q��¡"����"�!����I���y"E�|5�y6��w��P��6�?������Sß�'X�UJ�тp�\iE�[?i�鉆D���aG�'���'��Ǳ~���?��ʇ9�fd@,	�>,�4�Ɵ{�J�p�o��:�v����+2%P�q�I��0шd���	�◿I�y@���d���3�ǕB���G	>ړxP�!���x�f1��IS�M킡���p���iݛ6�'��	�?Q�?��k�1H�|��Q�X
���$$���y
�B��͠��,0�q3f�V���F7�v(uӮ˓+` �z��?�;_Ke��˛E���@7�[;����?9!KR�?��������'��uPT�v܉����<˄I0��M��K+'���`$�
j�'���I��Ӭ(���{A/	V�H���Q�-�Ry8c�͋̠m�J�)yG}�K��?�����D���D�N�).(�JLM�'(a|�Z�8�X���S��X�噗��?��'�~Tȡ�U&�v��7��8�y����$�����O��|��S��?��d�:Z�@��ܣ!�$�I��(�?���3�Sa�ϒs?��PB� �A���|B̟���hS��8�k���)j�(����0K��N(d���;�#F�~@i{a�;s
q�:]�M�&eи!�����T�< 
r��l[�m�O*��<ڧ�yM��Y��$��R&���F�yb�H�M���G4|d��'��O��F�D���[���᠊,z¼��"�$�?���?���V �T�Eғ�?a��?���y7�߈1�Vp�p��(��-X��:^���M	��j9k�K!�� ����L�_��|�F8A���vbZ�D�L5,�խ�4h�� ���68(���󩟶��I38~����K�3עh�#@�f��d'?�"�ɟ���C�'	{V��r�I�����/�|�҂"O򡢐k�,Cb�Y̅�!��D�sR��r��4����<1�!Ȏ�~����O�F`؍q������U)���?����?i������?��O�4��SeJ:2����'�3���'��:z$[@/ͽJ��0�(@�9	uD}�FJ/1��<����n6�=�*�/7�욠���7h>����#�M�R�w�'��B�h}y�BߎLB8�%W��?����hO�"<�Á��.�*c\V�Y�v�u�<�#�F�yi4X��
�<�P'��t�I��M3�����bŊ'?����@ u$�Rs˛ 1�M�o�O*��� ���$�Ov�S��y��!�����[G6
0@d�΁g� =�j�9��0�Ys���剏g��yԈ
)�
�ąUI���wA	�B*���-H�C
6�A�㣄:�(OD�#��'����T{�<	 ����S�ob��3�D3�OP����� 5]�R)L'�i)��'����_73#TH�H7pXf-[��6o�S��j��R�M+��?�.�N�Ձ�ORl�"��<<���V�JC����O��$��ZId�H�'ش&+�oK<e�O���/F���MY\mط˛�G�n�q�j(۰-�-f�ja��Gϲ�RE*֎0��s�B1��`� ����U>r�H%�'^i���ɧ�&AZ�BZ�B\x��)��!� 8Jd"O�GIT^��[!�>MȐ�H��	ʟ���O�8~�� ˂q�H1Ƞ���8�$XE��!�0��O6�D�O��$>:�� �2i�����"��Eh�(��#���"���-DG
 2��V��c>�Q!n��a��$I�~��T�&5�,�bl�]�^����=aҀړa��&��<���9���지 �L0�h�)'��� ��/:�(zP�'����^tP���O�=Y�A�(ɛk��@��r�,9�y"�ǥ~G�|9�I�3u�L"��G����Y���t�'�	#�\���^�3z�Z� �4-�¡M�k
�=�	����Ɵ��Zw��'�I �R<s��R�Q��r/ŘW�1k�
�4 �╣S��3 ��,l�(Q������i�9��b�S	��B��C�6U�!:���9%d��0���'��+شv���pTB!ʓD!�+1�ӘP�"	�,
C�d峄�������q�d�Q'�<�"@�<Ÿ(��+����&gb�AP�)�\ '���ߴ��=�$�G�i72�'�!c-C�^T����ʆc,�Pۂ�'���Q4}�b�'��ɋ�h��t��QCP6-ڮ ��y"(�9�j1{�k����:��4OB�	�ًv: ���1��Q�	�,�ji�W!�7A�!iw���q�R��Q�8ړ`��E�����!�Jtش)� ���H�k@. ܭ��(%��%��3�u��f�,e�e�?���4�L��ɁA�y����Zd02�i��	<�O���j�O��?}��'Fݟx{�S5-
aZ����Wm�X ��ݟ��	�=W��6�Kq�Y�S4-l�!rb��c"�O5�Lp�Ǎ�B�b)��l����O4y���T�Y��C `ˍ	��h�V�շABq�K?AS"��9%��&8@̈]�e�)?q���ş���_�OK�$�'�����w�d�f�-jU!򤚧.C1�f�_ Pf�����چ�џ�ʋ�)�B5�7d
t�Qa�aK�v���'Z剅� ���Qğ\������|r�+H�|L�Q��,\,�Lj��9T������1J�j��e�t,�|B7�>QǨ�ɰf�f�[�k�>
 ��ѽX1�jK %��pI����0$Ń��-�ӕ~�a��O�mh��^c_�s� ^����4�'y��=%.��$�O��=Y����JTE�{�v��B�y���=Xգ�H�e�^��`Z)��d�\�����'���R�݉�!#k�͢q��vp�EO� �
-�	�<�Iϟ��H|r�O�6�b�̘-rez�Jt��i��ɚ�d!4���"f#�s�
q8�N׵"Z�.t�'���z%��2v��mz�dBh����@�љ*���b�j�&E�()����ĝ�!odӌݢf�L�I=�4q*��^�*! 2�W�oN ����O��lZ�M��R�$��zn�!���ȳ0lP-����.BN���2�		y�%�i�ik��@��\�$�O���O�˓�b��d]?���H�H���ip��Ae�
���M��ş,���ݟ<���|�TF�vu�dpfm��4����큙qт�@"��2�,��/�s��y��C+z��p�CB7&S��b�Ѩ G�[�$�8xL��b�����E+W1q%�A�����F�%�d���Oz��'?1C��30� ���L71&(�O����)n�Z(�7���Ҹyn[�n��O��=ͧ7���%_��Q�X����H.�?�*O�U�q�㦡��ݟ��Oܔ����'@���.`aV���x�����'��ݑITp�&��75��%��	�Z��D$ڠO���*���CƣO�ll�h�ǀهW���� t��Ũ<�ڹJ���NȒ,�p�A���0�cl�|�,�9d���`Ûf.�bŁ�k~�����?��|��)ޕ2BjlZ1%(S�t�hŕ�}�!���|:)U/`�FD�u$5I�ў��I��HO�""c��.�(i	!�;i��=ڐ/V����t�Ƀ~������x��ϟ|�I���B�:(PL�K�-������h6�<���&g�) �@�V��|2K>���A(
!��a@ f�2 3��h� �a���Z̴y'�+#� �|ZL>15�L1B����I'Y��B���Z{� �IJ�g̓�za�gL�V��]ԈK6C��a�ȓi�����,&n� g/ql@��'O�#=�'��If`9k�/�
U�t�	�j�#CH���R)�6zT� ���?1��?��	Z�YZk�X.,-h�ڣn�����Q�De��d���H�oZ�+�j���剈o��i@��5��m[�k
t)�����j������rߦ ܴG� A��+�O.5�%�xB'W�>�ty:BiB((`�A(�0~�Δ
��g��6m.��OM`�F��Ҕ#S"[�hP&"O�5��!ć]��Ӵ,�>�`mQP�|B�pӈ�$�<	�������'����G�`([�$ױ@iq��=��'q��bD�'�r<��:T��0Vz�����\��vIїK����r#!�D�f�הs���
��V1�(O�bc�1���k4���H�E�R�E�E�ЀZt'�1"�@��T���G;�\YT)���M{��2扁e�����L���Å[(`8)�dKt|B�,ZT�ٜl���f!�@V�|F{�OԢ���' �D{�+$Mze�G),^��'����'c�����O��'Tܶ����N����)6$I��о;�$H��?!a��/{��m� I�'qrZ��5.ު���.r@앗j��E�W�G�"2	���Q~KєrE��Pq�M `J����]/���U�!f��Љ��g��.������3#G�OLe'�"|� ��)��Y����6�<m`Q�!"O��[iֺ!��}�%�"wY�����h���91�9{��8�DT�]mn|k6%wӤ�O6,Kf�*����O^�d�O��Nڗx�0��t�U.UB|�C6�Y�|�b刦/ϕ}$Z5޴g�4h��h�w̧P�4Т�����q� �1��DHGF�H.d��n�wG �X��J��M���Y�F!꣋&��~G�Q����1PE�� ��iV�Vg74��Pk�Ǧ� (O�4���'��d�?�OzuQ�%�6fh�A�2��OPX)p�f:D��"`B�Z��Ӿx� ����<���i>q�	qy�
*[��"u�T� ��kv)Q�/�|8�O�T�"�'�b�'Tzם� ���|ڃ�	e1�ɩ�ωnj����'��H5�Z�Yj�5`G/�5������� �ơ�A��dۦ�K�2�P��q�ZW<Ĩ�K�/Yɺ �)X��OL���-��u FÃ\K��Xf*��\�R|��%Dz��	�9�`��K�� � ��d�nC䉂p��q�n��H�gJ�)�`�&����4�?�/O"��E�ߦ9��埠��@]$�����Q،�!�%����4l@V��Iߟ�Χ<�����bA�b�(ap��0<n<�(ϼ$�x��N��mY����냢|���L*ʓ3�|X �H��Y<�!�mλ|���e��-N�z�a�nD��{�.Wh�z�7iJ����<�wi�ڟ(�I>!�з'F�j�E�K*6h��Fa�<)��ڏIGLccN��8֊ݛQH�_���hO�	���(�o�0!@����(m�A�$A1�$�	�Am�Z�"|Z�O2Z�a�Ǟ<d��8��K�a�t���OBD�g�8��i(�AI~D0��IXt?Э�,%��q��
�z��	1|q&=r�똗���ӨI�/iQ>��c��m��S
7�8�� �Fh��&&�Ŧ�#��l>Et��*�bPp
8(�X��.D�dP��Y-vsX��2#]�}�2�S��6��J�>]�Q-�>*A�C ݜg{��E(��y#��\vy����E��3�?�\`;4I��@��(ƠL�y0M�<4&AE��8q�iIt�4D���L��`0��%(� ���H�u �)���j�2��t��^ƨ�O<���'N1�1O�@��ɃJđ��+�5
���`"O�bB���H咐���^\E��W�h����ә0u �Q�R,\�L���,@'�a
c�#ya�$N�i2�(r!�8�0�g-�O�ȈFC�F�N���d�$dH)~@�ti�@�G�&��SvO����O��d�<����&�0n>�`��~�ؑ� �ә/��,K���(�����I�cI�">�#P	RGBI���̄�p�!V�D�
_$1Q��W.[>�IS4�^�@�p$��o�'͒����?Q��TE�	z��)a��ۉg| �	�M���D9�O�<Yƅ�8!m�mXpJ�X�����'�nʓy�CS��7j�X +�+�r����'��ܲ �'��'�����h��͟lz'�G�U�^5!���.Ht�͢�g��4اm�u�NU�G��4}&�sM��l���n�' �B4Ӈ��Z�b��B�«V�F)�Ug���V.�1Ĳ8�h�� ���B�@-�'e��� �N^'$fmڕ�2W��y̓a����I����'���G����E�ԕz}����kђ{�!򄄇 �6�� �M�AGb�3a�ʨ:�ў\َ�i�]����p���.�"��$eL�N^j���O��$�"]�E�7�O����OR�d�h�Dن"��s����)�X����ͬ��#�L).��aS��En��D��6R��+�?s�ry���S�&�T9A�n�`��A:�+�R��aiXc�h� 3�!">��
I)�8{�a9gM�5D�>*jj�!qΰ�	̟F{r8OE�R��-Zw�x2vj�� �,-2�"Oֈ�"㏙M�Ҝ��o��m"��'� #=�'�?)/O�eGD�	d�Aۂ�D�5��m�WY��F�O:���Ov��러��O�瓘`-h��C�4"ହȥIذF�P)��h�>K���"��l��	���.,�Q���7��6��)�p+ƀu?�ɓrC#_��E"1�
����Q���,Z�����S��D��|`��xB��+:P�(�뛀X���d)ړ��O*�ӗ�� |�t�(���T4�yP�"O���,/ZV��
߶9��U[GT���޴�?!-O��R`�u���'�	U"K���n�Ɓ!��M���D�������O�$	>s�VdK�*Qf0�9(���'�LhKO�{ؐ�Ѐ��:T.M�,�g�4#>���U�!t0h�h��>Q�����_=�~!{�o�$3�L�#M����sJ�c�'H�͠���?Q��T�C�bDA�g
C�����#���!�O��KdM��$O ��d�G7A�,��G�'��k*�2�뛄+��ܫU�	�9�`��'%�I�s�'y��'��ӖD������8��G̓f����/L�ᩢ� |��nZ��lZ��X��
���� �_���}̧3]�X���y��sQ�Q�y���ϓcP����J $5�1�$�M6/�)�c)ʧ%t	�A!�7sϤ�Õ��a�j$����������'��� �4ڀ�g�rP�El��.����"O�1�R���Y��I�L��Y� �I��ȟ��A3m�i��� FM�
?8��T��O����O\`2F�~�6���O���O���O�!���0\��JF��y��Uk�n��HnnR��� S7����
Ь6�T�'x��➘���ה,.���b��T��[���->IX1ė>��;FBR�UD��'���A¢��ȢP�L��t�7�*?�u�FП ��X�'e��
C=��˘;�pC��L�^K!�W�}��誀�=��咓+֨W�2��|�����$T1� �[�/"F�TaW�?6��(մb�Z�d�O��d�O
�)�O,�p>�`���b��Y �.\�xt|S��95^P��G�R� �B�G�'\�"XR��	�J�>}P��FF�u(���+��L@r�b� �a���"��#¨@$pQ��8���O����N,5e̱���ȕ-$�]�f��O��=1�����Hԍ��L�;4B�L���د&�!��<_��S ��a�;����?�M���D�Y��9�O�r8�8�����<�n|vǙ2K��d�'6pĠ��'z2�'���8���*Ң�c��*K�6q����:6^1�lƶT�d�3Eg�$2�~tQ��ɟr@q����n�*T�G���gLt!&��K2�q@@b���PÌ�rM�#>�C�ϟ��	V�'4|8L8Ɔ�)�`qR�L����0?�e�Բr�̭{AK�*����~x�H!*O�������q�"d�!���"�X���	џ��Izy"_>=���<��!ƸV4�$Rvk�7\e���$��e?��Ĝh�'�T �*�,׮�&/�P����ʠp�'����IT�t�U�Mw��Xs`")~���Cc2�7�O�I�b�P�@��O����:�DUş����|��gL$6(p��	7>Rpo���B�����9�j������]m�{���a��r`��C��):���[2G���'�Ȍ*q=O��]џ(�	�?a���<�*	�7�8Ec0��
*qĴ�_���j���	*t���	;�?i㏓Knz��B�>O�1�hD�H��ѪҫG�ebw&�ON��4�'��@�'p`b�'�?����b��F#r����p��R'�ȷ�Rq�2�'�,�����?�,T��?�b�'�����M�2	�/��XtB�MB���cݸ
�,� @�i��I�U���'�,�˟H�$�O����	X��H�$���Ky27C3G� ����o�L���O���������"�ݐ��ܴ>���c�iC�d� �qqk��Y�z��gMN�q���<OjY)�z�j�o�Lt-�O��d�O�:Q��$|��b�
60��dӎ�qo��2��Ӧ���4����y2d�_"�"/>ǆaJJǟl�M'�ޤa�6C�G.B7����l���ܴ���X?i�a����u���7�A��@ Gvv"
�'l.���^2z��M�e�ܴj���4�?����D�O���<�o���� D%l��X_�h���4�?i���?��?����?�-�|�S�8,U�b��(	j�	fȮ*��7��OL���D�O�˓��d��7�4�[v��3��JQh�2UO~o�ɟ���j�F��~�"�XN9���� �^ ���Z����O֢?�I��kQ,�F:Eҧ@��feX��#�D�O��$%���<A��z�v��S���v��Iq"���f�:}`ĺi.�[���I�	|y��'��I�\�(�`�[7;�P�&�A_�!�$�3.@�����8�rDY�nэ.�!�D�y�HLGeBӮ�y0��7Iv!�/ĕ	RÕZ�R`bLA cu!򤂑9�6}��i�/J�Ĝy�J�(c!���) v&1Y��@�x�ژ�# �YE�O�d�S�G"oSH�ˁgD��5�!J1(�ZpF��#p��K��W�
�bTA������Q%�=��b��̀>M�q󄆟8ŊR��p��nI�`�O܆]A�!Dj��4����>y�mM�<1�9���\=wj9�c�ҭ���+�☔r^=��.��d(Ȩ뤁�	�p�a�(��	�F��D01{S%f�}�r��
C$th�i2�&E�/*�]{��sp� e�K�m��,�/`�i�G��LSI�%�]D�^	�`L �Z��gK27͕����JH��+�YE��� $ƚ8��	D���D�W:M�]�'
.��C���'�ИSq�N�{ް ��upq�ʓ�.`�P?�"�
��şfv~$�ȓ`��i�I�&���OF�i����ȓ%��:�̙�.�xH��DG*�^|��=\ �Ӱ!��) �u3�7���n�<0gH��{���#�
�\��̅ȓV����֢&'����M�?0�܄�~���!�`N��7*��U����ȓ@l��;�Ⱦze�9�q�A�!�h���"���8b+��M��"p`�.VL^��ȓz���*P��88K�-��*])����S�? 2$�#'D�"j�2�E�b���"OMb��w�ʇ�Y>O�}�W"O��1Q��M1��	>�<�!"On%"�*'z�\��D���И�"O���G���E1v���x���"O�QBV�7���*��P�!�"O8MC���ؼ0	��K�@��C"ONQH�d�dt\e���:e���"O2�#���=s�d�3��U�J��`�"O�E���K�?��A��]Y�̉"OV�FR�32�!t
�v�,u	A"O(�Q�#@X��D��)Qh����"O8�ce��P_ltk��R�z���"Oִ0�M�N�i:gc�:8����"O ��;�r5a��/u�#�"O�Lb�Ѕxr���Ŗ9S�����"ODhڳc�D?Q�W�E���i��"OL�	�����@����4D���A�"O줈1�X?E�X)�ǹ%�*�a!"O^x��!��S�&=�4�L=Cs��Zt"O�� J@���15i�24�����"OXE��ȫ-`<at��	��kg"O1P��6YG�Ȼ��]��p��`"Oh[�B�g��K�I�ܤp#u"OHy�����8!��g�jtR�k�"OxP��ɶ��=�Jm���"O�h:�AF�t�� (�
�1%`^2�"O6l���5f��`�)ҹ;'�Iq"O�
�jε$,�`��Ҍoʘ��"OBq�s"٥���K&�O+F�b���"O	��D>�0�����{E"O��e�T��)B��+�ܖ4�y�M hɊ�0� _5`(P!v����yB���G�b�� ��]���P&�_��y2�ӧ߰����˻c4д�uA���yrm�E����3�ܮ[IJ<�����yB�O�"�ѳ�A\�T%��6�/�y�I�
�v��"jΜR�ȵHe�X��y��I�ke��iG�Y���9Ń�"�yrꇸ.����f��9KԮ�Q���y�)��[�.e���8GBpeRS$E�y��O���: ��=?��L���
��y�(��B("I	E�05Kv�I�(K�yR�[�~�Uj��]�-4�$����yRM��Y8䈢��ŃSB4������y��ʳ!<�@慅P��`�ϝ<�y�lݞx���&�!C좌9"�^��y"	�S�ƈ����3��E��h֙�y�蒧]\����+��<��$	��y����h��N(z+�1����yBAʜw�hS�!&D��1['�y���v�QC�o²���KV��yM� u���S
êU2Y5@ �y���G�J�����QPd�@��́�y� �r7�q+����7�E넩���yB'�" �@��%�(b������y�+P�^�,8���SR STN̙�y�H�XB��lCO*
x:����y#F�C:ʩ�5ll)
�̒��M��jJL��m�sw��!�)^>���Tr��1 �ɱ*�yQg��a�ȓ��t��U;� m�@A��G�rP��:��`��F�]��͉�Ƒ9}�@t��\e�u�&u͸)I�+�8Uk�}��S�? ����hL�>�.QJ4ͼ�Cr"OR1X#*PwJ�L2ӯĲ_͂M��"OJxz��#\�"�r�КI��ls"O���g,��� ���aU9%���:G"O6pQ��L%R� ��ⅵt�NL�r"O@����О�(��܂Z�v8�V"OX��V�F�=j|��F��@�
�c"O������R����3��mCc"O� �ڲ(�[�	�54�T���"O����@�
6��CL�52<��"O��	vΊ=a�ȫr��43ZAI�"O��b��{�~)*"!ѲQu�0A"O��jd�Ģ|���э'N�к"On�1JS*f,NX��+	/�1�!"O�0��\X�H�HL%���"O�/��g<:Pʂ�-.1u"OB\HBN
k�|;`j��<;��[�"O6���n�u&AbPxx�e"O�i�q�A.uR(ȣU�2pP"O��`��b�2P�C�t0Ա%"O�����H<hR�� R�B�"OV��P#��� �H(T���p"O�T[�J٩qh������J�`ͩ""O%�I�w��iÄ�%� �
v"Ox���*���CF�6x��0�"O^��i�1���h�[+WsJ`�"O�C" ��u��#'K�� v"O���7��?��2J�7��T�7"Op<QakNo�|��
� l��y�"Ob�R*ɧS���ÄH�n���kB"OP����2I}R�z�`�?d̰C�"OR��'g��d�a� �< T��"O�Q
�
0zA����#%4e��"O"��Z1~�Z\k���
j�1��"O�z��(?�8�H��Y���8A"O�0��K�ya�|��b��U���"O��(6.��M[v�qU� �y��<��"Od��F��=	�C��=X��Z`"O�$��b��Ir��������"O� � ��|�zU.�=
�B-�"O��q0c�~� ����;K�]Hs"O�i��P=/��Z�@�+���"OA�g臖{��Ip�FW�LP�"O��cS{��j6�����"O�ty��L;b댍k���wx��"O�Lqg
ٝU���K�e&��U"O�����\$zR���@���3)�x�"O�Ż#�D)W��T��bF�G`��g"O�0�;V?ĜzʝM1ܑ�5"Ort�U.}�H@�E�x���"O��3�Y�o����9����"O�(�S���1�}rC�$A�4�S"O�8p��:dy�}����.�����"O��#���R����6B6z2"O�� &Î�|8.0�5�W�6�}��"OJ<*@K}/q�!�H�"OL�8ƀS]!�P[�z�RII�"O���F�
�n����C�~y,�CQ"Ov��ӂ��eཙ�"U�zs���"O������>e*��$�H��YD"O!T�H4�H�R�B^�==���b"O����=30�<��Ր
J��"O8	�N�5@�V���8!�"�r�"O.��i]"d��BFA�*���96"O� ~��1w ��c�V6>�8<�V"O��;5�<t��q�s�S�J^]��"Of�*�F�4h�`GԂR�hT"O�e(�� ��x���e��T :%��"Oz���@".V���
2AD"O���D��uS�x1���,;�"O��q��e��a#I�-S8�@"O�!#q炅h��0��˰%��"O�p��D.L��������A"O��(cO�K`6�Zl_�l�HE"O\��5,��S �Qg� 1���P"O�e���ŧS���s�RY��(��"OrHC�8@Thc�^�N����t"ON���˙�'�؝�����0C"Op�Z���KPR�&��1YU���""O�!B�l�k.�s�ņ��$Y��"O�h0��i`�0�eï:uđ�f"OZ<B"�Q9E�P=���nh��P�"O,qh�D��#e�隲��YV�qJ�"O5j@���01�q�ařWT��7"O�,��DV�CN�\��ҨhFT]X$"Od$�� �^�.�R�[C `��"O��8P��"�Ԭ�7��%����"O�Y+A�\�aF��Ɗ�&�j�v"O���-O$�b��U+Gc�)c�"O�� )ڗ<���$��P����"O��Y4�E8ܕQ��k���!�w�<9�t0�ڗ&��)��0P��q�<!���/��v̔��J��5��G�<��+=4�%�SHؼ;�8bq�]�<�C�٨2�^͐��ɏl��RHDp�<�!��z���u��7�̉�`'F�<�p��#-U8���,�=<���cΉy�<Y�K�iu&�`
�;��˄(
�<�+˕WG�ЀӊC)f������y�<�T#�Y.l2�DΏ��s͑)]�!���/=�إ���׳$~��-��!�$�+>��a��Wzv\��L� �!�[,Y�"�q5��~Gh��,�T�!򤔂�X�p����ِ+�!�$=F�l��i^/rp)���!�$G0k0�*�
�]q� �(O 	�!�dƿ%%��3�M��`舘p͐��!���U��U�d�õoF�L��+��Hj!�d�~@��B���C-h�b�T�H�!�d�5Y3>  �A� T���J��~�!��6a�T�V�L��e!p@9a�!��3
A�ɫ2l�'Z1�Ǳ{!�%~��ඇU�f�P� �+ �!��VaM���AD9�h�e�̮#�!��	T��m5"�~#�}��&S���˖`hcc��ǂ���)��y��I/B��&O?{�,{���yb��N���Щ��r?L�racD��ybD7�F|qR�Se���'LĄ�y�M?'g���QIӛ�6E����yrNǬ]V�BO�0[pD�3 BE��'�P�&æSz���n�Z�كI>Y7��b[� ���=|K�)�R��{�<����k�t��3	$�4���r�<����YLN�:��ݞ�-��#�S�<�g��8X'^���M\�$zz�����l�<�S�7k!�<����
�����g�<I�M�b2�3-T�����h�<��O��z4D	�`��u��H#��c�<� ��0k�������g}jA	�"O~(����2A����@��;�Т "O�,څ��B�����@\@wf��3"O���B���(�D&��si��XF"OAB���!l�q�^�ubR@	�"On�Q��@��������H1 "O���U��G(�I �ȕ7��ɣ�"O��ֆ J :1��KI�;�>Ģ�"O�I���Lh�|Y��&<��A��"O��`�˘�?n���#M��?&*q�P"O��,�/8�h,�*�r%j�b�"O��{�bH�2����A4bN�p¨�7j�mZ�\v>=�D��9��_���V�|�"�ɠORb�(8�O�	 X cX��0���Vɦ� !֮LHҩi�EN��(k�hR0"���I0E�S��Q�����
�]��#=��+���Љ(@i��!��S�����S�Hc�A�D��@x|ܙP(��X�C䉕����d�w����a�ɂTG�7ޠ�̒�*�1��9[���
I������A���$-�>�(��Ƶ9�1ZE"Om�R���AA�{�n�:� Y'yyl�T��l�<?��ݩw �r��8T�|9���P�I�MЧ%���)�O�@@%���}kCn�:E����%����]H#���vd6�Q`�_�<����)QO0Ԋ�d�%m��07.>_�J#=�WΜ�X��s�Ȃ��
���ߦ�S�L��`�
�4�C��73v��ċ9{��̈́��tѠ�Ӹu�L`�q%U�-����^�ZTu�ʎ)���H�-��i��#}��O\ÕkO�6pAsu�"��G{r�äGWp�D��M�\AxZG*Q�?}~X����CY���l��u�%���y+<;����Fx"��';|X�+�T$��p�$�&�|�Ǐ՞r�ND�M��>q� ��}�g@?A*N��' �\�2���4���D�?� p�Op�3��~#XtB,l�4�Ѩ��3*�5 � ��Ɔ@�/���2��ĎP�|���0W;�Q���N�Lrg�x�t��o�w�P˅fsʾ�qu�B(� ��@��!Z���3��+�*���қM���a�	3
>"}�10��ЗB����%H� S�E���?I�`��[�"�s�'��q�\b?!Ku�T�p�4�\P������H�µǁ�tA �i:�u�� Jԁ?3Z���㈷d�>�{A��H�1�-̰8��yI��'��c?m���~f�¬E�Y�4jֵpt����lE4!�*�X`h�%#�\��ɵc7FL�����L��[�[�g�7�֨)V�4Z�A	�8+�`���������O����!2b����77Jt��;��\��N��B^0uO�=�h��+P����O�X��q6o��f�:@�MO8-��u��D�-'�>9�e��+��4y��F8'j��"ɀ���'�I0����./ �x��	�[aq����נ�@��P�r9�8���9������p����\ܜ�Z���mFx򪔳��I!��>�z��B��J8��E�4B�*��c��:�M�%�I��{��,�<�Em0 m�4��ʑ)X��Ɇ�C�T�  �*[s�����<����u�E#Zd�J��P��`�C�N��Z5��I��؈������9���}�=B�ҷ5�f	) �Q�S��r�.�O*�ȰH��=��C�U�t�7*T�B���!$ "i��R�F�>Zc�D*�8��!���Q�O*T r��}Yh���\yQ��$#1�d%@�̧_z�т%bř��']���T�<s3��(C�B8v�)��'@��X�01� ��*�a��R������'7�y���HD�� C.B�:1rd�r�w?��92�
Ջ��?E�q�B?�P�F�<6��ӫ2D��ǣQ'��9�s� TS���%KD�>��rfd�3�O��=��d[�L8��-K��\(�U�F"[׶�Ɇ'�>O2�K/Ol\ͧ�(��&�/�P�E�&W�& )5�����'~&!+1���g�@�$>Ot��P��Z�Fxa�C�CF��	�A��	�J@}�i��$Aud���1$,>����~��J3b�"׈9���#hh!�b����dІ�ēQc��B�q�5yB?Op0C�D>%�!Q�ԣ!\u3��>A���4��b*.&��*ǯ�ĸ'_&��D�ؽe���*�鈄<i&��hBO��1I��Mj!-`�y!�{*�Z�jp������R�~I�$ "���F���� 9z  �ʧv}��KDLL�TRGm
�=�Z�i��]�0X��P�	L5T���7��sޱ@�JJ�/4P�B��C1v@;b;}"�;Pb�r�VRHː��,O�Q�e@Rhi�@\2gT��wU��[T�%�N$�d��$N���J8a�.N)r�ɘ���M��h��	�Ya� ����?��ǝ6\���=?�A&���(E���CW�-p ��v늍a�I.����5[C&]� R��O���Dj�30��i��a�d-D,H�@QJP�&?���J����~�O|Xбǎn�p�0�ծ{�P���4K������,��|����4;� A�f�!�M뗋<"�P �X�t�Cȉ>9H�!PqO�P?K��� �x��eV>L�y���'�<Y���>1�BW��x�i_2ֶ�ȋ��Odk�/EF�t��1f�7�YD_�D��ָ1��J7lYC��IՈ!ʓ~)%iv/ώ=���6�W0v���*A�&w����'<��	Ħ~�˓�
\N|�sL��765�f��
t���b��L�xG�	�ukC�.��|"��;B*��+��ɠ".�K�霡�x�!����Rڜ(�ꞑ$_N����B���O>��OD�H���ĦS㮽�S�.@u �A	ϓc���W� � �C�'���(�M�vE�̫H�0dj��֭b�!�hG�!Y�����F:�>`��0PU�bP](�B��
�L�{��D��JL�y�o*���
Y��+	�d�b-3�/�l|q� �O�J�)�"c�B����7'��X��#1�4�)Qg��Lc��y���>�(�Bw!�2��'�x�'�0����.�쀣�ŵ`ʎ���*JxQ��M8���бv�b�C	�.��ńh�Jpip��fd�	�NhPMnZ)n�N��W�ʜL����iQ6���$HԀ`�4%B�&�)�H�j �^�y�ǚ���H�i=#F��c���&*x���R�4�&�2`�-&��l���Đ�H12GAOL~�9�A�h��`��9D����J�t���l�n7jx"r#!i1� DǺ���t��7wb��D`�0�*#G��3�X �f	�a|���u�XI�"���eK	ע�٧��z	� �ȓ0 B���j7ƥ9�+ĩ,f�*TJ̓l��<�ؼC�ͰObd�9�gO�,�á	Q�<1��E&��@6��RSZU�sgVS��	R�iݽ������O����iU|d���_8�	���'���p�'�3�l�p���rF�a������@z�:�Γaw`�cY<��=���ƥ)�����4�cj�0K4�g	
|�j]��Y?O뎟5<9s*�9�`	
���KC!�dQ���ESG���k��p�G�ޜe����M5D�v�?�����;�x�;;W�=x ��`ǀ�^򶱄�/��
�&R4o�(��T,Q�	�Z �x��HB}$ �P�"D�RN�6���{��R�W�� �%�G^<���
�^���D�x��ܦ���+�"��%�&C�ƹ[�� ,(ZP� 
	��i1j��q�;4m(Y	��h�4��
�~��Ӂ.V6d�r �/V\i2&A����	,���`D�'�p8���f��u�/r3��އI(��瑎y�r7M�W# ��2��z`<�3�Q�hnQ��JkI1_P��k��ܺ#�\�)w�ۊd0��m���M[�y�O-P�Zu�[~��LV�� $���bD00@ո[HNta�M`X����fW���kwM��!�<H�W*C�`��o�`x�ԫ\����?��޴R��4��'zB(��-�3T,e0!�߬=�\�Ǔ<��Q��ɔ>3�i�w%��PJ>ap�+U6:��kR�R	&0��zb�6��O�b��������G�,�� ��B��A?a�$��P{����H��(���:��}≠CѦ��q
;L��1�'��dz����^P�L��"��K���:�-�>m]��nZ�	2P�r���Ǹӣ��� �>��CZ��Dc'c�Ӧ�.�@ȸ�KJ�R��E�'S�
t����)xNM�J?}��i=*�����$��$��B�-�7(6ѡ0�'�=�v�s���xM"%�BŃ3}{�0�gf�GˠȊ�,R"
�<9ѳ�)B������V��@C�|>$�`�CY�lSY��'�V1⥤R��M[�'L�3F�ǻQ�Ͱ�Ǔ!!f��D�#t|��M�,[�<f���(�h��(V4�s�b
?q�]"��/eQ �>��CI4����'/���1g^.Z�*P����L�l�6��\���1��M]���i�6/Ӑ�>Yp�	
���!	��@�*`έE����'����_� 3�,�� �u�v���Р x	4ߟ�9�iN�*�<���A�"��ɒ�a]��ū���ċ:u�
� Q��SR���~���QE�2%�q�6)� _����2�X�*�Ӗ	i杙=,�@�ڭ>�`�#GV��B�	c	���r?�&)H�)Y�F�1AH+���@Ң��"̅�I`���z  %
hB\)��!����K�u�P}��F3AFZ܆�ɇr����R�.B��3( H���=$���÷k�^��ҍ�1�<�A��<;�P�Q�`]��F}�V�2r��@H�1��l*����ē"���VFWy���iWJ�5ÈIY&F�����%��V�A�W�Tv��wn��*��3�	:�L�c�8 "IS�E��]�Y�BG�6=Ee�"�Eۄx�#�i�dl�U�Ix�HP�I��=p�X�DK�&�e�&�$V���e�HG`N�x�F��~C�!��	�sv���� D����UH���p�IgZ�C*�;f�[��K�O�V %x3�
�C�8UI'H��4���HeB�w���8`�C��~� �T�#֯+���Ҩ����'D@hVK_� DH�{U(LAp�\
�4HMj�i��4�r�!H��CC<k:(�
�)Ǡ[Y:0�ӑ&�Y㥋R�Z�3�I f��i	U��,�"%�Dk�a����p����-Z�i����!O0)jh
S��p"$�@c/p�rb������PF%$qQI�DE��\��/�,�~�V� ���ad"�K
Du�2�WJ`�4 I=��l��HD'M��s� N�`C�bb.��|�0	�w���r��+(��dʕH�=.��l�w�ց�p=b����jݩwd�)� � ����3Fd�K4)F�2L�)%�E::�0a@��d���$��2�^���-S���H2%^�m�̰*�'�丱aV4�����x�f�3,O,� w[�b���ʘ0.옂�J=0�lZ�1sP"˕=-?��+'�Z�֕�a��@�����S�2B^ɢ1lM\��X �>M���>9�M�qjY�X.7��e�O��S���[���`!�q�D6n�D(8�A
�u��X���y�S,1J�d��#�
Mu�!
�<)��]�U���a~�R#'1Vi���>:b.)ْ� =`|��+�/��D���'m
��o_�"���I��.Z��(ڐ�-@<v�*޴yɰ��A�ȕp���L�w���C�("5ў�*v-�|%��E6P �0�@�B�3�J�[���YEg��C�,�y�9s�d貓�Q�u��9��Z�w��l�,��=h����1"P�Rk�\,��,89�)%l5���Q�R(O�p����]�P�Po�|E��$'X�� �]K6I�d%��q�.q���Z/�P���'֢�c�'&4�Z�T�==�1��e��n���gN[�U����կ3���>O��Y�L�}*1��m��.*����wd�\{�JP5j��2�oΜ ����y�-�V��oW�P9Vf�k���O-Q��a�hE?9b �?�h�l6 NP;Pj�����K
=q�r�%�Ͱ�=�Y��F�K��Ey�l�9e��̲�#}1X��J�&�P@�ל5��㧢
�T�H�Sƛ2 �xX!@V�*I���?�EJ0��𤓆q�l�s�k�#^β���!�x�:ic�W?68��$[/�R@�E���Q���r�o�3~2�I]����g�:od����c�Qb3˖0h8�m�	�'c�Mb�%v��tQ��� � 3��4�Acq�R'E��p��L`�-�y���`7��w�,� �3$'\�8�
�+61��.`m���CK�@�ёG�S������s�t��&���)�a�H8��	�Jrz�ӗK�,3����	�S���Q�]�&YC����A�F5��Fz2(��NX.U���*;D��q���dC���J�(��@��afQ2�I�:X$��`l�n x�j5s�Ԭ�A:O2�7B
�7 ��0恽eKzh� �'���xW	)K��Y�\�"~a��H%�8SQL&��(����y"f��O���bM��`�"�&��	��Ě1>��d���C����$̎=�:�ʱC
�R�fܑ��	Va~��!k�v��aڰ#� ��W]�N%�0#��»(���sF��	ĄW�K}F 2Ì��ȑF~"�^ f<�]��b�=p9`m�@T�#	�$��*[�<�r��Pi�t�֠|
��"Dqy����OQ>�"�G:r�2}C���/`�t�3�I:D�p�$�9���F�V\Q4���'D���#HY��Rq��dִS�`�L'D�T����'����g�����#D��z�`��Q��o2��� D��[a׊� 샔G� \g�܈�`*D�|��J�͙Ẅ#/��Y`��(D���A_���R�fU���Z�(D��۠gK�b�Ơ�q)3w�Z8���6D���W�^�P�` !GPB�@"N4D�x��c�(�4-Z5gũb3�$�>D����Ӯy,u�V�M� Sp)p��8D�DK�(' �VOCn)jWk$D��W	ܨ'΂����tr��%D���@aY�V(ja�0��QF<���7D�T�eE'thPX��Ü-Z�`%D�5D���ꅕ	��ʢ�O-6�`���/D�@{G��L�� �X1pf�Ya��/D��zW��L��pb���5r\�"�0D�$3��F�U����Ad^fjx�b�#D�(3�)�~�@ �B�<h���$?D�t���oe t�B���P�9Wf>D�t�a�
C���/�l�F=�0�/D���3�ou��� ���tnbMR��*D�ܹGO�?9�J�rCA
���7	)D��F�?:��Х&�vHrgi$D��H�B�F{�����66>L$�"D��A���>�HzB���"�!D��p�0,�
|�g�Ua��o+D��kSU�.�%�� ,�按D�*D�X;��J} � �O�"�zu�5�7j��;��ҁ\�xU���%�ĒO<�21���}�B�ĺ�|D�"Or�:�B��-�.�Z�Ǌ�{���"OZh#qZh�X�P��ʍ~����"O� �5�6n�%qe��?Q��Dx"O�i�P��D#:�c
T&!�L)��"O����  8�^`q&i�������"O�X��HxA�$*
4�� �"O���ĸ�Ӡ�+�z�A��F�<���8f�`����$����B�<y�BK�Y�XͲV,�!�^M��m�U�<9��t�����,��WO�P�<׬�[�N!�p�H_'td�R#M�<�t�	�]r왂<�^b���K�<�&ȓ=g�|�r �C�$��q��I�<���W+6)��	ԃPq��̎H�<	$杗2��a����=py&��u�D�<��aއ68̀gL�;]:a�BJ\A�<��f�-ZF�]� ��*P�H󃋗w�<ab/ġ}]���ǉM3�z,[$�o�<y���8z��y3m�8�rmS7�Xj�<�`��AML�6��C�B��Dh�<ёƋE�b�	�NK�,4�P�H�`�<�k�0/����(F�F䰡�!�R�<�a�-�&�(�/�:t���G�I�<7.E�԰��Q�U�vX��n�<��e���26L�"��SI]g�<yT�R�%��5�A�K��2����x�<��)�h��+��T��)9#��\�<1`�{��:��I�D�@`m�A�<y�!L2��0;�B��%��hL{�<���9{|��q��{���"���w�<iC鎊]�����蚖[?Ĕ��Rj�<���Ƀ`���۠�����pg�m�<�U��^D�}:jwM~����Kp�<I�'N b���	a[\yp�o�<��CS�t��g�K�4�]�f,�U�<I�F٥\�~��K_#!��U�<Ʉl�l'��U`�9��Z��DF�<��a��45N�*���(E���J�W�<�7 �&��=3���0s�"�ٕ�JR�<�SJٯv��\XE�6"�x�*afUP�<�%i��BS&��I�3'��Ju��M�<ф��$n+�'M��H�'C�<�� ȂD�t:Gf[E�HӍ@~�<iG��NuV���兑0-ܸVƈ}�<	V��*y���s�H0a�b|�<q�ċ�<����wF��Y��$�N�<�A����W���v�jm�$�^@�<��Tu)����C^l><�"�f�x�<�f�ǇsEƠxY����Zj�<�WB�:o�&T�@��1'l͘�`�}�<��S@�-8S�J�
Bl`����<��i��9C��@�1�v�+��Rx�<aFh��yB�(�)H���Bt�<�2��g�^�Q@�ϡ9V���A�f�<��a�,�QAm�s8(�Z��~�<��L��Х4b
�^�Dh���Jv�<16��q��8�ҋX�7kF%����}�<q�d����W!q�v���o�<9AiԻs��p+� *�&��#Ri�<�� 'n�$���U�~0꠨�o�<1�c�'N�j��S$~ ��h�h�<����4g���]`�y����g�<	��:#V8��ێ
@��q��O�<��e i��AEd
0I�xQ90�G�<��)�U{@YHw�.v���{�Xx�<iE"�.Xn�svT�j@њ���t�<� Fڴ�۩DNr �PG�e� ��"O�Ŋ��[9$ؕ��Q�j��Ż"O�uB�&�6�$�ZA˞
+�-iT"O&��aJЋ@X1e�މ�V@;�"O�P��gG2#VMB�HʉX�:LAp"OxMcBbP	K�xq��ĪH�X}�g"O�����{t(:d��� �X�O�d��r�L��>`
�5��
�:�!���Z�a ��5^����;v!�)t�)W��y��GO�8W!�$P�D��&�(p��Z��H�$�!��=<�a�ILG ����)~�!��f:L���_1)pX�u+�5!�D@	2H`��a	]g�@�`��&x!���h�ƩO&W� Sr�M�!��f��H����8RTX���u(!�-/JՓ�U�lXc3���- !��6h��6A�y�rP�
 '!�dX%�d�JH��x�tE=L�!�DO��l �.#2�<�!�fґr�!�D�rR�c�K��H�4Ł�u�!��Ұ]�3��OL� �����Ew!���=���XqgЇ1/���ECߊ(�!�DX�Hg���+&�	�(�+#�!��ŗ:�����}?��QTDץU!�$H/
���ٓn�)YL,����9�!��<M�"ӄ](U�2�	�Β�Q�!�dU =|x��7D�ЬTްv�!�$�8g9j���Fɳ�.�(Rʍ�B�!�䏯��D���6�|�X��-n�!�W
. ǄG�E[�iiR�_?K�!�T3��M�DVH��9TB�:wH!���~��0c�m	t��E#@)!�S�C`����~�f���c��E&!�$�D$���7� X�xh�A��!�䝢'�č��]�^�,LSd�ښC|!�$κiށ����2J�~��b�Ū&x!�D	�3И饌�8��1��E�$!򤏕�P)�S�d��,��!���G�jX�T�~�Mu��d!�䁹W/XMQ%�G���%�2<'!�$Y6R��A'��/J��9�N�5z�!��ƐgC��OůI2"�sS-��b�!��$�Q�R�ӀX>%SN��H�!�D���H�)��OWݔܛ:�!��23/V�xP�nc�Ydm��!��0#��=�]*�l���3�:Y�'Fb�r��hl�y��2����'��L���ϯaj�%��(�19���q�'��)0�E�:]UX q%B�EW��s�'�n�Zi�2^ҥ8E㛥A�<d1�'������J��	vg� *��	�'7��yw(T�0���םe¥
�'���p�C�Wޘ8��N�Od�$ �'zZ��n���1Ȇ�4r�<tq�'��43$j��u+xq:�|M�
�'����R���I#�t��J�57��h
�'!�53�%L%@"С��0I��
�'��[�R�"�$S"OQ�b��	�'�R��Ղ��Y�B��/� �� ��'�"�KeʕtdYx�OTiJ�8
�'x� e�	�r���&b݂e{����'F��X��#�H��E?c����'�ƽ;�!�5�)fѲW�4c��� J�j2꓆t(ʈ� �-&�(Ia�"O��9"AK�d\�k�)��k��p��"O���T�E�J�F	��)}��'�#�+CǸ��@"_�.o�ȸ�'g�	�6�٭"�]�'�Z:|<�a�'��y�4Lq��R�,M� ]� K�'0m{D���b$Ѥa
�
5��'f��{�n�E��T"��U�t��}�
�'�jjh�$$龴���ס����
�'��tK����o&���؎}J��'�dh����y���i��=(���x�'���]�L�1�-ܣ'�L���'ܡ8�,ӂ{���c�O�l\.�j
�'P��4��K��j�B+k8t��'E(�ӲX
F���gl�\�T���'K"{đz�*���%I�d)��'�@�@�"Y% O6��1�R"mq�'�����#k��\���47����')l�҃��&I$���	�W����'Ʈ\�C��Z�d�S'��R��[�'��󣖰*%8҆��Ir��S�'��)����12�� ��u48I
�'�2ј�	�\zx��tB�>e-2�'(�%.쵩�"%Gd>qҀ��2�y���m�ʙ���[�1��zA���y/O+�\��1`���XAH�4�y�@܀T,�!�����^ i�j���ybhӾL"�h ��ڭCV�9�y"�W� 8I&�قNA�p I���y�۽ �`�;3�X+A�����AJ��y�L0sO�ps�eC�Gg:�X%��y���$�L� ���>�T��D��yr쐘n𴼹�I�m@��4�	)�y�Ş6��a��a��^0T�� C�
�yCSQ������(Ȣ�	����y�k~�l)Y�@�.$w�P�%���yB̗*Z���e��/�p�Ń���y�[�>�X��	O0.�� �4"��y�M���쐺�J�C4D��y&�8\^��U��� uZ��
�y�#j|Ե��T�0�A�A�	�yB��E�����L�zmd�邋���y���(`����n{��[�H��y��
$kP(m;��mf@yA�\��y���G.��۱�Ne���� �Q��y���;�����!ZVȘ����yr�X�l�FpqF�ʹ��������y��AY$ ��QG�4ɑ�d���y"˃z�p��р̒]���3N�y��7\rr�	7`�Jxz�{u�ݬ�y"�U�o�"�V(ǰn؆��'��8�y�ל:b�A���lM��bO��yr�֧56=$$��vV-�����y�I�1d�a�(�,&��- ̟�y2NԇC ��g�ǵfOZU!3��y�X�#ݲu�q#�e@�p���%�yR@
 ���I®��Z�8%xp
ʠ�y2�Q�,h�Eb�oH�O��z�I��y�'p��m"f��q�x�4�҃�yR�+hS*��U!g?���%O�
�y"K�q��4 �gI�`�,q��\��y�ˌ����'..ԛb�8�y"P!�du���N�\���Pf�Z�y2�̹{�tͣ6JTT�r��`��y
� 8ib� ]� McT�g	� 1�"O�-�Ʀ��x�:�.�&n
�yp"O�H�P��&1�����F4tH��"Ol�t��)O'V����*.���"O^�;F�P�+ظiㅕ�}Ȁ=#'"O��Z4�9���c�ף0�6|�Q"O��ŀO�2F�C�־cڸ�b"O����0�L=�#��KҜ)`�"OЙ4̉6;qvĨ�ȋ<k�PS"O��9p�B�X�����Nh��"OHr���9m.�1�&�lY��f"OV�ǌ�!�B�(&��Lxi`w"O�U�)$ظek`eĥ~k��*"Oޙ+�N� 2��$��fh�t�"O`I;���B�-R���]X���"O�M
T�J�6@���Ž6B�(ـ"O���B�`���*Ł�8��J�"O�x[��M���[���=�"�I'"O��Z���T�M���C�l��K�"Ozl���^�-���	�i���H�"O��3(@�5 �YC�L�RwdL:�"O�e��䇽y,r��B($h�c�"O�hӗI�[;�h1��A�?S�ؙ�"O�X�e*�=0bx V�b?��`"Ob%7��%���	��Ȧ,B�u��"O��#@�L�>���1�M�`F���"O�8`�E�$l�����٫]hpI�"O��Y7E�;aN�;7J�~C��[�"O4Tۅ�
 |)+�OU>i�@!��"O�5Ja�/s�,Չ5A?g���Z�"ODm0��\��p�`�=&Ѩ��3"O&LC�I�7
y���j�б�"OF<����>�D���T�Mݢlr�"O������c��I#��85�b4cT"O�C3�F����ƈC(����"O���%�T��K�'̝&����"O�<3�<_N0#E'ی��\�$"O����P8{=���&@
E� pz�"O�`0G�9��$,Jv0�d�Z��y��+��Y��ϗ"<�H	TH��y��ٞ������p�$ѪTj�#�yBo��V�]�-�b�6M�7c�B�o&����G�Xh
l�B��`3�B�	�{�ؔ���G�ø�wJ��,��B�		�qY�g�9�����]��C�I�8��YiS/�w��3��85C�(
<HP����͐�⚋9R�C�+v�dY�LU�T����2�C�ɛF|��f �<��������C�ɡ��*%�I�r�H��A�ӄ-V�C�	�Sݘ���IE$Y�4Q���`T~C�ɴD����pE�gwpy2,�-��C�	�1��a�|BQ FR,$�C�ɥ꘽+b�(�3#�Jt5�B�ɪngFE�쎪Gyp!�NǄs<B�	�Dpj�"�%ɵ�,��Ha��B�	3i��x�A�S�\4D���TB�I�7A�T1��؄8H��,��C*B�	�L�֑C.��W

��ፙ�|&B�iU1cC,�?R��=�P.ێZ��D�
�'����Fْ/;��K ���&��4�	�'�Xy��i��%Y�� �#MEZ���'�@`����o��:^h)tD��y���Pd�&	�0%�h#L,�y
� �����2}��z�D=:4�C5"O�q+��(c�lj6%�!{2x
�"O@-+�ß76&`K�#K�ݔa� "O�x��늆/K�����&�8|А"O����Ђw�~����ץ[p�<z�"O'~W���JM�e�ɤ&�0I!����i�ˉVJR��#D�2 !��-m鎹����\9nT�a�ٷaE!�1r�����(.N䡗L��!�B�Mz4���S�|ܙ���ȭp�!�DD�Y�贩���^�Q4�7V�!��;����?zu���ة:!�$����ڂ��X��7JQ,!��'�phx#I׭,j�����!?!�´73��D�7�%*�����!�\!h�2H2 �)Q�H%�+��{?!�$�b��9�.�w��Äi�IP!��]�m��a#���"w�L�µ'�N!�D\*"�5��B�.�>l)0�8C!�$D�#�4t���=
�4U�B�>
!��U�[�F��G1,PxY�u
�5.�!��{f������~���A�!�D�<w-B�`�#�Q�h�㚅Ot!�D�&#G��8�/Z�mѬ�I�C�	tm!�]P���6"&��ݩcÇ�!�ğ�]Y2U��eƻ��E�C+���!�x��Se�=4�T�um!�d8nAb�P��~����Ҏ�^!�䍫X��#�)������B��Y~^�z���;Y�(1�*V=<; B䉳�j�G 	w�L�;� 
�T0�C�I�-+�*���s��RA� `��C䉢q��h�Yt֪U��eE7z�
B�I1V**a��T�n����	��
�B�	�N�!�����V�����,�2RB�	m�v�R�DV�<P��A	htFB�ɿ
��@�%�
f8�C%^�z)PC�3=��yAH�L�`P�
^�k
 B�	3@D
	�T�B�L�@���/j�C�	�������*�8�6��,��C�ɍ8@����̹_�B�̓E^nC��(Vb����͚vy�}�TAJ�n�6C�	!'���w��p�"Hb�B�3rΡ�8}��E"�Y�DfN�%�	=�!�L'�!�@���"Gh��!��.T�!��K'9

p�B��D����#N8�!�'|4�2�	�:]�ʄb��A!��Y�j�갎ޡ3�h�8�߀9!!�D��9�D��˂'jd���.M:R�!�d�)(��D6T��7nN��!��q���յjY,9C��J!%�!�Iu�)CW��mt�����Ǐ�!��b2�	p��yC�0[7k��5�!�Dɒ7d
�����y7���e���!���K�(ْ'�>o$�Ta�'� <�!��?���RBM�_
 d�e&�PU!��|;��WG㖤����$v!�d�z��V#ӕ^�@��[�Ҕ��'�6�����<k������!����'�4��B圸����#����'�D����Q�7�h�p��*����'8i��bH9N�u���5���'����0hɦO���`��?����'�;��2d�Jd��)��Kr܂��� �1B ��0t��(���"i6(�T"O�-@�ަ'� ��R�b���"O :3��)6�P�F�M���@S"Oqx��,�2P3k}��Y�"O����ݿ&� �������q�p"O�u 3ʐ+�a���#'���f"OX�{U%Ub�F� �C�C&�8Q#*O�dA !V�sk��PE,Z��S�'7(%H2Lܖ|�\A�g70�J�'��hX�ف(j��I'Hԍ*��L��'v�9 &�9e#4k�";�I�';\���R�s��)�������)�'�����<{���ӡ����B	�'n�9�Q4/�nܻ"�Ϟ}��(��'G�a�l*A.��
ri��_/4��'Yذ�KƼU�|�&��& ��U��'e�Z�h��g�А�u���#�'m�M�Q/��m�P�x!�d��	��'ӂ���M�n$܀P��j!:}��',�,����R�u8 �ɀ|�<s��l��!�ĥ�ò5�Ty�<9Q�6o�5a`�P�e�$�HgL�s�<���Y�5�T�a���$Zx� �iEr�<�"�E'�:� �I[!�`(�Bk�<��ʦNft���X�K��A��Me�<a����%�]�Emɗ,�nx�"*�_�<Q��?��URr�� a�1`�_s�<!fo#��(Q�E�ܸS Lk�<�͕3n�l�#��M|��8�@Hj�<���W�%R@h"ԦO�Jh�!�cQ�<!�i^#`���s��;Z9��7I�F�<��]�|���d�XXY����D�<����9�t��g�=�:8cP[j�<Y!�di4�b�ǵDO���aXb�<	6��I[n䩄˴HTZ|��e�`�<�PO	@�Q��P�
���@�`�<��#��i�Pp�C'B��!��H]�<#	������ ��? �!A"`�<Q�]27�\@�U�9\��<9�ng�<y!Č	"���7��=FphIt@�d�<g敆V����@�_�9rR �%��^�<�p�L~=��#�X<~�i�!a�<ٕ	
�}�|�Q!�$#�I��,�T�<�rn֗h��@�Dh�	P���Sm	{�<Q��Q�.��*�e �ok��b�
n�<a�
 _q(��B��?nQ HIC"�m�<)!�o�xT�6n�8�<,�p
�g�<a��e�uys	̙H�����L�h�<�D�F�J͙`�PFh�u�L^�<��;z��L��M5)��ԋ5�S�<��S�|�aqD��\U�� �w�<yf*4%��p���¶}�A� �Z�<�r�Ǯ4� �	[�;^��RJV�<��ς/����@�Y�ހ�ck�G�<1�����D�$J-E�� H�C�<A�J�A0.u�烀^)�yr �}�<��/����R��D�i�:���k�z�<9E�E�c����lO1]���{'��w�<$��X<H���8Y٦a�Į�w�<I�cDYShX��
1R���̗k�<�mƪA8��ʡ�΅80�]	�O
i�<i�T/��!�Ff�Y| Q��f�<1�7NJ��a󫈢A�ޙ���d�<�7\�e̘T��锝�0؉��T�<� R�ɐ��$�ҐĦ�m�0г"Ot�q��F�3��Apr��:Zj]�p"OL!!�����IYłϯ��[3"O�ܻ��*4F��I
E�F"O�0�0�5 H�"!={;DI���	����.��'���U?�@T�&��aq➠.�d,��M�ZЦx
��?��2�d41FjN� ��H�;*��,+����Zp�J/�2�V��P�����I�a�
��R���Evj\��Lr�)���|
e��	�"aAc�:vw6m��kc�'����>����{�����~b��E�XP6�9�,��c>2�Ti�"vZr��%�d�b>:p�RY�C�4��LN���|B�`�Z�lZĦ5���W�1� @8�c�WS>�$��<ȗ慮��������O�>��'�B�i"�p�!�P�s�	/�
q΅P"��(��Q�"Wb�����W ��2(&9��'��[c���r⛨ x����K#^�Aߴ0*��rV��S�v`�`늱��13��.h,dK�.D�
��s�%"�QR�z�c��Q ���ف�f��1�r�'��<�Sk��Ms�-�"=�hX�"f]L���~?����<�p�O<�
�CvQ�dr6�I'A ����d�O2�l�M�H>q���u�lZ�o�jT;��S�-�F�Vg4͚��O�٨-�
Gq��D�O����Oz(�;�?��4e�V���Cy^�%)5�L}x��5�'1Vr���Wrȸ���;e����
 @:� N>�ޓ�p�i��B�t�Q���ץh��p96I���*���a_��S�Y�V�٦g��L�e�$0Q��1q8����F�?m�'��S��E72��r�xr�'�n��\}� �{P\ �éYT\�Т�Љ�Px�i�Z�d]�\�fѣ��Q����� A玲Rٴ���|R�����$!�9Z��x��qRcȅ>�z!I���h�@�d�O0���O���O��$�Ox)�2�O�����(��7����V�d(�G^�[�8��P���Ul=PC̫Q��K2G��h��-@Ӏ� �~A�tL�7\�(J��Ze*8�.}����%�8Q��;�!�O�8/�2.���BT,`�j܉O�1T���o�֟ؖ'���T>�[�F���`�
��N��u�g�5D��k��L>*�M�DJ�>��E���?�5�i<V7Ͱ<QU�T�N�F�'@^?!�T@V�{zL��Q�����q���y���3���?)��_����T( C�Y0C��2�rE@�i]�C�l��$���Uo���E�H�@�����R�'1 �w�B�fOe�v�9t�b� 5!�
~q���Ӭʀ ��e��j/c-�M��!�B�As1�B���uӺ�%>�l��dXf�!�,-(b8�핋a���������))�ɫa��,x2�ˈ&�8�PK^�*;r�'ў�8�M���iě΅#߂�#"g��C�Ќ������~b��>'l7-�O��d�|�$((�?���M��λp(ј&@Z���0"��E�Lzt�VYj|j���p��T `C�pd�m�5P>=����
�a�h�6�؝_�J@�"i��m觪Κ���m�h7�Q�޴�Q�6�s���Gb�!:b�����{6��q�N$9��'��6��Ny������C_�K�B,��A��L	�S���~2�'?�N���	P�m��M)�&���AA�ҤP�Q���ݴ\˛F�|��O��.T���@�P)ږ?V`�Cb�~B�$����7k p   �   4   Ĵ���	��Z��tI�:F�����@}"�ײK*<ac�ʄ��	ڤ´�xbjR�7�I007(2G�U+DUrF.KW$ts3���rv�y�Ʀy�"�Æ�u�FR:=֬JA�,^)���a�O:pC���0B*z��b�_�}�E������-O�K0	�O�
��O��+�Mݛ;�@'H�N��ɀ@��5M���!��[���$���T�Z��5z)�t�Z}����;_���n
<Q�wn�'|w�,�����a�����9o�&�C�b�:k뀁SJ>Q�Ɉ�O�(����.2[�9�A�n	*����R�\�b�4Oba;��������|�3��s�v�NU�[T�M);�p��q�Q�n���'T�m��}��K���{!bO�G���$hM"��k�;����\c�Ĝ#�uX�'�>a��d�j��	: ��<ɳA�9��ɃγS_��Y�EK75dU�f�V�IO�Fl���"�d�-qNp+孂3�y픳b�1���F���2fFה�?�A�R�r]$�Њ1�ʩ@�OplI���;��z�dE5*(v����V�B�	xK>���@�m��S*󤅀b��|���P�m�C���Dx�<ْ�Le��an���y��ߡZ���'���[����\��nv��5G�}\
(� ��*��0ˉ�
n��T� �d��ȶ�(�)N-&���a�, K��Mp1�X�sI���,]}�Qϟ�i�̈�@\�I��?$�B�,�!̓" ]�Vˇwf���4jP+(�k�h�O��)�������� B �A�2�O4my� y�����']��3����w&N�i�O(D�O���O< �r���t��a=�����_�f�pc"#O�B�q3qc\�/.�Y��/�"��[�*����Į�(FR�q�&�OH�������@G�>z"����[�Ģ3���ړOR����Ԟ	��'�v�����\٣��/3<� I��G��`I>��k�����<I$�Q�C�������j ��{�\�R�'���@ ��^1fU��
!l�J}���OQ�<�d�@�hPC�# >�P5z�"�p�<���<�q��T�C�(���]D�<�� ��� J�)W�	>E��N�h�<Y��M�$�tkr��'���SA�i�<�4�]8�wY�Y��� ��^�<��Ņ9t���F��R1��bf��]�<im�	��)Q��e��yJST�<���4Ys���ޑqz���g�~    3
  j  �  �%  3,  w2  �3   Ĵ���	����Zv���P��@Xx����W������K;G� �$��=� ����8�҆�
zn�(
��U5}e䥐ć�Znb	BR�B3c�XA����(=��цOM�;OZ�xa/�X#��b�j���)å����h��ܬ'"�`���	�(h�	8�-�L�}�ʗ* ��C,	�a5'��l�(���DJ�~\�t`�e��R~8X�W@�X��[ֆ^4�I䦇-k�8,0P��M�l��ҥ��:�]�P*A�F��iI����8���	�Ls"y���A�`cZ!�f� 
$��T��c^ If�JJ��$�揂%OHp�ȓD��*C�N�#��@���n�����b�JٱeE�j����Hʚ~��)��E����J ��2	H%��D7����Z����H
K�dP�@/	����ȓ%v��Xd.�*)��x).,�@!��CqҜ���2Z{8qh� ���Q��Pt�1"��Uk������u�p�ȓ$.�t(ԣ?�zaE��id� �ȓJPּ`Siwl�zV8y�(݆ȓr�89��+�	$��}rWGJ�5x:̆�e���`"D��.�UJbM��X����ȓ^^��u`�V͐%I�t(��Ki ��s�H�fJvT���S�EAD��U�l�B���P�ŀ< 0���D���Ԃ/�zf�;a��ȓȎ��IW<s�|�+�-�62?����I,S���*�)�&v�9��P�\�4h �e�d��P��6dN,��I���?��)�;����T��"/�Hd#�ėg��2��d"����I� �.�j�^7���JP�@G�0+0B*K��a�7#�y��է]����oN�����޼M��}�#��9a?f�����ٚ��	HVyRF\�tw8��VE�����S�����x��V�%3r=b��#_�܊�}2n�Z0'�3vIn�3�mڝX��X�%�>��n6t|8VɈ)9��Q{%�&/�Ņ�9�\Qz!�6os���bK߷ �J��U(h���FſB�5�Y���?9��O"^�����T�L�c$�WF�I,�̠b&�_��%�Ab�A��6���W,1X~*ANm��f����y��Ŋ/�Yr3C�}�D34DM�WܬY�j�w���	UĦ�h����@y2ǘ?"k�DZV��u`�(��@Ƹ'���u���D��'M����ע[N5������1ax}ӖL�)[m���P+����@�?��D�Ɯ�0c9�����J�Y`z�K�a<�p=��'R~*����,����!k�0���cY�C��x���?L��"�Y����2
�k1r QPB�%\�!���
9#P�+2E�����"�Z�X#�~҅lg�ӊ+ꮁ*���Lb�B�bިxo����r�1�	�9#��5��ّ`�@��bRmˬy���PqH�]�v �HfU�͘�Y��y3�z	�ybU�Y�mz���Rۘ�'[���G$�0�E�S,*^}9�$ܢ.v\��N[�8�8��ŷs��,�f�վn`�Ԉ��/��O�9� ۛ.,TX�'o�/>��4j�A�3?�����'�|�KѮA���:+w�b>��ǈSP�*�S���,e^�c�i�9;�������qs�����'�*� ���G=���S�9���D��~�Q'?�L~r�	B1;��1�"�)�¤2��z�'E��H ��&@�	��\�h�
fDB�F fw�I�d�P2�lࢆ�	����ɽ 0�;��B{8�Y�'���k���¾��Cɩy���-On	���O,e'�ȱ'`G�f|�}j�H_q��� �16���)�C�5�tDA@Y) P�a�`ɼr�4�X��	=L�@!�Yb�%�$E�)'36���I���$I"�ĝp6k�|J�@��ĘO�l�2���6ĉa4i[��(���N#}a}B�i��QWa�3�* �a�hQJu0��P<5��8Q��2Z6\���L73o�'t��>��d �Y	�х/���ՠ�J4Of$�&L�(�PP��q66�;B� ,[*�~��2,	�<�`�K�+�H@��P��N�ɱ�iPBy2��c_�=2���&�꧃�$��u�29!�G	��g�Y�O�qzFeV���$ڤl�8 I�VA�G�$��G_�J�0چ�4��qG~�� �(���;E�E��eI�
����\����DIyޖe�,�����
��'_���P �= ������>,���@JO��<������#�ߚ8� <����?j��
"��$R ����'4|P(s�^ 1,$b?�� �ٷ��8��1c&��:t�U��Ϝ�$Pɧ�����N]Fe�n�2b�b,��j֋ �!(���a!*ޢ\l漗'|j����8r���&��Mm�|nڧy�T3�G�Vd���c͞{'��'-�'�,BWEܴ_aڐ��J$�D�	9� z��7PP�wOkդ����w�0Xrm�=��RE�?O�@�? \@��ʕ�/#�X26�Y��z����O�}5ς�IN
9��4�
�O�LdR�$�0=��i�#�-;� �Te΢�=�O�F�r)6�I	0�ɻ��D�4�d� ��($&���=�e2S����<pe�|�Q�A@ؼ � �7 &��"�M�OD ��+b�0|d�Y
�~��ē-��� ��ZP�§��a�b�_#H�J�5��D?iE��
>I����-��р�2쓖�,[S�%���Ӧ"Z��)���1�KR�$I��(��Lsf)�6ɤ$:�׸[V�"�4'R�I�cQ~��a�hb�L�=�Ͽ���[�
�Y�G�a\@���KUyyRo�?}ȆpQb����,Oĉ�5JF�Y�b)����6����E��#�O.E�'Y�f��1�̏J~��O ~�R.�&_����%���`���_ܓ0�Q$>�-������3J��e�A]4]���zV6퓴3�<*䨛���<2D��J�3?Y��b�� �Y�2�f�0r��8[C&A;d+�-��)wg���6��I,cw�%���4�IB6���ַQ\�3�Q�"l��| n|���8�E�3Gw�q�f"�~P<#mX�E�>Ysp�g���[���ռ�+�m��]@��յ*"�Y��u}���-�Ts!ܲ|/��M�OV���w�hN��oe!K��O&�D|��Qgt�r׿T!IN~�V��}T���%��jК�@`�$KJ���G�?���+D&�@���ږMX�ē�19�O�7PrY�0o'gTd�͓Cx�	s-��Ksvqp*Oq���w��&f�B<J�E��-���H�>�f��B ̳4��D�ad�QDf&,O�e[Ӡ�X2���6qr��{��>�.+,b�i�jə,�U� ONX��è��D�/a�>Ab��00�l�ѱդ����4B�p�`�\1�����V&=�9�3��Nv��7�]^�e�A��3ם�<E�DnW
5� ���D�.���j�̙w�ax��l��O��z�.�]��;A��<%�Z���w��+��S��L�Q��/�S7?i�ORiz�b݌/��E�NZ�S�T����'*J�Q�BóTB�=��kʊKp-HC��*D���A"�.�&��Cؒ��{���T�D;�T����ؔ��ըO��C�Z�@d9���m�� [��O��&R*���$
�Q�Pe��'�B��D'��"��i�S�կD�b�hL���6�\�	qO>�u�R�Ga��u���vd3�O��q��:��d+CE�4h��f��K{qOFd1V`��}џt1E��pM����MO�o�����<����4��*�����-�ҍD�s(��	���e�'͂m]�2�V�\�z�)�N�>/������~�+\�4Z�x���^���' Jz=��$S��H��b�2j��Їȓ$��5����:fː���d�` �(JF���0%�(�OL� !cO٠E@@���H*�����Ŷ��Q�G1����ɃX�F�BV��}¡�U�R�*7F�J��J(��$��QhQ��)�xGN���>��"ſ7��)Y���F�`<@�ZQ�'Ŵ�J���;�$����H��'��8�h�(C�ԹKPa�4Wp�y)��c������n^�5�V2:v�U��ԛ?k�6�݋ ?F�HBϞ�
��x�o�O�b��i�C\��gA�;k�r�j�
��yv�(##���\Vd��.�V�Щ�e��b���9v�̣/�D�c�B�}<�ݠ'���#�Ю�c'�} #���~r�� z67M׿O6��Ȃ�јth�4*����c�a}R,KG:����;rl���t�t钿��R �i�m��	�)��O�� �iФ�5�[�O�Z(�ǆl���d.#����,Zx��0�;ғA_��	��1��S��MìO��u�իH�H�s�e���O^|�\��F @�yY�A٦oL�[,�I@t�p�$iFM�J�>��&/-_*��l�dM��T��\Y�Ġ�CU`2�Ӻo�?��*�d�Px!i�/{4i[�E�d1�Ĩ���W���O��%4�Hӓ	z�V�&S��]�q��R�X���'�0��n�NЁP@#�u7�d?�|nZ�6�: YbA��#DHbȕ�z:
���K]�ڴs�i�?i]�I�T���ag�j�IK2`����M��l%����F��
�?Im���Xwڒ�m�08�KOx���2a!6�j9E|�%� FG~�'ɜ0��Ӻ#񈈘g��1 �T�CE�M1R��{&N9C����%	���%>�ˉy��7r]��2�ފ��d�h0�~��ywVe
�4��)� w�`}!FC-S(0* ���Ma�=�фS��4�0�
��Bb�	��΃�0=	�\�F�hӲ��"T���3+v����'��5 H��-��IތX�#S)z��)vϻiTR@{�	��!�䂆i�(�P�,E?iٖ���B�n{��
�����aQ
:H`(�ខ'�(�R�$U)���b��z����@M�4��.4H�X
v�F9q��(KW�'�t(JUܴm�b��GE�^^~����o������On���ͦ7,p|� ,�41��^�y��n�{���b&�ނ}/HL���4��iE{���E����l�;r,=�G%E�A�YR�"V�*��X!�5M!>-�fW�oab�6���Q�HQ���2Q�az���*X*��)��I�P`%��?�w��0����h5��AX�̗:�*��!��_ɆQb-�5����	� ��#�X������Ͽ_��	�"OVI�f�҉<�h6lִv�J��a�
�������Lh1��:!_VH�b�©]<i4hޤV3ʨ�=��	��A�J��Q�Q������I�LbT�ֈ
�R����bL��FNXڴ��T���b4��>\��UI��F�v�~`H�>f�
����O��n�j���4!n�a2����'� t�)��_���:"�S)9J�míO���C�Q���P j>@P�y���i[b�9$�KY�Dl�R'O�f���!B�T.�� ��]��$�Ua�
*�"I�
�/"� }��D�L=�v�&n�����'oΆC��܃N`�P�i� ����0#Hz�y��\*и�.2��o��PA.٦6�p���v����?�O�ᢣ�T�>�"	�@��:0F�`�P����#��Hdx� e��+� 9�nհ^��'��f�0kV��/� -��&��q�����gL+$�L8G~2� Y��B�Kݿ#�!�fƑb����El�#��%���F%�ڵ�CE���09`�Q��eS֦M~�T��C`�CV$���6�I�N��r��f�09��L*�^� �4r��Yg%���.C��v�Q'X�trR*�./��r�͔*K����ÑS0�q@C���L��`i�*�<;'Dpaz2�Y�K��r'��x�8e1���^S%j�H�2�6�L���r�cZ�����P�d7Z>Y�w	3�4]HĹ��� }��{���<x���ʚ�K��pZ3�*]YN��$�O���U��u#��Б�܁/��0��@�}Uq[1�:}�6mA<Fߠ*���ß��r�Q�#L�k`i�8�b�*��9�I<?1xJ��ǷCO��c�Vk�0���_�$��}8�l�/���d�A=^��v��W�6� ���8,&���S�n�.C�JæQ��#>a`�-�����O#5�F�M.F��ـ�Q�.-|4So11P�ab�=(N6���&���#"��\�k�F+e�����
��	B�x�Tf�=а?�U��)o˖P�d�f^ĽyU#9���`�+��M̻��A�W��)K�Q��y��]�PdT�ab\/��g�]f)t�BV2 ��yb�M8&�t��F
F`kF��Ы�L��!��W5��bM�2�*�˰A0�x�qW�6�"ŧ
�l�!��?�I& B�mr�k�NU�xB�ϻK��O���"�ڿ78�� LЇ-.�L��O(�xu�۫,��&��<�J8y�GJ�g� �:�e�'.�ȕ���7�$�z��'��D0�Fv�1!3��Cf" �a�\$q�Pbb�#�8b*�{�HD3å���� �1Q�7�w�.	�l�l4��H��C07H���'<����O�A�ơi��ES�h��`+HO~�g��~B�U&c�X�� cе�箝�?t�d1 ���Y�֤ׯg��iSD��\�c�'O��׮�v�+D^�X�� uܸ���l��e;��G
����W�}����OD�#�x��D<5\���"�	� �@P����%���Ұc��)��O����i�,c�^��8*;:���@�-|Z��10�@�6�<����"_(����0�7/s� �'aT�Qmr��'�����i�恙S��?K�<�0V"�O�py��e��j����>���� ��M5�(?�]�"D&se��)�����gcB�ɻ8���T.;����V�o꼉��<>J�7gIL��8�V�]-m���C#vE0}ZGm7LO������b>�����O48Ȱ���O���!ʣN���p�"O,�!�Ҭ������r�AG�D�;�ҡ!chI,ሟFk �X7?�|TmܲAؼ�+��9D�`�FM�$8����J�i�I ��-TtMC�{r��x��E�����לq�jL �F+D� �"o�&�P@c��%]|���Dj�hP� Tx����N̓F䮈ZՉ� 3F�20.7D���#��(�iJeAB���I�U
6D�P�� 7������-s\@q��&D�Tc腌WY��
�	:�ZP��,2D���"�G��&�r�h�j�p��3D��( ���e�」=E[��ad<D� @U���2Di��J�dIJFh>D�8���������V�]��}��)D��S�hջK��ٙdϵF}�9p�-D��j��[04��1�c��$TܐW	?D�h����	y�x��PoL�w� Dy�m<D�4��a��O�IQ6)'�.�K�:D�"dO��4
�����e�$re�&D���pN߸e_����D�/TӐ�Q�%2D����K�bH:E��GS$^��%�B�,D� 92.�Od@�J ��>��	���*D���퐔:������c���FO(D��p�&97Rx��I��T8��;#1D� ;a���܍B@dQM��Qq�c+D�@�P�L>?��%�C�W�����l�<AE�Ϗl�T�vo��\QD�y�<Ag�$	�Ѝx�l�"G�Y��^O�<� :H���..�<M�#&ЇW�t�"O�B�-�-���yeX���"g"O�u2�5�Z����L�N�n� �"ON�炑�lnV)��+ �%je�"O��ia�w��5���Qa	�L1�"O���Ħ�imԭXT�T;n�4�$"OB�)�DȮb|��j��G?d߀�*�"O��ƮE�BF[ Q�}I�ˇ@h!򄁗hj���'˨8>f0uf�(W$�x���92���ɋ\�^	X�.��xd>�jGI�O:B��)S{���!�8%<��jGn�B��!E�A���	vB�-B�bFTV�C�	 R� G��ȥ;c���`��C�I�V��x�)U�P�7�W�m��B��?��xC�L>|^���T�nB�	R��h���էR���
`�,`B�2a^u�Q�ea��ꦪѹ/�B��LB>T�D���>�0�s��C��O���&J��I �����3U��C�I�`AX�q���'M�TҗȐ�)��C�	�"��8f�Ү��ě#J�cPB�ɶ&FB��ҁ�?�T�c��K B�	$W.��G"G	n�r�r��	w�C䉎I�T��cʂ`�8�bt� L�|B�I2a�$���E�"}I`��MbB�I
F�.���[�B�H)d
ԖK�PB�I_}��LɃ>����m3��C�I�,�HԂ HQ�>ݮ(0��(][�C�ɔF�P�"�1��R�o3�C�I/$9�A��D6Z��ٸ���v��C�	B{]�u��F�3�HYv�B䉐����	�<e	�h�jq�B�Is��%�AO'ĝk��׆)ΪB�	%z�V5��,� *o��y��5�B��<�D���ˊw,�y!S"ӐU��B�I�L�014��9�z!�4ל~gdB�:GX�)��->'��C�+	�FB�	 >�.`Иp�� 95a��z��B�'?��q�0��"�$��gݸ��B�	i�ڜ WyO���ZW�C�I�t5j&@K��,i9tM�8dlB䉆�b�Q�b��
uL��g�F�C�	>
��:c�)!4,�$y6�B�zW|�����I�CJBm�ZB��= �nL��ͼ1$tx�C�;rBB��-u��RA��i}��2�*�?+lB��$?]�d���|ك�W�L{B�I�p���d�`�6�[��Y
u0�C�ɞU�d���ƛ� 	x��){�C�Ɍ%��؛� ��(�$���-�(2��C�ɒ%�(�3����Mi(e�$�ԗV,�B�		N Ԉ����"��r�d�1-PC�ɩz���3�+#���0V�O�G~(C�I�)��JQFĢ/�u��\��B�I'y̜!�cߥr���B-܊j�B�vvD��@ը>�*�3%�E�9>�B�ɥ`N~z�Q�:�f r��P;O�B�	>e:4���"�p%nu��(�`�`B�i���1���* Y�"%=7� C�IG��Br��&���˔��eC�	��iv�6E��(���'�C�Ɏ3�Y��]�?q�x���D�g��C��2��{�a�\��Գv�";�C�I�9
m�g��~xl� ��"5��B�)� �4�&ɟ�I���haM5#k�d��"O��aSg�@E�0x�K� 8�q"O`E�� �,!7�T0�4`#�"O~,����K9`!i�o�3-W� ف"O D�r�HjR4�s�ŏ7h֑!w"O�����*C6*�)��
�sM�E�"O|šs��0��1��-�\ �"On99Џ�0Z=z�xbk�H��� w"O���r⃵$�h��R�H������"O�q뗧��)/T�H1�=9j��aw"O" k�8b\C��DK  z�"OƘq�Z4�"��g[1��|@�"OXU�R$jI���ݹ�PL�cj�+�y�Fʤ2xݑt  A>���*�?�y�՟_,�XYT��.y���U��yb �$��M�c)A* ��I��=�yB�g��h�KƐ(N���!�y���2 �8�欟�N�:�@��y��4KP�w��#t��틥�%�y��� V$�1��ѹ�P�$BU �yrk��F���;�ȵkX�p�#��y�a��=��cS���V��� �yR��tB֬J��أO;�!"� ��yk���m0�
@�G���P5/���y���$i��QLAzBԳ3B�6�y¯��x���$��:��QC���Py��	�2c�w�A� c(��!EHJ�<�P �� �9�B�+;O�))���_�<�&i[. ����Ӄu-H)a��Nw�<����e��
�L��@9KD�UG�<QF �|Ȍwk�O��0�A�<��+�)
�Hp�O�I�8��&�~�<��)ȓ@I�r��@ &�](���{�<�s�9;ޔ &�֘J�̰9�Ay�<�!�ӓ�:`��'�-b`22��x�<��E�$t��dHE"$&�yb�@Sv�<�cB
M�fԒw�֜"�$�z��{�<��mÑg� l�u���ּ���y�<ɣB��)�H2#��P%��_k�<�w$�a��*S.4��@h���d�<Q�Z@t�:��&]����$a�<)cD%E�4�sGɧ�P(0僗Z�<Tٴy��gX�N�����U�<aʁ��~hw)<p	��e�<��aN� Av@Iu$Z2j&Mї�Pe�<�Ä�N�t������U��KB�YL�<I)�<\XM��-0w�>\K�_�<�UG/G��ERu�.�zT��{�<�����36	اE�du�(@%%y�<Ɇ	Џ6�	&OP�w��8Z�a�j�<���#M�X��TM�)p �
6E}�<���60���*�F��1)t!��+Jx�<y�ͭ6W�`�6(�'.�T4et�<�!"-�Ё1a�=|&�)#t�m�<�c,�C�fQ�ݰY���B��j�<I��Z���1`��}q�ȡ��{�<�F-�
�H�������x�<I�B�� �^�0l�h���1��z�<qE�X,�(b���4�!u�Zs�<��ߍ;�]��!;
��,ٶk g�<)B
�!��!Y�ʁ�R�PL�։W_�<q�A�%t����/I;\Z����q�<i0�T���� ��ƺa� H��+Fn�<�!N�9����(ݮ:��p�$�@�<� Z�C��D=!-��J��F �`U"OE��'R�/ػ�鉁L^�Z�"O�1��,ߔ}0����PY�"O�œD��+� 9����!��G"O�a�zU���αA���6kWR�<�B�=6�qҥL�~2����,�V�<1��C�DTT�@��6��uࢀ�O�<��E�#�h��8A�<M��`�<q4`�� ���6AӰ�c�c�<1Uh��Nd�4ς�p��̓�'�_�<���xQJuI��%\H� �҂D\�<��Z4Y�D�0Ӆ�A��ف��U�<�3��'�*"R#G�z��5�Z�<9#bA�?�I�e`��#"�Tp!�L~�<Y���?%�4P��K����&b�}�<	'k��J<�IiW�Ϛ�@A�x�<���W�HB�k��e����% K�<a��)C���lʞN��(� � L�<��CC&Q���D6g^4�v���<9u��j p�pH��b����TE�D�<هN�7A�|��Ȑ���!��OZ�<��EQ6�Zl3b�P2� �RF�k�<��)BD�`�DHo� ��i�f�<���%C��5�6��H��9b�g�<�SnN�p����M����HG�<��Ț �����U|6�� �K�A�<ٓ��6#ۺHc�g��@n�����~�<b� Ym(C¨"(�ii��O�<���؞F�9yc#Ħ^l����a�<!!��1���(T$�ȶ�KY�<�¯E�/b� I��RyC!FJ�<�WbS	K�:�j�@S�1�$	s.�K�<����z� 3nۡ_���RV�a�<U�O�=<���� 7Xx����H�<1�AI2H���d�Q�v��\H��E�<���s� ��P���V�Р���u�<��'�,c� 0��Q�q���A}�<B�A�|;*<����q��DSƬ�w�<� �̓Wy�B0IF�_`,�*�|�<�i� �v�e��dc�1!fO�O�<A�C��|>��m�7i>��%I�<�,�X�����`~.����^�<�0��8�124��v5j�X���W�<�W�a>����i�(���
R�<�4(ˋq�pꢬSc�E$M�x�<���l1>�X���+5�I�H�u�<	7�X�Ty�Rt�&�&�P$�{�<qV��n�t��C��%g�Ce�Vu�<�ƅO&r�P�+r�"iv�J�<�+�>/C ���k��v�Pd�I�<�'��t��f
��w�aW��j�<qS�,J��L��ES�B�!EL�K�<����q6��y�(�*|p�-K�I�<���rhZ�c�˘�Dg�Qz�k�_�<��*KU�"��"�W���Hu��]�<a���:���u�^��R�<�X�3�j�3��P#_��H��Ds�<�#�V>TȄ �c#B����I�<y�g߽0�0�3C�Ci4Ĩ���B�<����@:ds'�9D0�p���z�<a2�U�W��@��/dMf-8T��u�<Y�@%��Q�ާXu�M����K�<Y���(�(R� ;��g�@�<�@�la�⩝ � ���@�<� �m����<�tYy�Ǌ�7F��p�"O:ժB�_�bΈ�FƜ[/<q+�"O*�Z�(ʼֆ̙��A-T)H��U"Ob�
R��������4|PYC"O��@w��f��,Y��-e����`"Ot�ArE�)p�n�PL�p"OD��f���,����*@� �~�)1"O���H�W�^��2�����:D"O*� ��N]2l��%��3�l��"O��A� :�N]����l!�,�"O���d�iAd c�E��dVQ�D"O�ESv�L)�Ua�ڧl��c"O�+��8w\��(G��e0�m�"OT 	�  ��   "    �"  �-  78  1C  O  �V  �]  �f  am  x  L�  ��  ԏ  �  Z�  ��  ��  ;�  }�  ��  �  H�  ��  ��  �  N�  ��  ��  �  a�   o � B � �! T( �/ c8 �> �D )K rR �X �^ �g  i  `� u�	����Zv)A�'ld\�0"Jz+ �D�/g�2T8���	#Ĵ�#ۊ�?Y�� ��y��%+|m�֠�&Κ!���ԓP��WB�^fХڡI�'@xV�P@fO)Bu�] ��F�+��韚z�n��Q�ؓ>�j��U��LdP��Rv�<H1��Ȳ5�Hr�U�ѭ;`.����Uۛ6�\�{jS���!r��9r ���B�H��B86���9֨B%\��E�'�3[eҁo�؟L�'lr�'@�f����H�*��B@�J�b�'�:6�շ7]���?���E ���?�$ϛ�8@�����P��p�f���?�����?��&�^ nH؞X�����p�@�"��n�EY���o���@�V*��d����'�,<�E����'`���R�C�eSt�J�0gXM�ui/!�I�<���2$�� �� �5E�䁱y�^�S�l��R�r-��R>IpR�'�rw�(�d�O�d�O$˧�y� �0%�6�Q��`���qgĉ��?���iJ6����ߴ�?Y��i:��Q�w� AaːE�4(��/նJYʀÁ��,�#Q}b�'@��'O��ۇJ�
�.a��O�?���u��P�<��(0��Z�T�#"K�?j���W��g�01@��,�?9��i1�7��lQ̧��^w�:��$���'�@��#�#�pT���i0Aq�O\=xp��X����Zc� ��U
�g�oڄ�MCAi�4P7jxk+Q�
N�ӄ�����q�wJ�h��9k�ir�7mF�A��%Z�X���b�
tb�m���\4Ÿ@�*^D��OL��8�5AS�,�A��M땹i�r7��g� �
ӂ��Pw`�C��v�b��eF��t)��T�R��u��/WަM*`ʝ�.�n}�4n������H�?yTEZ������ qa�J�=U�ˁE;�?A�'���O��D'I�B
�*��"&��L͵;�$�v�[\���E�jW��'>���'\b�'��1Ku�Wjq>Lғ�}Ӽ<�5�ƨp{E*h �Z¢5�A}�� ؚ?aH�۴u�p�z���'�t��Rm�,���Pe��0<Y���AyB��<1�d�x1�s������v��џ8��ݟ%����П��'H�+%�V�#R�֯NʚI�ֈE���'�� ��F�.y�'W���f����l�c�O��|��@�	*n������O�˓��閾i���iy�I���?8�`[q��!������O���"!��j�M*p���lZ�%��⦭�-�P	�����ppQ�#��䜧e��qrdǫW�x�7c��%!f<�)�95��ś�mU���:�"΂'���+��ܦ���q>�cB�E t�A�+�<��p��$���O �$�O@ʓ��O���$l�1è)C���z_>�k��d�O&eo�	�MS��j��3�,<Ѐ��/zd�C�Έ�1���p��bӊ�D�<�2윃�"���?a���$[���m�/8 �B�jħ20�谔K4'��`K�!��Pň|� �|��g�C���P�"g`Z(�4�M�9h�����QJ �X���V��X����w�<�-���`m��E��V Ȇ�.޼�qLI�\6M�hy��U��?������|�.�/*��Ҕ�Z6@�H$�+�)]r�'��	�@��O\�"`�CR��
��O����9�'p�
kӂmk�i>!�Hy��H�J�Y�NS�0J��S�֊}4�d�� �yB�'���'�H��������`p.��G�.i����^Av�9 �ߢA�*�Q��U��X��B���<)���~d�TD,�Xb&��Bn$D�$g�XC�&��Q�<X`���X�'��L���T�];'�ՠYzu:����?��i�
"=���W+��Iǧ�2U���]
2uR^�P�Iş@%?�@���xH�EC��v�
<	7��O��m���4ț&\>��pG_'�M��?)#�Ґi�ISt#	!hD������?�%r$���?Y�i�j���K*O~�!��˒!T��n�r=�G
��e�y��"F#~�X����'i�ʸR�H�'�i
�G.~�j�rrb*Wr(�E�Gʍ[����W�4S&�ߒg���O�0SF�'U�o{Ӕ�$
K��m`��M�4�M�Ӆ���˓<5�8�����Ӻ������j���q�%ʛ3�$ v�%��'�ў�#�M��h���ԩ9v�»�x�RU`T=D��f�'��7M��g�L5l���':���O��͑`�-0�Ҳ(.����#*.���'خ�*a�E�No���.a�,t:#&;�ӟOt*�`�B�(�*3W�3xH�'D�AUI�;w�T�1B%0$��ISR�l��� �s$*"��#Gl��������F�O�0l�ħ�O8P`Iv�C�6�h$)�4LA�dJ>���䓗Ob��&!#�����]�u�N�V�iM6M�ɦq��4��!tq�gB�3�~Q
5*I�bi�iXS�i���'�+R�3�4��&�'&�'�R7�!��S$!��J�L�2�P��7�>�|���h<z��tIY>)�3�m�n�� C	J?4�y�I]J)��i�]��ge�-�Y��؜]��9�O \�#����y�N��fê�cgD�Y=b��G�$�u}�@ѣ�?Y�����?���K��(Vk�m�(����(?��8O>���0=!Eďj;0ZD��8_�X��"ߟ@��"�M�ֻirB�v�.������)�|��]���ySa��w��Q��DСq�K�.�ĸ�	� �	ٟ��\we��'h�i�U0!e�w�<�f*ݥB��O��Qb���'�D�f�P���f,�B�!�d��'�������h��J����A��'	*����8wĖ�Z�$C#S|��0�[�KY!�D��K�8(��b�0\��!��A�*@�'{6"��͵��4�Or�[�F��UO5�>]��F�UN��'��9�'g�2�� ���#����0�RoGvQl:� �� ��~(m�+��bX�xrU�'N�<:��i�t0�Q�6>�0Y��B8j7*P@�X'L���@�[�7��E��� �D�O��9�	���hSn�y��Ձ ��$����@��X��`X�sn@�G�G�K"ܘ��/�	@���(�Ol�cwb�!��9@"������u�'~�I�+� ��Q�'zA��Z��"lI����i�m�6da������?)Qd��?���;u ͫ-��l��&z$i��Xm�)]�6� T��OL�-`�r��]>���-/�|�Z�(1Z��f�~�&5ز�N6`�tm�PA��?��Č�� PVaDW:,�ђK7?�4�����	b�O���θsߦ��D���[��!�$�$k���bC���
�&ƈxDў��	�HO�*vGϥj64��Eo_�S��������I��I��HZ�J�ݟ8���t��ټ���0���q��8R���ٜ�@�8�4dP�@7f�20H8�*�B�����y,�䢐�Vl�P�䎒#c$̑$��2
�(�Q�+A"KEr!2�L�$���'t���s�Ra�ֈ&���8a@��lR�4�?Y�$ֲ�?	��,O�dȨ3e
<�E��'�L�$ �CO��$�鉃-��#�����\�C�UP��'���b�@�oZz�I�?��S[y��9ިX����;����(I� Q��R/�R�'���'���������|:��
�SH�u��,N�tܪ���M]�TўU:u�W/!�(p(ܴ=j9��	8$Ѳq���=���;���k
��Q�˻���� S���U�'�8"�dpF{�郤%J,�&�õ.઱��됑)��3�(��EP{�b�;T�jj�`��_��=��y��+~�@4{�oܼh�&�ЇCŬ�����|b'�X0:6-�O8���rD❈�@�,��Ua'w��$�Ol��r!�O,�Dd>��cFʏ7>(dD����kܴc�`vcՄ5�����ƙ�`q�j�RX��<w#՝5��0(�̄ ���F�iC������8C����o�BE���`�Ԃp���Ey�Y�?���|���E~�����( �@�,A��y�LH�1q$��W��o� 13����?!0�'�4��o͏P�e�Λ�w�;O>�%M�v���'o�^>�J��ܨ��@�9lԭ:�Πi4���c����. .6��	H�S�L<U��	�t5�g��&������$?Q�I�x����tAǇ;����H�/!Xp�暟��a�O��$�"|�r(?���{�↸}� 5&�Q�<�ᙾjʸ�Іhװ���*�J�'T�}����[,� ���8�ಯ���Mc���?��R��|�����?!��?����y'��<[t!`�`Y {�@��$,[�9��ap�
kB�$,D:A�l���t�	"�u�O��W"�n��U����<����F)M��f�o�$�����-b�����A��'�u���w2r��'��P�&�����?�:�`�|�J��?!���y���/В`��
K8R�Y�B����y��_6R ���Ԥ�~�9�B��?��4����@�ɞC�i£&[0T��1S�Y�{��u�T�_���I��L�I�T�[w�r�'3�	�Hq"8hv!����Y�C� a*�	cO�Ax��m��+�*�Is^ ��=�+aqHEΖI�l�˳D]e^�I���6`�6���mv�)Q�'׌K i��*�z"�����BK�+`�H�iNN'ufjtۂ����*�1j�O�9���4eN��v���~�|��f�M�V�(�� ��$k��k�͜�;�����X8sgڒOzXl�q��$r�����4�?���e����NǤ<:��&�Ҫ`I����?��dޚ�?Y������ʿkH��5f��e%l)��Gp�I��.�
AYX�F�W�2����< ��Ey2,V
sY��D�e��]��Ѽ2乃���):���%D�N���xdS ���Gy�����?YД|2��Ȳ���M�92]i�,��yR�Eu��,��H�Ԕ��"����?���'���K��K�q7�X"�F�;����J>�ү�����'0Z>�R4CEןtg��f-����	�8HT��矘�I�����䀛~ОH��)TA���O���I�p1R���Hux�Ŗ���S��0 
�G�X6k�7V'��"�d)9	<���_���T/b?xK��*)��E�fcWW~����?��|��	E�����'x��y# ��z!��جkn��t&R
��P�ɩBў�I<�HO��� %d����d�]��C��{}��'�BL�7F`H��'m��'��9�6*���Y&2����H�ƀ^� ��ܑT�4��0��-՜{���?m# ��*`"�ɏ���x�rC�m �j�-x3L ���P�hAhd�D��E%G�%�
�+�}�4hBݼ;$�I�z��F땭E�.�C���M���iy�KQ����Y����8TNDd;��t�4}ʗˁX������L���9.*�yGSd8v�h�mѢG��d�O<�m���M��@���'����O��D�`@�O�ABl���BK�[�	�'����	�@����H\w)�'p�i�<6o�M�U�˯"����viB� v̍���S�I
p| ��6|��	Ǔg΍� |)83��3|u��i	��" ȗ�3�tD{�'R�[Ѵ���O��;���9�n
�	ēO��m��`�4�j�O��eʜ�n��$�O4�=��dD)8k|-�d&�9P�\�P�C+��{��$H�;Ж�:I ;Gv ���ؖ{��'��6��O˓�����V?��ɺf*�"�N�:���Y�bѾ4$��ğTHRlH۟����|2�! ��h��إ'U$b�%�R^�RV�R�����C�NB����-�MZ��#&N)nxq�"�K,HKt��+6�`T \_�`re�}G4�>�R�^���E~b�B}P�,`��>���wo���0>��ɮF��G���zeX��Ԭ�g����� !��N�#B@H������Idyb!�f�6��O`���|��,͓�?�$oǎ.)Na"��� ���!��?��*���CJ��Y~"՘���8H��*���-�}X� �#Y�v�2+56���'�
=��[�]
|�t>)j� z��.�E�U��A(����$&q���$@��1tPB�����@T?���h���I�ӈI��/ّ�0��c�khB��3A�����▂��p��;ޜ�=A����`�QG��de���hő+� x��)��M���?1��:.� "OÁ�?����?)��yWז�hD�P�˕kl8r���0�0u�K-�`ظV%��3q$As���y���lT�$iF�Q2g	��)AG�'��b��B@%ġrvC�&tDY0"΀�V'�SC �l f#d��da��,�!U7��S�/�Oj�m���OH�=�(� H$v�����4D8���cK�y��͸5�����Bm� )���<i�Ar���S�Ԕ'�:I�GLke�9;�&�+i�f�ҥ���T�nMؖ�'^�'jrb�~���?�sD��*;�܉�D�`�F�ʡM��UB1��D
	E�d��	�K��f�&��Af"F� %d�R��ؔ.���B�V&�d!�
�!=D�D{�ˁZ��!@�=C�4iX�#j�("G��O��!ٴ�MK�����<��I3�ïvXF�����찖G�\�<)5���i�.܋B�
���B��M#��ir� 6��Iɟ���H�2=�Ek�&Zp#g�H+L����p���(�I�|z��^9& �d��JL���������cU�b[@����`_��b�3�W��SU#į3��lz�#�$�����بcuԉˣdȮu�\���O.%o@�>fG]�$��q~R��4%�.�v�øN�P��L���䓟0>�w��/-1�T�R��1 m 8�[7���G�O��a��33ԕc��YU��2��'��I�^���	۟��	B��Ua�h��|��E�Ef�3��H�F�Pr�'t&}�m�]ha����|�8��!<���?�(.���XSR�n�@S �'?yC F>������	�B��"�&kD�>��6�֪�|���lљ2��$?��-러��D�O&���O�,E�b��2��>l{�l�ȓ �LEё&O;t�Bq1`Z;U�8\D�8�'y�.1*M�uȲ�i��O����I���Iҟl�P.�.g�4����H���X̻m<�M�q�mP��)��"rv���A�.&���$R�#X���a�A̧��'��O�"m ٓ�Îc��<4,��1���!�Bܦ��p�ǋ��O��<�O��)q��6]9�ܛ�E_�{���P�'��I?M�F���O�=9T�G�J,��sD��� �����!M��y\�"]��y򭌰��	�RF ��H�����'M�6G����*� s��H �LSZ��P.�?�(=��ʟ��I��H��������|Z�����ĀuЌ
^�T�s�-a�Mk��kw�I���N�Ul��=��&� �M(%�JEq���X���rCP�w��=cQ �� �OG51ʣ>AgK:?" �wH͢IZ1�D��~�����F{��I�Wǖ�I����\J0���-��!^�B�	=Og�X�R�^'EΠ�P�	�!�z�O0]lӟ��'%�����"��Ԣ^��օџ��1��#?���'qPP��'0b<��5�����F���{E�1\�L @�ߛXg`1�NՎu�Q�I
:}$DyҢ_l����H�?.�q�:�fyd�=�䨺�g\�S�=�D�ۿ{_�iFy�E���?)������'E±��Z/lb�{��!].�'ja|"�J�M��$��&�q����?���'�x}�6�#?�vU(r��>��1�����Ty�Xoß���J�DB$'"��?K �4�ԉa�:��"�P�#��'��!y�����E�cdqӄ�!�o�|�Οv�f��*[�z�Hb���Z����cRB^5,~�a0�
N�N��A[�-�*,�&?��I�6!`��
�@��|fL�!a'?�U���$!K>E�$e[�f��V�Ho��YlB�	�2�hD�N��s�ơ��d�#�$�=���e����� R��AM��{�p=�_�)�I`�'Hٳ��
�,���x���|�UA�g�zM ���8��٥,ܢn5��
���R�XY)�+^�^��|A� j���	�pL̍�ĥ�A7|��1)̈́j�)�P3x\����G��T�o<�-� ����O� �x36M�1
BA�4�E�6Ũ��`�'��	
3m����O��=�����UHM+�͋�Eڂ�y��=���X��94�ý��^I���T�'N�ɰ	��Pd��q�T�Q��i�����ݤy�I˟\�I��X\w�'7��ȔS�8�kɳ?�<�b��*k|l�ZSO��Z��D���ro�e
�s�	/+h��f�,eL"D��ǅ)"B�Ყo]6b��YS��̘|�Hcٴn�6}���<ʓ[���;ÁJ�z�N�:���(Ȕ�C�)�ϟX8��+tvp��ϐ9�R���?Cj������"E,H��&X�2Ϗ�X���%��Hݴ��q�4���i���'��i���\Ydو�bߌ�L[�'�R�Nn!��'q�Iݾj��� �$��7)[�|(�"
"X)���T�V*-�R�+��-O�}+BbܭCߎ�(elS�Ɣ	Bp�p��d���uѨD��MO�9)�h)�&�,I�����X�9ceb�*kbxy�B+�Z鲝��e�v��������!T���?��4����I�Y���+җBy�Q.��\1O���-�O@�?��&mB˟@q%/�)�؍�"˦b�lysG	�̟x��<vDZ�S��R,D�
M6)�)�*��V�;V���O����#�[%t�čbăı`�01��OV5�Vn��s�\�
�G_	>D�b��#a��,IM?)z�f�;{l�ĳ�K�H0��!?�WOWϟ��	O�O�Uq�
T�@���)$��j�!�Dϳ<��q� ?z���5��-6џ������A�C�lt�XRD�ժg��'$��z�d��B����	ş����|2�T�DCX�ۢd	�4F��bE�Pp�!9'��->dP�r��/W�%�|ʑ���8T�� xJ��d���q&*tb�I
_@����X�~�@(������hF��1���SB���~b*]4�R�YVg�)4���aQ#���?a�O@Y��'��퉇:���&+�
(��ۆ�? �J-�ȓ($�`5��5F��+�BG�C�@)�'(#=ͧ�?/O�A�R��d��I�&� [�x�	ÅUv�(�M�O��$�O���V��|�B,��Xh$uѠ��1J�`E@��#t����FS�$�b����Yow�(B����H�<��f�Q1<i@����螇 ,�r'���q(0΅�x�$y���R6A^�6̣:kO
u��n�e.Ca��H��ǎ ��������s��⟈���4��3&�����
(&�b���J���=��y�	U�Im�q�	Z,l+@��!�䓥?!����B�=j���Ocrkӿ1U虮Z?�I9��r`��'�<E��'�0���m!�/L_|�QQ(�rw65��[P*��E	�?E�:�o@�|��?)��X����@7IU�6x�!R��	=��*4�׮H����ͅ��aJ)�0q��q�G	�-�'�@U���?)�ObhJt���RAfMJ���"z �17�|��'vĜkrB��L	8�́5f:bH��"�i>�K�U�T]H��TL�|rA��Gz���CyE �7��OT�$�|�$B��?����l�xm��F\�0�����?���y&t�Aǅ+~� ��@�k�x�)D`�|5~��̟��P�CBu�(p#�\����5���(#��8
��B��+-C�ԩ0e�2�5��E���S	1�� �B�V�[Z�\2�+���+��������S�O�R��e���p�"c�.!D�9�'HJ	cB(
��.@B�Wx�ti!��D�Of�EzQ�w�x��F�Jf(ع����7-�O��D�O�]
�^����O����O��`�8�F�0cU����=q��8����\	�2#ӵ)P��s��"��l��VX 1� �n��@���_��a�^+>h� �띀C�x���5�Y��r�C�aڝ��f�(�pա3��f�R��ĝS+άjb@�aΦAؐc-�!�$þL�d��sI��[^�#�J�U��	��HO��+���������s+���!G�"tH���+I�%vj�$�OD���O���
��Z�r�d��$�r4x ��	[�u+�΁Il8���� H#���ƦT��Ey��]'��i0lXA�( �I�B$ƍY�![1���Q�L�:I��7-H#���z��N�%�Щ��!/�ԻU���>��T��	!=�L�d����+��<�Mr�U��à�$��a+��^2Ra�ȓ��(�4G&%
�����y�&�x!޴�?�.O�=�J�}���8��.^�Q<�=a�_�{p��ز��ڟ���<r��)��Ο,�'rS<]"7o�HP(|����M�
1��ZS]����d�B"�����]�x��Ex&'�D]��bËq*=���O�F���O(R�`��jE����@�N����w�x�Ѐ@�yoȱ�?u�|BJ�<�ؒG�ȣX��F#��y�o��Or(Q+6-��]���$��'�ў�S
�?9u�ϹX�(�TɆ�<|��a�Az�IB��ٴ�?9���)��v����36|�piA��ekaQ�Ha�����O�|"u �V�ǊP�|���r�|"ʟV������n�|A蕆/�0�6�������`wIV ���8§=��x �
#�z}���D�Cg�p�'A,����R�ɧ�� 4��j�-آ�kD7d����"O�	��ȞN~�<�f�ړH��U�	�h�88CsE74Ε��W���@� �kӬ�O�m2�fX�Re����O��D�O��Ί�[(�!ɃQp$��.��dщ`�^,�<�P�4q��I`�Vw�'F�%pc%��PA�<q�,�5.T%@�1��&��|\Z��/�M�h&D	�E�O��4v��	��f��`F�3{��(��F�y���-�ʦ�.O���@�'Q�D�?�O�} �/P�ll@�0Iټ9��(=D���d'��b�(�(�%�(`�^�[CϨ<Y#�i>���^y��@!Y6���5ʕ<M�l8�/�&y*2�U كZ���'���'9֝��	�|�RDY�5�L�����8q� )I�jZ0H� � +y0*�k�v�~�����wop�##��:�>ةt�G�9=�)�7 �#�@����O~�x�����OU'��3���
�!J�g�
���M�W��x�4	Ez�I^9�1�U�pl�{w	T�.��C�	�s���b���:~��3�"�ΓOH}lZ��̖'�6�;��c���d�O*�id恇4�BX�"m�^�m�H�O>��Ô� �D�O��S��L��ϝ�NL^Ū���v� b��g*JMc���fў �ql�9.��E剈g(�MS�m&T�p����۹!Z*����ץkĘ`W��9D�֨ʔ"��Nk���R@L�B�b��R��O��'�����Z>N���C�o��h�qH$D������?7��CRA#9W�h#�)8�IV����C�Or���\$���R���"�( z��|��G;��uӌ	��S�|��.�J1~�i���/��2'e�k~�@ȯcM ��H�e*:P���Q�Oh���D�l�$4ڠ�W�XX�<��O��!7f��4�|�YbeOP�p��)NR�~�Ro�����©�v��	�(��������)}>�ǍK�Y3�}Kk�4S���Gi:D��1�G&v\-�����S��@�R <��af�>�a���c�q���#5��;�)Z��ɪ���fy�LPI��3ʓ|��`��U
y�a"��A.#�8�<pcLw��$�"/@��FT�3'���8�8��)����d�4VNT��A[�oj@��5|�@�OdP��'1�1O�0�&��U���C�[�<k�"O�l��ͤ�%:4�N�+�[$\�<���Ӧ_�:5K�r���W�<S�6���`�/M�$��5(�5I�/�����O 8��L���O���I���g}�P�S�,=X�$�+*����O���W'�0�уCw0�Y��P���,��)�l��tLE5~����aЎA��#>1�C�7I����`�l�0��O�*RS��"�O�.|!�PРXS��d,<F�F|2���?1����Oײ�
�V�N+ �%O�}eFHR(O6����1�����Q^Y��8�N�>E��}2��<YVA��� ��(P�-z��p���qy���]M�,=X��Y>�;CA�?M�I�ZGF|�n�c�z�{�B݉</6���37���H�ӥN��d�0z5��b��j>��|*�ş>SS
�U��?BX�-p�bF�<��#4fk|D�G� Of�"�bR%jSĢ|��A/K� !1G�O ��l����<��۟��IJ~J~��OVQТ��,%}j<{Sm޹$��t�P"O�(��GS�1��Pj�Lڅð���	9�ȟ��I�i�t��(���
(:q�B�O��O�$�W��6 >���OV���O0�i�Od���B�6����H
,k�&�����{�`�ʲER~L���<>C��!ȟ@���{r����H��SunI�0 ��t9!�`M�C]��q�!��9eB�@̟^\c�{�M5>���XGc��r�l�(�����d9�r�'�ў8ΓHܴ�h��Qoqr���ٶ#�|I��h!�J��^e^���`ǩg*4q�I�HO��OV˓u� ��IKTΐ�� �d֡��A�/v�h�)��?����?���?I����Ԥֲ�h9�H�{������T ���oޥc������
Q|l2&��q�'�8�s%�\�|�b��V�M+~�����'N{�����+R�Y����L3^��E}��˯�?	T��#Q,�8/�����_<B����e�'���@d���QgɌ$3��#�%.D��ئ��}D� �k��p�Z�)���<��ibBS���Պ	���	�O
瓗B��Dp��B�!���Hw�B�jsR�$^U2�d�O��$�u�0	qR�Ν1�D|At�
�S��(/�8����	#rP�rTMz\B#>��Ӫ��0a�G�a��!�`(�3(p	+U+�
�T�r&M�]I�걣�c�'�le;��?���D�ԣ*y`ԎF#y�d��b�%��D1�O�庣_�_آy"�+@aD���'���y٨�7�=Y��,C�0�t�'�dHz��'b�'�ӹ_��I�X1�PZf.h�D�.	��J��M4 �`̜.��ّ"��3�ܤ�cf��SC�''�Z,���Ьzˈ9#b��g��1�R��i�T�\(:�����3�K<�'?��Ų�� 7����u��/N���Γ8"���	��0��'��� B�۵(ܬNFt��I�M�n��"O�Fƚ)+X<;!-í,�����I�ȟ�Hk1G�j�@iy`�6h�u[�/�O,�d�O@�AS�F�b�H���O���O2�	�OF<*T����U쏙$Ӳ��P�K8"� j2�Ԩi�,$81��Xx�h�b�X
p�dNAq�2o����D>0��-Е�� R����S�p v�' Aj�����@� ��S��"l$�!#?��������IK�'+�d�*=���8c�^ך`�F��Zs!�dZ�^yl�*ơ5n�K/5$l��Cɑ��Sǟ �'�\�#�F_^;GF_��FD1�ŕ&����e�'\��'L�O:�~�T�9pT���
&Ef��r���(�4te�ؘ�S�b3'�}��Q�Q�0�ªD$bx�R�
�j�EZB+��+�ي��.9�hX����`���I,I)�Ā�6�����Ej$}�愝9�^��'���Oh0�Ą�-�0p�b����!b�(D��KԬ
i�x���	��Zʸ5R�G�<��iaR\�� `����)�O2�,&5���A	F�v�B)C�τ\���6(�x���O:�$�A
��KʲfΚ�J𩇔*1<	c"�]���A,H7�"�J%���|�z#>�1��VXȹ�<dȄ���蜴<�5q��	!O[td�%K�Bd6�X�#�j�'��<���?)����Þ\�$��`M�H; �yņJ���d3�O����a �*fPT���ހr�,���'Z��KռQk�E��A8fy;s�Zg}�!�'}��'Y�^���O89O� �B���@�Q؇�I]6d)[&�O��<	��i>�)RBA CT�xWNH�^-���H8�ɴZ�O8�����Ɏ3s>x�Ң@�o1�����'���nԟ(h�m�<�t"ß�I�?��4�?�E�+O�(U#$�L���:/�*@����4�?��S9�?y�'�]R��M�;y�V���I0gW8o��pO��hau����'���	29O$�ȟ����?q���<���«/�@��3OT8]\a��g��<h*@�I؟�����՟����.�@4����:>���"<߾�rk�HQ��v	�,���d��&��'�P,��)�~���?����?��eH�<~�`��&�oJ�@���X����&�?i��s����>y�ԓ���4X��t˓���)����Q!B�|���B�v5O�*��'��B�	����O|�D쟸ܛ�ę5`�l��_�r@r �K�<L�ɕ~R �D�Oz-���?�b�'�����M#a�Ճ}���tE�H��"Ys�	�z�F8O�i2�Ex�nھ{y0	�O^�$�O�慢IA�.V�X�I��x�'�z�>!�Ne�PsSA�ͦE
�4�*��y�#R�a�����Qj��*	4՞����:xƛƮ�.j�X7�u}2����6M�?A��Ua�m��ĳ@��2	Ǩ�j��<^�!�D/R~,�[�f�2|�4��@_��6�'�^������z�G�5\x8[�v�z!�ff��'���'h2�'���'(B�'���Qj"��@�	eE�N����2
�ڦ���hy2P����yy�Q��#������ıHM�Qx��A��M����?�H>q���OR���<xq����K{B�<*T���	F�'��8+�Y��抭CB��bAk��$���Iݟ�'�ؔ'���R�Q�Zm��j+8g�}��'z6M�O���?����?�-O|�Ģ��#�A�"�v�Ib��@Þ��F D�`�#�_m�Q�B�w��0Uo?D���&וT�r5���\ׄ%Y��=D��
 =��l��_>}�v:D�袱O�4>�n�ɤ��U��Գg�4D�x� e\�^��@J��Ͳ����`3�?���?	���?�0��r4&�����s�����_�v�'M��'�'���'���'WB���$��x�fؕZR�Ѱ� ����6��O����OL�$�O���OL���O
���!GX�B��T�?������bj*�nZ՟��	֟T�	ϟ��I���������	WEV0ɱ�� ϢD(�*�~�8�ٴ�?���?I���?���?���?��� 9�Q��@�2�aE�A��ecB�i�R�'���''B�'���'n��'��p��M�@����6@��n�@�D�O�$�O*�D�O��$�O��d�O���7��c1F��E��-z���qF@ڦ��	��,�Iӟ ����ӟ0�	��$҃B�>r��<�6���d�,�.�2�M����?���?Q��?y���?���?�C�\�"L2UN��Q�|�����V�'E��'���'�"�'���'12@�� l��
�*tǚ0���$��6��O��d�Ob���OX��O���O*�đ�?d�(r�U�Q�a��-׿k+�m�ޟp����\��ß��ꟴ�	���I[�c0��	n�D ��K�@ǈi��4�?����?I���?���?Q��?!�2���a?�ezp	��'��踑�i��$�O ��3��e�'>����*G�����մ&�(��4O@x��'���O:�ڟ@�	�<�CN2:�"��!Ŕ�K�� �W�����O�Tn�ݟ0��������$\&�n��<I���J�A��^�ƴ��V�M����O��S�˓�y�Ot�4�>�ɬs�(�QD�RU���
�J&8�?1e�i|���O ��3� ��`� �M�*�����F[8M�v�'�����O��m��M3�' 哙>v�y:�,ޠ���;��� G�ʓm�"����T7#�-��$Ğ�RF�n�<�c��E��H��{r$�����N�':ax��W���#��ȕ-Y���ս�?�d�i��m'B�g�:��<ͧ���`�$ܘ�[F�M�"`}ja蜬�?IԽi*6�O��z2Ie���= @�⨝�	�ݬ{<�u��K�."��_����������G{r.�%&R9zb]<��cQ�� x剄�Mk��H~��'(��^>e�I�,�~镋ֲF}����	T�:�d�;�O0n���M��'�>q{RCĝ��|@�&)���%j�*`�Ua�<?�"J �h�|�^w�<��O��D�O����7A I�㇈�7��`��M rN���O���OL���(H�`˓2V��B�>�4�(]�bY�a��:V\ E⋨h-��'�q�Iҟtq!�>�;Ko�S
�MCqȏ*O٤0����;� ���+��w<r�ش�yB�ig^�
��>D��|#���>�3�O|�	����B����(ܚWXNh���_�!�)묩�m�*<�@�r`\�w�a~��F�_q�Pa�j
����c|ݺ(Y�� ѐ�#9���d֢�J@1di��i2C�wTN}��-	u�>@��C Nx.�Qk��I�IХc��g~TBDeWS�~:��C���'�D.R@^%��i&^�i' J"0,��8@[�M�nQ���`�-/I˓��y�C]2�?ͧ�?y��av����Mò�f�eYG���2��5[�B�,bW���I6�HOR��޷)�\��c[�y�T�%-U�e�bq�a�O��m����d_�	a\"<��O��`�N&5����T�Č���"Od]���:.�ʅ�v�V�V	��3��I!rd�ؒP!ٵqVL�c�)B�4��'�*	�E;vm�s7�-�T�$���!�H�u���7�ۅBibr�ʙ�R$��h�G_B��ס:!�D	�p�G�A��1я�6ˮL���Du�����8�����m�#Ÿ�f=#�@�3
Ă�jܛ��ԎpF\�"��80�C�tȹCG�r���tOzy��'y2�|��'x2�H>L���=[�a��E�M�p�7ℼJ��',b�'b�'y��=��6��O��d�6�Dk�	��M60��KM�x�����O�O����O,��1��O����O:��[<ȅЃt� �a@�#{���D�O��$�O��	%�`��~��'dW.�F� C^z�Y�i�2�v��K>Q��?��K�?����?1ʟV��0!b/�y[e�^x�H� �'�2OV�%Kl���'�?Q�'%a剻� H�7k�������?(���$�O��A=|��$�O`�$����5��� ;�:�r��)1��
�J\7Rr:Y
(IAh�8R���?�;G�����kіW<��;:�,\��q`G�U²�'��'SҐ|2�'~�'���5(��BB�_uTP��
U7d�"�|��'�R�'Lҗ|�-��1���R���>(Zl�X��O�H2�i��O��d�O��D.��O�Ո���$�C�
zdW�"H�M�'E�7�}�@�8�Ԉ��.' jt�v����x2�� ��p�U��V�8F\�`�Vl�P�I�p��a逃5T��g��	�D 0��R�	�&h��DY�t������%PD6�z`�U���i"�h�:W�����P�	�p�Y��-��}���/Dlf%:�R�����1�X1C�BT{	���%�#�05�"�FX1
, (č��?I���?�����n�O��dj>e�sfJ3iX�`�E��A���mtr��e��I�Ykn�P�@˛vԔ@�EU�n����7�� �0 �D��S:a{�M[�̦*�iZ�������	X�K��'��Y���q��?���G��:��`���:O�l���'7D�@�o�6��TJ1�J�O`q3� 4}b�y�d���<1�X d͛V�'q��i���e��x����tg������O�)�I�O��d�O����S8O�h]��cT�1���-ݦ^2؃7ā�s���(di˵0�P����'o���ūJ)o>l5�ff�����˕u�:�k&����Z���F�ssp���O�\��8�K<���Y���Ia��#<����+��(7K��`��=���?A���iЈ+>&%�"���^��7��s�qOڢ=ͧU�DF�
+����"��$jB��<�d4�'\�@zs�u�R��O.˧���3��M3@��j����6'�9�h��ɔ+Ca�(�WȽ��z��9R����P�X\ӝO�Og�pcӫ �E��E-m�샯Oh�K�L�gT�i�D�� vH�&B9��O�i�ՇW{w<�k�i� p�&��O�ܻ�'�6��ئ��	k�O��� $a�2����Cʝse\9N����^؞��
O62�v���C�*{3�(	�G;�u^��(��3м��
�PHhb�X�;3�'�r�'.BD�0�"5���'{��'�Z�]��A!�
�{J��&┃H���	ԏ����k��HS��mr�'>c����6�rb	���pDK#L�#����ͻz�V��!�=%�4��O|�V�Ο��	>
W<$3§5/.x�F�>��Sb�iD��E"�"]B�<���Mrg�l���A�Ɩ�'\)���h�<�G,�9R�����ņp���y5�\y���7ғJA�����ԟ7�f@)�b��{ЬY� `�47���PF. 5'����O ��OZD�;�?Q�����W�%7J�G2h��򃕇rبs2�:I1��U 4K�yi�"zW���A��q�:���� vՒ�6��-T���d��"Y��y���M�  3D�V���yfM=h��Qd;�M[��?9���?����?�����'I�ҠIV�S�+��ey�L�z��%��.��`W�'��Ձ��V W��OlX�'��I+Zd��ش�?9��M�J�J�x!6��J���cA�p���F�d/"�'��ʁ�z��P����|�X�Ӻ��ˇ ի���g�0s�lV�'�8A��ѢdԜ���o��pVlD�2PS�E
09p"?�ԇ�џ���43]�'4���wgH�$"pUpb_z��D���'o��S:+0�	����^G�����n�t��D�H?�0m��zFN�JW�ʸ)l��T����	"{u�ș�4�?�����	�-U���{�t�iwn���ҕ�u�^57�x�I�DGǟHs��S�h�2p-����T>Q'>��F��?V\b2Á��8L��$�>��f	-mt)�T��Aa�$�D	"���R1��+N�l��WJ�����1��~��ZI?��~���S&��� ���"-dB� J���O�����$I�xdC�Y�H
 [���0Q��i��dx�င��*9G`賦GA'������?����?��Q-d�������?����?!��"7E�f�t��GN�y� T��Po��TH-Ohe��G�S&l�'>c����ӊOX��c�g��F�r���V�](��j��D���N|�>1��վRs�s���H�����4s�L�F�n4�ɄӉ�?����?ڴB8(�ƈG%t�H�1�)�@Ӗy��<dp�aȵsF@3�NN��&������ؖO��.�~=j4O�i�RtY�&�DZld��7�O�YT=���Vl� #F�5ҪM�?�
�
��ŀŨ�嚽zql s^���c7D�r�O�
p�~�2�nN�i7%4D��˃�}oN���*�|^6T`�5D�ЋTk�y��tc���A��[�4D����g�6t��
�j�$k���5D�H��	@TH�`;Zb@맀0D�� E�.ADi�@T�u�<u�ê/D��h��Q6*�hW=X�髶,D��;�k���*7M^����.D�@R�H�&hvLG>��\Qs#/D�LarMFh#���H�a~Ⱥԯ D�P��`[&n@d$JGӒ7~(`æ:D�� ��)����.ʈS�R�6D�xQf�^@	AtM�{�X�B��!D��*�w�$$	amQ��hZ7�(D�� �GA唘�*�6-���� C$D���E��s���R-� [��m�D6D�9���;,��A 冂P��Ҫ5D��f�7I�Ұ�aH"V�8���5D��r�IS�f2� �u��̎,�@/D�DHe�E��ꀬ�!���*�#7D�����o��I)%�!6*d"�j2D�ܘ�Ͱ8l.�X�Γ�.�AF0D����Ög���P��.!PbD£*,D�HA�ჇK�U�fꌽ>�Hp�!a*D��"��?L�X����Lx�Qb/D�P(�b�Y��t�Qi'� �A$'D�ܘq	��<��`,�9g����SB)D�`��n��H8+t푇<怔���+D�BWD2Sl��˷k�BA�q�I$D��!���:�4Z��1)f�Ү8D����)	�okĄ*(4B�X�9D�p�ÒV tm[��ԋ@�ֽA *D���v��"Zf�䦖3h�d9�+D���f	��Dy���%��Xԩ��K:D�8w�E�YzI��יGԤ]���,D��3�GH�AUe��)?���6b*D�Tc��Xf��á�N����,D�XY4��d�P�A�&d�~}�	,�Ir؞X�-I���ݨ�._�l��S�	 ��o�+>�smO1]����$1B��-QS4�Vn�I��tAL����$:�S�? �ׅ�Z��gо\��"O�� ˝<�~��ƀ>OO�L��>Aa�)�ө6
 �$�#H�@�/w4PC�ɂ7wjH����7^���cP6'�8�x�	ד&��]�WE�&<�0@2��A�B���ʬ��Sjψ#
<���_S�B��'D��(� ��4�C���,����#,O�mDxb�K?���+�59�L�����y�`
�Z�*4�B�,1�ZmyV�\��Yc��b?=C1��n?Zd��L�r�1�@�*D��Ӎ�RgH<���O8R��a��o7��>�0=IQ�D�*��w�۾�(���DQH<1e�K�6L�9A��]&$�XD�?f�!��YI�q�0f�8��I��M��$0ay2!,_��#�b���*���]?|��ȓR���a �>�j�%ɷ*zv�$�pX����ɕGb��[���Oʤ���ĂN�!��]u�l� ���c�伊FkJ��O�ن�ɇє��#�̲\��	ʁ��"HC�4$Y�@�K��H�F�X�AK�oX�E+�'����<4�(k*Q�j��8�	˓yj�\�ڣXM���R/Ƙ'�ip��'D��	VIF�U^%�����"����f"��Se���Oh�d2!�2
�p|r+\�<�h�'��(�ϼu��hM�V��,��}��5LOV���Hά,�u�C��4D����UO�("��p��(�U���S��L�Q@R�<A�A�.*Ĥ8X#I*oȼ����pX�LEy+8g�ڍ ��8JG�8��W�y���6��"��9<�����)����hO��L���+S>�$iP��	�
S�lS0"O��b�b߱}R�q�A�',_�cX�\Q��� �a{����J �'�'�d�1N��'d4� �	rCt����R~:8�@��LXk�A�	*�Ԩ���S{4$�@�[���� ō%a��*s@��#<i�a�7����(YO^�V^H �nX�/��``�'�$��R��Y��:���C�o���YC DH�I�8"<E��gυt�$I�#�L1�t�ӣP�O��	i(��3�ᓬ9~B�k0�֠"����NQC䉴Z�,�x�@�[m2�Ⴖt��c�`
 �4w��xB)�:Of��?<gr���xb��9�.�3%'�,l��#sG
?�:�R%M�{(<v/�_�zIg�	�l9)�I�~8���QDI�*�(�Ȓ�p�9�DͅG�0��"%<�qo۪/�4DҕJ�6���ȓl�b����\�!�q��DL�nΑ���|��.g�p�!!�>m@��ȓ2�)�B�_%h�:��?3�6���zFD��@
U�2�����O����f�����,۩���c0j[�b���[���ȑn�i��=�V�A��ń�&FΝGJ�3]7: ǵ���5�ȓ?�nM���B �u��ˡ(3RP�ȓj㔕S7�B���ڒ�ҝO����%�z�I%Đ�]��UZ����D���ȓw��ƅ�J���C�g��͆ȓC]��z1 �""�=�B�1��� �GbA�\�8�g��3wE
���g첍���,�,T���Lu����艙4F�0���0΅] D���`/ܠ%�J!L�fV�ņ�\���Q-߉J4�(�Q�/�䡆ȓ2A�8�Ff[#E�P��T�����q(\ᣪ׽^	:CӾ,�\��S�? (�*�ܦfȹ��Hq���P"O��`ՈE,I�v�{'��c��T��"O %âe����ap�˨;�L�k�"O�Q�f��c*,���	�'��c�"O8 ���+��0���XP���"O5FJӦI��(毞�QA�久"OB�2�I�cCHɑg��3g�e� "O�m�����<�4��G�E����0"O�h;AΣ,��̓�E3 �2ź�"ON��Lܫ	�Ia&eיJ���"O�ua⣎�_t�!a$�2K�P���O��r��N��0>���A
}�`��S�*�����m��d�7�h��ش$���0+E��!��A ]t܆�hz��rW��	��Q�rΉ�V�@��?!�)\��8��	UF����S�i2L�2cH�}�r IÙ�C!�
'`�)̝	sp1���cU�TDxB�*�g}�)BK��I���&>�Z�G���y�Iɪ
�p���e@!\<�xW�H������>��aE�[�zD��HOҵ�
�/FZԲ�
]ò%R�'�j-��3O֍Y�N+O��Yp!�L�-81�L��Tμ��KS��1�O�}2�nӱ;Ap9�5+$��uy���&��Q��'�>	�C��2\��YHZw_�i�'uT�1G�߅#�8����C�m�܄ȓ���R��čA��:���f���ѹi����ahV �Ak���=5.�õ������y�j��P�Lx�@��C��pm�2�y�b�>�tQbi[)L �"��V�/��3`A�$����tB-`z�Ð�?��%��'چ}Yv�^�KA" �3�r�0�� ��Y�AC�K�����J�oȰ}�W�E|�D%�fOH�i��&,ڵx T\��˔k�a{��Ƌq��%�ckѵq�U1%����'�EU���z�f�Xɚ�:� uS���Rӂx�����q2��� +��a���,����'P0�Ul��p��q)��C�C�Y�|�H�J\�a� 
0wZ$�e,�J�ӕb��.9&*H��Gu
���U�K��!����$������B�ρ
f�y�a��It
�I@/��R�����\Ū�ǀ��'<l����jۖ�h��@�|f���
��(����<]l��Z82D�Rd�^,v%�e�3͂
09�qكC�G���J��p=��f-\���)\���Xۆ�Tb�6վu:��֛Z�b9j�`��u*�ZSM��P�`��E��|�`ۥ*F�} ��V�#�!��+�r)�2! �b�� 9�(Mxʶ��Ao�+�{�ʎG��@���[*�z%�J~��<�R�^40��ո%�O/#�F�sQ"O0�˰�ذ�����~nP�ϓ:j�����lf���gT"��n�a��A��'��w*��3\���î�5o ���ytСl�A3�5�Ү�j9�h��'����;�#�N��q����7.x�q��)�><�z⁐�I"�C��&ƾm������'ل���B� }�T�L -��립� �P���IP��/�VcuH �B�,;�g��y�
%>�����(��r�X;��ɨ����p��  �.����J$<��&?��w�H�z��T����H��"P��'/�|�
� �����'mDI;�4o{F�:�� �2��$��i����~�L>��W��X�M�U������t؞����5?�EcW`N�"�)��x04��'��tA	��O�ѣ��~���B���<�dѐ-?~�nUG&%���Z��#<�S90*V)z�l��-@O��~����	^��!��I���W�(2�\�6�"c�έDy��K����?�+I�r��d§'^H����cjC䉩y����0��]�*�i�7[�dZ>�e���>ʧKr�U"B��%�ZŻR���j����SƪD#�X$:�$���g��!��y���*ljFIٔ�WOz��0�̞�>����	�Z'��&QoXB�� ��bQ �<!6EүX#��c��l^H��@�Y�cS"�SRe*�t@�Z�R`/���C�	77Zn�K%�8�2ɠ�E�>|L�7mK�}���AG���X���:ol��}�1[* 1[g�!9���¥|�2�ȓ*^�q�ܟ`t�1�C�Ϧ&;�p���U����f'�#= �|J�v��O<!�'��t	Ԧ�;{AȠ���!p\=�� �e5Ƌ�SG�t3����X���ѵ�H8:dx#E�7r^���~y�̙�㎖XȞ0��6��=G~2E��u��R��� 0��Fv^����$FE��y4J�7@����S�? �TVӳs�@����Y(-(��r�"On��w�L�4a�C�==*�O���*F� �T[���bdZ�M�?�` ��dUq�alqY��D��k�d���8}�ȓl���1��F"
�*D[�Âz���?5��#.ɢ\I�ј�fQ9*��ȓ�f������(�P�k45�a�ȓn��M�sj���Y�R��1b�2���(�H��H&.�b��ǄU,��_"Z��UŇ��ba'�X�r���c^�y�� @�z�9f�T�T��p��;�1�cy#�xFю!�i�ȓJ���Z�8:���	�
~@��ȓ2�^���ӕ		V`pF슁AV�ȓA��� X=+�y`$�Ěk�v���I��U(��)�
ዒiSiAL�ȓل�x%�U9�"t�h�mǖ���Z�L��?+J%y��3መ�ȓ<�x�dN� �������8��ȓ�8�E!t,Y!�@�i2r ���,Y ��F�0�2�R��X	Ez��ȓd$
�����+{���`�8)�|t��-L��I��N6U6�j4/Ki���_���D�n�.�CGe�l���p1�* ��@Cu 4^� ф�*2�ks���/y�+�M��6Y��ƽ�%%�-_^0k�Q?�}��#D��h��<E�=��ʟ��� ��=D�L!T�M4��F�ґ�����j=D��a�l��-t*Yh�bO�.�(��I;D���voJ)��0�3+�@��:D�܈�Qx0"�S�ʦmf���&l.D�8�"���d%�4l�( t���-D�\2w�s7LL*���	S���,D�l�p q���`#���P���a),D�� �y ���c��P�7�*D�xzr�5.|)�,S&	lzp���=D���g.�5�� W�U�D����?D�<�7'T4�� �TK��F.p:�+T�� ��߹wtN�ԅQQ���A"O��xW���\Q[�%Q`ݸ��7"OD�[�.��\���F�΃6ؾ�r6"OD�Y�IP�U���`���*Ġ%@"O���l_0'$2� ̲��X��"O��bu�O�F��v�ڄt{Je�J>D����D��=�hd� e��1�8D�\�s��t���	c0⸫��4D��J��Y'M�(%cI���3QJ3D�X��,R��@�M-��i2�4D��wB��'����ꛐmo>|��K3D� y$��a&��׍T�cF���l$D�<{�o_	�al׿�D� u�=D��a�嗶�$��gb�d�~���:D� a�	�� P�Z6�H�>�l�A��=D�X@�&��i�(p�P/C����" D��pg��p`a �޷5ą�j>D�hxU�a'�Kԍ_�n|�	[%;D��B@(��dife��^'q�.���#D��,,�B���#<3���m)hP2B�	�B.Z$�a�.�.�(T�L�B��/XP�\��m�@��JW�C䉪.��:7�^���t��/H�����3� ��1�\ G��?O�y5�K
;t���²}�\qh�����R�K�:�.-���v���?��F��s��US�
����R�J�B�)� :�ё�Ș���#l��/�*)�p�C;]�����	�M:�-������3c�(��9ӅJ�*��p�.�uX���FM�+�L�X��ş~�Qb�&��k&M�����'Ap�C�eU�}���H]"!W.M�J�����54j�4�u�t<�a4ғM#BiyÀ
:u� ��L�(��y�'��A�T�41 ��?��I�� �
P�H���H#"�`,���d8���cЏA��D��8Sw2e�U�cӬ �5���H2�a c�^�L<�}��	�&�@P�va�h<-
��O�F�@i6�ɥyˠ\� D�~�<r�w�������Č)�7'��r�p�[g�/�P��μP��l�%fq�=�e(�7,Ije���ΥEG��z2��!Z�r]��t��)�ӱ65��s����l��y 
�G �p�z��hy�B�7m��AY�.4P���U����,%\5�	F�
W�#���$s���I!;�pT���?��f��R.
؃��J�k�Ibm�Y}2�F$5��{Q��tМe���nchEP'�P�W�(B�I�1;� �=�b$ښ�~I���8���=���@�VT�7��^'R=���8s���ł@������A�xLX)�.I09e0��Ƙ{�qOA��c��P2��)-�'�e0�B��]�Ɲ�D�Pق�'���R݅`�ɼ"MW��4�bHb�\%+f!��K�ɪ��O$ӧ�OI�XJde�0):�H��h%x�m��aW�1R`���0�I*Ғ�Pa�:
p$A�&eӎV�:�'=�uDCb��ispoL�6(���J���P#�`�֟�����Gw�k���>9cX�SI�x#��*8��EC�s���:���7��i3����I�4�?�ꁒbL���QoŎ[ھPЦ�َ_d�V�y�`�Y�놖�MS�d�r��#?ɢ�twȌ���R]�<�i��O�l��1F~B�Otҧ5�������ӎ<����`�@C�ҬGR�x��Q�@\.�yw 3Ik$�9�,+��ye����~b�>q/�潰uN���H03A�M��m��l�,_�:]��Eh��KS<�
an��W@Hِ��>tt�O|�
ͅ���Ś�c����]�������|���^�abL�5�Ҁ5Rf�Q��`��%�'LCF�s+G�f�&k�Ry�0l�|7R�s�d6��*���C���i��'R�#�Z��1�i�t5�0Qp�@q�H˂d0��O֌)��fQz�� /C%/���aiݸb!��0��'��"!��;ІNr��h���M@�����H�C�`��	#&�4 c��Ƽ��Hc��������b���b~�Iu?�f����O�B6�~�Т���Y��q��T���
S^Y����)G�m3��1�.׉L�l�O�1��y
Y�c�S�r
l͂-�:C�x������	��~OT�����У�"3��%p"(��qƜ����NGR�X #��8Y��H�����	�5s ��Jl���͹.Ξ٩�"�H��e��4q_��;���{�Z;�	�l���G~R��J	�$���8)� ��G$5(�D����6���G3&n�ѧϛwr��6jC��0��I�~����S��ȼs@ ��X�&�ϻW�b�k��k�I����)��v�z�pD(*�v9����?
�y�ш��\�Vp�?1�c�*N���pP��U�y�dRcR�a�OG&s��qb6��3��'f�6��O�q���׸T��ѕ�iv80�Æ�>)T�F�)����p�X4mA� P�·�l՛��JǈD��"u{ �?��q����FkB"� �b5@B�o3rPhL�D�,����Ph�,D~g�d��H��E!ik�)ϗg�&�F�+������M�|ߞ杕iu����Rc���4�g�&X�Ro��p<Ytn� ���w�:Y���9čCA��i8XR�MRp�*��C'c�TEP�W�`��0�H�(D������صr~ڨ��,�&A�L�e���o��d� '@d�S���Q��Dz"ЗJق�C�D�3`2�Kǃ�����z+�d���ԚZ��!��`GK�hɢ�*\�*�L��� �Y�v��ǓuF�P84b�!�����xcXuoZ9JF9@�M�A���Bg�.k�#?�!HU�nB:�3�A(V*���֎T�[TBት0C�
��A#	��#B�_�P6@X	7����<aC�\�z!l�λHH�!�N�$ K�\�J	��%��Ih�$� ��2��&�*(���F��%��)%O�\���883:��5jK?8ԥ��ޕn�7�C,��>��ٟt3XB%�(��� ��qx�F-�2h�H���6�t��?!H$1�Eٵ"'ZC�	1~|@�[VF<D ��Y�V�O<E"��3V��I���M���b �PW���y�!�S��Añhe�^P� @N�K�8���T�D��L��?�'��T��.\sF8�`I�4Dա
�'4�b�A��d�`��fvE�A�N v���ň^FX��( GQ94�HM�R! ��X!gd <OHL�V)4@{�Y#�O&�c�(�j9���k�/3l�T"O�����k�b]��ʇ�>%����ė�~������J�O,�:V�@�����R���� ��n�P�0�zኍw�t�����a�ЧO��V�1�3}���6��x(���2�DP����<��x��C���{ H��`��t�M_>��ō�G�q��I+ް���V�I$�c���M��d�f�+(Jh��@j�v{x�ِa;O	��ț�)|TZ�Θ�&����i
�����W�Em�k6��;?�?!6�
=X)ޙ�7�]���v� "C�C�	2��d�e3H,��J�D�6Մ#��]�p<�'#�2��U�w(�})��[5o�R�Vf��y$L���I��o%�hꃣ�RPD��Bэ^z�����_\\X���W1V%��"�'��[=�^���[Š�-S�l���3.�Fz����`T��i�6`�G��9��6zs�!���G�|���14F�+q�0a�3�k/~E�#��<���Ǔ;/����P�pei�K�5�l�2�}� �lm~���ӀZ�^#?Q��6q�|��EZ`fġ1���Q�(C�/8L"T1�
C�)&���ߔ=-����,R5�p<���?���ڟw����L�c�!�� J��� �j�,f͵_�v�j���&�P����T�<� J���>i��8�b�����j�A����5��#6ϗ)B�z��1�F@3b �'>L��Z� ̈d]fF���	�^2vM��l}��Y�
� d0�����F�'�M�X��Ԫ�P&�J��$`D�;�ڥGZc�~@�WIɲY���dڈ= �XF��=�-����O�����%�~#?��۔P;�iB��ҡl��i�+�-~��$/���H6h�d� ��Ń# �a$��B���� 56PցH\8���sA���λRsf��&=�tpn�Iu�-$��nZ�1��`�2�̔Z��7�� b1h`�[�ڈi�艵
m�<�R��ADb��2,�;k6��졟#��6K ��B��1e �YvI[�	rBm��5���� kqh)�ĕ�o�-�&�
�tԒ� �"g�X�0�o��>m�ܠ�GWy��-p(3��׎�O�Ց��,؀3�֝(N�t��D.M�F�	���2Q��6탮uȤ+��R�{A��X"C1���!��|�b8����x�`Tʄ:bᛆ�\Q�<�c%�wL��S��+%��ӊ{�x�:ɐ/e�u�)��d�>��C��M8�2�IP�|����;eC���Wm޼�򢑨U�N�Q0(�<y��f��487Bɰ��&b2�w2���G�u}��� �9Q6!r��$���ß k���E��,I`p|Ũ�O�*���*ιji���@�*<���0�8�$S�x�x��Gi��|@Z�;��QM���t}�1�Є�{W�bF�^�1�MBӏ	#J�	�sMM&d���9O0�ֈ� �Ta@�F~}�d�+ K�x!w@D�o��%�3�M�`d�h�1od����E�D�����ܼ��O~}y�)�5E�xj�/�ҪECu�Ƿ�y2䀷�R�(#�R$t���S�O�d�s�	%~���B���63�9��F��qǜ��]�~[���`�q�E�Ő��ܳ�h�W��0qD�	�y���'�����9���M;���2��͠��lFq�p	4�x�;�DS$��O�i(��@�yX���h���xs�O����,�amhMʲ�՝pO�!�T�k���Ԃ޴L����j��X9��΀Vt���^�gm�I�>A���a_�u��l	0SMt�rA7$�ڰ�N�YI�1�L�7���	��jt��` 3��q�5�	W'Z���j�(p�!�Q-\�ipu�!(�<0)�d^U¤��	'�L���W���5p�6����c���Z� \�l��Q�'��ѥ� P���@�����2��Y�IZ34�e�Kh?�xl�)���:�9���ɩa�:7N�<���PM�=��D�('pd��cJe�s����#״
�l�����GY�9"D���D�X�����'�T�#�G]Q��q@����Q��4^�p��#�I3N���W< J��YFI��6��4�f�P�A�'S�5�b�@��x��L�%�yh�O�YYbh��DO$�"�(-|Ǟ����e�iI�LR���s䉿�?Ydd��$���!�$]~Zw�(p��	Rr�s�&�H 3�4n9�0FB�7N��A��) ��PF~2J�$s6�{��� 4T��΋z#�L�d����@�\�S�O��H��&"g�P�Vi�|^H�͡t�X���J�	D�{%(}�� ��/G{<a��.�v�v:�If{
`���d_!7� �$�Ԝb��%���;%)0��7gۋP���ly���yER8Ir-[+6�RaQg>}2GU9T�0S�j�4:/`Q�2.��HO�י�V�yc�Ŏ)�^���mLp}2
�3������h��i�ś`#@=Ѵ�P�K���rGȱv�X��㉝{o�:��+�x���K� `p7��9G���dM�^_|( {w�����)��Z��3���$%fmi�W~����;+�%S�c� G��P+�(\8�1��ORX�8�R.Ah8�ݎor��'!�}�^�	�I_H���$X=�,!��닠\$"e��ϛ@ A���J68��Ȣ�'̎�g �0Eˣǅ+5p�X��'�"]8BT�:W��C�/�8}��'�$�ж��;���ӣ�� *�L���'J��ᰣ��L���A�H�1�@��'W��4��	 D��@PK�˴���'Ȋ5c!K�I�����CO��б��� @|�!ꅡ0c.<3�$�c��	"�"O���pϊV��1����n,z�"O~�ăǹS?ވ�ゎ�a�0<�U"O.�sh
?a �KA�A�\e��"O�U��-���ഠ ;!v�`��"O8 �s��F� �d�%RmԵq"O�zGD�$F���Q�N>��`a"O��9��N��N��!\=*%,��4"O�Y��͋`�� F�{
�9��"O���s�G)ba�˰���r��BA"O�𰰮�u�b��S��(^�ʹ��"O� 	 1�褑��Y�Yij"O����̍6���p��L	zAZ��b"Oh�qS(G�t�H8"&ߗY"�ăU"O������*R9���:Kmb�y�"Oz�ZM�/~#&Q���ÑWg>�"Oh�)T��r.I낅\9
�x98�"O2�b�o��N�D ����X�(�"O2e�'�j�)�b�q>��"Oމ����&�:������ p�ѩs"OB��H� ��;��W�zd�+�"O~�YG�ЇV�@q`AF��x��"O���B�� ��C3%W��J�"Ol	�#�Q6t�$��C���Z�
�bA"Oޭ�ɞ�B�ZQ���</�}+"O�XEC�b��� ܸ(��� �"O\0Y�m	�iD@�с�_����"O��p�	m��0� �'L�c�"Ox����TF{��e�ơv9��)�"O�0�@�E�[������ױy�x���"Oj�{2� ���$�Y<�\Q��"O2�CAF�p���q�V�|���Zp"O^ *��Ĕ|c���d#����dJ4"O,�B�Ĝ]�z`8aC�'zF�
"OpA2v)ʳd���gA�!=h�
�"O@��.�Lc*0���p-�Ȣ�"O�P[u�ӹ'�d��R%��E ��"O9)$������U�t��� "O�ı�B3�Jt0�#]�N��R"O��1�Ɏ1~t��
�<jr��"OLԒr.Qy�<�#U� �2��"O$�*7�	�nF�)�����G�<YU"O*���Hj��X�Iە.�ިb1"O��JEG���i0P*�TN�A�"OV��W��n�P�kM	X��P�"O^��OX��.�'D�3[5�<)�"OB���'M M�̹ �M6  ��"O����큎"�TPS�\7b���"O�a��� -S!2� O(B��L�f"Ol �W^�-��쑧�� �@"O�� $&�X\XvAK�Au"O�������H�v�q֢�<a:���C"O4U!��섘�� ��S�ȩ�"O��k3��,t0���� x�P 9�"O�-+֪A��5���n�lkt"O*=3��ɮF*((���;�8պ"O��3 �o�ɘ��T�f�D���"O���fӆ:lybåB�t��L"w"O�]��!Md���b�cAX8��"O�Q�dQ�}l�cV�J8���S"O>�XQ*׾%��tq�ӹ1"�4��"Oz�ȕFI1 �d4㵃ã�RUat"O�{c Z-x(��I��^	$�`�3A"O0��S���AH3J�>l���ab"O� .���JU�\��L�a��~���)�"O�S�+B�fH��U��N\��"O)(&�n�Zh�2��
��"OX�('�K)D~��$��%[hAc"OZ0���#��1��\x���0�"O��i' �<�޵+R�gДM�"OP�B��K
6�B��R+=K�r���"ON��5�-C���:��4[��d �"O>l��%;�4��I%	�b�8v"O�ᰀ�g����e)[:{`Lp[Q"Ob-!g%ޝ	��}��!��a"O��V��#T�`�f�)z�9c"OH�� H�ujY!W��#.D�T��"O��2� �3A���`�M�!5V@�u"O�(��G�*^u��#�P3T���"O$9Z�OE�^r���&�5o=2E�"O�p��>
����(_<@�9�"O�� �ʏ-��1�D� -�d�kv"O�H�B�P/y����uV�|����"O ��_�T�\A�Ē
n��}��"O�E �	��ayB$�;Q��T��"OL���_��Œ�2��@5"O���kݰH2<�"���)�(E��"O��%+\ ��#�5�d8�4"Of�*�m� c��l�q��/px�b�"OfA ��1#�-��C�%�m��"O�����Ôa���Ø�4���Q"Oa���M�����;]/��"O��g��S��؉ �P: �z�@�"O�u8qc��@C�D�dhHy&L-��"O���q�Z��)(֍���ԙ�"O:��J� 9�-�I��2"OF|K������"�?<�8��"O�I�4�Y�����o�9{�"i�D"Oݙ�F(p�6�R�.��J�B�a�"O�ي����2p�^�9�^���"O�0���8l*p�bL(��A`"O��	1o/n��Zv*�P�����"O���e䙈.���i��S8���"O�h@�yڱ;&� 	�͢�"OD��@�W&e����2N�� 0"O�xN�
S��{��O�nɫS"O�0�o���(ܚ�j�F����"O��(�ǁ�$�z�'}x2!q�"O�A����6� ��ATTX��f"Ot�b�J�l�v�)U���.?�	��"O68+b ��&) ܂�쁻]B�!� "O�P�$''u.0���ڿh6�4�"OdM��E�
)=����$?^�w"O�q����P+��b��m
ސ!�"O�` ��G�8���:t^�}�6<CR"O��e ��� v�Wr���Bs"O��	�tV�]��AX@�*�xe"O0!��k^�zx� ҂g�l̈́�"OjL��&�4t�@��Rƃ�p��-p�"OlQ+ˍ�z.}�Хј(����"O��r�ƾ3r�f�2Q�0ѐ"O��ၑ#9K��0��69�^��"O��
�B�+!��}�,ns�P(B"O>8+����ed2�A`�[ ~T�-:�"O`P�1�ʤs����*~e>	15"O4q(��
�|�hL�o�"^ڑA�"O��r� EA2����>P�(�"O4��bm�;m|�̨Dh
�j���"O� >��&X*-����]�,�4�k�"O�Qc��	;*¶��1Ƙ�W��P�g"O~}�V(Ѿ]���zu+۲\��|�v"O4PQm�NlhQ��+!��x�"OR���+�60r�h��|��d"OF��Ol��TȽF��i{ǈ"�yb�W;SD�G&VG!B�Ő�y2eߗ?���0�>\d�r��8�y"�C�m؁��X�d@B@,�*�y����_�5(� �=U��Т�G��y
��|h�m��(�hpj�ybf�97P0u�a�_�#O��y��s�N�c�ǎ:�v	;�o�yb㌞Y� ���](LO�U@񂒏�y��C0FFB���ܻF]b�%���y��-9�$�� >�jL⧉R��y�DkUt��-�(2. S�yb�[#��P��%��ıv���y��ۆx�\M��D�? � ��l���yB��yP��kE�ޠK(�eb%���y�؟R~�t+7矪q@�h�Q�W/�yrL�8lFh�ɑ*�#�D��(=�y���w�+q	ΎC<1����y�ĆuO\(���G�M��U�7��y�o��5�ڱR�&ɀBa��� ��y"�4W���2S*�
O�d�(����y"��3�F�@���A�$9����(�y�OԈj����?�8E`wʆ�y"��P+��y�R�����gE
�y�lJ���9�m�*n��:�PȄȓ4e�)q�ͻ����#�}�@=�ȓ\j�)F�Wa�Pp���>d)FɆ�~Ւ`J�Y��83�W%!de��#�~�Zd�� >��̘v�Lu����ȓ6�d��&-<x0bCV�CC>y�ȓv� �RBG j&��s5��gѼ0�ȓX�`���D�k$�Esǧ�4-6��ȓ�y��*T�mFHɲC�=/x,�ȓc�~(�0��9U�%plޝ�b�ȓ���p�ɝ]$h�E�MW
�?�
ӓ:�bY���m��e��dA���U6�,3Iӫ{��Q(�ߌ:���ȓna*� `hA ?^�H ����]�!���8n�Nu�4n��{L�2�-Q1!!��7�
��q�H�@ιf�',
!�Cv7ص↦S�i��r�!򄛙-�����G�OP�dD�=o�!���3'�>��v��C�C��6NQ�' �l���·]� �;�G�'�hy�'��Ak��<�꽙����-&X��'�X��eY`��Dpϗ��v���'�������2���Ò��P���'	z���DJT�0��v��0y��
�'�0ф�C�6�T�)�̃=(k�q�
�'{عZs#C+U�	#�N�0���
�'��- ��E�A���66w4(�	�'����DM�Zɐx��KH *��-@�'�ĕ�5��{|Uh#��)4���'2X%*u�\'Д�����r�n ;
�'��pP�>@�*U��Y�h'�%�	�'ɞ�hg�Ӗ1�h���bŜ�Z��	�'�樉E��vZJ�` ,B���$��'�I�Ò�y��`2��ה�\ ��'g(\����7]��Gb��m�E���� .p��K����ÌW+�)0"O�� �2&f��lR;@uF��"O�s#�d#�9sA`P�A`�=��"OX��
����\��1!��,��"O�LiШC�
 FCC���@�"O�"W炇-��$���+	��x`"O\YK��]E���1�I�Q��)�A"O�������>���@�#�=%�r��f"Ox�B�
�{��dv��M8��x�"O�:E+J4�F���/ʧ=0vQ(�"OL!��+H�u,\X��DC��\��"O�A���9_ծ���@Z�J�ܵ��"O`�P�̈́bx@!� O��M赂t"OlIxEA�eL� ���np�"O !hD쟾U0:�oL&u�1YS"O$-9�g L�(А�KX	mx��"OL[V�+��ʅJ\W� ��"O��a�B8]
��UJƪT=TD��"O��
�*��s$�`c�(<s/"�24"O:(�Ѣ�[� �eL)�ډ��"OD��F�O#v9jmb�#�99���� "OPD���]�$�Ca#�#+p�X�"O����'#*|�C߻;�`"O�i��?c� tA�♓$��`�"O�wj*�2����7�@��"O���X�)��A8w��J�X��d"Or�R��P:�z��C�`X���"O�"P$A��� k��k:���"O4ؒ�^� 7	���D<0�@5"O� �M0TGz�@Hڡn**��%"O�MEEԭ[�2�	ud�!Z�v"O��q5F�=w8�@B�Z�shX�""O:�r�!/\5�q��G�v2"O�����/E�U)�(K5r��-�
�'��i[b�L�r�b��� �9	$���
�'��9q#T�qϺi{C$J�|f�0�'
r�XS���B P�`���uN���'��\ �E�?����A�l T��
�'f2ejg��:sj����Omy
�'���n��+���%֋G�x�
�'�p�3�[�~M��˂�?nL���'�=)�"�D&h��01Q

�'pX�BS@�:m�XR��?2���	�'�6ɨ H�p���7���Y�H|3�'EN�S��y��T��4&,H
�'����V�[���A�\� �	�'#������ �j��'c�#`<$p
�'aH�z�N�*Y/���d�
 ���	�'�ؐY�kY�,�
챁��I��=	�'����V��,ۭ=D�$*�'�z�#�/o����,T�m�`2
�'鼕+�E6n��1P�!�Vd��y	�'�0���#ݣs��a�bC>d���'7�=1��U�=4�1 *�`�ء�'�ЌX䨈�X�ZP�˕Zrl��
�'rH���;k
 x)�gS JT6qB
�'���k�i2OXi+�JG��܍�'��j$"�<�l�����.����'$x�)�"�Xe�� o�*��9��'DN@�G��?��\zPe�?.��,I	�'8��2 H�u��1b@e�!
�Ĉ	�'\�E�!�z��iɇ�5Z�Q�	�'�H�Q�ꈑX��0�n�-�����'�v�� NM�BB)�V��.�U���� ,Qْ�nli�GMX"w;�@`"OD�ra��y�$qs��N	W(�B�"O�xѥ�&&H�p@�C�2(�7"O�p����)ɲѨ�����p	�"OB�J�]�ed�����O(\𞩉�"O���㘯xc0��/!��БT"O��2� �6mn)���֥v{|�c�"O���a��L��8!Øl���G"O,���J]!I�
E"��W�H�Bg"O����1b�`��1�$=�qX "O� ����p������=X�du�B�'��M����G+@X`��±K�!��1b̚L7(�JŎ`a׋�J-!��e�y�d`��R5�i�j6!�d�,H��rf�5���e�U_!�D\�.�*���� ��d	#h��^T!����	�4+7j�������x!�$��@�
V逷Q��T0u��.e!�dݐ"<J	���X��ճ�E�CC!��'~�pLBuO�|
H�W�T(!�\+$�.ء��ۯ;s:�!g-�#!�D �r�г�J�\T�Ip+�Q�!��i��5��["W0N�����!�d 3#��*���v�`A'K�!�� ��^M�D/�Fc��>�!�I�3��93k�
6��򠉚t�!�D�kHL�*�H.<��B!ܰ�!��Q�@���o"0e	�!�"�!�d�NJ�C� 	q ��V��!�DW<b�r M �DQq�M�!��
GE(R2C��S�&@��(�!�J�]cP��nF I��m��!�D;E�`��k�+?��x� g�8a�!򤑾J喐R�K�b��@���/Q�!�Bf,�����p*�W!�ޑI�h�C*Pa����Ӛly!�?rQ*�*�
w]�8@Q�K<V�!��-��9��F�hR���f��	�!�D_3 �xH�7N�e����1k� ��4D{ʟN æ�M�R����B�r7�E!�"O��ІHC�WhECes$V�`�"O]H%��s=t9
�P@�"O< 0%�,&�f%�;_��!��"O�%�X=�Es��W��f�Б"O�Ty�����4��F�.��BU"O��s�Ȝg.�a���c��U{�"O��i5Ę��t
��X�ҰA�"O����Nn=:0k�Cw�۠"Oȍ���G�u�DX�g�Ͱ h���"O�C� �V����t�W��B�"O�0fm�$������J3�|)Bb"O�`���tz���jT�|�V���"O|q2E�IR�BFI�?XN4q�b"Ot�9�cͬ@wF�{���M]*��"O���a�;D�^x@@D��4x.�#�"O��q�b�7#%NUm���δ042D��@�Ɓ.�6�v��:��*Sk.D�+6Α>S�$<�X�u��mCV�>D�����Lx�e[R��^�DM@2 1D�H�D�6rF$)���Pt�;�e/D�D�`e�>]ޕ:CjAy�,-�q�+D�p��k�����B�(�١7�(D��H�bݦ4��0c"�[-3���$(D� #G
SS9�`{gB��x�#3!%D�� \�Jͽ5n�H� ��:u?
՚q"O��u�0:V�9sKʮL�9��"OP%�͔\b�D��lF�/CzD�'o���Rs�Qb�$���n� �'P�1� �\fꍈB�E�����'�<�YE�03Uh��PI�U ��
�'p)+B9�������y@��
�'���� �Q�
�q� )C�HЮH�'��8�J�.K*����^�?q*�+�'7FuC`�X�s>L�"'	�4���"�'.�e0��H	4�1�A�<(�ީ��4�Px2Ɯ1Z�%!vN�-�h��!c���=Y�{�A
�TU�]�fAU#W��uC��E��y��G�_X��r�ܣ`�������yB��s8���!Z�M�"�A�D!�y"d܀N!ل�I��Չ��؇�p<��)8�~�PT`�ːƒ�*�!�d�܎A�+XB�ȑ$�,�����㉴ NdxB��ïL�h�;q�E	��C�	c.��`�,x:\pɃ,)��C�I	�乢6o0˺��f ��)h���d#�I;F��'&^��0���8B�	�|�<}�DE�<S�ASp�U�6B䉘Z�T��f�j2TE-�\��C䉸J)�1A�͟}7D���,]�B�I�g��H E�H�w� �*�H��aC�I�2�F4x�)Թ!�@ `�D�]f�B䉰g��\x&f�p���q�زn��B�	;/��(��J�4�����Ҩ0�B�	�Ez��-�]X�ʓ�D�B�I?G\�2"Q�ar0�CE���2<|B䉝q?�eC��4�T�V�Ϸ6�ZB�I�"NT�	4ꟀdGd�А)N�C�0B䉤'[����`��;������
E��B�=K�N�A���(�J�Y�B�Sc��p�`Y?"�:�Ѷ�Y1f�xB�� |^N����X�(�ʲ�C�W�:B�I�D����&�#+��2���2�,�>���	Obx����R K\����)
5!��O =��У4��sj	��%�)�!���4s�t����-|؅��m)G�!�DV�
셂'-�4�~h�e/�.�!��R�ފ���Q�"B�ٖ.�<1z!�Y�d?,ܹ4枩Q�u�GOD�J�!�ٰR���D�9K��)q�ȁ/<�!�D>Suv�QPd�z	��R��E�vf!�$�!M6BY#!`�7��#P��$9v!�ĞA�����H�N'(M�@J�-u!�$.%tA��!	|�rQ�^*�!�$˧$�r���mFN�3�ȋ�YW!�V��)��-@>/�� ��-j!�$4�l�ۗ�ߣ2����Ŭ W!���0m�y�)�=� ��%�#Q!�$�a����"R�m��XR��Ңr�!�J�b����_�"�lI"!l�!�͡Bl�큵Iճh�l��)w�!��_ܙВ$2@e�K���c!�$[5o�>[&`H�@H��DE �y!�d<z���� �C�x9�~�!��֛%�
�sW.-(p�'D^�)�!�dܿZXRE8��K���@�˶y!�D՘W8��(G�\�	O��AUW�K�!��3��ħ�*CRm�GG8_�!�Y�=`@�ڴ#�;I%�Q�Ʀ�k�!��  �Te��t-p����T�+Y��"Ob���
�	7z^-��&�w�h�"O0�#�� D�Ѳ�0Q��i��"O6�[� V�	��h�k��U�V,�u"OޡCc�!��v�C�A�9�"O��p++36<5�F�N�\� Z�"Odm�ag�tm�Q�HZc�B�ˢ"O dX6_�-� ◨	�9��qIv"O���޴�䑲_M��Qr@"O���V�Z�2*.0�DF,�踺"O=�gc�~ަ)8R�u�5� "O�E0��$4]��Q���3���{d"O.uX0c��3�x�2q@���r�R�"O���%e��6����6I��]-�y�b@!O��4��F\��Mr���9�Py��G��D�����M��rfS�<��a!c�a�Ċ� ���Q�<��L�i�2�g�.�Za�3�	P�<	t�� ZX�����Ԑk�bD���BJ�<Y�)�LF�hD��
y�x�"&#�n�<�ЮObl��K�%��@�͒glCT�<0*�(R�Q)7��<2q�@"�
W�<�DH�PT �;�["~�^�ڇF�Q�<9V�A�TX`K��ޤA����L]K�<�#�G=uXK��C����!	�$�DB�	-/$�q��$����C/�Q��B�	b@�C�&��?��<�v#��oB�I�`�����\�> �@2p�C,f�B�ɜs�YӪ �;~�Mi7�C7}�B��JF(J��W�<��B!�B䉐2�Q9���Z:"�,��s1DB�I+	(z�Ġ�.:����6S}�B䉓&<F�� ��.��|���'��B�I��R�B^�#�ܙ;rj���C�X�Z*���j��A��
D&qC�I�<#l�+B�{��Z�8Y��B�	�@xD!s 3F%�����$>!�����d�6/
,S# �x��7"!��[�0��P�&6#P�i!�s!�H	��1!6G[�McN�@M��J!�B���mkЎ;Q_�@ J^�o!���!6���K0�%VF�e3�B��{!�؀P�YWd���z(�76U!��D��PD��C;cP^ ����-2r!�D��6�t,�7�³y_��PM*S!�1B��ȅFXA����7�ԃ Y!�*�B�&�  ���r�Čo@!�ЏG��K��$>���R�O#!�d�uN8pTH3f�͉�-\s�!�č>r�Bj1ZZb���*W�Qr!�dY9Bn5ӕ�ulڝ@��Y!�d�(z���`O�hS4pA1NS# e!�$�ExM[��'jH�����b&!�D�x,	�!�(8@���NE�w!�d��!q(-+G�ߒ[��M�5�ѸN!�D��e"h��އo�&M1�ꎵ0�!��fC"���^�!!�HR`��!�@�M�D��xr j4�ۥ*�!��\75�R�*"�<g]����&�5(!�-H�Ó�ìmY�h�҇� ;*!�$E�R\��M� Y�x@���>�!��zI�Ƞ)�fG^���NB16Y!���*vF2�Oʗy4���n؏@L!�$A1rΌ�ed^�,�E��o��]�!�� 0�f��
� ����4Q��ZU"Oz��C��^ij�V���)L��R�"O,�2�"B;|�UmZ�_-��'"O�q�R@�4�����A� ���"O��0�^�Y�D̈�N^(i���y�"O�1╉�'���ʏ���x"O��ا��=7T2����^�@�p��"O ,3F��!-�PY"�íK��|�Q"O����hV�8u>12��V����r"Ovl�`�Ag0��a@p�XX�"O���	�"���AH�\n�Dx$"O���'ҳ]6�҃厭B�$�3�"O�Xb�eT=J�����C�<n��� "O�9�0�8�^ 	#��=��mu"O��cAVd����t�|���NF��y§�~�rZ�� � ̮ 0�`�<�Py���3~Ҝ1�0/�<p���b�$TW�<ɱkW
)�������Fr����h�<Y�#V��*}B�	EY�VLz&��e�<I�j�4Q�a�%p��sK�e�<��(әL[>Y��o��I�j}C�b�<A�
S���CB�-kY��R�Es�<A���{C���D��>E�\ 	.U�<fj�=�bu�:.�8 ��o�w�<)�J�9f��5C8}Q� o�<q$#ْ)��)Q��Ѱ[{:x9�	�r�<	���{�zx��F�%=Tٸ� o�<A��J%59,@��j�~a@ �Edo�<���	���<���E0]]
P�6M�d�<����-7<.C��	�W��쑗��c�<yt7ssr�I3ES� t(%�*�K�<��-� �|��_�C$��R$��\�<DŞ�ni���� �����l�!�$���
3.��V�`u�g�W��!���J�<�b�C˹(`�f	�Z�!��&:'v��@�'�U�3��$5=!�d��h��*)~��Ad�/E!�$ԳD����@KN?;��ږ��	0;!�'Y�1�'�'�]�.A��!�D�����҉ʭc�Ta�6� Gz!��]�7�(�� M�������,h!�W$>�z,+��άm�r�j�(R�X!��Qh���*�=4�h�Y'ݺ8�!�V L߲��Bײb��$�eK��!�d��1�h�2�lG��\�ţ�Mw!�#���kUO�e�Ԁ�#L:yd!򤋻`ۂ��f"��f�会֡�!�X	'�0*$-N-h׊�{`�
�P�!��ƭ:��mQB�ث-��0��0}!��y[���P�O���ⵇDf!��^{�f�{Sj��Gf@� b'�0\!�j>�4�F�ª����Ֆ0�!��
=tp(� ��P�x�t$1E���Dp!�dF�U�ȡC�fJ�ႧB�<e!�"-����$��h�
���f
)[!��Q�(W�P�ch�)*�e���S4SP!�DP"OvXad�� �G�C�2�!�$�0�`Q9�.�&a	h  �o3�!��ѧf��	F̆�^����V>nt!��>n�y��j����&k*c!�ǽf�����KS��x��#g�!�$9\��@�(�y����	�~�!�$՞$�I�M-^�h��NO�Y�!�āZ��x*�C;\�~T���!�!�� :Q���+?8`p��b��s�:�"O�-�� �@bxy�+P�e��A+�"O��!l�z��CI�%��"O��T��6ܠ��g%P%y���B�"O�3a*��yO��Uc�9���S"O�q�F1"�"�H��^��S�"OntK�"[+^������_�2�!"O��(���5	�Z���c3�Ʊ0�"Op�a'.V��# IHm�"Oz�cN�
X�X��H��B����"O��
��$���@1��<��1d"O$)��L�2:��&H�]��*P"Ol	��ˉgN�,*�C�$@҂D*`"O(8Qq	�	$��-�C	g���	"O�S� ����"�\)NO���"O��S$�ԁW�f}��!	nCD���"O��#L��u.�E�W�F�O�P�6"O�aå�������fF�X���#"O��S��;6$,0��&P�H�����"O�ɪ��֌?�DAY0�� ���"O�D���?{�0��B�o�z9��"O�����H�2��.��Ja"O�-��6H���ˍ)6�|)��"O�J1��}�1�3`U�,��qB"Oz�Y�R#r6���d�>cP!�w"Oѳ��H#AZ��I���p\��p"O*y3@��U<����[i�$P"OB$A�ǔq� �d��	T��"O��Bb�ތ<$p;�	K�'9�AI`"O�@��M��N��a7#M�!��pK�"OPx�DM?�̓SaB�1$j�� "O@�	�FҤ9�p��%�� ����"O�%�#��GT�Q�a�	�Tn��rU"O��� GK2MZxiB���gb�Iaw"O���cm
�n �������}K:$`A"O@�"�k�>�M�5��3u-r��"O��Iq+[�<����	��qj�S"O�t�A��&x�q�i�(86ޥ��"O
 Jr��)W{�@��`�P"O��p�	��
QȐ�d�q��"OD�i��ϓzb43��F`
`��"O�A3'��,s����0g��8Y��k�"Oi�V���S��p�!ő�:����"O�؉��#r�x �A#�0"<yCE"Oh�h���M���@��$E�TX�"O~X#�l�  Y/cr`�"O	�Cȍ�G  ���3
=��"OV���lN�k���<]�2"OƼ�"�I;2ed�ڇ�8$٤��"O�՛�ᖧ{����4 ��h�ج:�"O�,#wF�n9�a�u(ٛ:����"O��7N]4zcB ȕFԐK�,D��"Olij�U:%�y��'0j� D�"O6IՈQ�S�ȝ�Eg� vL#�"O���"l������#W"O�a��� q�uX�g�5Z��x`�"O @�����.� ��"5�JԠ�"O:��W �u���G�c�b	ҳ"O@`��o�<Y���9s��z�du�0"O���JU�7�G�|N��q"OID,�	z��ԫ�`"@P�"OV(RpC>:h<��	�3G+��8�'��#�@n:2eڤC�%	�����'�m$i�.S⬩g��	�آ��� ^��"�#{m�0!ψ�i����w"O���4�B3<^*Щ/�$E�u#�"O,�0`�L�u]R��צ2��"O¸��H�PYB��G�֩)�"O� �s"�8�f�8PgɃw����B"O����ؐ�F0�/�+��!��"O* z�AN�jd�-�r�;{����"O0ЅcӴ��U��t���3"O�`B�%�6���B�.u��,��"O6D��
�)2-�� S�ܮؚf"O�Y ��P����@�j{�Ae"O���n��<��M*�Jج4zҨ�U"O�ժV$�&�\�,v���"O2�ćAeh�p$�A�PY�ҥ"O@�#�@-\P@�:f�N�*>���"O��e���T����3��Z9B}��"O�HzR,�r�Ry�0��%"�T T"O�	�c�G�*�
�r�N [!(�z�"O��BǛ�P����se32��ʰ"O��)&��:����׵8���"OX�RV�E�4��P�6(��("O��yB$��f����Q�[1s�t�
�"O�H� -� N�pH3�	H��E�a"O�,A�-׍%�Teh�$�G����G"O���n˸v�D�{�)^�`'���"O���%�$	Vedn*����%"O�ɉ��;JhM;��/�Ƒ��"O*�b�O�80ŪS�o�a 7"OT9r�d�|��L�siD}���s"O�� T�ˤ2&�%���)�f�"Oع�5 S2�Q��Kz
��"O^quK[-4R�/�
s*T��"O�QV�ʀDY�h�N\n���"O���#Fʹ��mT��^QY�"Oz����~T,��&���&}���"O��,m*<�ŋ@�Mi�C�"O�!��胭]��\2�
��\���G"O�0�%�C�5�l!!OG�UXd���"O��9���������V�ڽ�t"O�����\�mjW�6[��=��"O��bi� G���F���h��3"O�l�ά;�)aK�d���"�"Oz��M-X:����d]��"O�`��l�$#����ԇ	q���"O"m-)s��IǓ@�����	��y��Q}ϔ�	s�P�/Lp��2�yꙟ-�J(#r�D���EC���y��!D�AA����,[�J$�y��pI��̔��dT�r��&�y2@�+$D$P�m��	xu��y�nʵ�P�'��~�}�d��;�y��M����1��,v��<�s�U��yB/�( ��e�E�	>��pa�0�yB���H��x�#�K>:�&�;�����yb	�����(
28��[�Iȃ�y��?����l�#pb4���ĳ�y���JѢbھ����Č��yb��A��\�1�\&��s҂��yl�:|Q�k�a�+x���Q��½�yR�Iz�)�'%�$ ~�2�*Q��ybA�&T��\`Cl)��Q3����y��-z������R����kٯ�yR�ڳ734�"Qg�/}�tq��f0�y§2����V	�f��8d���y
� ���j��@���[bK@3(Y$I�6"Ot���J�|r���싺=TT@1T"O��z��2A�:��aJ�)c"O�tA�������T�U�\dL��u"OR�����(T�Zxۀ�ν.Z,�'"O���� \h�I���)w�DAQ"O�	���Dd����i�t~<��"O�hR+D�~|�R��-��3%"O�A$��E��腦�y�����"Ov���9,�������+�"O���PHA�	���*\� �����"Ox�r5�\��(�V$T&���"Ov,;fa��l���]��	c"O�ъ���p@!ٖ��/f H�"OFl�V�[2���#�>D��x9"Ovl�Ā�f�p�c�W;F�9�"Ob���F�2Dt��s(�*1���"O�����~A��⨌�	��)�7"O|d�� }�Ⱥs��=�B"OJ�H�Ini�Ǧ��"ϊ��"O�R`)W�w�z\���\�_�B0�"O6����]�`���ZjĨ�ء"Oց�� Ĭ4j�����Į4�av"O$y����[���'? ���S"O�kr�ƃm"Z3���7ʬ��Q"Oi��ƒ\[�a�\!;��P"O�@ ��Inv������d��)R�"Oz뷩�,n���xq��I�B�#�"O�|�q�W�v�T���0'�(�R�"O<!��BV����Ւf�:�"O�|�ů	�.2�(��R��U1�"O��剋ZL�m�"F4 �-�"O��YV"'Ӣ����#x�,9`�"O��d��$j �A���h�VX�E"O�z���-a�D��C�Vyt�"OXe c�׽v.�#D�=q���s"O����YDI1�Cn���G"O���5��0$E�P��ZG"O�|@�AVUG5C�,��*�0L$"O���"Z=(�j�Qf�.j<tyC"O,�i���1o�V�ٓ��6���"O|ekE�
&� �y'b�#G.�xS"O4,y$���4F�8����S��$(�"O@
W�݅+�2ac�f�2^s�ä"O�L u��Mb�]�k
9�8�i�"OhuS�O9i����,��`��3"O�1�C,]<\�P֬։N����"O�f��$|�p��k�iƍ�"O���`Q#;w��bd�/#�\���"Of�!Ĩ\,N�=�@��]�D3�"O}@vD�n�X`��Q�=T��3E"O�)X`�գY�tl�àӁSN��"Ot�p7n�Y\���O	� 6�X�0"O&���[�R-��փύ3J�)�"O"E�u���Bh"�p�"OLj�o�gn�O+��Q�"O��)Qc� |�LYeA�9g93�"Olq S��?YP|#� �%�����"O����I�>t����ԉ'HD<Jg"Oa9Vm��-U�E�3�\_?z���"O����K\�?jZ)��CU<t0�u��"O�ͻM�>ol�����4�X�i�"O8�x`��;��b�D�F��Jr"O�誕k�=G
!6���HH��"O� ��m�)��	t ��8�"O���f������%"қ'j��"O���S�Ar��nP)7z,��"O�aqb!��v5���0.���%��"O�A j�-5��5rW��-vE<|3�"O�x�t����,A�1�</6�:c"O<U���!-ѮYC�a�+x�ɔ"Oԅ�1	6YAT����%'���v"O>(��J�Fo�1򧘨&svi�"O��
�LE$<�8a�m([2���"O�Y�EP,�r�R�-STHl��"O^ᵭ�� ���!4�K& CA0"O�}SA�Œef����Z��Xf"OL����P�DP�Kʤ[P��G"OJE3O����z6���G�U�F"Oޘ���ڄ>����AV���r"O`���%C?����玬~3X:2"O0�K�O�XE�EXq W.3v8�´"O�1�r�(xf��d�şi���T"O
(SU~�TUK�h�3RfPeQ�"O丙&
�&G"�rWH��C]���T"O�5Y�GW(��Y������3D��ӡ���dX��#���e�����1D��Y�b\<9h���Y��#V�0D��b���:cONa�φ3.�z1���.D�ہ�G��a���W=@�:�?D�\���
#)�i�CI�r�cQ1D��3��[�[�h�&��N⚤�ae.D�ԑ�(��P��q����rM�\��%.D������@�����v�j4x��-D�SP撖*��QS�I�N�.4�'�-D�<I�jB%2�:�8��TjRct�*D��{t�H�\��k�\���a��=D����Ɔ�&��8e#�	LrH����7D���39�P]�ť�R�N��b'+D��#�F�B��עa�Ѻ�#+D���3�]�R�i���&�U9��)D���d�Z�������
Z�A0�%D��ee�"�6���E�\2P!D�dH��� �~1����(�����;D�ԳT*�%��X�ff�4A� 81 4D�H��̕6Nv�HՋ@���/'D�48��%{��+0��+r���B$-'D�����)d"PʄEރmI^Y��)D�hZ!Z�<�҅D��Q6:��!�1D���"��uE@�*t�&E)��,D�  cl�, .���F� � 	y;��+D��[+B�:�4}ۂ��:B0S7�=D��ғ��^,��Fa�.-!����&D����;Z ��x4��j��"�$D���
�!$8���K���R�?D�8���P�IS��Rj݂R|���u�1D�|*�
t��5�s������m0D�L�*I�	����c�@��+.D��:���me����U<
�D�#/D�l�F�;	$��ؑ)B ȸ��i!D� ���
w�zx@&Â�c�l���=D����CK޽��)���R�{�&D�,�#M0lNd��v"���.&D�����?	@= d�!S;N�b�� D�d8t��[���B�,�l� T�3n3D��aL��Iڎ|�ëݾx+�`94�=D��^:b8��kI�8譸A�;T��q0M\�`A[b�M6�&9@0"O� ���학�&U�#
-Q��<#""O����]L4H��^�V���"O�b�͍�il0| ��	���C"O��;�ʂ�^�xX)���zZ.D�"Oz�Ib��Zۆ$�e�_W���Q�"O����n)��G�"
x|��e"OI;�$!��:5���aA����"O�1��&�6t��8~8���"O����m����jB�OM�qF"O.�ҥ�X#2Z�h�Z=�С"O$`�W�Em"Dԗ
��q"O����\9�j<����U�����"O]�e� 		���e��FQ�"O�%(�k��9�����2-���'"O8iz3���&!|�J`�ʿ%���"O�ASL2Q�N��R+�=:�����'�h\����8e�*}ku�M�E4����'���ED�U��DS���n��	�'���eD�����&`	���'���H�GNo@z�$��d`�@��'vT5�t K쪕*��X�|���'��P���1#��DxšTyM�u��'�D�8�ڔ8��(��m�r\J\��'Z������{9fU�B�q��R�'@�� ��A�G��u��BH1�'�XpCF��3�`��N2^���'F)��L]��a��\j����9��;��݂!��5zu��,�2�ȓ6J�y�e��z���k�K�)��%�ȓj�x`��J	�l���3�dM�~}Z������;��{C ��,��لȓR������]������8F{�$�ȓdi.Q*�'��C�H%����f+ @��N<>\as ��A�����%!t(H��!|����H�/��hE]�\ ������$m���x�k��џKk���ȓa���s�DI��BL�9��9��l��-آ�ºO�L1���K6I�ЇȓD0i���	�&|`B�uF
Ňȓ?y@�h4(),}�4���9]� )��$0�l�A�VҀ5��H�4 s�ȓy���҃���(A�h�&Յ�x�.�Ƃ�$,6��jZ�v`^<�ȓ&9�x�)��-D<���͉�	s`���Iڌz�K�s���Q$�A�}�L؅�d(L0�@�)*�CӮ=:��ȓ@�vJRĀ�h D[�J7$ߌ���d48�eU�J<t(@�@T�p>��ȓ_h���q�I9x�>d���G3��H�ȓ~d�r����u��l!�( ��������g�\q��K1@ǧ;�^���PHL���u@x���'�m��b�B�CcD�ۀ�U
T5���c�,uY�)��g��Y#3hJS���ȓJ���G*Ҹ`զx���A�?����d�}��K?R&z�j�"��M�ȓjVP Rˎ�a�t��pR�U�����~%�e8�`Щ@�r$ub��?o���ZI�D 揑�H�袥�4y`��>���*Fj5�0��%�	4��q�ȓ@�����P	ʮ]!Я\�u7�]��2��3��@�]V�S�@�M5�|�ȓG����p�(L���&f0&
��ȓ���h��CJ��1#`��(:��Y��S�? ��*a�"g��}������>A)R"Oz�OīC%��(`�F�~�^���"O��v/��b� ��F�1��݉�"O��P�ᅀ3>	ʗ'bw�t�4"O�j��+:�ݢa��2�f���"O�Bef�o� {%�^%*�S'"O����+/#Z<�K�D�"8��"O��ɕlçWq����d�};`$	�"O`:��x#�������g(p�#"O�m���=>"�J!R!�x�""OD�Y���FTH$C0�ֽ��
�"O����WaObhB'��=x�"OT1ʴ�\-*莹��h� ��Dq6"Or�ҵ�ي!UJ�)��B. ��H"4"Ot�GP�Pqr�S�*�H6�1D�pJ�� Lp"q�R
0���j�h1D���J�X���� �o��A!�/D��!E,��Plxj��=W�����,D���CխV���c&�C�`r��.D�����S$#��m�Bl�x�R�Qo-D�"adέx��LC�h��$s��.D�(�T2H�&�se���T\�4��M0D�t��&�(?��X{)\�<���0��!D�4�W�XMg��b�i���[�-+D��)�@
�Z�P����P��ý2j!�=���q�R�t}�R�R1GM!��5{^��q�Y�Z�1���S1!��M$tBXi�D,�%d� zt��	�!�d٬aS���\�=�JA�4�[9`!��3_V H�A���R@��ɢ0Q!�ݼ"���n[�iVڍ�%�
�,@!�d�=�m��l�;Q?����A�4!����Wh^�Rg�$jh��m�%!��� >����׀L�t]Y�	�Q�!򤂞�bY��İ
�2�r��:)�!�D@�l�$1��s{LU�ϗ�*!�d"h[��#!�wB�{P���!�DK	
�Q��CZ��	�J�> �!��\$@�t�:��F*|:���#�sC!��Y�;^Zt`�1$ �b�54!�D� >��ѨHΟ$J�y�A��;!��,{i����ZxeiEA��!�ȋT��3b���~��f��!��@W�\yQf�8Q��C��?J!�$��D��MC�-�/W�\�Z�:�!򄕔<D0��W��wPiRá�6�!��0V�͋R�	 �* {7`���!�$�6}_04z��E�,v>��ΚC�!�$ŔN_H�C*5���`d̡-�!�M�fJE�!hM�;o� SwL�9e*!�D�
~22��w��;_T�W��17#!�$��D�����+m��nϸj!�s7���1H�o���X��֋\!�D�6l�i�M�.��=�r��=!��I�"�4	�����F(!a-�i�!�$J ?H� �B {}v�z�*X��!�d�=\ݓ�c�!^�52��0�!��]�'�^-����eM<�"� �G�!�֚|E�$�^V҆�K�KZ�~�!�X<M�N)��Ԕ) *���D�!�DNY�Ds�C89�%P�C�J�!�DżL�����^�_3̈j���H;!��3.�z�	Uf��x�2�@�Ǽ":!���^� ��Cq���1#Ƭ�!�� �-�t��~�ج�F�t�l��"O�-!A�ʃ �,)q���5>`�"Oz����;��y�*�\�F<�H�<i�*˶_�0��	vv(���l�<	&���n�ʑa^�c<X��NA�<��M��|l�Z�mB7|qщM|�<aQ��7I�z��=J�f��&Yt�<9r�Y|n�����q����#�n�<��
NV�R4�\+gj��k2iTh�<��S�H	H� Ș$b.���f�<��j�o�r����<����Ee�<���B2P����]��EJ�&�{�<� j�H��ы��P2�q�5i�{�<E������f#2N[N�(*#�C�I<?��10VkT�!�4�D�7?��C�I��p�hsIЗ@�ĈA
�>�nC�&7~`�R�̊~�d�X���*a=fC�I�w�������E��k�c�D�vB�I>Oq�Q7)G8MR H3��8!�
B�I�ێH��U�j��a�D�Ќ��C�I�i��#K��.?�!ħð',�C�I
3XLR+ԲY��9Y�'�J_�C�I�`��t8���(y���0bfP�C�I�W?���1+
P�H\*��[���C�I� ���RGG�,�b}aՎ�>�C�ɥe�N�Q!ՍV�����`اw��B�	 �X�E%��U}$��EX�,�B�#B:t��V�i��I���-I~B䉯]�Q�֨\,�A�p�@�U�C䉒U|lp�b�D�=���gB^�27�B䉱�IcP��G%�љvfݫ9Z�B�������/�#�*��E'��*��C�ɩz�KB�p��(�$荺&��d�"OT��S#մ:���Ce�kF�%��L�ȓx�L��cƎ=/	$ ʑ(2�M�ȓ���Kњ�~����бGǠ���d�K@�1g30�� ɪc�湇ȓ���R�hH�8@b�	��פ�� �ȓD��[��ޓ`�`�eaH�5��ȓb�.��d
U-I�y $/�Ht�ȓh]D�	�Ɣ�_+`8�U�ڔ�Xx��'�,�( 	�0Oᣳ�(Ck�%�� �e�q� �y�(T��c_�O1֘�ȓɼ �Q�JjpV@V��0vg�܅ȓg!�})� ��`�yH��Ӫ1�����A���z���!D��x��C!8�nE��4WF�J�-�Cw^`� ���T�ȓF���h7��@�dU�3�0T],��ȓ?��0��n�pJR|S�j�Ym�9��@t���	2y�0���)攅ȓ2��1�s�� o<�BcȚ|����ȓz�hѣul�����4nВ6�ȓ �2b�	*Dy�'�ŋ� ��5Y����㘥J�$�����)��Z��IEưh��[9-Pl�ȓ+���E�[� >��q��<�����#k�!8cn�KT���r@ӵZ�ȓ ��l�#�b�Z�$�Q�A�ĩ�� �����~��D�p�˙r�2��ȓg��䋥#ׅ/S������I�$���Q�rx���u�� *5mܝuj�نȓ����&\g��	҄*��a��\�ȓ �`�����),�<�@��0�ȓEg~q1��,!�a���E:z���S�? h<H�b��p����@�ʬz�d�D"Ot "��I�N�jCB��訅"OIh 
39� �́x�D�$"O�� 7�1��$�E�FTq�"O���f�4�&�[�@?~��%�%"O�x�iK�"�i�Ó8PT�v"O�����#�h|��EP�����"O�%{�J\C�	�EI;6ZA)C"OdqHd���xb7�Q�|L�SU"Ozdκ4�rD��I�C��A@"O`U"$�@v沱 ��M3$��F"O��:�bƒ ��{$�Ӆrl$���$;|OpAwg��_ʊQ� BKk�D�"O0�HE��.�v��`�	�ԥ��"O4q
��H�O�`E���	z���"O��0jŦF�Z�3 ɗ�ԉ�"O�Q��� �ژ ��
$���"O�E�U�+w�y��ÙC��8sc"OȨ3�&C<'2�e��������7"O��0%eD�Ii��p�E�v����w"O������9�t�x&�V�;�ܸ��"O��k�#Ѽj46�r��V�o| q�V"O~t��D�P�Q���QgT}�s"O8 �BW9�&�{uG�ySV([�"OH{ӌ��8���3'��Ox�"O��iR*جk�,3�ǮKW�̸`"O��J�(y�Z� W�vR|Tq�"O�`B!NWN�U�7��=츑G"O�T��-*��d�B��&�>���"O�uK�/�"6��5:e�8�)�"O�Q��f�0&�̨��D�8eZ�"O,�i��H"��e�+�O�A� "O4l��C��h'<8�fJߩ1鬝{�"O.�`���>1�"@p���W����A"O��*���&����ↇ5_
��"O�Y+#s����ɋ+�VÒ"O��WF,�r�O+"�T9A�"O�(���.&z��U���&���!"O�I��I߰��!p�g�,���X"O��7$�_C��z����"�
�"O�8���<_��T���H��A��"O�y���1jXAH���˪��"O`����5r��;�ֈ��'��r�̔r�Z���L�S*�Q�'�(!yp+BPB�����E��\��' ��g�_�|�E3�Ě.�p�;�'ҺT����H�1W�M~ ~U:�'����a�K��1 @l�?vv�'9�+�ϕ@�<���e��]�(��'�h����-r`0E��-$��I	�'����-�D��@�rd��V�Y@	�'�>$(F!�P��u�Q.�G"�a��'�B �%F��]
a�H�&B�dh	�'A~=��JM*@��0�@�Y��'�4��ᗐd�؍���=�(��'pv�� �<x�=���1�q�'���A�c�iǠI1�4u�$E�	�'��R�M��%hV�.w��h�	�'��Z�+�8072<�ՠZr��dj	�'hv	�4M�/.0I��o�5c�4���'[���@�I��\3EKMa���C�'V�B���1/�݊w�ʵR����'¼H'双�H�a����f�x�'&\!IGa_�1�`[�l��+������ B�A��9cHL*1b�Xqx��1"OpD#��ǰaX�����Ui���!"O���e��z���5O2Zh$���"O�"�`�z �iE*u��4{�"OʔQS�!�>�Cv��H�iR�"O�P�O�X>���Φh'���c"O����H�:2݂4kQ�
�*E"Ob�6k �1�镇6�|��"O���d%\�{���
h�� u"O�h[���/uq�1�f��<L@`"Or4���W�dL�q2�әn耘B"O��)KIt�ذB0�ׇ �T�"O����.S��l�c���X��"O�*��6���瀅9�^i��"O´"E�C-e/���w*�
jæ {p"O��Т�d*$�r(�)s
B=��"OX�Z��l�8�7�5b�5"O�q��aB�+�y�2�±�p�"Or����9��p�Ǥ��C(��(�"O8p�/�<O4�A��ߡ�Dr"O�<q�Z�d�܍@ �1�F�S�"O�x1Ԁ�/��"H�v��- �"O����G1'ݰ(q�/�]���YS"O���ʂ��ĉE�8RR� "Ohp�!䘋i��Q�.�M�� �"O��҅މ1�*9�L���:�B"OpP��ȱW%z5�Ø�D�Y�"OصS7��x��%
�:k�u�"Ot� 2'ͤ=r�ɡi��ɼ���"O�t��Y�v9ӐG� �Z��"O�A�X�T�:�(��nb<e{�"O�A����$�����ɥg[�,�#"O&�����w��a��!���"O�	���T�!Ԗ�eG���h�"O*�����8� ĐcmH=D�.	
p"O�ܪUmo7�����شo�Q�"O&�iD(�0a����.SZ]hqE"O�8��B�et�qT�Q$�z�"O�e �M�F|� ��c_�BzI��"O�� �hI�yz��ðD"vֺ�� "OVM�u+�J��iʀ"�;W�ԋ&"Ol�sDm	Yo6:сY�J��`��"O�YcNSp�3�I�`y�X�"O�q[$�$$�$����$LL�3"O��@2Ɗ���A�VH8�.+�"O`�s�$�8gD"�z�ҹt&�x6"O��3u�($��%r�b��:CVa"O���qaS1)_V8c�D�X;TD`"O�`$%L��T0Ӈ�̥C)�5��"O�0��l\.ޘqU�H��&�q5"O����I����	آ\�f,�R"O�yI䄫*\����2Yr5x�"Ov �U���_�\|�.n�洨C"O4��-kD������у"O���$�ܿj
��h��U����r�"Ot,�FI�1<l-�U�HV#��"Oj�ң�Ɂ	���C�gC$#t�hh�"O�)�� T�HAq���J�XQ"O�����˦$��B�aN�C�"O�YUK�}T�aAoFB+��1"O<tT�n��zVND�,��4 Q"O~ �Aϊ9T�, �M6�)x1"O��<�#_;��HҬ��IjBɅȓG�N�3''�:��:Q�2�2���S�? Ԉ�&Lc2,A��V #%"O��Rȉ�l2����S�r�"O��XыX�]�ƅ �G ��٪&"OV��c&��J���fF�uܚ��s"O�5s�ɇ0	�x�C��*`\t�V"Ol���Y81��#�!=���"O(�� !�'-���C55pӓ"Of��V��e�����_P4j!"O�-�0e$��)aկ%/�X�"O����"N4�HV�ù2J9	1"O�"��f���5�[385;�"O�Q��L�����C6r�jtK""Ol@�Ȝ��dTCr)N	C߄��#"Olĉ�BX��^=y��Q#���"Ot��U˘�1B��CE�%Rj�"O.��Wb!l2H2�"�U��y�"O��	$KW��%Bp�K�7z���"O�����jF�U1�*_�[��V"O)����7>z,5`ϋ_��,�3"OZȡB�R�E��p·O�v�b��w"ON!ě
O䴣���Ӿ�"O2�C�D�1o�p�(��t'T8A�"O���q鞊9��i�sG�a���&"O��WۮI���wނ~ �9�'"O�|���'�"}�'���Ej�X�"O���J1v�P�	��J�\���r�"O&x��B۰���-\�*e9E"O@�hF��� `�����# �����"O,�I�����@P_)p���"O���#�Qbx�J�`�qx\t�%"ODJU'0o.]�g-MB�tCe"O���*�<AV�A̔��P�z�"Ox���H�?o��r3K=�Ve�F"O ��,��,m|"w�M����"O�9��>G��dmT� �L`)�"O��v��f{*��K� �b��"O���qM8���ٵ	�!M����E"Oȅ��*�(B���q�'
$wt ��"O�YCB=/�lQ����w_b1;�"O>uHVeП!�RY��E�CQ>%��"OjY���՜}2��Ir.�*ljX��"OP,��C�3D�HH�l�7v�^չ�"OD�S{Ҹ� z��L�0"O��C���V�Zi3Bٺ4�^��w"O��Vm�	u`����EQ9�2��E"O��ӵ.E<=��He�KC�21 �"O��;4�Ň|Z`��ƠF�30"OҜ��!�<V� �ΐsL.m�"O6���_�<������DK��y�"O8З8T0��C�66@�(P"O<!I��îvˬ�)���?RH�d"O~�e�А)���#B?"6�� �'�� �0�> ���� ,x�'d0L���$�l�;��d}y� !D���%��PY4U:e��=��8�G=D����=kr��\>(�x(<D��Bb�U�2���K`�ښX�l,�2�,D�(��oA-�tu�"�Z�P��=�� =D� ��֥>���%`έiDE�2F D�Pz���j��Zq��cFYJ֮>D�4;cNVL����Ț"��� +;D��q@�{((D3��G;��D���9D�1�g�_g���D`D<s7b:Sc6D�h��*,20��&�@�v�$��4D�� &#���cC��I/6<�n��"OnI!CK�fS~As!o��#�8���"O�ls��G��	Bi�o✴��"OxY1+��� }��NG��pX�"OH���]�ez�h������e�"O�X�v���S��F�"�NUJ�"OP���ۤ?!�X�.�'r^�(d"OD� S�дh&��S���AY`��*O|����2��##�G UP�k�'F�X�5�E�j�H,1qm�T�Bm�'��8��͋[<�"Q�΄S��Ts
�'�ȁ�]r6-1��P��(	�'�\��q��:7̄bS�C�Y�0�r�'+�+Gd�!y 	��V��c�'��J��E'"y���9!��HJ�'ҠY�/�g�ݙ�m�(R���'�V�{�
�+Lo�X8pj��MrP�'�"h����=3 �灈�(d$
�'��t�q�%r��-K$�����'�Xa��Ռ5��eP����s�����'��x��[	O?T�[&�R�i�6tZ�'���V�&4[�.S�h��H�',~�rE`�5[^�(fa	\$R���'ln���R�b��&P�2!��'"�U�w�]0Vl��	U�1��8�'�4%��/�N]� ���җ&;�@`�'�Ȅ#5��2��!�᭜�a�'f�]�2ѲUN�11��/���B�'"�Wh#T:!J���,X~FP:�'8�|Qc�
�8��x��aA�?�Fq�'�bx�4��	t��0���/FήxY�'��03
����{7%F�@Ұ4��'��}!����/=6�0t�L�@�a��'ͦ�plg�R���
4�|$��'q �Z�i�#��8F�X0X@��'\�-M?@���x� Wl2��
�'�,��*M�W!������ddZ��
�'�ڕ`Rk�L(fA��)��X��u��'���L�1@�D͙�hHzT^�b�'oҜb��Iw�Jh*���|��q�'�:�Jv/L  Ebi��v}���''~�b@Z/��ɣ�ˌw�h�'������y9���J��)
z�'�@�AO��y'���N=��lz�'�`$���ԧ-4��� �71����
�'m�٪��W�>y�\��Cζ&sR���'�����'[:H983I�
wҜ)�'�@��� \��Ib!ƿ�"���'��"`�� ����5�Fh�'�ʝ(SÍ�2+�H�`5&��PS�'�~1�7r6J���CԒ��8�'<�R!.�IdĴ��ۅax���'O�q���G��P�q�	c��8��'n�qr��G(,���L�a߼�'��8�Ԇȥw���&$�Q�4ZP��Y�<I�A� �LR�h��`�(�b�l�<���&�����K�*m��A[h�<�9��|0��ȋs������y�<	 �V�
Nh����<.�%�Ût�<aǢ�Cs���۸-�^<�%GQY�<�!/�0I�~=��HV�g;~]��ϋ_�<��9J��$e�3"r�ɲD��e�<)GW�(l�&!�_��	Y�B�x�<�v�Ңt;ؘA��^�n���0��M�<� �	8�.M%�Ҝ��+�4I��"O���ȓ���ir,�L��'"O����(A{j�A��^|]$��'"OZ�e���]NqQ� 'I�Zt"O��iao��P�Da��H�ֺy�r"O��m�5��KΚ�ʸC�"OB0�-�$O�� ��Y�R)�"O�P��	U�.��a󉔇6���P"O�E�%a��V�J';�bp��"O*8�b�$~�0�gH�0k�d��"O.m[�h[�D��W�K���d"O����@ �>�<L2g�>,p��F"O����D��q��if��vz��"O~QR�\�u��P,܍^�&( v"O���IH�f� ɉ��-�
y"�"O��хf2Cx��#d�8��\q�"O���#���yZ��M�]r�e#v"Olp�R�,`�Ȇ��Vr���"O�Y�5��q�������1�~4��"O�P��F\�L�H�#�͚1v� P"Of,�a��(*��*�,�	Ղ�g"O��zT�ҾH��Ĉ��� \�B"O$踠홸k_�X����u�0�Zu"O(Ԁ2b 4�tupe�5��L��"Or ��f���:��
����"O�ÀFY�j�h4��D@e�l�"O�!Ñ䊖5J09�ȩF��e"O6�K �1lxX�a�H���q"O
�qS��B=�ܪd�;e'���CGܚ�Px�HϝU�P���ҔyIv8���ө��O�#~J��Zܸ�@�ʀ����OO؞���|2�/eV� �O#�,XS���3���5�S�O}����CS$����#P��zN<�M>���iI�4������H�1;D��+�ў\���?D�)�,��;u~5��N�D9�L��	b�lJ��A:|l��V*�:��B�6i����F�!\P�ѓ�C	"RVC�I�����3a��9�,]�l��#>q��	�(v�a�U�_W�t�!��H�kQ����I -��<��C <��p��+gՊ��g���'����R��ǆ^"�$!�K��C铢�$5,O�$�u+: W�!9�c!�h���i_ў"~n#T��p�����
cZl�!$ϝw}
B�	,�FyP�'49�L$�'.K��c�E{J|JgI�����V+�+ҼDU��Z�'l�?��$`�:^,�Y�a��b��H�Qo���O$�=�OW���U��	�䠐�	��H�}��)�ɂ�#ƚY�rL�Q�D�x�@��i�Q�Ї�IY��5hcM6���@�O���h���ؠ*V�E[&n��:5�Y� f�!�,��<����$,:��roB�.��O��=%>]I�ű8x|8ҕ��:?1�M#�5D�|��%�?)5���eC'���s��/��hO��+(R��v��q`:���p�B��4}VЫb�l��;��!c�6M�>!	���c�	���-Yl,z2-տ�hO?��B/9�0:#���Et���L��RI!�1C���UO�*4fe��lI�?3!�`/�y��R-#��)�@�KQ�(Ex"�~"��t����tdW4�eI�!�D�>p.XQQ��H!���s�U�	!�ƴe�R�������]Xc"C�1O����ZR��Q���Ӄs�&�	���'��{R�æu�'�l�e��)ub) '�?'RH����� h����J������|j���6O���i5��M����/w�d\@�O�"T��jp$��yb*G/1�$�#sd���
 ��'�<�*ش����"|�'7J	�Jm�vx���$Ү�����&��Ya��W�^*�$� �
2~���"Ox�Q7QўlP�	UQ"���a�O���]�S�O61X�m؏G궜���jP����~�]:~z�H �hE�m�T���y��9P�"��Y<J��}�#끉ܨO"�禅�d<6\8@K�;\ +t���d�'��D�>E���+s���Ó�^]���^(�ў��ᓿy&��(e(_�O��PaOmX��p��	�[ X��s��h�!T(֖7�c�D{*��6�§A�J��3����%�V��"��"O��Q,�.�6l d� ����"O�9�
ڔ"� 1"p��	b���ڄ"O�#�Ō? �X��˺R�l�8�"O�8�� ߶{�D�3��7?��D�"O��)R�|\��:�	��Ϟd;T"O�#�gū[����Ǎ�,�D*3�D,�S���tU�Co��$wzp����:!�ғ'`%qÔ�qZ�Ph�n;d�=E��'D!@��E�e��xi�I/�zl��'�L�J$ +�ݡuK���ę
�'?��B���p�~,�@��� j
���'iz�EgϨm!,Z���޼(�	�',p��tJ
�q��C��Y�8�+�B'׆�O�a��T�Ŏǃ}�p�!�-�.Yrv�ȓ[:
� ���$<�D�!C�(L��Ez�O5O,b&#�=~�HyhR�;���"O�a�D��':��ɺ3��%h86�i2��Ĉ%��0d焄N=���D`0	�!�D1>8���
�{���Ku�#�!�5j�x��N�Z�V�3oߺO\9I�'��	�'�v�S/\��̺~BX�MkҤ�J��5�ϡT|&�2s��4{Q�C㉲VN%B��=q�d"�ْ}/�)S�4�~"1O\��2�~���Իe N R��0haAS9O$ �F{2<O����'2�Dj��4@������6-ް��	�v�����i�|mZW�:�j�,�`h˱y( ����@�6<�����ē' X�0���UP6-��#ǯjx�ɰ �%$��y T [R�� +w �����;�I��`�?qO<�_�i޼���/�i�����O�<��I��d�C��$Un`�.D� ����'����<�����,H�T�
S�C�#%>1�$M
k"�zB_�T�'���C�`��:T�d�Ϙ�Y������$�S�t#��|(�@� 	OI,yb�#����<y���?vU��j3oٴd:6H�g�B!��c��A��AJ3xq�2�G�O��	X�Oc���F^5Qy&I�����'f�;���j�|k���zi2��F?�O?�IX\��9��X168��� �J
v��d�����V�U0��Ce�;U�qQ�E�)?O�<��d��D�(�%�^���Hl��r�!��P�R������4"z�i@�ט_��	C�� 3E�~����Y�]�ԥ;��,D�ԩ�%��b�V.X��Aa�d8D��Z���0T&l�����q�����-1ړ5��?e��G�t�e9��� i�yaEE:���\�*p���f!Cׁ��u&E�R��P��?��R�>����V�ذ�юY
'+xeiB��C}��>a�O�#}J�݌|���Q�K�-L�A`%ݙd�EɧL�g��<4E�_J���#��Cj,4�SLi���	e~2��T�M;�?%�*��ԁ�yb�'�$U�"ωE������Z%�r9������ fYR��U�@��b��C���!�'a�	�Ui�T�@��I�@����P&'W�"<�����k@��W6���cA�h�,��ȓ}s<ub��;D7�(�ML�=�ȓ#.�`!KQ�~�J���J�`|9�>��'i�>�	����cf�\�34����Dz�B�	k	�t�)~�,���eŖ6͑S�'	Q�ءv��)O➠cf�]�!�~l���:O�cڴh�z�$��Z���P7|�8��ܤJGx�0�7D���
E�2��C"nO�:�n���*:��M�O�-��'�)cUr�-����(���'2�䙁DR��-�Q�����z�yb1OF�E}��TH� ��49$(��Q�X3J�\ �'g�W�r� Ci�v<�j�\�'r�'�O�<If�ZDib`S�P�@��  �Y؟��#єI����qt��U�IB�@�ȓ`���Z&��4�ؘ!�O�<�v����q�'�)��ʙ)B��Ń��_P���c	�'�
��1l�5��dЖ�1G	`ݩ���.,O,�a��Q�(r܉BTo@�)~08��"O��d��S�eY� �*��"O&i���N> �훯?���y�"Ov�HFǐ~�@�H"�`�@)@"Of��!�Ҁ(��M���A3~0��w"O�d9D\Fښ�b%ҏ7^�QH�"OJ�k��x���`��^���+&"OȠ�`��%[�:@��E��?����"O�5��c�0.זq)a��,�v��"O`m��M�=0f��7�rÚ�Q"O-� �)%����L�%��T�"Oޡiv"	Dڤ�ci�C� �+"O^�����i�2����Op
�S�"O``��@�8�^���f5PY`yK�"O�����?�$t���dN��"O%17H;�L(�d�Ǒy��p�"O6У�DM4K�V)�!E%��L�e"O�|�����\�&�ϭ{���"�"Ot�+Q$��F�0�P�A,�\�Y�"O�E�P� /"rP�Ps��:��eI�"OA(ef�K���St����hAp2"O0XAD'/
�4Tۧo�2{&Q��"O�ٱ��ǯ5���R�^:^�"O`@��@'<8&\��-�2iTҕK�"O���vL�;��HJ��Ь�h��s"O��0�H�S<�2�]�a�pы�"Oh���1��!�oב?�j1�"Ot%w�()��uho�8{8�!r"O��J$
�&��Y�5˓V�j�Z4"OxZ�e�-�4��3��d�F���"O��ۑ��e���t�!m:��V"O�HY�I- � ��'�ǡPS�� �"O��I��ۻ2�ҍ�_�eADd�e"Ov��&�:�ub��9=�I�"O��� ]�i�*T���N���3�"O��$IQp�<aQ�����-:a"O��Ѐ�FSf��4JG 3�f��d"O~�C�%֫v�аE(ƽ�d��"O�\�ϗ��8=1�ff�`�!"O�{D+�갔��j��+�}'"O��rT��jXӆ҆#"��X�"O,\᎘[;�,�P˝�:u�C"O�E�5�F�V�:��q��0?����"O��a��'_!F�Q���ވQ0"Ojɉ�ƆpMQ[y��-q c��<� �-�c�L5K��f ��A,�V"O\�	sm��u��$�	I@|ؠ�"OxL��/G/P5lM0R�I�o�"Ob-	���v�ଛ�Ϟ<A��}ɳ"O�{4�X9Q�����-X�u9^���"O�=��M��MV���ץ���q"OL�"�$Ì�N	�fD[�h5ډ�"O�\4�E2^������M��Բ�"O���"
0ZE�r�3���ʇ"O�LX��X-s.q�@�+j�zE"Oj���D���AjWL-Ud�f"O� ��c��2��"��޿\J��V"Ox���G��2�30��6�=��"O(�c���\hmb��ƥR�F"Oj�!��,�n�x* �jMzB"O� ���ªvOrMx5HT<� �"O4���AL~��K$�رf���"O*��slI�X�&�#GYx�:4�R"O��ڤ+ߺ6�ֽ[��Ӡ/��9�"OP�����\�z1#3��<g�L�p"O���� �!EbضX���"OZ�b�fؠ��bk�!G\|s�"O�)ˆd�N,����	_��=�r"O�ڧbS�u���ӧ� i�����"O���DX��v,b�����Q"OP!� J�,���d��{�����"O�H1kԢJ���V�U�A~ �F"O|A�&��:	7�ap��:S}v`H"OB���
+H���GkYml&4�A"O�p���+ �b��A� Y�(ʵ"O�=���L !t�)9a��~��B"O@�J �	4z��E(׊I�q|%�A"O����A3E9���q����|�"O��l½5�D蛂��Q\$�W"OL�
P�J0`'vġ���Ei�%��"O���J]$�|��s.D�TFi�"OL鸂��t��}�oZ�^q:u�w"O�q���C��{mN8JY�ye"Ov�"�6p�<��&��L�C"OB���F�)#_�,�t�T����"O��	?pLd��d��C���#"O�}��f�
5Zn�� $��=�@4"O����䁬.aN���T�i�*	�"OD43AkM�mzdТ�NH��: {�"O�Xx�ƕm�D([�,�
�M��"Oa��lْp��l�@ܜ
��1�"O9��?|b9��( �n�r%�C"Ol�*�&!_�h�"A����(�"O��:�o�3*����<����w"O<�C&oL���Xj��U1Z8�D"O�Ai7�R�EDD��e@!}~�#C"OT��d�O'XҤ`s�ȑ6
\�Лs"O��A���V�|��w4T�	"O�:$K�5w�
�(f�V�GU0�Aa"O���4�� '�JC�Q���	O�O�����K�o]d��((`�aI�̸'���)Ƨз+��}X��ϔ����'�<tr�^<Zа��gn	��m�'o�\凘�#�����2	�T�(�'�(ۆ+w��iqv˄2�,�j
�'�y��#CpВ�H��ɹt)��'kZ��VM�4@�xeeQ�&<�@�'4��Y��{�P��m��| ��' c�犕O��bo�7��1��� �<�o3X,��t%�:����f"O��Kwf@�
�&�5*ǽ8�����"O��	�OGc
��-����"O�ȧ�A0v��$�$��b��RG"O@e��̿/P�)�"
�2�"O��ED�1%�
|�Q��m�L�"O�`iR$�2�昡�#S=58�=�D"OXtY���!��x�Ƙ"�iQ�"OР�C��C�Bnɜ]6�h"O(����*	q�b5�	Ȋ�y��? ��a���ܜu�
e8�����y"� �̝�nE��l���y��?�����'�A'�C�բ�y�N�w�T;�  5�$P����.�y2C k�܅�R�/A����"�#�y���,v����+=W�!s�޻�y�'EpD\`���=� &c��y��:G5^͒�횈|��z�h���yrB�<99���JFx�D8{� ֍�y��9S4y�B��pJ8�b�f�=�y2�I s��zub�s�8�G
&�y�`Yux9��B)e��X�b��y�m�qiL�����cK$�J�Y��yB@-���FDX�^����'ޞ�y�C�s#�mᢗ�
2�1�D��y���qK�c��Z/�>U�	ܭ�y�9z�!𗎍�#І��r%��yb�N�M��@���_$n��1c�OV�y�ʏ�Z^ޜC �.q�ְ��I���y�c�2g =�� ��7�0���y���>�N��&�5�������y2�8E����E�(;"��Rg��yB��:��(Bu`�Q�
)�%�y�d �:%�w�V.?�-x�ݻ�y2"�ΰ�w�bp��ˇ$ٲ�yR�Y�{���6 �Z2V�"���#�y��N�AS8A2v#�$UeT,Kn��yf�y������J�2	Wm]?�y��Heך-�o�6kz�\ �Ϗ��y�jۜ�8E�/�n`�0���y�*��_�$�b�@M:Je1eJ7�y�P!'4�ٔ
޺x�-��Ξ��y".�'�v���.��|��K�I�yRI����=�&�Uy�f$�uї�y�k�1�P��UH�
��!�;�y2BV\�^���V*:��`�)���xb^m����R����U&,!�-_�bȩ�!�<�>�Xs���!��}��잤Q�ڱ5j�wu!�D_nZe#W���+~�<��IX�b!�da{�t�V�Ƥv�Q�j�#~>!��K�@�=+�G� }`��p��;O!��Sh�i@��L�sA�Px��_��!�?,�||HզZl$���a��$�!�$J��bY"��R괵jU�ʼ!�ӧc�#�K؎@�֡!c !�D���D�!aJ0K�Fə��M�k�!�Dݬf��,y���G�t���մD�!�D��_�N���)C�
iwN�B�!���LQ�!� A��e�oQ7#�!���v�c��ϱ1��`�����!�$�(ƪ��a���.���L4n!���-r�p��E�n���) �A?r�!��2rH�Q���_�x��d�Ņw�!�� p\� � nǞq�D�V�<m��Q"O��y�&�3_O��k�Iǯ^�� 3"O�ETgW(.���3�Ƨg[̴�2O�����Fh�!npX��0D���A�2E�tҿ-� L2S�8D� g�L;ib��#�đ�R��͐Wc$D���SN�(m�~؁��<'��}K�J#D�īW�!��<��NT(S��q �4D�LB$�&CF�е�P:bk��*�B6D���V�$t����j�5)�50��!D��z�훕?Zf(hbm ($8��>D���4��앋�F�*(��%���0D��1�Cf�9j@Eۦybt��"+D�\��k�-����Jx�� )-�C��.4������&+�0<`䃽(�C�$(��I���̏Q�,<`��&cz�C�I%M�l��a�Z6M�:�C��'B^C�&u����<#|6%S�@�AC,C�I�Fk��02��KJ����-RhC�	�-�Z��`-E�2C�%@� &1Y�C䉛y�ȻT��}��1��J���C�	�5`ݑ�+�t�jŃ��E"/u�C䉋"�X���_41�D�֮DG�C�ɓHׂ@����=�`��P�®C�ɧ_�T�!AĚ�<�J���J��B�I�P9R�:����rkX��ehP�-��B��b:�p8gFKX�uƀ�bl�B䉚%���Z#�ʏ0�2%J�hߴD3�B�I�I
�Q&	��}2��5F��V�.B��(��}rq� 0�ʼ�AG��D��B��0(�������T���ZV�O9E�C�ɘ79�4yQF '�F�z���+n��C�	�)�hj5AD>�θ��� �^��C�	�.�,8���'��\� -ݎ(�C�	H<�92G��Nٌtb�CV�LהC䉽Zc�0ʧ�R���Y'
:P6C�	'{A G�]�f$�X22)�+�@B䉚Y, ���P�L�>	�O�J6�C�ɠa�J]#%��&9�vp�gL�s��C����b*h8�Ԡ4S@�C�	�oإ�F�3HL�薡D��B�B�����C	�>�0�Vr�B��~��E�t$��VO�B�Ɋ0��J�,�)O�Qs&
��o��B��+#+v<I`T�"s�"`�8��C�ɐI��)����W~2e�1�щU��C�I�b ��A�/`(]�"只_�C�I�!��ظ�6����ە3oBB��pD�$�qB�g���)6a��QrB�I�0�&��k?M� ���s�TB�	�9n�񒅜�8L�Ѡ��ă#q�C�I�ϺYuL/o��ia��]��hC�	�d��5�&n��BAgm�22 C��==��*w*�'c�)�0���
'�B�	�P��bP�4���!�~�C�I����gkA�4�����ҪGj.C�=g"h���;;ڦ([gHŴjPB�ɤ��a��̌f��$�b�Q"O�)�qnK&�$<�D��;G �hK�"O�8b�2X�ʠ�� V�NQ�"O�p�$$Ai�h�Ey�䐑S"O��񩊛r< |����^g���
O𼀤턨T�L!"�@ROG|A���>�y"F5 <��@��ةARl�f]�y
� �-�HYC	hPBҧS�CF�!Q�"O�B�j�	t�I��;:���"O��E��v0L�1b���~\ɖ"OB]�r��qX�(c��?�y�"O�A*�KM7W洐F�P�,��[�"O�ő�M����H��K�*�B�"O6�p��wD(����T��� A"ORm��C(z��cM�]��ȋQ"O��c�H��Z��D�)}PFi�'"O<�5��u$ya*�
f�̱ �"OjD+��[�B��Ͳ)ħ3��� !"O\(��f	3�p�0�7>`�}��"Ob�pQ�I��8)�F�ŔA\�$sv"Ob	3��ޑ)0�y��r:��2"O� r5
�u]tT�U%կVz��%"O��
3�J*v=<E{v�1� ���"OjX��U	ņ�	�)�n���"O�=شF�2E`(��S�x�@�"O&�R�녥Tu�1(��ޝ2�A*$"O�9f#��*b� Jt�A�acD���"O�Y��ٸeg���P"�c� �Ye"O:�����=���*���"O�yڠHX� М!��BQ���5�G"O��q��A�=���V�4.8Z�j�"O�La�/A�v�2t��?#&���"O`����|���	:y�qF"Ou0�GE�5�(�#J\�$mBC"OBI	��RC�X1r�̽ѕ"O�����R,D��,n^��"O:5�b�ƙ8�I��-�
�@"O�@X�( "R��b�L�ƅy`"O�D�JG�yMlI����f�ڕBb"O���V�
l�r5K�]�X�"O��R
�)rG�����)1�"O�\qC_%,i(xË���̉�T"O�q����(Q]��XpHI=\�$Q�"O��S',E3h&��H���"<L�B�d&lOhP����d�uF�"!T�%��
O6MÎP?�����V"L1�`'CG�!�D	�\
�T��/kq�u��Mс��x��	8_U¥�& ������@� #C�	�r�L�#��]�!�f�@��A���'B�#=��&�Y?��݉D��wO�Px�&�V�<�RB��b, ɓ�g`���,Miܓ0@�z�	Q�S����
7�XA�o� �Px�茊ue~`i1N� ps�a1�B�h��J�d�2�n+2�� ꂇ1�m��I��O�i)�兆'���jD>&
�x@0"O�m+wO��:ڬ�1��ʜ3�dء��xB")�S�'s�i���pƪm�FnSEw���1���c� �a�R�YƋU!��>y��'�HH�Á^�(Չ≗"�8��	�'Q�x�B#�-Q"h���N�L4>y�2�9D�@�cg�	[r��I���@	L7,O�xGx��=[�Td��.�/>bJxI�k*�y���OMH%2Uiɍ)�@1+g����Q��b?���I�Ԑ\�&pF�Q�U�1D�|��`�V�P��f��t���:C�,�	��0=ђ��')ʶ��ՃQ�^?�@���OH<9�I��K�;�i�����4ቈM
!�DL��HR���8G�(���_ay�,'�4 ��ʹRLA;eh��Aq�Շȓ
b���)HNzH�͉Ba'�������G�h}ydkP0t`Z�R㊣~k!�� ��)a��W�N�P� 
�+6�A��$�J��� `��J�����[-`�02�<$�P ��w��J��.,���¥�
��yb@�RR�	{��Ia�ő$<װ<���A�*aBʕ�g�Fhh�b��!��/IF�$��wD�f 50��'ўb?�a�̚5	�=A�oͩ$�c�$D�k�/�r�<�2�JT�T0�u����<ٰJ�+P/P��$T K{�!��?c��$���+7qO���G�/�}p�P��'.6Б��t<<f�I�e�f}��',<̩�5V�.QY�+o}�C��^/oL:XGx���j�?-
b�]�"ܸî��H!é7O�������'bHӱdǓv:PYS�fRM���8�Ir8Ex��I�>v�ܹc�mÛ>o�p�I�7;�6�5z����3�)§Q���d�R:k�jE��� �ȓ�V��jŧQ�^�!쉃i#� �<�Q�H�l$���EO��X:��	-�"̩u�Ֆ<�!���L�FQ�֠C�;�,8̝�D&���T�PxG�?P�B4��#e���r�%X��p<�˄��'�����jN�	�渐` NJ�#�'kPaz�	�0<Nȅ��nX<<�Ji��'�j]J���()@�ع�鏱!<$`�'b�!���(h_����A��Z�;�'`�A�6FX�f�����ф���q�'�DٶIX�ޠ�p��9��@r�'vv�J�)W�b��*@���'�ʔ#C�A?�uh%�V�>�xx{�'�xC�!�?BY�[xM�xI�'6\)І��
��|��J�+q�NH��'Z6��1i��U�g�� F#X�2�'�|�w
��kOv�␥D�F�*���'��0ʖmF
!�l��5�����'q�9P�D84�z:0MN	1D&�x�'
=����>:� FF��f����'�L�I-"l�$��U���yp� �'zք����W}�Y��R}jQ8	�'�����@�/[B=k�A@�M~꠩�''<���� TڙS0��T�I�'��X�+��
��$"@KƩV�8\��'�1;��L�qO"̀��)F�T�
�'g��&�6i�4y
��ȑ?�PU0
�'���jb!K'S�j�:��\�"On 
4�ҟ?���r��
(�ԡ�6"Ox�0���>8P�%��]�f֖��"O`K'�ޜ;�(h���{�җ"O$+$dH�3�]�c
 �f�T!qR"OFd�V��>Vb�X���U�%r3"O���ृ�������V9���"OH���=b���QP� m����"O*$@�1 ۺ��L�)D��	r�"O��q)I,/z�L��k��`V�O`}��&���0>1���^�)0�A�7dB���J��1#*��	$R�a�4��$:���@�t8�tb�:�܅ȓ(<��ԃZd�m���v����?��.�:Tr�`釵3��&CY^�i����HkĈ6C��r�M_'u�!�d�	3y0��! ���@���-T͎�Dx��9�g}��
r;@|ˑ%\"IV�őщ���y�L�^-��Β E�z�I�⏲N��5� �>���̊}�q���HO e�\�+<��S�Ȋb/�z��'w� �2O\�`@T��@iWk�eGpc��$���a���w�R$7�O��@&k��'3ܙڒ-�>�L���	<�h�Ie��|Sbc�(/ݔ`�[w���'����"d@h�Q���&�=�ȓ\�8��ʛ�܊�Idj8+6ZL���i�RuSGB�04�B5+7��
J��yP5��t�F��y ��(� $�R3z۬$ ��=�y
� ��z�],A2�w�ԾeAV�)�(�)t����2$��xAF��d����Z�ߺ۴�d*Al�� ׅ�����9taz��B�tzf�k��ʝ9�B!2�Ü%M��p��Z�i�)�'�J�.��$�f���v�=lOZ����z�-��LFT ����d��2r`�6�ޑ���� �+&�D�+~qx�
ݘ�D��gϑ��@�`-X�u.^ݢ
�'��� X�:�X�3�*��bc`��#��c�Խ��Dy��<��� 2OYⓌ4{�N�
_�e�G�B5@�=�˄�e!��PY�d���\7�x�)�X8Y1��K�z������H��\1 �R�Q]�|�ǮX�߸'	^4���Mȉ	����(0��0"����W��� ��R�x~����$���*�o�)�4��!�F�Hc�/۩�p=1�W7{��9[6Q�2���/[w��,��ƭP�]���óf�6i�T��nB�o����M�~Ć)I0�����:� J>!��6G�"�q��Q,���0Č��
�ysl�%.�R�+��G�&���7D�*�aJ~:�0�t���Y�8L�˙��8h�"Oʘe�6���L�:�,4q�o��aP>eð +}��sA�C#����O���+��'����CάS�
����O"}�(���:���m�&K�x�
��8s0t+��'1��|pB[�fL�S�C6S"||*c*Ȇ&v�zj�0�&`��ζQ��e��ˆ���'[p��EvĘ����:�Ny����`SA
��0�t��Pm��&~�Ū��P�]́��'VQ�� �wS�̍�S��0��u�`�;��4*�/�#ZE�@ZA��O�)������EF�E`��D��y�N8����fC�93 L�ڴrr�c�!MDr$�#�IaV���~H>a�
��F�8I�AB�����"(EK؞�AS�??I�e��.t��"��@X�ɑr&L�B�O���T��P�r!A({r�"PG.pf���6�4��:��#<�Ӷ+��@���ޏDԐ�C@,:*=K���!2�!�D�y��슖��?7'��#���G��DyH�{����?�]�Vq�9Z�6:&JETa�2�:B䉧c�z�@~�|I4GW9
�����	t�i�r�.ʧ?LZ\h�e���ւ!1
��e,e��qhU.a\"�Q�B� ��t"�d�(m̱r�R�\�,�2��ͦH�y��\k����e\�1�y3E(��'��m@n.ʓt�����3�a%��/%��aP7Nn>-K1��(q��QdC[2f��=���.D�(s�oöeN��G�<$��1�o��eȆ�I;Z����� 26' �AƤ?��c�؜9�(�!�M-*d����r�<�&`I���1ɗb]�i<VD���Ĥi��9��]�}+�9���E�}-@\�����~ybjN� `Y�D�W�R�2���<�0?AP&Rp�(h�-�^�jw��1hw��'��]�"�U/��>�ÉH)�te1�%��)��b�	�o�'EH�H�k/@H��~2Ԭ�S% ��e�U�""�!��Ko�<�q�.1M� z7MB���ˎh�<y�/��_$T�MS�mĸ�CABh<Y�(��6Խ����{�2-Lקp��|�pc=�IO�Ol���㗯��ڱ�ޏ/"�Z�"O�\1�@�$p�L1W�N�_'8���"O.����#iN�,��X.4�2"O�)y0�q*Fܓ��0I\=�0"O�`�T�*":�+&'Г%�1	�"O<��a V6y��=&�z F���"O:���M�:n�~a����oԔ�"O�$���L"�a.��iI\�ۇ"O�@ 2*�7�p�@��`��*P"O�u��k�;��5P���E����"O�Q�3cW�Zu���Ӕ|�U�D"O(�x�!�	Hz�*0��3���r"O0�K5
Cz <�
��UZ�.%��"OFD�P��*%>6d�p�	O�p j"OD�C��҄6���KЁ�HW,�e"O�YЖ
X�*�֡��/�3~Լ��"O�Uy�� �z��N�<?Q��G"Op���X��\{�K��e7���"O A�%�D $ ��+�1��#D"O�d5�*.U����i���h���"O05�É@<�����~���"O� �9�thE7zVH�hv���J4R9`�"O�Da��':��Y�@�}-���"O�x��Y�$mb�	V#J�@��x�"O$y� �r�8��U�EEɢ"OV�c�%�sΜ)*� ,�fɨ�"O�P��$��Ft� ��z�X��"O��3�ѵ)~�+.�p(�-$!�DP8+ڱ�@��A�X���^
i_!�2 4b���.�PdP13f��t8!�DA%+3Nqb��o�`�����. !��2S�:@���r0��_�}#!�U�",��2�%FC�|0Ó�O!��Y� ��B4�}�
��C"�%g!�$ů	T� 4,ĉh@jq���o!�D/U���pq��:2�I"Ѯ̏D�!�fsDq�A�-aIC��!�^" ����,H;*�HU���hy!�G�D��5#�a���M��O+$�!�d�)R�}��'���.�P�Z�N�!�WBnl�Ϙb��uR��&!��,}"���[�	��"��h]!�$���¨k�!�X9{���8{=!��P��T�2I��U3�J�l!���8�ےj��\#|!C�$T�!�$P�M�`Չ�ݩ0az|��R=�!�D�5~|�ub�3/Kr�ib�>�!���sVypUm
�!]�1j�EȪc�!���,?#PR�W��j��Ī]q!��7aHz�!6�&?C�Q+B�V�=�!�dWJ�z#�a!B�J� 5�!�؉z�ڀ�aC��.&�*@C�0a�!�	�*��-k0$�y2�]PE�P�b!��H�:���[��#&Ze�`�Y?#O!���<F��@���*ΠKv��5Q�!�dC�a�x�16>$�Qҍ�|!�D�'S�!`@��A�R��mR�s�!���)F�H��MI�H����lF!�ą$n��aE&\�H��+%,�4�!򤌡y#�-`�eM�I�~�)R�	�!��S~�nl3���y�F򥌁"s�!�L�2����8a�t�7k�!��R!���W��zh�|1&��Tm!��۞&��HӰ�ݧ&�\��j�O�!�D^�g�(ђݱ��آ�4[�!�d28�8!�D,z�i0�CJN�!�D%v �2��$d�0� �tu!�@�r�#]0>�"*ӯ�:�ra"O���2�ÙKx��ȣ�g�P ��"Oj�����alx@�� �Gh�"O�]��"ʒw������N��%"O���D�qp}�&�7�h�"O@�q��=�v�z���e�@y�"O&�st�I'�Yc�A��r��6"OJP�ʇ�gbjA'� c�i�"O��Ǉ��w������->Ʈ��"OR��h�DM$`�Q�S�JΞuB�"O��c�'�'R�ܑ�,ۉF���2"O���$��1:ž�h�aݶ6�
Pc"OڰA+��"wƩ�d/�+8�lT�U"O�l��#��1��_�s=�"Op��e,�%k�bـR�Q0r�
��e*OVL�]��p���<]�����'����$n[�G�6 Ѕi>]�bl{�'%2噱.�����P�_
����� RPP&�֋���)@΅(�^e��"O1�#��#��u�d`X�'�����"O�r��. �n=Qa*�(�8H�"OY�,)u;��r��Aft��"OR@����k� �'ƌ\�e��"O�t'NY?��$���E���"O��`@��|a���P6��)F"O8�[ѯ&
r�8ւ�5*� �"OD�yQ�N� ;rثGoN�hw��I&"ON͂v�X�de��Qu�Ĝ%}):�"O���È{�8�9��o�2t"O��G��z1.��#ŉ�ϲ�	�'R�8�Sf��'�)b`�&�0��'��GM��Z����~��0s�'nB�H$cėX�!rFO�?u�.��	�'A����Q�_�y��o<Dq�'�*p�ᗌ}D����i��D{�'��`!6=D<��f_�o�(9a�'��q��B��&}pqA�E��`-4I��'I��c��i������v�(�'UL�{g/�-�T��� �����'�6�A1�Tڌ�`H@7$v���'y�)���=�<��	�&�i��'��5SM �3K�Y�Jj��\��'T�1k(���ђ�e:��T1
�'��D�L[��B�`A�	�R=�	�'`:�kE�@��1�Ѳy4� 	�'�x�k��4ЌĠ��� 	�q	�'�d����\�5(�c�>%��R�'�^8�S���Nh�������'�`E�"�J�sT����Y����'�����֝e�dر�+DIt6D��'KP�)a�J�oP�H`�Ͱs@���'��sC˹`*�p:WiQ�k`eH	�'���1��єh2�u����W�4��'J��
�m��+;FH;��F�A�9��'^��a�G�����0K�|1P�'o>=�����p��5�P�85�Y��'�HU��'N�]�B��%N�=(Rb�
�'f2���eݬ<0�	�#��+����'��}�p��Dz�s�j1.��D��'��a�B%hR(��D#6a���'��M#D��2s�B���
�(��@�	�'�^���a��H�̑�c)��|�lc�'@8x�ъ[��a��!�RP)�'CФH�m�;w�cC�Е�|p�'rt�.Z�_����"��?�$��'ϸIA�A�)lȜ�r/ؙ����'H��a��
"~��E$�R��
�'1��	�
+"�40��H��v]�	�'��tSE4=����B�83�N�{	�'�(��$�� 	@6� )�'��y b��-<������lu�'��԰w��[6��`@�<w6��'��Cwg�S}�	���11t$�x�'���S�=9����Ue�������'Z�i�7�L�|"���T��9!��L��'�pp�G�>jJQ�ꎵ7ր��'Z�8pQ�X�O%sC
6 Z-��'���yu���9(����5 j��#�'b�݊��;��	� ͔OmPyC�'k��z�+�]_�1�AE�#V�����'��0s&K�V�R$����+FC��q�'oLܩf@�&c�@Յޒ2V6�9��� �X���4U��(��,S�vX܀��"O�Q�0%�N��u���#]4��s�"O6�U��b�<%�s*ۂG#�l�"O"��
�v�&4�ɘe�>I�&"OlM۰�Z�O��=hr�Y�@�xd�4"OP T��	{� ��D:T�|Tq�"OJt��ܛK�&mC��!�R��"O��S�DD�x���r!����h#"O�	�똭<�!��#��f�ft�&"O��#)L�"	� y�B��'Nܹ"O>89UME�}�(ua$�ű��P�"Ol�����((��v�pq4"Ox-�f��-����C��S��;�"OD��h�61b��׀�M�\TYV"O�p�SB¦;nL�U�� #����""O�	;�
�9y�vԹs.Q$y�0A��"O�ɆkU	dހ�b��~��43"O� V��,L�������k�"O�d��j$гJF�7���e"O��Q���	�<�1)�$#�x�)�"O�H��JΨ-��؊V�
�1~�ŻD"O ��V*w����֫�S\�ۀ"O���gZ)x�%��;)L(���"O�����AJ,3Tc԰/0���"O.5+
Q$~
(@��$�j���+�"OXdyWGђ!�Б+�	��B�
	�#"OjEs��k�z̨�&c�,���"O��(�?���k#M�{��z4"O�1RW��ՐэK�
� ec "O|�U�ExVXJ&,TC}��b�"O��Y�ɚ��\�s�K�_=�S"O�� �m�yA���d��*���"O�"��8E�9���Pi�L��7"O��ٰd-9b�X�� X�,�&"O: �G�-_ڭ����"�p�"OR��g��P��4�&�\�NF�*P"O&Kr�N_�JLS�؂>nnM
�"O I� ���x1��)\8XX
���"O0��	�B��Y �)�7o� �4"O�=��&� ���h��'Y�̳�"O�%�g�n�`�y��_d��p"O:����ϣ}18�i�a�;32���"O���e%E�
�p���"��<
�Z�"O�5������Qx�kӒ&��A�"O��h "s|$�Ӗ)��7��Y`"O
�i�@�UQ�l:�� t�X"O��Â�UA (�E0����G"O�����1tR�)
�̈́e� ��"O�%)&l͍~"(Sp����1a"O }(�1 �����C�2��}�3"O\-�ꅗ#�
M�bbJ����"O8HQ/�H"4�r���8b�y#�"O��CE��]~�{G�:Up;"O�"R�G����g��gOz���"O�!�!�S
д�WЄF*H�zG"O$���D�꺜+�τ�W�F\Q3"O���%I�j�~�۰�͋Kؐ��*O��I!��<=�XJ4���[]!��'���t�ɬ[� i࣢�)8a$3�'�.=a��ٚZ�:�CdaG	3(u �'"������	�xȓG��7[&*�'�J)K��?m�$���$%�����'�l�[Vh,���٢m�>M�d�'sVpAo��S�F�C����|�
P���� v��Ӈ�г���Y��X	U"O\�Y��@{����E�N?�P�0�"O� �$�D�Va�Q@�3�6�a�"O�����~!+����-	z�R"O�(�6�^4P6�	w#�0���"O�][s��
c ��w�j�2
O����O%i� �;��4i��P6�hO
��C��0FAhP�'8L�u0��O�̂2�*l�y@�'M�7�V��!�>��
Bn�O�����n�
��E�ē(m@�mY7^�d���@�S�OQ�{c��@�c�A��fJ�!�޴un.q����iߜ|������Z� �� ����+�����b�8�N):CnȆ(�|���D��d�`�D�Y�.����b
��y�4���%PrtL��x��K��O�����f�RO��Bu�.d���tY�|�5GUj�S�OL��A�އg7xy��B�t*�\�ܴ>I@����I��j�ne�0]����S���6���"�5�D�P�΋5��9� �5ꀕp��Dͺ`$��ᓌ < ���"/P�	چ+2�� B�C�n.$��� m�p�|�~:e�I���������]	e��t?��N?��㞢}:Ai�z��=�$�8J�x�U �'��X���<�)��x��4�gN!w`\¥KX��|��/���0|B�c��d���A�U ���1�h\]�ws)�J|J`���.�Px��V�B����C�X��-h�$���`�)�:(N�*�(
���E�2�ʇsw��GPjyH����J>s�J�A��e�v(��ɹBY�v)?	�O�?���	&aW�ۤ�Lb3�EHG,���O���S�v���ґ�J,<T|�Sk2�zc���Ln�S�S1xS�蠀�޺w1rU�3A�
@�O`�G"�)��ON&���`J�rŹ$
�^��R�x����R!(�z�L ;��{WL�_A�V
D%[N�c��i�hR��y_~��i�"� ���$qH��ʇ���T_�'iDR�*��䛂�˭@\M��'w�	:�ɍ�?Txe���/G��
�'6�(G 
	m����A�B��!�	�'4eJ"��UZ�Q��2��x	�'W�sA��!* �PI}4` �'|�E�h��Fw��ѭʺnr�\3�'�ʄ�0��Id�}�UmX-X�����'Mr��c@F>K�<��FH9g\���'����lD�@��8�,V�\w�5�'��D��wΨ�b���P��D��'�0�S�!\�7pT� qD
�C����'��x;�aa� ��!��)�=�	�'���kQEõ
d�qP�+(k��C�'l�SK֡T�B������ �i��'K�����1B�TA'+��9@���'&���C!zU)��	U�q%,��0h9D��q�>�����k�z�a;D��C��`�~ C)�����I=D���eđ?�`�#�ӶcT�mkek-D�tr�Ŋ�Y��Mb��n`�H��*D��㴨ȜC����� z�h0���(D�����!JL�m(EkA�/Cm(�D%D��&j�T"�#Վ0��!D�`J5L�8biy��̷s�2� �!D��0��J473��K�
?�,J��?D���7K0| F���E�86j����>D����+��D��RFJ6u����A=D��@�GS�n�"�ۂG�!	|�\���'D�@�J&C��k��Þp�����+D��Z
����a��BC��0���-D��
e���P��H��u*<sW�,D�XӁH�B�H�(X��	*D�h �·F@�l���e� ���)D�� �T��f�O�εs�*��u��'"O������ ܐ�p ơ;
d鹁"O�Qծ�^K�4ZU���=P&%`t"O�i�k�4����W�\:0q"O�����3-A��x�B��_)� ��"O8�����F#���LZ�)� 1�3"Oݹ��K=��S�k\sX�"O
 �E��!:��
�)���� "O.���IÙ]���  ���ɲ"O��ٔ��t�f�ş[�4	�B"O��j0�
G�$��Ԫ�<�豢�"Oh���-:@@*@k�E�"O�	�E��a��&�1s��y�"OH�V�A
b�Ł0�RZ8��g"O|�%CK�%A�M��-��o�����"O4 ��F�vfh��-�*W�X���"O�e8a
�kG��I�g��͛�"O�B$��<uQ���0h��w�B��T"O����䈐 5B�5W��=;u"Ol��q	`w(XP��k�Ĩ�"O"\s��������U����"O�	��M���je&��,y@�P�"O>�0�0z�뱂�� T�("O����Ȓ M�i�R�D]�~y�"O����!C�>�����9�t��""O`��c\0C��	�DU� U�@"O���S���?�L�%�$� ��"O���.��M��0�ď�'c>���"O��/�6�"U��	la�<��"O�H��Om@���mJCN� 8'"OJ؀w*��"H�|���ΧC:j0V"O��s�h�Ѕ��	.͊�"O��ss
x�(QI��[����q'"O*T���
8���i5˰y�J�"O��0D[x5��I@�O�?
F�{�"O���DnH�*�(���/@12׆���"O���A�y��8� Z$ �6�[�j1T�X��L�`���_|�p���"OִH�d�W��	I�A��s���Ig"O�%� KX�CD1�r����4�0"Ol�y���k�N�Da��}��[�"O�`�!-�Y�0��
.�,��a"O��#Av̋���m/����"O��Y�y�-
��I�2~qP�"O~�I�#��O�Eh�)ɣRj� �"O ���eT��R���'�Bvz��@"O��� ��8hP��gY�j�Z�"O�4����:e��2��3_�(W"O���!�T ~������X}r��6"O�(���:(�H�
f1E�9��"O�8�6 (�^��4�x	$"O�4����S*�����( (��"O�Q�Ô�8�@u�Wk��d �){"O���Ђ�>Ej'+�=l�
|�"OJ��BGY�H� �B$��c��d9�"O@ua�$����|h�,�0���q2O�`z��F+?�h��f�W�z�tՅ�ch���&�1b���j0(H�I*����mA���ɖ6.N�eғ��kˢ���)�N��\=�z(J�fфJڦU�ȓ��!!0�M:�N�� ��)?}4!�ȓTJ:Ű ��\���3��R1���r"�h�K
�G.8Lp�B�7�
ф�{X��;�CB��f  �P�^#v��S�? h�� -Z/7X�Z �-Z�9�"O���E�[$CXD:�U�I�"O�� ֋�2�,�k��2}�P�j�"O�1���`��l�W�M
:�6��"O:��ņ_C���、�*�$���"O��)���!�R]��O$��!s�"O�-PNP�L;�M�o���A"O��ڗK����j�.�%͖�"'"O��J��ŀo�|x�D(Y�6Z�IV"O�<*�$:p\J�o�|��C�;D���J�6/��٘E$�#y �㐬9D�|x��hF��yQ�X�R����8D�d�$�Q�2H�yÓ�ܻS�$	�UO)D�|�EӾ���7�:l2�`2�;D�| !lD"H�%OŒ�۴��<"HB�	+%�^��C���j8�A"2L�N|B� A�h������=;ר2|rzB��1q���D�[
ql-Z� �ZB�I�?�����ƕw2�=ӦO�"B�	2]��XKRK!���$�E�l+�C�I�w�
)ĥ�:A��A(c��-]�VB�I/F��B�P� YJ�����x�HB�I*�tőA�

&�ű�AY*Q~~C�ɏoҺiB!��{Y���5��6N�,C�	���P�$O��p������?F�B�IU~�  ��h�BE2#�Ĳ^r�B�I�X�^D0�ԏm��Azp�Æ�\B䉃Z��y�Մ�)6*�e	iL*=�ZB�ɬ8�f��х��51��k�H�BB��0.\8���P��h;'�nC�&K�(��JE�2�����ܭ�C�	�:���S랞1�u2�b�
��B��E�J���-ѻ1���'2�B䉵.����/>=�i��M1rB䉤88��&cR�M}��-ҷ;�dB�	�������X�$��T��b
6PB�(7�8s�ʧP3���+G�Rl<B��)Q��+�� �:Qg��.�HB�	<+%��ф�ʦ��Q�:x	^C����MS2�<)����BnV�{�B�ɚ!]Xг��º��sG�?'��l�鉊?��R�#��y6�	;�V�X��B�	NXX��TF��k5��� )�<;�^B�	�Af������)����î��x�FB�	�$�0Ⳃ���a� ����B�	�%�x��W#�5_��u�Rdİ(U�B��b�#5��>k���cd*�g\�B�ɘ�jP�u��g3�����¢,�C䉑��( �(�'
[�u���w�;D�L�f�yl����<5R�
$D��;�&=^^�8&�֤��*�"/D�����ؾ@.l�H��T�8�8ȋ��,D�H�a��q�b�`fH*h���d�<D�,9�	Na.Y�.ǚB�$��;D�PѶ�.��b��n����9D���7-�(�`%��ƀ-���[�-D��DA�5.(2У�T��� v�*D���#���=���#F��g�<��(D���C5z���B�%��%�E%D�����N�d�x�k��^>��
 h#D��Z%�fl��WI��ߞ�4�!D��ڔ��:l��ib�q;0���� D��R�I+'��A���O7:':yg�>D��Ȃ	��Rx��-oh���\�!�� �\JF|���Ն]�Rj�"O��d�ce"}(w�M�fG ]��"O:|���
���u)(}1�"ONLA���ƕ���1t��(`P"O�%����(���QSĐ�l�h�"Oڵ�bn��Y�I>�$x��"O�)bwMC/Zr��"��.i�h��"Oڥ���4q�e9�(Ծ^z�Ġw"O:���)���xIe�S��<]�G"O@�y�A?~�X��aoêb#�:"O����F̹GE��#��'H7H)a`"OL]I�A�j=p,�%:"�$+"O���䅐��U��mI�>���$"O 虇C�?Ra(�#o !}"���"O�5���#��qB�7^ �L#�"O,A���+%��K	��to���$"O���w�H:�^���*� Mr�I�""O�%��g��=N�ɐC���l)"OԀI�D.C����!�%YׂU3B"O>Yb����X�(B�a��2����4"O�d!�	D�kKZ�9uBѝL7^�#&"O�)�/�3�*���Y�
� �"O���㆝#R��9�����~����'��23���p��ʄ�oYbi��'�fpA��+a��p.��l?d@Y
�'i�p���M��t$Z>#0��'f�:d�g��y��b��[�'#l�	\�F:�i��KX�9\2��
�'�ܙ�A�M�4�|��8*W��"
�'@��@�=�\Dkt��� ��<�
�'��|h����y�=�����Xh�#
�'��@��:if��ȝ>	�B�	�'5��آ��(B��0��j�dX��'����r)¢�Ec�!�Kb\d;	�'uX�
���1̘3��كX����'����/�3dpjSG�yD��w,rӺ�*cc�
'9�������I�\X\w�B�'؛��ǒ*fx`W���9Z�`���/+|`8S$�f�� ������:�8	�5_���pE�I$�5a2X�w�\��̚7w:�%e��A�% ��Ǻ{��0Xڍ"�ԊO�z�I߀o?�II��ݨ�?-�M;r�i�V���	\�I�I\<9�\tt�ytj��[���<)�ph��)h�o���k�&Ac��ǆj��O��!\��(O 聐��ߺk�4�:XTA#W`0e�a!S��1�'j�'zrX�a�'���'a��bҁ�0� sr��Yߖ1bP�B���
C�?!V)��ȕ�<#��)���(O��2Vœ/N��:Wn��U�6z�hJ�x"(��� �*lD����O�~�N��t�<<�|��a��9yx6���O
�	� �%Em4l�2���x��<+1 >��	ϟ��	H�S�ӑa�������V|e��D�m���I�Ͽ�ŀ,_*��'��r4xa�J. �26M�����'�\��+b���O��'e��!��Q�{'��c���M�F3�?9���?y��W�z@��RF��Jp4
P���3ybM(�����ugN�^՜�i�/�J�T�0&�����'jh=��YY����@�$,>��*�Ĝ�� �� �ם8��]�s��4�Ke���^e��yR˒/�?�F�i �\��SY셺�뗦}!�Yt`-�Ĩ:�$�O>˓2He2��ڕBZ&QYu���$,���hO���ܴ��$��<y����$��Xr�܊��А(��|o�ݟ��Iԟ擼u�D�����(�	Ԧ�Wa�2����o��.���ˉ:Lq�D��*�����#i\�}��jć���i�����w�4���f��X�a'��6,���L�5shz����)v��!�'���D{g��LѼ�ElY)b�	GX�� Jς�� ���&"�f(o�"��$�H���DGF�HA�DV:��ύ�H��������?�3��4c2���10��Q�d�O&�nڸ�M{J~��'�޴9��ղR`�v�t��͚.(�L5�s�'rr��DL҆���'�"�'�d�]����I��AP�-R	��(C���e�*N	�6B�L��t�slT�m�6@b�^�-��?�(^�v
�T⦯'�����GJ_���{w7n�z���̊=z̬�P��YQk�\x����P!p`�
AO4E3�H�@��DIӆa��X��'47m V�Işt�IV�,�ʔG�D2L�!A��99F��D�R�<$��U�
U#�&B�Ȉ��+�"#�ƚ|�+u����<�p�V|����� |17�@40������&;, i����(�	��؀Peџ������#5hI���L�M��I@���%GX8hRiR!t9b���-8s)�uH���$�&J1��I�'Ɠvf-�%F&e'0 0��� Y���.˃i��o�7�qi��ɗw�.���֦�j�΅�U��j'���?C~ms�OF�|���?I������'=q����#��xu�E�<Pj��3O"Ћ���M�tA�AH��B���0� ��M��ii�'9�'W�'��X T  �   -   Ĵ���	���)*thŖ>"�����@}"�ײK*<ac�ʄ��	ڤ´�x�c��7�	�M�������d����F̘w�` �dk�k�a�(�ئ�Q3�V�uGC�6A�� K4��(����O�I�*ͼG��9B�E5�hX����� �-O��Å��|BH��OP���&ļOa��hUgK�!�
yb% \(3� -���)��<O���������:*� �J�.�2f�LV �bǏǺ[��SO/�� �%[�(�Ĥ1)O,���9��a��/���>%r�KW$	(��g撔)hŹR�b��+W,	8��^������>	t8�:������P"Ũɪ�]*P��
Q	�1�ɔrq�]�1Q�����'�P`�"-KM}*V����R� %����s?��L�0��~.E�ѯʧ�?%�'����DQ���9O�Ac@�H�`�Ah�D��x�G�pf�عu�xB�K3g��0I>)d �	e�,D)��s��@-�>Y���yT��.���#��O�,�PğK\�'����6�ݟ��D�r��-C ���D�DPv���R;_��O�Ҡ&?_
���<��h�#2�����{P2��n]�TU��h����Fh�$��U,���7��T��C�f ����D�'Y5hP��-�q*z��u��,��������wމ'��	P�I*�O����䌀&�8��bܺxD�aD��
'
�Sx��$�7&u�+O^��I�4������d���@���/FZ8c`�� 5QN�����C7CM	A�X�'�(�D"�8 "�|�c@�Sz��6fx� �Ҵ��X݄d�U�FQ}��6}��n�	�[_�$�;~��82W�Sj���L��?�B����vl��9ŧH<G��ě�x4���<F��	o����1��P���1\�+7I/��dՋ��0ِ�|�E���TH<Q��Pv� ��f�=y]f�0��([|a�/�J�Ʌ+�>�� 1OD�Hu�ϙaf�����%��H�tiR�p�DC�I�f�~ �  ���T�aJP�?�Ʌ�e�5	j��,oY�c�P�h�D1��}��4��N�8N	��B�H�nh��m� �N�p>l8m��=z�=��Upp� r�0Rj�� ���"�r��x���wnY3�$��e�ydVA�ȓ�0�����o���Y���
%+�=��A%`�����y� �Q%�(���ȓ(����uƐO�Bd�Q�Q?d�ؤ���N�C�Mi&9I���;A�����6�黳A�&X��EC�B�|�����8#䉈u��j ��z�h
�Z�ұ��^���
#��;S�`T�m[�4|l@�ȓ��� ��;oY�3�K _�VQ��B�N��內!(��El�:Lt�$�ȓs�y(&b�`ƽ��Zt�R��ȓ2�,Y����w��pQ�DL欄ȓGi��Z�(ϒo#����o�$-&ńȓob�b�`U�W��4R��T<�Ņ�~:hP"�U�,5��#^U�`!�ȓ>��x1�̛<�4`T�ԱQ���ȓ�,Ț��-����#���$���.�]�`�A	y�Tă�oG/oJ|��2�4����Be�@UkT�)S)��Q�@��a�NCf�EkD���a�*)��a��4����ZV|�w��
���k�9�F��"NP)��F K�<��ȓZ!<�#v'_gh���$4Fࢄ�ȓLքDj��?S,r�x���wX�8����9�Gk�P����O�N� �ȓ7�$ R�F;4}�%Y�<��k�1����UXx0�N̑58��ȓH	,e�V\>9>P�ֆ�Y#����:�z��P�u�����݆Q
V��i������u�����
����S�? � "�Gʔ8:�Ӥ�U-a,D	A"Oq��Q�N'T�SuH�x����"O�њ�2R�r���iځa���R"O����H/i�Q #�?��ef"OD������O��+vᜟ1��8j�"OH��dێs���E�Z�����"O� *W�U�Ht� &؞e�n�w"O$1����M��!����4g�J#�'XB/��Yl��o*&f\�`eVK�d0jǌKu5�B��?ѓ�K �?����?�Aځ��H�T*GO5�xk�G�<g�(��4�Q�0�̛�lI�r�:UI�rJ�EyR !TZH�C,F�ʈ;��Ä��J�
��=�R�@`�K�e������#/�H1��ϛ2@�'�L1B��?�$�O�����#LƘ�����"Q�*��O���OV��?e��	�<��*�%�.Eؙ$gZ��?����^�'��� iW< !�@_�k�0=ӂ�ׁJ0m�f�lӎ��B����eZ�M����?����z�ふ�M�pc][�֥�ׇ�1Y�z��C"-'��'l�:&(["zE�3e b�Tm�$�d�I�6BI��啱ITA�F#�;_q������W�8����0^gx$Se��<�����Ƀ�bZ��gFǶW�*�0�55�	2���2��٠l/}R���?ɖ�i�N�������G(4$<(hwẽE�b�1��D�O���$�~�,�{a���0
�XȴN�xY�'�<���O��@̦9�ܴ��0�*��wI�;uV�s��^6Un��ҫs��4�?�M�����=�?��?Q���u����4�<S!ML��4Z�약|��H�e.��1tΊ�Q��	Z���|�g�	��Ēvj�(Xd( [�*ع��[cǆ7P��0�FDL(V��Aj�0��:���Y��e;.��Q�V*��%�؁�ݴh��f�'��
1�����da�V�gDU�\d ��O*[�f���iEby��)���	3��/ȋ��E�'LPo��ӧ�c��IoZv�\�"���S}r��<��<kEC�E2(T#\c�p�`H�cY�$�O<��O��;�?I���?�Q�{�zQ�� �f��5h@F�4_J1(�I^:=bh�@�+S�/ e��cY�H�:Fy��$��!5��c�Li�TNC�[n�xIR�e �8�+�+z��|���A�@�YV��W�O��b�D�#R�9` ��R���AR8F���'�O��d�O�c��;��N�C�c�Üv�� �c&�	��HO��:�'ş�N���m��hX- ��s�I.�M�6�i��I]2�=�ش�?�ܴ~^~٠�eS>��D�%���o���7�'K�j[1^���'�e&/��%�6+�	#��{��!�ȭ+��<#��1Ʈ	�`R�rkQ�",uB���ٻ"��I��Ph�]k�l�=l�^ ��N�`���k��ŀU��/	:E�pqi��a}1Oxq��'��7�R{?Qs��h��/
+���N�q?��lQ���Zw�1��D��O9�=���p-���g�����:0��)*ੑ6V�h]�dK��"����/y�T˓`��ŀ��i��'��8p�ڠoZWc.����Z�<๱h o������?!�m�-����)B�y�`�C¥i��d"�����I��)��jD�X҅�G�_�'�� ��-۔W+^���V�q��5��"d� M9�`?lvM��~چ]���
��RT�6�d�+��}�<%&>�$>5pS��H'����PJ"�����'�� �I_��6֐*��㧄��VF�H�򯏅aў�S5�McT�iA�'�vy�� �n<�R�B�L\łQk�O���(�$<�:�P` @�?      Ĵ���	��Zt(��?�����@}"�ײK*<ac�ʄ��	ڤ´�xbjR�6�F��t�gf��P�\��h"R>D��@Ezad(uJ�ݦ�	�j��h��(��M/�N!����E�4X���s�����ҕ
l
7� U����''Q*x�R�}�$�"��:E��FU�$M�t�T��tf� CLD4�"�N�h@�}B�D�<�����#�8�jVy�Cۣ����(c������!dc�;6�B�bT�Z�%��I	��ǖMn剨�?Y�۸E�$���vχ*r��� ��:T�$��h2�UI�O��3�_�
!#P�X
8Z�������-����S	O?�xG��%��]���QC�B���+U^�`n�>s%�O��Kq'O���ē��?iG,ωInD���Θ���,ܭ�j�`�V� ��'���@�)ey���O�`��G]"�z}K@ܕ[R�P���^7�ㅛx��K�X�N`@O>�U��i�|�'�*�`'e�+�f�I&f�4t@M��]��5)CJ]�	�n�����k&�����n���ݤ*��Ya�dų$n������U��Y����_?�A>O��#`��?���S輸� CT�a �m�G�E����'�n���u}��v>�xq�Q.@���̽Z���IIxp��h͘"_f�)���c,L�e�DG�#8��)II�-pJjasg�G�\���l�$��fD�������?Q� �8��|�"@O=K�H��'��MP �(�PyeO݉k���&��X"�|���9�?��+B�0��'�X#�_�B�ҕ)BgG�$����<r����P��O���|��z��#���<� �P�Ņ�V���J$��O�%���v\VDr�+w� �\�~�O��$����%�<�BL:��(H��� �&�ɛF��py#�>�M��hy��(�.6x��HT*��D���Oi�}�L��}�-��ѦH��X��H��"O��K$�  �\ܓQL>#<1j6}�+%?��]�Va <��yUb�'��ܱp����'�������'k��Q�  �dC1H�����h�]�Q�ȓ&i�  @�?b�RVs���V-�68�8Ё!�'���'�R�w�M�	����	�C��ײh�S��C��
!�_  ��$%pG�ߴ%���º&nQ��
q�6 �
M�O@�ZcZ�c����O%�1K���2�@��%!zj0�gd�/0��́����^bN ��$�P   �  �  p"  K-  �7  &B  iH  �N  U  �_  *k  Ht  �z  р  �  U�  ��  ۙ  ��   `� u�	����Zv)C�'ll\�0BKz+�D:}"a�ئ�pgm�|"��f��Aj�
s�$��@�� S���e�J��"���x3��caJ H���������hW��:E�H:Mb켨�%O�r9fի��7<LU+�B��)q'��UײJ���N�yL��I�Oکˢ"S�D��
S��+o��M�;(�|@u�m��!�:G#Z�@t���M�Iɬ�?����?	��?�p@I�\�\8 U�TFպ��+�?	�����9�����O��C��O���O&��*�H�8�i��Ô)(�S@��O���O<���O�	�O�(��i&J(
�@�^�D:#I�,~B�8a�h�>��@��:4�l����%�V��0���d#����Ʈ�xD"����LxC�\���r�L�?)��) �z����y��V4i�
(�d�ϿL�<�Y֡W��?����?yԾi1��'���'��߼�An,>���F�ǫ	~��E��Ɵ�h�4vO�&�a��8l�՟�+�4e��X��i�e��$�+,&҅�E�_��t�ä�2"��z�,ғ/a@iiӂ�/Dn8�i��K��Ms��u'� 5'����vxhq�	7d��Qt�g!2�5I܄z�� b��l��?M��`�0H�G�,0�0������$�� H��n�r�,�a�ŀ�0� �4CIYU�� �.�?X ۴{���v�@�q���`D�8���@%�O��
�Y1��\~���ΦY�ڴN|�v���G�m��n�)Yκ��T��!�Z�ɝ�x*!b6aL�/k�i���^���y��$fk�6mP��jٴ�J↭C�B�Ma!�W�n�~�����>	�����zdN)�޴9�����YƵ@o�*݊����'"�z�ʂ�Zx
Q��*<�J�%�Q�,���'��~Ӛ�)�^���M;-���Bj�O��'@-Q�x��4N�&}�cVg�O"�+z�l���O��d��c��1��R27D�n�*q.8��8J�`�I�V���0��S���
%D6���ꦝ��h8F�i����-S_v���#�#&�ʰ���=��[��	+Z�:)��)��A@���&�Љ]D���O0��/�d�O\��<i��^��2�,�X�(LR@F^�5bP4���?�ScE��hK>�'E���O���d1�� ���	zk�Z�%L�J��[���5H
�M����O��.����lhs�� F(��NM�<-��'��p�@	k�r․m� e���>�S�n���fPUSx4A�(�8 ��<�'�d0!���"En���+Z�T۔���D��O!BD�p�ِ&��DZ�/�9e��H�O���t�'"7�d�Op��C�k�K�,phQ��1S]�'#��'R�P�8�|Z1��X��1���*��H3R�OW�'[�Iu�IoƟ�Cش���kJ��y�Cd�$
YP��A/�?����'���3#˰��某�	ݟx�'�|Xb� K�_� ��a�j)K0��bmxL[��G,(⵹C�����S�?���3I�/k�&}�磂�I�Tib,��Y�e���NM*(�A%�"��]���Zs�DFɉ uD���w�(t�J�L�L�p�̇�s%z����i�2˓d=����?���O�`�P;,���C�
G�dX����?�*O�D?�3}�%T{�:� ��%�t�sP��?��<�6�{�ȒO�I��˓�Fǚ;�wƹ� �#g<(�����<A���?���lu��O��D�O�}������5��S��KC!Н&�n�P��1L���P&��hx��A��6a�)!T'��@�~�@�ʀ�z*��:@��bب ���7���TD5�]d \b��A *6 �* -�&�o�۟�"�4A��`FxR͉�h�ʙ@���9�M��?�)O �D�O���qO�xr��ȁcWF���W�4bA�u�'��6�O�nZ�M�-�ֹ 3A���IşY����d1���ʑS�p}8�O�ٟ���8G����ğ��MA`$ZWke��Iɖ�V`kV%~�ˈ�JT���`Ė�43���J6pЛaj��$�R��`�2�'j$It��"j��Ƙ��O�;p�`�h��ۋ�:x�J>a��[ڟ��ɵ�Mk�W�U�lS������G�*h,Ox�b�
�O�O�9��5+[,=@d���,4T���)=�Iu�����}��x�'�P�� ���� �H�7oYզ1�	�M�aH,T͛��'��	�?����,7�)8;
 ��@F�`�t�BF���I�Kd��AEͅ3}��:ܴV�����D�U#� ��j�p�p��i�h�	�6��h��Ilk-zxV} ��C�3~M��,�����?l#�ܱ����"��)� ���c��O�0o� �ħ��OX���2C�#�F�a��)�|�rJ>1���䓱O��q���I�]��Q'5b��T��̟<��4!��ƕ|r��3F4��`R�T�bS���W��+��6��O~���O���'H�Q�p���Of�$�O�n��F��SCjTj�ʃ�#N����Q�ey*;�"K�~���'��=�ߏ]�yc4�Q�t�0�c��,8�>-�&�.V���K��<���K���IW�xF,h�39�l�ed��}"@��*�8�����,r}B���?ً����?I��85Q�˾}�r���]��d��K>a���0=QGϩH�He����V\�7o�����M��ir$k�L�d���)�|2�� ��x���R�,�<]GА��C��?���?Q���n�On�Da>8���:"8�`�$\Zj �e)ۮ7CdC�	�T>p�5/Wz��}Y ߞ't�����&�l�5�הO?�8�F��؍p�M�'=�v���M���k �&�  B�+<�VM  �/D��RѨ\%!�Pvl�1r4SE-���ɦ�$��@�@�4����O���s�X�n�`wdH��n��Ed�O��DX9NJ��D�O�%Z%��&Įݼi�C�'�M� ���?�0DÖE��t����'M>��E�>�܁����B2~x�6˚�%+(J��,+bm{1#�m�@)��ɗ�P�D�O���2��GG2;�H�&�ߠ�:4'�@��a���2F ��e
���a��R����q
6�	^������OLQ"��ߑER�:��T�gz�PS�'��ɻ'�0��	i�'/���I��x��`UEEetB-���
7F�%B��?�F��?�p�	 b�tb>��UEH�Y�-jP+�L��Z]~F�2�a>s��K��n�ɸKd4���7Z��+��af�p�ရh�b9c�@�?��E4d��Ժ�A߭zO�XA��*?�E�C���IY�OQ��!s����� �L�D*�B�b!��DFJ8jA��|	ӫ=�ў��I.�HO��qA*&c�t��*[�	m�)a�N�٦��	ȟ��ɩ7�a�$Uݟ\�I���	��#����vo^D����A.�]x�����m"An�<�L�`�{�$�ϸ']��H��ϰ�
Y0��T����y�c��S_�r���P�y@N����O׈p�(�G?I�Mm����]�3I�����̟0Z�4�?�c��?ُ�,O���ʖ ij���/L;O
��J�  '�㟀��	 5��t0��O�vT ¤�;���D�O��oڮ�MSI>��'�r-O`��@���h� �֥��t1Sbєtڜ8�+�O��d�O6�D�º���?��Oٲ��ћ?LdI��j��mqJ�2���.R��%����}ś&�B2�p<Q��7.2����]B����C/l4���`	H۞yw� �����_&�hO�(X���2/�,tJ�M�$A��Mh��4�r� �O�,�b��/L���w��מ��'�1O[�6ON�n$��4_�G @���|��`�2�Oh��M���M��۟ #᎕�� �
�N�Y�e�d.��(�	'v��x�	ş��'9���cG�j4:�I7��(��6υ����J��2�F삣�5U��L)B'd�'3��;�
�0��#��P�f�P6�]! �d �aK�u~��p�Ew�qȅ�(OR�Q��'ḓO䢢��x¸;��ƩS�\S�"O�I���dEfiy�F<�r��'T��dZ"Y�r�@%eq)J!�9'�=�I>1��7&���'��Q>���H�ϟxbs	��*�LyÇ�
±�FSȟ������I[�S�L�`�E�"T p�h��ډ59 ���!?�#ll���Z�"� L��y�TK0F2�5��4��	�Ot&�"|ʴH)mT^�8sĚ�l��x���q�<CQ<o���Z�ӏ
A|ŀ���a�'B�}�CN�<�)gLܴ�8htm!�M����?��}�仕@ѱ�?����?Q���y�-�7SI Ti�FA&S6ڤP�'�4K�ra�V�O����F�	M�qʏ�G@�u'�O��5���yVf�ᔃ��y�l��ѩA�n�ᙖX�yJę��ꋬ����EZ^����'n6�Չ�w�4JF��-#�I1��LΈ{#�|B ��?9���y��F[&1�!�J�W*�$�#�y��MU��ukC�N���1�?���'H���I�I�j����M��-��(H� %��M*���,V���	ǟ�����8�^wHb�'@�Iб\j�ٺ@Ɍ-z�0 ��J�$�@:�eW�,� X��}���͌?(��&ʓJٶ|��'[��6�����H@�a����ȋ�+k2(ţ2n@�@kF�遼lu��U�xr��z�vx����/�H�!���6��[�H��ޥ-��8� aU*�������=1�y��98&�A#�?����׭��w���|��[�"6m�O��$ƃl&����G�m��%��NB����Ou�լ�O���m>�R�\�J��3E�Ot�|��5% J_��Ѧ�Z"L �%}����C��Z�Q�TцjV2g���KB�It x��c	bq��m�=;ԈpA�@��s�]i��7�Q�l�0��O�=%�L�2ϟ��u g���W2^��o=D�D��؀xt���Po_aX=�S�;�OB���7�0t�e�j�e���7ب�O�<z��K�y�Iȟ��O�����'��#�$Y8��L�6�@���'��d��_�$9pc�G�[&QBI��M�ĎY3$�(��!.�^hi�Q&�>����-�`�F�MN��ܼg_���4=X ���s>9�"�eB����Z�X�`�������K�O�$�"|����3����+SMА�7�LK�<	�2Pڄ`�!��'r�j���j�'�r�+�d�L%p"M��2Z��c��J z�, qY�p��쟠{1腸%��	ڟ��	���̻W�u(��F�t{@b i�Mp8�S�P�t�.xa�
���5��#�L���O��������~�+�� �h�#�G�;1~H ѧ5$ɬ�*3i�'B	$5���F�Z�T�M�1���0@����1����D�8|�\��6g�<�|��LӀ�n��������|�'�b+$|*U�K"Z��p��C)~m��'ia~�`R��NG�(h��c(_�?��MΛFo����˦����?A�B�4�O� 5|�N�,�@��MJ ��Y��<(���'���'+���h�I�|b�c� 1����Ö	��]���M�-�5z�M�/���󬙖
'����D� ^���L��Rg �K�d��R�Ż@��̀ū�;eKPt����Հ$
u-�o�,�O�(nZ2$C�EHU�.Bh�Cn�+���$�O��=���D�m�$��X(>#��;�Eֹf��{R�D$bVT�D�+۰�W/Ȍ+��'$N7��O�˓8N�-�a�i�r�':�8�V�_#C�B�c��?������'�b���<���'zB,�8t�(�i��x?ٛw��`�*��`�5����tk
Ó|�F�2�JD����á<��Iu�؟+�:�X`"�'޾i�g��O�T�)�O��D����I7bh��I>�8�ZC��u��E�'H�|����&��n�?E��=y6� ��Gu��a���'\���bfͰ:���e����'/p��.oӬ���OT�'_��m0������i\2����1g�/Y���?�Qj�*j|�V��j�Bd�ׯ*��i6��	���I4+K
(j��� e~��[:{�T�ᅵpP�*���5玩��I�d����O�8	
��=X�0u��i�Ot|�"�OXm���?���il�����AV�:U��'E$)!�*D�$9�NBI���Q��ݙm����Ra,ړ�?i'�*ݸE���5e���VT�E@�	��4�?)��?��hY!h�dE��?���?!�wY��§ȁf�t�G�R?��5��:R� ���q��%*c�V�Ϙ'*��n�7U���
k�F��w�F���;�,յp��M0cD��~h�d��Y>�#�L
24�:�pY�K�\�r@��7y���;?��O���)�%�X�ul����H1.��"�@1P�'J��2R��=��u��D�? *��?!��i>Q�IZyb�K?K��C��Q*~T�C��]^����OW�B]��'��'%�꧉?���/�d�B��<2z#O0`���ǅ�Zty��X8��"��/E��J&�4�=в U�.h��E#=��2S�ߟn�E��'�v�'�z�@#@�
� A3A�r"�̓�Ę��?i�s�n7��O(ʓ��Ҧ�k3�œSG��=z&��9�!�D�[�LpS�µ<����E�:�'g�6�C��'��Q�'"3OPXH5i�
$f,�*�& �X<X�w�'��d�0$b�'�iS#�B��~P�]7�h����A��k0��s]�
�6�Ě\i�d	��d������Q,p,� v��`i�<j`d2N�A;1n )Q�6����E862t����)y#�'���+o����/C(���D��>�O����KJ���Q����fsCO�%9�bL�Ot��
�_J��j�	� &*H�!�'A��d2����H�'���p��*1�` t��/.�|��Z)��y1��?a�-ʔ.�|��
ۄ3_J` t'�1&����r��OZ����!�L΀!H�ԲQ�I�)�N�2���u��D�@���nLd`��OW�3����y �� j]"�)eh˽A����'ӼDj���?��)}�L�Wb!h��S�ư?ܰu���)D�8��N�)H���1d��2�@�p��'��jX�>�UFH
rF�L���1xo�0�B�O��d�<��3~��q��?a��?Q�Ofa��ႅ����P��j���WfRr�X���W�
��IvP�ɘO������b?ѵ_,]���P�}:�
E�#n�jA�&��
Q^�`���S����|J#!�0g�z�ɦg�
AJ0+��_+F�pΒ.6�.��6?��|�7��O�=)�O��%�<��3�	�B9�$��9�yR�ւG��Q��F�y��y�/����De���$�'���c�.��c�J�;��r�L5no��sf��y� �I���I̟�F����e"��ZRhۿ.j!�5��Yj�I�D�;����A�"n#b4����uM Fy�ᏽ&�8�1���z�
��%�L�r�{�ӎtL�l���̺l�����Z�m��UEy�)^g��P�͑���� $K��D��?)��d$fX�Z�F�p����"�$�Ąȓ�(X�m�L� ����($��Zݴ�?�(O�$���j�+�e	����T�\�qw�J�d�$�O�L�l�O��Dj>%p�G?V�-p�g�z�l��#%ݔR�2��d�Q�^}�x��!ݨ9��Xv�5~�Q��ď��i],��PQ3O9F���ͮw^�Y�� f2�xjA)�vWvx�f[bEQ�88VD�O��d ?a�̨R��p��˖�KW+�K�IW�<�T�;�x=��HT!(�"�2�l(�Ox��I$r}���.ԬH��9%�"IL�ľ<q��
!���'�B_>I(��H˟�s mY�.���b.�t]X���ş���+���@�F�|�B��4
~�Tr-�,�+� Z���;��}�2F(���'1.Yڃe�dH�L�c�pμ9�r�ѧ8+�O$��0�Ft��0'�q؀��Oz-�e�' �O>����ڒy���I���^ѻU>D�ܓ�C�������h^R� �ia�;ړ�?i��z$BC̋��)"pjV$0�(�	b�	k#���uF�,���� ���|�7ȅ�t�69�2XTrђA�I��l;�j��*'�p(T�U*��\�|��Y�.�P�ɤlBe�4I��g�0��řU����� ݭx�\��N�<H�aX�I1��)N�!F�O� �D�a�]Pf~@���Z	h���Kt�'��	4�>���O@�=1ůO�EV�9��π�-Qx�d
��yҨ�7 E��O�U�4 �3�I��$�l�����'a��5:3"��$���%8U�c���W�j8:sMZ�
�b �I�`��矄�\w��'x�	._.��x)��k�I���H�ϟx�R8եơ1���o�/ (]���	49�Ե0�% ^���*)U��9#F����� ��b��A޴U��-hg,�t���삆v��b����1N�k�N�����4����+!-�U��.t���}�R���N�/y8U"����a%���ش��+a	���iI��'y
%�)Be�mJr�
�ZPv�[��'��<"\��'?�Ɋ(= |�� h?�7�
�r�6��S�Ž [���D
EO�(���%O`��!��;��{��ͤ~Gu�ܹ�ҙ���_�$��6@�F�E��J3ړN��������D���ɓ�т �$�����N����\�~���;/M��� �ވr�|�?)��4����"J��p���Of��R5!a��O>0��"�O��?����@��1P��iW�ej�7kk�P�K�0��x�N��U�Ϟ��UCC��i#0M)�L��_b�O��܀pN�-�<��橌���\)�O8�c6+���-�@[�t�x�%�l��)�K?� a��	�484�0��`t5?Q@h�����f�O��Թ
{b����͝����m�	.�!�X�Mo�=���!3\�y�W��qqџ@���	�3�"��5�L�SrT���̄O��'j��<z��	vB������ğ����|��Ą%5��J��L0]��$�3��_n��#�GO�d^>{T��:R�q�|R��8=N��?'A�əd	hE�ijv+�!�drÀyX !�#�+f��ʱ�-�2Q�@��R�O�����ށ2��[0"ԩo�`"��'<��)R�h�$�O�=q���
}j���/߆eb��	�y�ʖLr��1�
R�|H�u�ą��{���T�'�剟b��mP�3\�McG+D�$�f�݁;2�	�4�	��,PK|b�O��(�3��`83.[�{�"�qwC�Z�B3�hÝ��)�M�wXȐ
�	j�'�BkR�͝I���	f���m����l��D�Ŭ�c�R �瓟m�LY�U/`�H�H�j�S�<�uR��T�<T��y�e� $W�Q�l�O��oZ��MۋR�*��a<�� F�D6���F�3*��>�	O��1� ��)s`A� ��Zi�O����O��87`���V?q�Ɋ ��3hĐ �� �.��m������<�N�ӟ���|r����؄��Z帰ۑ�6-��p�$�ȭ W(�0B� �v����$X#�\�XQb΀k�^���͆�=h"���)�	��U�T��y�m�bJ�<�!�LS(z�$<$�d[���O��d4?�@�
<U �G�N�"љ�̄d��z�0�qBB=���h���
H��X9�K1�	W���Tg�Of�R�+�2>ش9`��a��ACU�'��	�]�n�sߴ�?1����	��]��$��^�B�-�@�tq�曪! ����O�dy���9Ab1���"�BC���w��Ձ��;���:4ƾp3D��XR<���PZ~���-�|� ��3=�)���
8Z�Q��Ǚg�L�s�O�-ذJK�:N�Yф(���Ъ�O�H���'��O>�T�D'<�����K<7����&D�,9H�4���Y�ÌEg	�-#ړ�?)q鉶7R�c�kL�,k�P��ႍr�4�?����?��N�K�А����?����?Y�w:*��ӥ�S-�=c��M�HW6�*ƥ�(<r}@�D�*`��w��!՘O��'�di��$
�{��B����>�]M��k,zԪ��5b��iH�Cխ֘O��'���)B���v�f����C�f�(չ��|�(C��?����y�*�X�#�ݐVz�%rUoG �yR��o��-8D��V*�ȷ�͘���j���Ě|���K�����
�X������7b<~���J�B�'���'�P�?�ٰ�دM�	�GLQ��5�4Y�RN�2��j��Y�LZ�M#�,�k�j�<�T��W�-��(Y[:%S�A�1�B)y�o)�,��U�_2?q�f�����OPM&�$�V���*��A	ICA1�J��[���'p<6�g�'�����
"F�bi F�Q$U>QB�n*D�L��牪Zva��˹v��@(�Ʀ5�	EyG)]�26��O��d��`SJe�rkD,T-I�)�)*:����O>
"�O�e>y��m���H���L��u����%*@'h��y?=���%猜v{Ic���X/Pe:�F	��f1xv!��Ln���S'.�xغ&ɾ;׶XK�n��ɓٴo��c�ĳ'��O�l%�����E_�qT$�M����s�:D�(3����ݼ��6+։+x�А��8��^������O��JU��C�ޡB"i�
GV�0J��|���C@�6M�O��$�|R����?y�dj�d�S�@�����kT"�?��=��� �(V�*��GBl��e�(�t�'Tx8z�'A/sČm��JR����'�V��#	�,QG�娦�q6����Z)8	DTJŋ�+`b�JO">�� ^W,��DZ�)�g�? ���&`^��&�Ȩ"��8[E"O���LL�f �C%I�P�<,i��	��h�����k�J�"DH�BM�^�xXY�p�z�Ode��B�n���O��D�O>���7M�����P/Jtx`�Z<=@��ҕ�~��J�4����h�',c�� �� 9���M�T�`�J�9��9U3u����H��Mk��\<@�rQA2Ê����(/�>��Vdޝrpe�'"���CA�2�8�x��	(OԘ���'m���?�O�Q����;r�Ó���Bʺ�9u�+D�$�pO
3���AL4������<A!�i>��IMy򍞵��Aq�BP!%/�P�%�,"-���Ύq&R�'*��'�b�]˟����|ze!I�V��`"�,���X ��.Ab #��R�����7aDMc7�I�cF\\ �K]9��A9E	����Y�
��Bmt�BAbΟ[�J"?��өYNU����[�z&ό.
��L�I�M�B�V�'}P%iQ�.\�~P�Ś�P*�;�'T��!�|���r� tB�M�K>��i�R�x`���M��?a'G�;V9J1��I<({PD�$�?1��
�������?��O̉�c��=/|`��
�
V���_�<B� ���_/u;��2�Ŕ0C� �k��Y�'l�(��BS'OS
Q�5㘫q��%"���,v�L@�N6U`r��uB�6eU$qi�B$�2�j�y�B�?)2�|�jg�q��1A��U���+{�d�<iD�aY2�k��/N���0dk��hO�i�ܟX��鐾T��1SS �=��D5�Ė4do�th�"|Z�O�h���1Fx(�FK�Jưd��Ot@W` �v�@��%�p&����	;��D3���!�@�����K�Ix*�%Q�������d^�R_Q>��.�7s�&�ԥ�*��` ?��K��t@ߴEp�>=�'^4���
�#j�J��_�]���ȓ7g�x3�
I�-	|-��d0���G"/�'0	�HP5��2t����Y�t|�m
۴vUx	�,O�!�-�|Fy���
d�f;��[�1�P�zg�U��'��)[ӓ*Φd�P�jq�Ԏ�0|z�p�<�&�i���� �k�̜�ʇ`�\P����D�I b�P��=�3�<?�����4r"y�1K�0ǜC�I��~��aƣv���񭇱2�|�fp��"|r���wr�y#+HU�z���瓻yA	���Oz7�ܰo�X2�L��!�@Tig֬cU.�0!�O�W݂0����Al�(!��YZC��!k�B�D��'��
ݐ�ఫ� �6�[���[���lڕ�6����D8\��09����E�eRg/u �p��Nn�����Q�����I�#�6(�C�~�����a�7�~��'L1�%d�R �T!P�(t㢹;&Q�8������j�L �I�@	��A$T ��OL�=ͧo�	�g0���̍[��?V�j�&0\(T�i2L� �'��ӵ!��t�S�����ƚ7[�r�b'WJئ�������83��٫2}���2Oc�}�Q��s��ɛ�.� �9 �t4����k��,���)i^�A�e{�����4��l��EdSXt���|��G<q��H���57�H@�a���<)G�O��� ?%?]�'��c� �8���D�H��Mx	�'�Tp0ҋ�xw�0�
��FR�����'?L"=ͧ#3��#˅\���bJ�=>��I"�,_7�?���ƈRaDѧ�����?a�?��N�O����b���=8����`XV�#,
\�1�i�D��������uc��g�'�5Ѱ&@*<�&���(^"�~� ��W�+
� Ó����%@Ϗ����!~U~����L�x��$~��cO�3�}���c��Md�$�O4�=�'+�U�9�P8� F�xSZ���'F����.W5���W�-p�`�j!�'�"=�'�?�,O�IT��* ��2Bb��z:)��Y]CBD�Ѡ��\۶��O����2���Op�S�j7����*z�Te�E��'r됩��'W� �L0�&o�n�x�c���08Q�$q���(]�Hͺ&��0���"Ŝ�qA�¤�A�{�Bp3#�&�id�I�M*P�d�}��[Df������w(�,U���*ړ��O&8jק�c{�@Uk�:pz0it"O�(�#GTcUZ9���QUk�u�R����4�?�+O���H�O���U�~⢢����0�K�o�p��� 䟼��	̟���؟ bP$�l��|���X�p����D�m8��ڊ!3�$�i�$Q9Dk�\ɋ����Q#�F�+iD�D"Q�xk����m�X�ƪC�9"�r�#Z�Ce^����Z���'!1�d����+b��LcƸC=l�KEU����I( ��P򃃅!8Zm:�nǏWz���pyrȒ�j��<��%S	�8r0���	�/l�@墒�b1H������5(f� @��*?� ������d�5��Ђ\0F���
�QFdQS	��cq�H�C��c�X�
�9yd�i�1O�ԛuiط@�����Hu�@�	=S��y{��T�Ć>,����B�+�>9�@R�y��*�?)��������� &�� �\cC��֊�8�(x`�"O0M����n�x�#��� pP�`퉿�ȟV�2��}[H��g�19��1��������OhD�	8(���i�O����O��i�O�`����p:��g�+|*ΐ+ 
UH�f��~�\�#��"�����\8�U�m�x���C	+mu�d!5HW�I��J"m.F�Ue�Bζ�p���$(�J�?���&�X f�B@��j<?1�M���L��u�'���K6 V$��d��#�`�{AE�t�!�$��>�ȷ��mt1ke.ܓD�R,��|R����C7qqːf�4�*"�;v�兔9d"M���O�d�O���O�]�T�Cu'�<I� x
T�G4Q!� Æ@��5X>����˿w�~�U��^f�p#>�)X
%�d��d��9we]��j��F�l��ze΄�D6֥:��Y�3���2�3ʓ. <u�	Wָ�j L6[�I�@�s�Ҩ�I`�'���xw���TprM���?�da��i8D�4�&���c
��Jľr#R�!�h�<ї�i#[�$��m (���O��I�)�W�^t4�.A�d8C�')�Q�'��'���E��$���'�1��Y!��%{���.
� �kC�ɦKz���ު9/��F!<@  �1D�B @����dھ$�)_�zr(E{�� �?��'*���'?�IZ�W�%{���#!ZD��&/�:6��Q�G��O�.8�'i�qs'K�{����' ��
�� v���@F��,~D&}����> º���<���?�����D�OL���O��	�v'��B���1;�AB+�y���	`�'�\#=iV%2B��`��	J��T�sS	��'p�m�N<qS��O��M����ቁ.�VŸ����zr�A  �ip2��Y�DO2	�2�'���'�����:y�<�[h[&b%l��A�/8(��I4�xӦ�D��)<���ڟ<[��?7��x�C�'����5���wLϛ7<�I.wq�<�"�����	Ά���u��'���O��4Ox2mSp��p�� /�⬂ëC ,�'� �:��'�8�$�p���u��	�<�$#�V2�abG*�r�^���G��?IU#͟���.x콛������O��i�O��zI��F�iiBmB�]�V��&N񟐸Q��O���\m#���Vɟ|!B��?7-N1C}d�P&C_#<����0d�Xŋ[k9�7����0��O���8`j�Ο��I�?�kd�Ϻ2�b"� �|���W�����t�$�I����Yw�R(�OV���ڟ���L*����@Ύ_�� �k^�/�:txQBj��	�ԙnڲ�MSa�L��)��0����7��Y��Q�RM�a�i�B�8Ƶi�(��t:O@ �~�(%l��?��	�<��*���2���#��ҥ�޶xmh	W���M��C����O�7���?MmZ��������Q q6l��J�)B�$GňbF��ȓ!P�#dP���@���\	;�an�����Vy��'���iԎ
��5�@�2��>�v�z
ߦ��	����I�P��� ��V��՟@ co�w��#%��5W�.!+��i��X�l�'��\� �'��Y!��O1�����I�Ws�+r���$�Ob�O��x��7���i@+�(�RN�5���'
r�	R���jb8��Q�r��-�0�X2.i�'��'}�'��	ߟ�Pj�)P`j�D�*K��y	����M�������O���O
��?a�O.���'��@����`)\��'}�-�FLR=81b�*�V�&i��'�0�#S,3��H����GM���'��신A�qnD��a�N���5�
�'vX�� ̄�W��+��*[��8
�',�@/�^�(
�g��V�����휈C$��� ��πtp�Õ8��)�T��s:pBF��#Ё���BB�&��#� �v�Q�g]� ꂀ�F)H����C�DԔ q\��âƌ�@<�ZЯ�����Zk,c�4S��֛I���yJ �I����E+F�yn��=F�A�)W�H�a�E׹wO�x���Z�i���{N\-4�S)$��C,܏m�p���� E*"!�BS4�f�a��N���6�ãh�9i�ȗ8hVm���t#����%�V�]�[e�~��D�i�� �'o����E[�����"�3Jz.��,O0�=ͧ��'��5Y���"��	p�C)=����'2t��J�<Dm�qpƉ-0vL���'M���6ʛ)�豢UoG�q�H�0�'0�xB6�΢O����� e�rUA
�'��PiM�5��"a�߻L�ڥb
�'���p(�2P���y`%���R
�'��� )�V�BgH_��jiJ�'����p�ߧ|'�)سd�m*5�	�'@ [,��Xq���2��>MR�'~�]@w�����@�3��b�"���':�ࡳ��2��0�"^;8� �'_�c��2i
�HR���Y��ik��� nԱ h�)l2���1�Ԝ4��D�u"O6L32�ȝ=fz$�!ر��T�t"OM�'��1zzp� PA��,r��S"O� 
�n�6 ?����,}`ح�"OZ`'\�(1Ub˜e�����"O�D��ц~����ǝ}<\E"O��̔�<.��i3 ��K�r��"Of���h_�P;d�U��E�w"O�͊�G�G�^�pvF�/���)�"O�ݢR�m]���a�ԻG"On�!7�ӽKx��熭R���"OHT`E��\Z��#�I�ά�d"O>1�F���j����t��}����"Of�"���m�b�2��>a�Dx��"O�����AO�����1�ܝ�g"Oh�6ʃ*e�2�C�'����a"O�|�@�I�x�R�buǆ/lm 	�"O�S�NI5/S�d��3?�,�D"O� �!��<�t��t�"u$(��"OإyFO�-jިh���T�lt�&"Ox�(��0x*���!�%b�$x��"OL@ٔ��X��`���)p&�b"O���#`�-3�0���G�'" .�B7"O�5�FK�Q���o_�W*��2"O~��&M:v��u�Үɶ;��'"O�9Pw�
/ft<�9q��C���"O�Ł���&J�8���&��SE"OLɁ��.M�p���@'9�j)"O��!�-�\�Ĝ3�Y9*�`��"O4��>L��l��bn�U�4"O��Tȏ���"Y1j,f��F@4D�8a;#�D[��,_Z�H��J5D��Cl �B?-��k��D����>D��`J�!�Z�!mE���6�;D�lB��/CN>Ř@ʆ�o�el8D�d�d��iu��p��lH�����8D����'�-+�ba��@��
.���:D������-�BИ��E�4�e� �7D�po�k�� a�+g7��7�7D�!���M� AsF�P<	J�|�7$4D�xC�"b=��#��Êo��h��$D�|�Ul�!
p�띦H����t�!D�\
 ��tuJ�su��~}s>D�����3@<����b.b9i�(=D�|���>S�m�f�C6#u`���<D������N����53-L)Zae9D��Ӆ��6)�&؊��j����h8D�S�6o�yѷ�� a��T�7D��8"Bٍ��t{Rc�?
ް�( (D��q�-P�v���!B	�/�r}0 �'D���4��K沀kѦB�o�f��c�3D������<`eX�!rf �b�k�
'D�����IZ���ɢ��'�����"2D�T��L'���xd�ڧ6�H�굃1D�tQ6'@�$�p���nَ7{X{w.1D��#�);���L�*t`(��b�<I�-C]�jD�sa���iJ��Z�<��\�`�2��t�B�1��P1��Y�<	��2^�����%]8��w`Dm�<)4aKQ]�1���	'���D#�i�<�g�0]��K�nօq9�q+��}�<ɢ��)#��m;u�ͦ<,V��V�^�<q#
�<M|0}�֢o��a��_f�<� n�!5���[𘬀EH�x�<� �D)���j���T'�+WL4z�"O���E#���
��A�E�_8�͋"O�$��X6���K�d�,	4��H�"Oj���GG�$�H�1���d>م"O�u�iڎ.�
�cr��o0�3�"O �R0��-D|(%�jώS���I�"OXr��)D,�Q����:�5"O:Xs5�"t�6���i�`�"OP�� �R?gI�8� O�H���+�"O*�;$`[�b����f�Z8(�"O a��o�]Yc�\*w�ڼiW"O���֮�%!L̫��� kZI�G"OD�R���$b9qBDH��6�R�"Oh�`$��'<R\ه�4:�4�+�"ON�3P�<v�0ii�,N�:��E�"O�A���$}<���A0��\	!"O�T3��?�0�;"�u�`4�"O� !Q�_#4��і�3�����"O @��ܦx=��b1��6T��4��"O���E�� 1�~\�S�/ѾD��"O�a��n̓V�Fti��=W�N��""O�<���~ ��	�`�j*��#"O>�� N� ^&t3w�%�a"OB8q�EqBnM	�G2z�f [�"O�}p_2�I�gO�KS����K�*�y�)I�*`�4%Ǝ>���F� 6�yR*���<`�F)D�8@�c/�y�����0G$DK�E��ƈ1�yBN
2J=s�X�5�2}��b���y�
(g2�0J�?0XԀw�D#�y�AI��l�W��_�@�ʈ��y��%kْM��E�iA���%���y�+�)H��u�Q��e��M�aU�yr�])A
H��!��F���WBB,�yB��'�H�c�CԬN@���9�y�lU�ZY�A@��DR�m�e^��y�B�o���b*�?i-n<�R$���ybÔ�3��Yk��$^!��y"��>�y�	B����m�!O�l1����4�y��գe�b4�W��GI"�X0�E��yR ��B��A��@��9��F��yb��k0$�	��:<�t(��Gŉ�y2`Ԩ ^���T8��cI��y�$Q�c(J[G$�j�F	S䨋��y���s �2�0h�y{�bվ�y�e��-P���v&�*Q�pK�D� �y�͂%��M#&���|́Rʒ4�y2�C�x�����\kyClΦ�yb�38��%	�*]h����5�yB�@�Z�As�k6P�J�����y���?��F&�?dl�C��̲�ybj�J1��q�GЄ6�>T���ը�yb� }�q�!j�>(�~
D�^,�y���5A5����-�  4���y2oz4�q��@��a�(���y�c�'KC����ls�C�g�&!W!��72���8w)F`S⥲���eO!�$֗y�+�2����`�G�|�F�ȓO~�C4$׊������@1\���-9�I7�\��Z(h�%&�9���X ƌ��|��M'K'�]��Ow�P0%�&b�ZԳ�Ŏ<G�̅�@c(�Y�eD�<�d�6B�.��<����pGi<f��Ţ=ی���S�? f�E�	�Z��L2��X�`F�x7"Oе#���#(T��"j͵<F���"OxA���d���I�?u(h�s�"Od *�`Ģ2�'�H�0�ܡp"O�U�q�W�F�<�i��9�u�a"O�II�ήO��p��\V �x�&"O�	&n�����n�=t ��5"O��27�M�N�L��7�#�HDȐ"On���N��I���u� EӁ"O�|����<y��5�TDK\��#f"O�	�"���	m�ct���8�"O)j$��&���Pע�zn��0&"O�`@1�ҁ?�<���J�VΚ��"Ol4���8tt�u����	o�N���"OR8aGk�X%�%a£��D�����"O.|��Qwn�I��(>���"O�ʑD��%�d�	�_H��Qe"O
 ��� �X$������uLBF"O�����D�I�ܨ�E�w�,���"OJ1I�
]$(%;2Ȅ7T�axV"OT0�g�%*���d���-<�T��"O�t�G��0<4i�l�	p	V�ڔ"O�@��K(DеpT�����"O@E��A�]2Rm 
��w�mh"OPt��a��a&���p�8�w"O21���]:�`Rf�q���"OAӃ'	�{�X�%�4/1� �"O6�A�
ԛz�U�Rӎv>�Tj�"O���u.F=��q�r���SR2�А"O�Ѱ�ìfТ���CcI�E�E"O� 	'��ekȔ��j9�I3�"Ot��@I,w�Uxl�
T�$"O*3EI!]�n�s�*� ƌ�V"OH`��_�>��b׫\�/��a"O�|Ӡ�E9���FjH�^����A"ORH�sDѳ5��4a�	W�E�.�yR )ff� V�H�G��8�f���y�A�.�b����LX>�A ���y�\f� c�H"��0#���y!-C��*B�t(��AW	Z>�y��S*>�挋��_� �+v��>�y�U�Rt�Q����4���Z��y�'��������4E�?�y��1��H�� ̜�`i"4�Y�yb�H\�|)[w!%*M&�9B��"�y"l�-'-R��UͫOꦸ�a���y�
�3�ra㱋��I��К0���y���D��͢���=N�|5�ɀ��yr�۽xN� �cJg�8b���y2�t�h�`�A�3n�kqnڢ�y�ݢQ;r��dޙ.$ᑪ��y�ǀ�'12Mp�%S8b�����9�y��M?�Kޏ��(*����yB�E&pGX��f�J/s�l<����y�KӖpc�t��eڿ@|]�F��!�yB*ēQ�*���lHkX�% ����y⫟�sUεɁ��k-� p��_&�''�8��+�(�t��p�E|l�\jK>��ǢE���H%]�$2!A�~�<!�[:OM�ê߫k{%x��P~�<�4�@)V��MBS��e�J�i���w�<Y��>�6-�����ER�q��s�<Gˋ>!Ě�3"jČH���{cc�N�<�M��?�8kQ��*o�	� ��q�<��bB-w�.e0���E:�jg��X�<� ތ���'ǎ���a�����(w"O��є��7?*|�@��/( `�"O�ġf��;+���3�>%rh 2�"O`MPfݨb J� J;� � �"ON�(V�.}���I	$� JQ"O�Hq�#ͺ.֪1�EI
�$�N�1"O�ő'�=I�����I!LW*e[�"OఢP+F=M�ȹ�&�5n�f��1"OP�J�W����&L�r��%��"O�k�jF=O�87KEe�	Q�"O-`��E�8rt����hb�"O^�8��q�U8� Q�6wB�
�ݝ3,P�mڥ*�$���F�x���QE�`*�,ԹqDĨx�:Y슜@&8�OX8�$D l%�8���D�X$H��Y�X�d��gH��-Kf�M�t=E��' .0�C� f�TA�P�E�>zF"=�1F� W�����j�|���GϦ� M6 Y�F��ق�@�bzB�IF)T���.-�����30{�6-�:T�r}ӧ��"^=x j׫̛��������%c
�)�t��?��U2"O��j`�2;�ʘz�l�2af�1I�,��f�(!nZ	sOmR$�f	��'��̃e�&�<����u4~�z�6�O����Z�Y��XB�`� �Y�zW���g�)4�f�c��V� ��'���P�#D��������j��d_�d�fy)Ă1bY��-Mp}H��|�'	�:o��YIQ�L0s�Ma�(�o��0Jχޟ��4玢,M�T(cɇ*wg|y�shw�f�P����*%��R��o�츳e�M��5֡	�
mL]��-��,j��G��hOujƩR;�H�j̈w`Ȫm"x��efOv���֬8����"��	6�`�l�^_��&�O�Aԭ3��t`Pᑧi<�iJ3/�]�1�U�['F��SܧI|LiK1+�a]p�g�2��1���~IHI�W�9����(S�~a|"b�=,=��Gأi�$,
f�G��y��£y��<�F҂ �|i n�8}1�|k�O��`K���H��\��h�?d�}��O۸0���]	��:�LZ�\��$��!�J?b�t,�H��ˑ [�z���+?Ǒ>�X?m�� �k�q��p�珌^P�����>Z�,���Nc��J� �1*Ȅ5����2Q0 r��(p�
��L@xL�# w��OVT�7��<9��b!g��в���hU>3�͑�AV����	���@�V?��%�Ŵ��i "QT��؆.M*R\M���F�����Ϫ-@�=�G�ɝm>��R��fX��X�'p�0��ŗ���� � ����O�a̧���`C�F�<�M��jV?��Ą퉘)Z��(�X��p�Uΐ�u#��jC����|���7h��	�2Xq� �s&_!�E�ӰM�B���OA�4ZEq�`�w��-8�}���8��Y	�o�E5>�j��۬�g�4�xr�Q�K�� s�ˌ\iH0r�O[�G�����p���#�O�PX�I5G���(�/U:f(��QWL
�U�Uq�ϩr}R�a��ij�c?1B� ������B������� b k��+��"@@�kl�Q	�r{R�(�L��.ꖱ�1�O/M���(��r���f	�]��� �нR;Ҵ+�P>��O��;WdV4�P#G�v�H�jN
T� ��I�R��F�r�9��CJK���aR<j�^�j�Pl���`á:�&ġ��Ao9���E'=u�9 K�B�:�b��^"+�Ex�h��`��q &P�Dtt���d��>
�,�����m�⡻�E%*v:�T��	zY!�/�{�^U���N��f�Đ�t[����8K�D9" .�p6�I�' �X�#�!1���mK���'���ʀ(������
d��TB�*b�ZG�ވ+�.��E.����1Z��i>�رV���)ؾen:lS���P����'�T�j��X��5n剜����s� ru�&:��]��!
�:1P��J`:3T(��g��?jhBW�I�D�Fs�b��4\&@�4Ş�K�a���Ӻ�ɧ1�\���-�I����q@݉U��:t%J.BR䬪&��4Ԝ�U-���剰{S�'�r�&oEպ�`�y�4FB�\���y�ֳ`�*y�C`<}��'A�T��Иf@�Ij�#��z/qO$���h��J��� 
������U;���& rS��˺{��T>�B'=v�b�#*�
H�FT���Gh�	&��P�=�OԄ��m�
�?QaJ�.����fĞB+�����GU&�Y�D0�)�缫p��lP�3	q	�V�
�7dV�'쓔�X5~�ȭ�t��,����d£32
8�p-��b�)���J�W	�ɕ "��r�9O�pQ�	��X/MzpN�3U���r��&m"�XA���4g8Q���?`��h��t>NMq�Ip��Q׬�����$s�p�K�.�|���V���U'��,�1����4�`��OM�y��,켈cr��2�nĹ�숗\�N�J�܊w��O�	�La�]	sH�m�NI(7E�4Uś�!ܐk��Fx�O��49!��49RTA6�ie8��g�����X"jԑd;R}�R�S:�h�D�>�|��'�R|���� F0�A��4�v���杛T�4A'�>ї��w)0�k�F�(f�(���Or%����7)���@��4z�B9�vZ����[P�L�ʉ�>y��E:ʓ]Tݹ�͖���k�A+�ځHŽ_lH��'�ZY�d�˓�l4@J|��K.�<�rA�U��������T��W�|�+3U޴���d�/5v��%�Џ}b0Q�E9�6Y�Vk�2����/U��O��O�8Q���2K�	`�Mـt�4 ����b�Eɠ44!��'O<���H��"���T�H=�6'�3Q0Ƙ�$@\�.�?!��IF
!d�N�$k�h#�#իRH�[qҩ,51O�Yul��L���i�']��PD%ޗ��]0���C�0���a�|�snץA�ڙ9��H\#>�Tc�+T"��3g�۴�As�%U��f�@�{�"�~�ƌ1����4Q�ՙ�b�墵����72�����x����U&JK؟�떋ȵ"zlkƊH .J��"���O�])�w�X�MQ�q�5�)���������_Z"1"�)A��2z]�ȓC��� �&�&
L�����-b�8 b,@+�
c��${kx��*n�'����ja`��:����iA���"O��$�C9y��F�96��)H4J��+�8���B��P!ԙb�j��d�ax��H##1�pq�b*|��u�qP��0>qR��+ ��{��	�@��9����l�dnB�4>F<�PO�nL�� �"�4e�I��k4�%/Q��Ia�m�0+FCap�C$G�21�XР�n-D�HsFʖ ���#l��z���K����<���H�}�'�DIP`���~(�M��?ܘ�@ӓ ?�N�?.LN�I�7#���VA�0�@h�Oχ�x�	8*��Lhd���	�D�0���:q`M�.yMH%C �d]�n�LJ!K�PʔS����u稛�
�V99���7W$������yB�A�++x�Sq�\f���"�Cs�u�����M�Ƅ|�S��O����Yޚ!�����:�P���[�r'PC≗&��� ��ԥn�Z
UkZ`��M<9��>�!/�H\��5�I�vPX����ufPQ;�Rr=��d�dF֘CA刟
���z�r�)b�(۱tf� sb
 z�f�ʰD�2L2GkN<R�&��ln��Y���7#�S� �	_V?)G��8�>�����A��Ћ-�s�����+J'e� ��/�Ӻ���(!����'Q�Uz˖��M'@YaR|�B$b�j���S���O�'6\���#���y���,�����i�%^��<`�y�"c��S�Ϣ;���H�QmB�O���r���IQ�Y9b���>�����'�*L��e.��5���\��"u~�cv�r��#.=��O��7���Tq���П>}P�hq�J5�M��gL?z��Չk�ԑ2a�U�0���_T�4@z���>l�ց����̸�F�>�i�����i Xh��(ӓ=X�O2��OXqb+�f7p��II+UV�p�֐x�)��*�㠥N�l��	"�?i�t�4햟8�8�Ҥ̂<�<���̐~S�c� G֚�[�V���g�=��O �d�I�;�c,�a�dH���ƘU�X�mZ��M�O�F
Bn(�����~ڰ��&�"��u� o�%h�H�S����%���2nh0��;_0�%���_"z9+�Y>��'W�=A�Q�|�+w>Q���sB�<��c�$
�H�
Ȟn�☇�	�CҤZl���	1h�|y$��d���B�
���bŇ7a��xE�K!|� ���-ʧ*����4)����N�Nðaѱ��5^@�Ot�3p�'�)�)6X��́0"�'}�4���3?Ra����<H��x�SC�9y{p0!�+&��O�dۗ���|aYE��@jq�g�X�=)��:b��SA��.C2�J�副�0� `T u8�������N,C8z8��h������ K�ja�����%Q��d�5F2\+Rub� _	=f�]g�X�S�$·&]7�r��e���~+	�U):�`����y7��+;j�!���N20�e&>��x���njd!F���:̈́����X�#骀�J!B�,��H��H�9���N*� @�ؒZ����P�i�>o˖t�ք�8u�t��OL��ay��QXj������b`��a(^��E�IH���'�I�g������$�Ղ0G�8=�5xb��Q�(3P���<�H���w�DB�:����h����Jq��%i�0\��Ɛ�H��YQb��294�SצP�2���*�{��(�KC5���D��-5�		T�ղK[�XkfYRT�H�V�� e\,��ퟕv�t"CI��M�`
R�͂+�~YhbQrTH�P��A��(�E��=p
�|����@�zb��je14Xdz��"bKѡZH��u�G-t����ҏ#B����Z�;���|`h�C�;ʎ�C0��3��ȓ	��$��[������-�$��U,  qO��+�� 7��#������#�i�Q�2;D��0%�V.�Rģ_�$^��k��.3R��d�R��dI�K�vZ�3��$׆m���w)�M��L(tLO�:	�m�$�\�rxж�Ĕbt$��(϶R���q%�';�M*pD_�Z�rl�"ᜳ=7X�Y#�Ѱ����@�h�8�w���p?�gAԵ������������ޑ�D\���	�H
x؋E� �`�cM̅h����o>���	ցV�]Z�ʉ3j� *��Q��y�E�I]����"F\<E�pPcE8g� x���ݰg�>\��`�������+�Xz�����0��;kj�x���ŀ�]��# ^ ���'�4���#�t�pY+'���*Ox�����D�dCf�C(m68h�7�Ϙ]�\l��,H�}
��''���陿Z���J3�W;E��p��U����N�t3z�Q��G]ܣ>	t��!R�2�ӐǓ&�`��V�`H#g*[)-9�h1���(!h�r��2&��Ж��a�S:�#s ߸�nxB��T�
�0�c�]�] a~Ҧ�Px�B��&�L���ʖ:i丵c&��<��1jF��N,l��B�KZq���Fd̀��Ξ*I�8�b�4N9��b��L�B�,!�ȍ\���M	�6.ў�:W���C�H8p�	��f�BiR ���E�M ��'� ���Ls4��XP$S�!@p{�	
�(��3A��e�24nZ#.0A����H6��k�bZ-ѓ���P�bK���TӶH Y ��	�ȧhvD�j�fRK���ؽ0@�}�b�҃H��P�)���{M�A�<�0�'�ʁ���'� �0�E�	'U�_>�0 �0PԘ��˜�JH��,2	�h�L|�a�AdE~�%瘠a�杽E�D�6�J:&�Ф���؅*��DB"�
�"`�S�w�R��(��t�G�"���b�O@�
үK(/��H�5>����)�'<�
�I���Q�h��jZ�(a�̂'K�.�Gy��	��S�`��*�H)b���7k���F� �]�&IV�DZB�v�
��`�ȥ
R�K�)ܸG,Q�7�`�ʓ N�D�lV�6P���R��|�� �0�[�Af�hIM�xˑnC>D�hN_?)��H�| �0@� kڹ	5
ބM.�1� �$I!� O�$�d�	�~����ꎩ&������B�+�����>�n�k`-?Ϩ%�f0O����➙F6󮞉>7H��"��W�D�cD�e�|bB�1�l�c��-pb�[� �4��[�ɸ2���4[��@��>)�n*0���X��W�Z��h~�ʞ/>�kT!�A��X �HO�xaG��W�4���@
��(�w���1T�	��TRP� �>�u��A�<cU ��EeՈ1�JSI_�Ȇ�ɞn�*A��,�sD�� �K�.�H��b�8����z�&I�.O?U�����|ɰo�(���2O_�<a4+�
en�$XR�6�l� &�zy�hYXH��5
�kaxb�(vդ���X l���)\,�0?�&�@�Y�I�oyL���,��uO
�{�#��5јC�I*)4�J�B� 2�:Q"�M�GRJ#?I�)DT��?�I���O7n	2qj֐,E�!e D����C�Ka2��	�T��Q!w��<Ʉ�����(��$�����H9#���#t�v���"OZ`�Vj��ܽ�G�DC�Z|��"O0�Ӑ(ݏ~�Q ����"O ��`Z�f�4ypՅ|�jm�"O�Q�$H�L�R�C�J�8h�	�']���H�Q�qzb �1U 1��'{2<��\�tM!a���k���'�DUp��B0����c��HS
�'0��01��cn�ҕǈ(=��}��'��L�% A�2��h$�b�Z���'}T��T��l�V��	c�x�3�'�2��!h7�L�K�,ܲnB���'�4��$��
z*��!���i��u��'� ���b\�u�2�&h�~�Y
�'j��`G=R1�m�`p�C
�'VbTc�/�4t�*�;A��0��E��'�� �O�a� L1Fd�2�'�D<��4k���c �$}�����'������aK���S��{m� ��'O@�B��Ǌ2����� �r|4���'z��:gf^I�x-aƯ�b�*��'Td���г>�V����k��2�'�\Q� DqZtx�g���ε��'*L!*���J��9�&Ȑ1�Θ��'�0z�LɽrJ�a@N�U�1J
�'8����O8
�䪧T4q���
�'�J0��]U��h��ۡ�"��'�T�c�
�_��,��&��4��3�'�z�d��2��Q �CM�"��&"O�2���9��=�ab5sMPd"O�ɸ�ب,�
Aw ��Y ��`V�D�< �0*�K�5��e�V$ �#��'��C&b]�ue|�HD�/��Đ�'��ỡi¸ءC���)�����'"P�q��2��)����7Z����� �Cդ��>�Zu�a���<K\i� "OT��%Z 1!�%� �Q�*1��"Oݚ�$�,h�m�G˂vd43V"O4I���В^(j�ҁ��5�bM��*O�UP�O!C����͒h�B �'x>i�bG�b�Lx,Sb���'�M�s��+�����&W-C�5��'��(���?^H������+�B�	�'��4�b��jo����*��!Ɉx��'�<�3��	lJ ���0P�Z���'�)��jT�nt���Ԭѵ˪0��'�9��J�|����2�
 _�ܙ"�'-�r���W9��Ke���S@����'��*rJ�3uH��c�bvF�	�'*(ܨd�̗ ��vbNTP�J	�'�t�9�H��pV��s�〈L�j$��']Dm90ΐe`* �!��2��my�'Al�gEłY��H�WD�.m�)1�'��`�6�E�O��,`��$�^8��'����gL+4=(��""�Hc�Z�'@�5iq&�p �q ]�F]~Di�'��@��܇3�2<��e�V� ���'�� �AHT�dWd�h���wc�x �'�4���m��@�\ٕ�^r�ȵ)�'�Ȓ�\�u�T��
Y8�"�'z��!@ʤ\.&���K�N?����'7~8 2l_1K'�� �ğE�̹��'�v�SkD%x��`�i\�/u��2�'C�Q��!�H�zaK�=^��X�'��A ��~h����#�;8>	[
�'��0��F�O�`�xw���:h��
�'~�I:�-#���VhC�	���
�'���6@�d����ը~�IY
�'y�E1�(2�01�C� �+
�'��%W�L?m��C7�:��-�
�'?�\C�5+r�qkZ/4�j�'�D	��DS���A��6h
�'B�(�t�1I�0K�	b�	�'G0Uy��,Tƪ�:o��LP��	�'���)EL�2��9��	 ~�	�'8(Q9p�]S��:�+�$�Z���'�DBU��H~����["d����'I��J_��@b^,Q]���'y��ڣhX�T��(�-Gm
��',�	u�-"��8 O�q�����'�����nW��=9���w&����'Lh"f͓R�4}㶏 �v1&�I
�'â��c�Q�& �ĉ��a���B
�' &�����y��4�%I3W��}H
�'�^)В�N�|�x\���Ȏw\ԁ��'~<H�2QC��#�CёY��x��'�9c��R�ځ���#M��Uq�'(�;�L
�"$��Sp�ВJl�	��'�����靻e;��c�aY�Q��`��'�t{��2"�"��6+�/IN$в�'\��ぢD�T�xFlS�
yHA�
�' I&iջ#��a�e��7���	�'�����O7b
���u��?'��H��'��98����M�EC��ˌ�`�'�\�b�eYLS�Č,nѐ�'�P9`����@����)��[�'�nx��Y�EJ�#�TZ0��'���s�"�/u��YpY�R
T@I�'�z`8����#(�&��T (���� ��#����M���ч)����p"O�I�eo�p~T�jFk2��I��"O ��a&S��n`"��1X�\�2�"O��s -�=��](s#��<GhC�"O��a��ՄQ��Q93�@��2"O2	A�k̃r�`��ebڕPD���"O�l��F)_��4B��^?ԅ�f"O��2��*YX�+r���4�cS"O`)��܄l�DP�&�U�|OfГQ"O���BI�,uq�-Ҕ��o56LQ�"OQ�!�Z�Q�F��'a�-\,�% �*ON��Ҩ Nv�Z5f	x�ʰ	�'����A@$֨��� %v�m��'��xa'�?-�h��E& ��)�'��I���_&a�@��Đcu� �'�@@��u)<D�.ǂc�]��'{p]�w���3���!���#]M�x��'4^@��5Ft��KbI�$%����'2�m� @6n�� B'����S�'�.pV�mC֜K��͎N@�u9
�'C�P��f͈��Aa�S5��y�'�b9E�uz�r��72{���'�`y{�eͺv�2P
1GB�	�'��!�Ȇf]>|Ȧ$��^ր�3	�'t|����W�hx��G;EU�{�'i8�81G*e!:y�HK���X*�'�>�*u�9B�Hѣ߼3���'8ڝsg�Y_p�h�	�.��AJ
�'v@�
vgS��I�Ǣ2,;�s�'��r���u ����!7R���'���9�ҷm����ȟC��x�'��dsǂ��q��T�@·A*�Ia�'s*)c(HHh����m���z�'����+�f1�%�R*
�!�'���' p!e�P�Rꔤ2�㙨�y��B!G���Rj��M�}4㍃�y��^�8�diU�S�LQJQ�p�S��yr��*k����AD���F��Q�ͩ�y2�0U�BH[Ȕ�X<D���nO��y���a?܈�c"%2�h�LF�yB�I�Sj^48 ۿ, �	��EZ��y��� �|�y��mY��H��yÍ�#\Az�Mİj[P���ƭ�ybe��y��gϠ�At����y��̌FP���.d�J#��4�y"�5:�dM2r@ݡk2�����y�c\!|�
�9慘�"#Ȏ��y2Ȅ� a�Q�]K$�9�'P����{X�ps0,T5<5�)�2��2��4
�.D�,���^�cl.q���:�B���:D�@��B�V'0� �cw,!�6D�(�%Bغl���Q�\%���5D�� �Ƨe�ړ̓��\��$.D��Z���(}q���h�y+`���*D�$4�&Cg8�ի��B�QE�;D�$(W�J��kˡH�4�cdB&D�ԛbH���0󮊿C5
�K��>D���d+��g
�Y&ǱP���&
<D��Bm�J��ḃ��HN��/'D��JE)� v��I��l�T\5��%D�DP)�+��a�B�A��� j"D�X���}�6L0�L(��L-D� AjN|J~�S��"'B�qa�,D�48���zuR�RQbS�^�����(D��  Y:E,���4Y!��7u�z���"OI�&�W�V �bjH�+��� �"O}��͔�!��y��kU.	���kA"O�H�fm�(+�N���)Sy��"O�tqF.�=O�p�����[��tI3"O�,	���;^��Gn��ȕ�W"O�9����ٔ�T/4Z �ے"O1D�P��f�����?���0""O���,��n	,K�'E�d��}Q�"O~Iq[��B��U���`�"O�}Q�Ȅ0o�j\�5́�h*n� "O4EB�Ɩ���I��Q�o����"O�P"�n� ��������"O @hՁ)H�\]��i��:p\[�"O��(���%3��葨$\�h�"Op�+�*]�6�Ԫe\�"�>%��"O?f�v9b�I�[c�Ҁ�!��~V�@q�ƧCQl�p�N�>!��=PZ�Q�W�� � ���M��!�Y�`M pꧠ�{a��v�S�p�!�d�*�����*M
YQVt2׌ǰW!�ܘn�(mb�H����a�?!�dĨ
Zⅺ��H�*sڬ�%��^!�$�5:ž�7c�-Ql4���xY!�U�M�ve����.2Tz�.@�3E!�D�G��݉t"L�r�$D�s܍(U!�Đ `n$l���ʆ��
��¨X6!��ѴSx� !�+֕6�|x�d�7!��O�9o����L�-�\��AD�J!�D�5ڢ�d�; ˒�q&/Q�!���[�A���'��q"�GB�n<!�d�'\W�a�S�/t���q�U�v}!��0j[��h�S�u�T���X�A�!�ć6nZ�YI�˕7G�B�`1�S�h�!�䙣KzE��ʸ�9{ȓ�,�!�QWT�0a�i^�h稰
!	�d!�D�y��$�u��D��!�š��5+!�$�~G��1&�ٴ �Sn+K!�Ă�>�Bػ`H�g�F1`"��9<�!�>d�P`�.E�60s�mYC�!�[/4^�7�% l^� �̋�!�!�K{���"�U�s��5ZWL�q9!�d�9���8V�ܷp����v�G�!"!�$D�j�&�� �#�	@!�A�cр�
��˲#����g�4�!�D��/����n	q||�$��#�!�DO�m}�`A�.�1r�k$(�	�!�ėK��ч#Y+T��(;S ��op!���p�P�XDj��A�Be{��_�F�!�$�q�&D��!L9>�!u·!�!��Ş�yC���-B�M]�~�!�$Ų�0 t��-0���p
	9v!���2j�X�v��VxR�/o!���n^�|x#��V8xB��3E!�$�&W"��Ru`ךZ��H�K�#}�!�$K3+ ��.e~.�Sw@�\'h-��'��X��+^�J��V`Y���'j\��`�qA���K2�a�'�"�C��ċH�"�CG��'5��h��'�r�c�\-
�(����E�(�~�:�'��J�c��~]�A@'�ˁ0A����'1�Rv�ϟ:��#�^ƐY��';n�:b�K�Րr
 =~�P!�'4�H�@Y�|�e�q��)&�<�	��� �p���,���P`	;1����"OD8YӁU�+&��12��IB��B�"O�I��M۲-T^��b�GA����"O���>]y�P�&��
�"O�]����m��=�%�Y�t���"O X�'#cB�0�T�߬h�+�"O�:2�Q �ƨ+s��*8�� "O|����*%�V�J�,�8�����"O�X0�S�D֮�ʱ.M�P:v�Ѱ"O,�0��Nc�x�'�F�c9n} q"O̝%KY�7@[�d�<]�`|Av"O��*q΂��))e�C�v�
���"O�! ��� ��Q���2�&@Z�"Oz�p[R��8��8�j��۝�y���l���l��}�61�D��yBN�$Z㚴��g�M����CC�5�y2Ʈ+\͉�
�}�8hp�H��y��Z���Xa�w3>t#�R��y�O�k�.� �&I��I��y2�У^BV1�W�K��L��a���y�J�" j����K���@kҮ�yrJL?8���04c�9om�U��!ڹ�yrNZ
_5��eY"mc h;uB�3�y��.�X B�ek�+�iH)�y"Cժ<���q��iuh:�y�DXrDZ� �l�1o�T�15��yB��
^�Е�`��0u�4�%�yR��8����dD�b�	;�N�o�<q��-��#��E��"�CD�m�<��M�Lnh��\�"*�8���a�<	G/G����1�g���8)��F�<�aJ�+ ��H5���J��C�B�<4��%Z���� d�)X(��ȓ2��؋�	9]�YA�J��x���C:y����(G�	��hĽsf�ȓ`���f�5N���N;@<��6�>�UH�!S�<c�7hT�y�ȓ��X� G���U���|� �ȓpiޑCC����!��
8��4�ȓ6��E��(���ZP���ȓ$9V�{�R8��}�	[[:�ȓLy����&nĠ(�O�1p.�x�ȓ!��r���a�D���r]&h�ȓ(Z�z `��f�E(寏.g9`@��z���t�I�jr��+F��)KX,��7�b�`�GY�`E$�3����g�q��g�%�f��>�FA��䗉m_��ȓS \y�� �O�t�;6�͈I���ȓeB$2���)e8$k����^��L��!�v%�׏�=;�-"P� jMƙ��V�T)��M�jo0!�"�� =���ȓ4���"P����R���>d���cl�"��H�Zy�Rm� r�Fe�ȓ(<���l�2e�6p�c�e�$���f�����S9w�X8@"e� 8���ȓIЂ]��Ć�~��S"J�@����\BѢD�8�h`�Te��u$$�ȓ,�Z�(u�54�m�ɞ�x�\��R��{�ކ�����E �轇ȓ*��ԧZ�)#$t`�H�op�u�ȓf�j����$3�� 0%A'*�ȓ}F����l��k��K����&|D��>�0m�W%�4;�m��MמIc>�� }�0 �
b�����T47�l ��S�? &dR���TQ���['hb�"OL,S�)ͭD+�� B厣m��q"O	A�M�s ��Xԃč�ܑ�"O�\k@�d��(�a�ҭ�����"O���׆�!��� Bߜ �<�I�"O`�!�kK d���b`��$i��"On%F+N�c,MC�A/�숒"O�d��'H�R��SJ2.�F$S�"O���oH����Ö�U�<MS�"O@=*�oE� ��d���a����"O �&퉄�fL�N�z�^lp�"O}�r��:��r��V�����"O���S/�d���ycg��@��	%"O~A1���?6��E:�&I�
Ȧ��"O�BH��d��Ψ�(�C$D��00#����y��[�7���W�"D���� �,Y���$�v��F!D�0��B�4I4�S5M�5F�Uc,?D�0�5� ���8�K�?<@Ԓ�D;D���'$@�M�lxX$.H�xP�S�:D��Aნ�k2�)U�E�\�'�9D��+���z����]6D�@��Ս3D���}�4��vg�
lD��@l3D����n��첇�D.ypJ�P�.D����dV�6ٖ�q�ͱ"+Da�� D�TP��K�u1��˽sB�:�e=D�hi�j3{���j��T%��,ZB�8D�h�+$S+
(g�T�i�|��&a#D�|K`�S#S���pe QTn�d;D�̘��һZ�U-�	�Nyj6�7D�����`������]�A�,�E7D�D�	�6/(H"7��9t^�e�2D��0Aü^{|��4��E��
�b1D���S X�>%x E�E~<�gD1D��!տd^Ejv뇅Fp,�(ց.D�(X����ƽz���O��<iW�)D���v*�&w�lEp$G��3��:�#D�@ Pȏ�����/ɻL��q��D>D���B�A�������
d���E:D���S�U�0q�,p�I�m𬔠��*D�LH���~sH�!��C<V�4#�-)D��[抋�o�����_7)��+#'(D�`yc���W�LI�� ��v�7�2D�H�p�09$n�`����^5���0D���O�1fL&�A!��?�|t+F.D�م@@:@>.Q6%Y]@�p�9D�`��"� ����%A�k�8D�T�f��t�� y��T	� D{ �6D�<[2)�	,���#A �_�Pb�+6D��Cs��y���A#_Q?�|�%�?D�|���&	z�I��MT��(=D����NT��SqەvlT��(D���roS5����u/X�Vw����d'D�ԩ�$�6"u.E�3��|PYx�@)D����&Ԅ�j�@O,"�at�,D�P��M�e�<��&�7x��`�&@+D��xJ�"yZH���
*x�v�-D��!��q�|%���+E�����S\�<)�oT�t�������)}k8��Q [r�<�2	%FP1��ѩ��q�<�V��
��5��lW S��P0�-S�<����8x�e�@
&p/&X#�H@u�<93X�/I�}� ���H�p�<QF(�F�@6h~�ꀧ`�<� 帀�7V��5�P'X�@�����"O�d��Cɉ:5��[��C,&�ʥ��"O�( ����]g����̞4@���q"O�D��N+:��ׄ�x_L\P"O�wJ�4蜠�7Đ$��TJ2"O�7,\$k.N�j⢔�~���"O����a�'2�y��Ń̤��"Or��B�-xL�A�*��8��"O�QS3���G�IQQ`\%���w"O� �#*�OY�A���{�"O*�I����T��$��,��rp"OB�RO�e=�4���@�X�Tȣ7"O(��j�62�09�,��6*J�*b"O�b�#N7a��T�0̀S�,@0"O��)���q�F���T�
��'"O���@�:k� �ӀVð�	"O��I�ʀ<P4F��!�/��%�"O�@�B�W�	V�@�EI�T��!�"Om ����0�.͹��L'Ijp�6"O���d��z.�+?4\��@�"O�X���]��z��fʍ�� ]P�"Ou�D�U����iS�XH���02"O��a0�C� �-3���-	��f"OZ��ѭ߰|�iwZ�H�tq�T"Ox9	k�
--L�1g�%>|��"O�4Ҁ�����bB�Oz�ӱ"O$���+!��Cȑ_hJ ��"O��q�ʆ�x�⩋g�]>XW�EK�"O�����4y�e�G�1JҰ"O���W��'�D\��љ���I6"O��J�D�kZ��˧#���Q"7"O�M��?�")��A�L�9�7"OV���eEo�(d��N/��A�"On0�"�
1 !�wB"X H�i�"OV"�GK�Y�@)v���8r�)!"O�ɈRa��]t��� J�ȡ12"O #/�5���V1��T"O �0CΓ"U�8 ��"n.�0�"OLMPq&T$�!�'>a �}�4"O�H1�µG��,�R�YA����"O���搖gS�a�OF!�rň
�'����r����@r'�ٶi�(�
�']�|����0Bn8��e�\]!��+	�'�ƍR@*��h@A�Ԋ�:R�lY��'�8c�ƳY�J5�t�P�Kb|iJ�'�z���fS�nl4BN���'��1���7�Ez�%��3n
<8	�'��DyeaC�7'v�D=d*`R�'g�|8�D��1�2M����/Ddݘ�'�lX�Ri��>@� �k�\��-��'�0��������9ԩW�h���'���1/�p`L����*�jt��'>��d�.'����Q/��'�X���'K�d�Q�:@�`�x�A��j�#�'�!� CY�YIN�K��;|^ \s�'Lv��vjۘM=s��L�Ը�s
�'%��D#_�e�v5�@�\�i�<��	�'�PI��Ւ_���"0 ��8V���
�'��H ��u��U��^<4B�@�'-��"N�N^麆��������'+0��d�V�*Cl����O������'N�u�� � u<X��c�z�h��'ߔ��=@�P	�ÊN�����'}�M�o��5��\y#����y���� ����E	�Tݻ�։��"O�``tʍ&$�0���b����"O�uAǃ� �|�i���������"Od�r6L�`��mׄHa"OEp�g�5w�"8G�ǈMȦ�p�I���*W�$d��'c�W?���(Q�P���5D�+\x��"��7M�%R��?���*��=萣�7e���;FC��Xpݢ��$����L�]X�U�Q���Ig�H�Qr�G�E�ʬ�ql� ]�0��OU�2G��#���0��xaÊ^�'T�T��y��F�r���ħ~R�,Ӆ{�8��e�G$�.�B��)"�DM�KV,�,�ІM`��ߚZO�|®b�ޔn�Ҧ�qP�U�)��g_�/}��0�-����cS�8��l�	ܟD�O��Yc��'&�i0Z)U��%���*uc�	 <A��b'��s�*4`[����b�
QE��XF#��0��˧��Yc�fdz��Q\=�IXtDK:	7�e��4egJ�k­�,:�f�`$c&w�hgfź)��t��/ŌCu�s�q�Ծzn�+p�=:�r��'�?��in���#|nZ�"�8e�p�V�;#Ҩ@q��7��	ϟ\���~�CƧ��F 9:��P$����'?�e��!n�w�I�?ͬ;lϬ�j2�ĳ'�z�*�� �1����'NB�z�^!9q�'�2�'�2�a�����]��l�`bmѕ���#��<���B�j��<ar�W
UМD3Q/��a��\���(���+�o�	 "�B�+����B�㔎�Tv����n�0��;ግ<J��!鵡�~��ǐ^:�K�΄v}BJ\*h�T�Ꮓc�q�qb��������O �$MǺ�O,!�e*�>-)�	S9B�B
O�6�R�`��XR�L�/u���
�'D�I9.��4kU�f�|�O��$X�l��l׉d����芪p4j= �!*'���S4D��H�	՟���[-������I*�P�����?K����%܅j�l�[����'4�|���"&%��E�Y9R�L3�e%ʓ3#�����Vv��H�@�`�H^*$�؈xcb
�H��tʇ�Y��u1N ʓ���	1I��!�ԣ����2e�`U ��M������Ot�ʧf�.�q�W�,���䪋�-��/Vj2�_�8\E���Q)|�!�b�'��7�W�Օ'a�	�!�y�j�d�O��'�<9) �8j`��!Ԧ4�T2�G	T��'{�85�<�!��e��ꢇX<mv�;S슒A���R��h}���`��#u0�i��IF�H *� �Qtz�$N8uc�`pdLF�Q��(I3K+r�q�i E� �`fj�Y�N�&�L��,�O�lZ*��'�M�g��"�~hS�Gq��0��G
z����?��>)CO���u�'�� �H��QK�_��(��|j1�is�6�f��H��F>o��	���]�H���O�|(s������͟8�O�N=���'R�i'N�����s(l0��R�!d�}�w��EdRhP���c������C^n8i�@�Dv*ʧ��Yc]�T��Q�T��A��-����4l[
�eL��8��t ��L�+����
~�)�}��&���×j>^15�G�D�&�o��8<F�D릍�(O���sӖ�J��n��"s�A<�f����Ol���<���T>�y&�L�{�H���m�M��5�n���Lp���Ot��yݹb�Ų!~,��%�E9f R	������=����?   �      Ĵ���	��Z$�t)�;-�����@}"�ײK*<ac�ʄ��	ڤ´�xbjR��7�	'3��z0�J�D�z��`�>>fl�r�(�bi-�=��/�u'� L��$��iW8��I�K�OF�	�ΏN2ƕ+5�e�]H�
׽7��-O�5�Pő�oج�O��0��E��ؼYW��d(5�FWM���b����N$Q<m!��F0�剟,A��	T�;3s��-�h�����(��y��m��� �3*վ�K"�
~��43H>A�-X�Zм\3D�Tو$5+�6��H��۵ba�`�<O��5bH���$��|�#�?\����$��%K#��"���"�#�'�
�ዋQ}���ݟ�ÆI]�	e2�G�ii�=[ ��gupE;�f�9��W�?9b�'A�	�G����9O� ����*r>���AC��`b�#�Oì����Ì����@H�;��|�/5L�ͺ�o��<Y7�ש}r�@3ٜ��E3�c����+�F<
��OY���0�'
��g�4W鶡`�ٽV9�i�FO��lt-'����d�2lF���y2�/m��9�I4���a�*�� ���%2*t7M��<�ר�>���g���X��聨-OG�^T$��2e�k����랳S �a���#J�O(9�ī[C���	�� ��B [4K*�P�;���=((}�'�d���,~B0\�`	�S"��!D�<a�,���F�����
4��(RUD���,>h+OX���^�nāb!'�����D�hF� � Z0h�6q�I�֩U0��F�DJ���U�<���%,l�@�؁&&N=�a�X��6͍y��%{���(N$tQ�IM��P�w�O����T�O$i��45I��80�˔X$��BXh[p �=� L3Q~�'j�a�e%-^�M��FHǈ(	�O��J���Ғ�O`��� \�DP�Vp�tX�"O����	�  �����I_�'Eи�H���Y�JTYq	�f��'�~b�Qg�0%�0@,��&̶���hO�N[~�HYI�P����R1%	:l�����D��}��-m�֟��	T��CJ��'q$a���-��8��$.٬�Ȕ�`ӂ����6��%������Q3c[p���	��`������?Qj�(��?0eD�Ą����cJ�q~RA�bP�04X�됿/6� Y�Ƕ|�3�ӸJ���� P   �  �  o"  L-  �7  >B  �H  �N   U  �_  Ck  ct  �z  �  1�  r�  ��  ��  �   `� u�	����Zv)C�'ll\�0�Kz+�D:}"a�ئ�pgm�|"��f��Aj�
�����N�2	l�bi��s�5���0� R�M�g�Ԙ)��UǺsI�����C�
��&����!z��5�Z�hqn��eK�I���4��}Y��_�y�ڴ�����Zw�����O*⅖�v���3CN�`3����>|���\��P��'�r��b��A;��9�{ӪX����Op�D�O���Oԉ�7�\-6ei��j@T�������O������ٴ���O�`r��(�$�O���a
�Px�D����e)�;��O~�$�<����?���W�΄l��ܝ�� ݎR?v�Pb�I3z=8'Qx���B�V'f���P�sS�D֡}�h8!����26>�Xhu�ܖgv�r5l�7Ϧ���>��'��O�25ԯ-�x����r�Ъ��&k�5�DfG�P����'H�O6�$�OZPo��D��ȟ��	^�t<��`a4wU4eP�ݾ^�x���'�$7�B¦A�ߴHٛ�'Qt7m߈+/ro���q{���>$�	6��?k�j�E��
i�p�`��dG��� U�ߵs4n�*�Je�r�lz�eJ$�\7���*��ǉN\|��I&(�t;�
�,>�\��7Ğ���4?ߛ��O^���N��=3��B<@t9q�W�<�n̋!���y)�F�G(�n����xi�@��$zT�r�֢I7-�ئMR�4����KūM�>0�.�(C􀀹EA�w���:�L� ��~�^Ul�^@@�{Vg �u�F٠�́
���QN�n�H@MGK�tu��G�;�RQ'���t��ܴ:x�AeӪ� `G� _5JX�V�X�@��(&'� *������̇��u���cوwbp�쵩��]�"t��G�2��ڦ��Ol㟨3�����*�D�z�I�~B��'G�-��D�OP�m��?��� Uˬ��%I��*zR�'Z��(�R m����ذ����t�'��'��'F2N�Y"P��"m�-"�7ͅ ����#ҧkNm�ed ���0�4O��R�l���*�hkӚ��%҆F������Ă~u�$i�"F�U����D's�I��D�<���a�=J.b�q��3U���'
��|b�'9RS�d�	:p�h��夔�y�� �Ҫ[���q�	ӟ8bp��SRD&���"�MϧQB-]2��c1j�4g��E[����?�-O*}K��������n���yg�%q�p�t*]TB���ӪV��?�G� my&��+�����i�����IP��.h���`�� �m��.�� �O@)��l�"b4����O�y�H �Q�#�V����	$唑[r������?�Cҕ�����O�%n��H����_ͪYK�nЌ~Z���h�Ft��O����O��D�<ю��LS�f;�+T�õ��*���hO���ȦCܴ�?)�ix�:Aj���V9�)�/�;5\
7��O�ʓCh(�'�?����?�(O֬*c�=Fr��g�M�ŀq-D�Z�I\�h�6�a��r1�\s*�p��d�-_���T/�K���l��y���]x��i#'�-q��EarL�5h��˧U�"��u���p��25�:0����Q넍 a��M5^��B'��O �I:&�,c�(�>d�q2&o�� �C�����IdyR�'���w�Q"���&$t��C���P�����䟐��4]3�Ɯ|�O��T��y"�>qJyʁ���r���+�/�"�� u���I՟��I��u'�'~B�'.>�#��[�Q�М��i� ���3v�U��;[�P�%f'<O�]/�N��`Z�,L��u�P0!�x�;`eX�n�1�FY�fG֝S��'4$�S�oH�Fv�5� ǟ�����'V2
�0�DJҦ�K���=�_���HR�,�>UsT��,^�%��XyR�'���{��9#l!P����Q�p�ؓ����?1ְi��Jz���o�S�d�,,��7��O����-�b�ad+Z�EB8�҄θ4$�$�O�����O��d�O`���̈́�Oo�)��"��x6Yc?�h�d���\��]j͡�z )A��T�$|�1mʡ'�Ƥpw&���\8��F	%J	�y�A�Z7wG4�@L�oH�;O>IL	����M��I�'B���ɱW|Ȉ�/O6��3��O�O��/�S�}��8zu(@0M�d�+B�i�T��G{�O(�7Mǣ&�0��q&T�1�8���6nZğ�sߴ��b�erY�T���?]���k9~$VI	~g���Q#L�|���	��؅���)V�������Mf*�;��O��I����8t�* b��C�5���Ǟ�X�WF�k��xc)Q%{S�qRԨY@e\���~�2A?l[�`a�!�p�~T����~�dC�?I�i����b>e",I�_���ӳ�΅3P��)�D�O(�O�#<9�
M��j�X��i�����I�'"ҍ|�Zm�J�I�Fĩ �"I#(��P����*^��C�4�?9���?�F$��T�3��?����?�w�-��.��b�]��Z.SQ�pd��
�Ј"���l*JUS'������qO<��S)w�P���� 6��TX�ω�K��
�
��M��]�C*�i��lÄj�|Z4� )y�mϻ�6T �`?:e�w�V]�"�ٴL�y5h��	t�矈���<���;uŴ=�����W�f���h�I�X��ɦ?J�0��?_O��@�.u�^���OF�o�,�M���S��&�'�d�O0哰P�����s_�	rS7!@|	��zGtR��'|"�'9���U��ݟḨ|�2}H��cO�J�Cip�4PC�G<qc�n��($� \:���H�� c%?�`P�47vv%�$H��[7��4(#B����C��D@��2�^=:���u���/D��:7�T�#���3��#gZ:�#B�*�Dܦq&�������i�O~�؁m�9='�!�ѧM1m����A�O&���'p����O��S�UP��(}D$`��f��M� |t��!�{���rJ��|uH!�'�:���dT�`1�mN�-XHx�3CЪY��0�c-ƫGH�A� �TR�9�6�	�$L��d�O��|��R1i@�59X r�F8q���$�t�	y��̣���[�h=�pH��C�a2"I#��s���T��O�Dz�Й_N��p'��F��(���'c�I�qv����C�'O�B���������;���X�D�b�v���?9C��!HR�mS[� ݪ��.�n��p��s��ъU����TX�T��jG'	���=-nbp؇X�^_n�S�j�HA*!ۢ��}v^=���?���eR�e���������c�l9?�QC�����I~�O��Պ/@��T%ö;m������!�D̔3�*]�g�:_Jƈ+2?
ў����HOHI����	|Jp���rd�B����-������o��������	ɟ��	Ƽ��YI�4Ѓ҂���@k����G�RA��4N5� J��Z�1-����䁼U�@� �KZ�D7 �1�JƋ0��lR�Z`��]��%�&���S�ۃ�$ 9�'!���
�+�u� ����YQ�c��v�'�pS�'�1���x �%V��\��d蔄V~��ÙE���0=��(��9Ǩ��k�Q6U��X�������M#4�i��'��T�OV剒q��0���X�½�w, �f��p�����������$�	�H�^wz��'��IS	�N2��P4�h�ެ&�tI��;0��5i`fm�,@���'� 1@��x���S�޲=/���d��RB�����1�����䟕|'��[퉍uz<uJgC�;��e��>Ӵ��o�O�(��ɷ\:�	.ϗ?n�4;n�a�\��D*��[u�8���m۔�AԎ�}�J�OjdnZu�S?0��ܴ�?�����]i;���A�dP'mx�����?�"���?����d�2�MQ�b��Q
<i�wnpӔ�(�I�uΆ]�Ѥ�;�:��Eb=B8(���L�t���� b���ލ��iKΦ�v%ۑNv�i�!��v��`��]6Z����I
{���a�I:v\����M��<Xw!<��C�I2��AG�>�r�#�炥x�d����(A�ؔ{j�%�a�_,� 0�WO(�D��w�<4lҟX��o��O&|I��'���u%\<DJ�[/^#��'GL9� �'�1O�3}R��Z���猃�/I\q��V���$�g;�"|*тC�q^�4���c+�qk	6}B`���?���|��	E�?�1B�lؓv� T�&��K)!�$�?7�V�s�iW(fڲ-ō�w'џ���Ɏ�
�� ��"&�^���L	C��6��Ov���O��EI� �d����O���e�)!�/%i!���G�,
(
��R�H�� C2Zh����8�"b>}�$l����y���5 �4�bVBQYz��O�h�����3q9|�Xf�M��%�FZ?-R⋋�<~�]?n�2�)�E^v)���A���'�4��*�O�c>c��K!��nIh@jȓ�XY����m7D�zf�B�N�b���Lͣrj8�#�#�OR�ęf�����|��V?_H. y5�ӿUS��a!��]JUr�G�Q""�'���'�,�]ʟ��	�|�Oܨ0�V8Y�`�%��ϕH�n�@��L�f)
e@'ߖI��ᩗ��Ӻ[����3E��0�H�C։{�M)�ac�F��E���Dݸ7��e��*�T('�T v&&�P�P��w��l��M�U�L��L�nyT�db����-��!�$R��i�\�C�3|Obc�0�'D$�6��d)�K�P�4.7���ŦM%�����[%�M����?�� WJ�˄�;�>����?���L�����?��OR�H
��E��ց�1a�u�����'0'TI���@:+�&��%ʦN�$��_�'	TA���!��d�":zu2$�c��� ^p�&&(\He�܀H:5{� H[�'��A�b5�'ժ�Jp`�lZl�¦�48����'c@�u�U9^?�<���'�,�����O܈8F��b�-Q@�T��O�
��
�lmx��i���'y��GdNd�ɞD��"�P�^�U���b~���I�ѷ'S�	O(���)6-|�j\Q�T�?��d���X�� �gR�oE�+5d9?��½|�x��L�/-�2�3fM֙%4L����C�Z�b�'0g̕�Uf��
�x劙M��%�'.:�C�ɧ���RRɉ���pŠ�VHB�"OLݹ�f̷35��"�Ɏ�;�0�;1�I�X��$	W^"'�O����d�<���'�b�'���! �) B�'r�'���M�dd���ʔ/E��ҧ��*� �	Cƛ�J��Q�G�Y&z�uCc\>���$T�*�!%ˠ�`�iI65��:6��nhب@#�;i�^�+�˼Wf���B#u��s��%3KØf((λw]�i���"|(�q�^b1kߴI���'e����'(1������yw��#�(�˛"`\�R[��If��D�B��.od5ZS+�s&�����OR���s�4�?)7�i,��O@�$Z>($������>X,�b�)c�>QI�(��L�	���	 �ug�'�<�,�Z�&V�@�ؐ�`F��K�L��݅M���eH!-lظ�%D��p<q��{�? d���+��8��PB�֒�2$�eF�8j�ܽ�2,5��� ��N?`f��퐣�ԒO�n[�f4A�"�Q���=oQ����Ob�=���P,]G�4[��m�(t0��$H��{����F��ų�*{���B�q��'�X7��O ˓Nm���׺i�B�'� �����fY�b� .%���ȷ�'{b�T>(���'��Fڶ&��"�k�w?ٞwOJɛ�` ���x����c�у�,w�TG&�o�ԒԎ^4�.� ��6N.-Kwg,�L��d�~��yr	�O��d
ܦ��	�g,|<�FH;"m f�Rk�n\�'�X`������d\�������T�"t�߅#��� {��hB&腨BQ�e���c��k��馱�'�9�Q�~Ӽ���O�˧I0��s��R���Of}��!�F�_ĩ���?��"T�����G�V>����V���7�gհ4jB�/�����ӗb���W+�|x �X�?�Lmၡ�8A�F�����И����?U[�,��C����7ɞ�4**���*?ٓ�O�d8�'�y���w��	#ꔱ}PV�:Ą|Q�ȓw�PB�d�����Q�T�8��QD{"�'kn#=�tbޞmo¹(�HD&��8�#�.~&���'��'Z*�1�
';�R�',��'��\�l��%З�������.8��h��gÝ^���)£Uv�U�r��D�`(�B���6}z	�#c��]�X�1�%G;TW���gP&9[��ڕh�W\Lʧv�l��m����h�5S�օi3)�!���J�M�ܟ�'E�I��@G{r��\
����a�5q�6y8�º�!��N�tG�0y���1ڱ����'��"=ͧ�?Y.O�����gCڈw˨Z�����G. *�l�$�O��D�O^�D�s��'��C�"��d��,K�:���Vn݇2�i���B0�l��"0��	��8lhT�f �� �B��̽b��!��,[b�mC��0t� H���Ė�cHtɳ#/���흒A��`7�'C"0lȦe�Iny��O��O�x�ƃ�@{�7!%Q�Q8T"*D��FL�G���bTm+Z$RP�(���Ӧ��ܴ��[	Cm����O��	=E28��6'P1�؜� �ʭH����OZ!JP,�O���g>��u�ع3���dG6x���C�u�Z����n���z늛,;�+�-��+�Q���a/D�Y�y{�� ;��g*�5,\��,�,��e��\�"�Ͳ�c�I�Q���d��O���:?�D5@�Č(���&�`+��^\�Ig�t�� �[�t�d�֥l~x�ై,�O6��I�4l����I��Y	�,J�����<	5mտ�?���ԇ��O^�K�'a�*%� ���oA��Ґڕs�'�ZeY���6&l��#��?a�*�{#	_5h�K?���bA�B��z�m[�RT`�8?�"��ؠ��.B(Jx\�ɓgG�`!xɑ�3�D�
>�p����˺[������A?��'7�>̓q�(�$~:(�c$��!,����qS����
��7T��@��+�B�G��$ڧ~u*%��c�6D�V��" �͟ �ISyB��(�x�T�'@��'�r2�8�R����-��i�>�M�%���� ��p��?g���H�O�${�1�qA�hW?�~LO�{�ZD
� ��zdpQ'Ȅ�I�� �$�I���WbF�{�N�����A�x��lВ��"ɇ� N�s��O��$�	q~��[��?���hO쵐�)�7�*<�EN��0y�D2D�T;�F�	4T�h�M�5k�13J�<���i>��Igy"�R' N�#�@��P䂸�����B2Z�a�B����'z"�'>���G�`�����K�%vu��Ɂ�'7�E�,l��iRA�[�q�	a�W�Q�������R���4cg
�WE�5Q��!A���0��:u&9K,��b�/U�3�Q�� �&�����!N�yq%a\�7̌���O��=1���[
/����a�8~f��0b߅@!��̈́ux��-��;H��k�>XR�'��6��O�ʓ���9��t���y)Vp��m��g�l��e ƛ�?��XP0=���?��Oy�����ދV�,���&ʛxg��W�ͽ ��PE!G*G�F�Z�*B�X����S�'����J�p��S'p�켫���3@���5$P�u�f@���?�������U�'.8]����?��O��A0�^V
*dj#��R�� ���|B�'!tb1���P�&l���6�*II��B�A,5���5	_�&�|cm]��?�+O^�LN��=�Iӟ��OP* b��'`�ً�G&7��7���^j���'R�ԴOW
dڶ�9(@7�L�z

ʧ��	�_&��͜�*/N�Sqf4I7�I�"9��:��A�[��A�����~�#u�S�_GN퓀���y�P)O\]b�`�^��I���S�O�lT[���n8�1��뒁P����'p�d{��p���� �B�H���d�O�Gz��C#\���r�E�y��t⓭G�T~R�|�e��fB$����'JR�'H�6�N��@�N�K�X��"NP�#)�00�4������#D%j^1�.����>�~r��'>��P1\D0��3�H����?358�c�}l *��ĥI�GҸ�S�? lR��'V��Y����i@ֈ���'���~�����OZ�=Y5K�.ӼUv��e��AS�N��y"��CȲp�&E�V���dջ��d�����'#剏
IlPQUC�)6�E:�+�L�}1Ъ�^��I����ӟ(Y]w�B�'�)��.Hy�eKΪ@�MC1�@6}PKT�ـ{�(,�vF�-#���lZ�W袐b��ɸ�z���DY�� $��
�+ό�2bn0CJ���ή;���Ϧ=Cq�F�tmQ��j�fT$@��iZ�2�ba�Y4(���j������V?���Iqe <%�ziyb*D�8��]`q�x ��_�b���c�+�$���%�Xeȇ�Ms��?�E�B� �ҥ	��*C�^d�4횓�?���n�\�j���?i�O�ȥ,�0V������i�"�i�ŒY}XP��l֎u`:=��^n�ax�f�'T�6�J0�'�b���d�6zڠ��+5d���QA)x���ٲaC�Y�ў(�F��O�U&��(`���B|Zm[�N�Q�K��'D��cu!�XwM!�LL&�����?�It�����O>9"R*�?A�"���d3(��W8��H�䰡����O�� C �'���a�#�'C�2�ۖM�.(�\Œ&�'_b-ɦW�
T��yy�թ�����G��V����D�C^/�b���R�\y�5���Y�Ɣ'��!�EO3sQ��Kr�ezv�y��~�mO�O�B| ��*�%�����~5�I��D�$0O��Ԁفk���EIh�0�"O"�@W�@��,��a�ۍV��
���:�h���C5�,ۜ1c^<Gy��'R"\�X��B^;�J}��� �����̧Y%>�(�o�75�V5i�#F<�ܫV@���RsHZ|;H@�c�f̧NU����f��D�5�z�i���& ]��/�-H.�!���S��EaRR�y�\b>�A�.N���#PAcҢ������:⒟l�E��O�D#�n�}!�.7�LU��J
�$10��'m�=��"ӧq@@5�B��+O8�Gz�O�RR�DQ�\������"�(�c�O�S���]���	矠�I��ħ���G"sd�S`\!fc����5q���E9R.�e t�X��gP 7�)FyRGV� 1�ܱ`싘q�R��7b3X9�	���J���!�ύ�AQ��e%��Zt6�Ҋ�*%$�X�L�M���˵fؑI��|1�c��L%�����H۴��'#��?�q��֓M��t#�LM* ��4|O�b��q�B�0��ٴg���8Ă0���O4�d�<Q��6�����и6� _��� ��3z�
a:$���@�Ɉ#	$����'w��)AqF�+I��K"G�k�����nW�:�e}D�݁�J���O�h��/8��e�3l0(�*�=D�l82�C�Hr��  �!D4�*��g]�@����i≕F���$�Od�u���X�N��*߈$�Ε�/+��?�O����F݉8�5&/�|�1��2��|*�'X��C�"��gZm:��;dT�����$Q�F�0l�����c��Y�" H" 7�P�/D#��(�h��9�r�'��P��R�J�qD�49(P���Ȁ��}Y��?���Mߡ����)���c&�4?IM^<^���NհZ`Q���e�����՛I�ϧ%H*qӢi��L�`%�RLM�%!���'�J�z��DXɧ�01��O�lㄽ���� ��Q"O±�qc��R#���g�'	Pl3�I� �����4(��QAڇP�=f(�$a��Io����䟸w�<;r)�	�������0ϻ0Gze3�C�$(v������4�=9p��P��a��8��`K�Ḩ��?���DۼH�F-��
�)���� 㐦-fu���ؙ;�H�OO@̧���j�W	n�!�P����)I>��N؟��|�<A��k�^Mj�NM��`(�J�<� +G��z�k�M^/s?n�8 �Iqy@>��|�M>A.��˦��Xv����
_�-�i���?����?q�� _��K;L4s�C%-=�aIboO)  e�FH�]����C̦y�0�J>;�Q������.����⋘ �	#w���!�t�	b�T�X��y��-�M�"��.P�$��h�'Z�*����Rܢ�^�6-4�ȧ���?a��i��#=���ο ��������@�2D��7~!򤔆b��� �8������U�6��'od6-�O�!��h 3�i��'��- �g�y{ִ#�&�C�b�1�'orĕ�D`�'��ϥO#\�K���j��8+bk�
�r��p2��;ń]�5��eXmM!3"y��Ċ�qV�y:4BQ��R��G� Z�XaP^0$�p�R���,��d*�2�2�4h�c�xRe�O�\%�D�E��y��ܛ�@ g��yфK;D���Ԏ��
�����J�@;�`��N7��Z���TD�Ov�Rǥ��(;������E\�֜|B/ĩS^6��O8�D�|ʳ�5�?��EXo
�� ퟷPVfD	�d��?��� �*f�K�,�=HpcTis�I9+���[��l`d�'|���D &o��'u&�P�焰7*��8���;�,�я�iQ��K�I/(�j̀Č�x�	�\P����m�)�g�? p��@O�1A	�p����Y�ll
�"O^Q���:s��QTL�:��8`q��)�h��5{!G�2WyL�I�]:G�@�`F�r��OFq)q�S"��d�O��d�O6�n�k�ؔJ�"6E��M�i!4%����0 H±�ڴ	b��M}̧4nb��*���;2�Ƃ9��-pVl������U��x��FìsL7Ǵ*JDq�Q�܌^�P�OVhU!Q�[��y�%� �����b�D�/����iȔ�v!�5���?-��� ;$1��� ��"D�� {�b�r	�'�m0���>,|����%nI�Ě+O�MGz�O��X��{D��6]�%"�鄛��{��P�Hȡ�������I��D�	5�u��'.�;���i�j��2K�$��Ӥ��p*��̽7F�(B�D
>~��sShC�$�@F~r	.�.��J��e�_���)��(�r�W	Qs<�1��4�{�@�qe�_:p����~�dL����?	3�i��"=���d̑d�Ҡ{a��)/
jT�d��;r!�'%�8sd)��br
\�.��'��7��O>�8 p�藿i�r�'�BQa�9RxMIP<�hS�'��]�b����&�8�Ţ��)��l ���?^X¢��8
ZѨf�z���"MK,�b��1pp,��C,@��Y�G$qE�T��&�(a�G�-��	�W Þ9jhLP���%q1Of\P��'�Z�O^�ˀ�>J����&�.=�V��"O����֍IX쩸��p�ܔ�3�d3��|�p�'r�h���M3 �`cҏ����h�i+uX���z>�:&mN4d��'A�e���
6!%?�P�B��i��
b�n����)�'i�XQ���O`!�	�S�H�D��'����3��Dؙ	��Q2s{�D��l�%f(%�����mh�z�O���$�q�Z^�v�;ҧ���Hʸr�n=+4��fHE��� �y�hP�x���Y`!9YL��� V��OxD�T��tކiq�����9
�`��A�iB��W��8���M���d]��Xɲ$'X<Y����-�8W1O�-���'��0a�,y �[� -�r5k�y��6�0=Q6bz.��X��G�RR���Sښe'��aWn�O�b>c��q�oY�TEh��v&J7�e�Bb'D��XroĨ!Ǫ6Y��h����<�T�)�'%�2飅�ɬwP�P��$w�Ĝ�� �:&b��qӆE� ՚w�q�W�׈r�2qd�L9�$�wH�$�#jζk
�U r�D(2��'�h�Ҷ�'���'�h�k�i�6}u
�0G� bƆ�;�>���8Bo�V��x1�I:}s�h�0��(3:Q�(U?���(�͇|��XB��+�z9�ӧ�7�dU�߇Ta���Iۉ��&���'GB�)Y"�Ҕ��͜(w�@`2uDғe��w���!�A�`� �[B�yz���5�$?��|FP��g'N�̈��� b�``� ��<y�{���ĸ�S>���*Y�?1�I�+|x���Z�RX�em�g��x�������v+.j�
���t�X�O�1��uӡ��ZX�i�6�E?�h�!44O8��}��d�q	�R<�ڢBԙcX��G����'/����a\ *q��C�q
�I)�~��'L�)��;���)��ԪÆf�T,k2J�e�<�U�3Sf<QRa�Jh+f�[V��?1��i>9cE�ycF�Ip� .W�&�ԩP�Y�:i��ɟ�&̘�*����ܟ�	���\w�"��4m��8U���Z��� �́�zZb�I�Ec��0	V��B��؛��?#<�`eXeP:�{뛪<E,a"ЭW�9:��X�ϸX�������*�a+��}[5��
[���ۇ1�t�Kb�D�/�f@�'Bη2DA؃��И�'����<��N���3�Δ�d�B�hh<�#��9�P}KO�<IZ�Ke���?a��i>!��Uy�n�fc��{��2b	���Y�_��ٱ7G�#!���ȗ�'���'_�D�'$R?�@ed��7�PX�i@(𙉥��"��EC�z�䓃b��H��$��D4�h15i7_�L8d$S98�b����H�P����C/�5"`��O�Kp�'�`�@�Ģd���FL�!	0U��'�ўXF|B��"rQ�<��n\Z׶�g���yR�Iu
x�5,�T��� 7����$	Ϧ��I~y�lB;:Ybe����S#3���i�`�w>Zi�$֑wY4��_;# ���O��DA��(	B"��gs�у'�֑M �C`/Q�Ma�}:&�ւ>J4%QBN�+lz�Q���	�M{L�K%F[�.��XA��+V����f�:\"���&�#)h}�6#k{�����	!jll�d�O|c>�X��ĢW$��� N���]`�k�<��g�j�rr�ҨVN�5a�!�;p:ن�I���dڵF\�(@'�m.�ڧ�����I��@��	�A��&?	8 ͞�?����O��y2�ߦf�-;P-ݯ~�����#�j�0�Hy�D�	�O�X9q!�;R���>A��O�Z"�I��s�T�9�Dg����߁���8�ocL�@2���.;�0��Iʸc��S@�|��a�X�`)a�'�)2���?��O�O��)� RH@�$Զ:�V-�����E:$"OTh�e�-�DT�L	�rU��퉨�ȟ��!#�|z��!��~���{G�U�M�8�$�O,��j�Bi����O4���O��I�ORq���T�xEȓ��7u?<����:�� K
<���"�!M
\3b� �㞐"E��k�l�
�H��@��hen��b�x���! ���{�)��F�D�wn�㞔!�Lp���-̯{�)�e3?�џ���k�'��ـ@�
,	!G�Ȋ|8�$�W{!�$�q�t�����|a�,�%�wqr�8��|j���Y�(�0�J�d�Va����Gr:$�jq�zT����O����O��	�O�L��pvnٗK��hjN�QP��kgi_)�� ���žQ��E>D�4E؁J#ʓ5�܄�d�% `]JB�9)����B�/61�����b�W<2AF	�Ѧ.�n��	�A��(ɖ��5
e�$��'&#�p��_�'x���s��&��T㈛) ��Q��)D����N�0~�a
7+ΓR�H���<�p�ip�V�0�aJ�M����?a�O�H�j#,9C+",ȑ������x�¥S��?I��g�0�T�P2dGȤ��H�� wtq�O�zeK#�$)@|y�,X��x�����W���AM��@�j�Q�+�huR��R�H�Q哒(܀AU*|�����,.!ؓO�����'z�7MۦM�	�|���?;*p�P!�8n��\��OK�̳#̟d&�֝H�O���Sb
n6�x�Fm��#s����|"�i>�1�4I ��"�aJ<��k�H�� St����rEg�b�d�O��<���?1��y2+Ŏ(��=ґ�@�V��`�r���~��	��HO�P��cɆ!�X�%�u�hĳd�<�I�x��OI�������W�m�@��[���Z���x�p�n�� #b�J�<���џ0���?���$�?��
�f��	2O݆����3o$AP��4�?�R�^�?���'��l��M�;x'(��#EF�	�U	�_:@�Vi�&@����O�@ٵ�`�T���?���R���y�"�=j5�Ct!٤ KFD�'�0���[���?q����?AP�'7����M�;E��Iv�F�Q���� �`�R�� i�Y�I�&X@���O0 9R&�U���'�r�O�r"NR{^�x �U���s�� u���$���'�.-ڰ�'P���Ue��i���A�UZ��}b���v�Q�u��F|6�}�HbQ@�O��$��%��Sɟ����?���˙�d����V�ۢK�88{�\��x��l޺��I��Xw1B#�O(��ܟ���������ħ<�2��'�+x�Hy`��z�t�ɦB�o�2�M����I�2�IW�-y� ��W� tzvlX�V�DoS�1̓M��kܴx����OB0O��7j����H�ɓ&O`�k$I5Cڰ1�(oӦm������YZ��Mۦ�Oɛ�f����⴩]
I��gk�> ��D����<<V!��Z�K�؀CE��9f���b&d<<E��'��]��I���t-�1GK��A��r��z%��V�'���'���'�2�'��I��Z(e=Pl��@]�٦񕉈��a�	RybZ�T�ICy�[�0U˔4��@D��;gt����O�Ms���?N>���OBA{2�
��"�	��%N*��ӣV����x�'���U��j̇O�@�F�N{Rά$���I̟%���'G��Y�J��W�2cX� K-7�B6-�O���?���?�)O���?U�G*ֿ�(��H�|x�q[W. D�l�Vm\c����2-�j���(D��犖Y�*,`r�3H�4���9D�D(�#V�=����`\�:5 A�b�5D��
��\�MN^K�C��A��PV�3D��I�Û�] h8�Sb�1԰D�C�3��t&�� ��&Φ�!�Sbn-��b@=̶�*e��z`] �BG3 e�՘c��-^F��b��T�3w�h� #��W���g�ĺU8���t�H0H�q E9�T��'%̌8U�-Md½
�a��J����TD΍Y	��2��	(9焄8��!iL�
F\�q����yRp� ��H��d�#cZ9d�P����3MD�s� :'>���O�hAd���A#>�dS$኎7� �$��4`Ha�N2jbl�Q��L�_?��� cf�nڍ2�IP����G��,�=�ǯ�LZ˓�hO��>��"\L�CB�=�����Ƚ8��C�ɸ"�	�4��	C�S�$GĢC�	�7����lΨg�6 2�NP�1k*B䉼v���1K��8bl8�fcS�C2�C�ɔX����I>_�>�B��O�n��C�I�<M�H���I��,ڰk���VC�I�V��Ԩ"�����/:D:C�I
��\�&�Ô`�,�X�mڤ|�NC�I��� �L���q��S�D�VC�GDX��H�N��9 ����LC�	5M� ��Q$娱���^ wZB䉜S��ͨ��B���XT*�)ZVB�)� `m@N�#$��p��KR�,�죔"O ����0�'��6�M�0"O0������m"$��!;a�"OZa!D8l���c]+*X|�'"Od��դT%-�J�zC��j1�"O��y#E����	�l�4HD��"OX�c�<,�����IF��P�"O���q����ա0̝��P���"O�$XR�Ή.��V+1u_̙ٗ"O���g�F 8�*i��	��WV��`T"O����\�h��%c&؇;t�}��"O���&Z���2�R�s����"OX�0s �0S��hr.��3�bH�d"OJ(�Dּ(�@A�ND�M�E��"O�d돨d�x���	m�,=X�"ONyP7!{����k!S�V8��"O���RI&~���:5J��w����"O��jt�N�Ґl����Y�X�iR"OR遡kW%Ay���� Z�i�"O��Zp�!��p{�I�L���"Oh���ϕ�Rn��Ҕ
�F���"O|��6Q��ٳP�ɒ�t|��"O�uy�].�	!�R�$�(��"O��{f�C�im�늿j�r��"O\x��lӻ1��˖)�zR>YX�"O2�+��L�J��q�_!~2�aT"O&�Q@ɞ���)*橐$x���"OJy�Q!\���Saà�HD"Ot-�BŎ4mr�'�_�dAS"O>�e�9G��("�$D?l* ��U"O���&��L���b�O�)m�,hC"O2 s�bW(?�vٻ�c�pbT��"O��	@b'�V�pb��5?X��"O|�
�d�hm��z���>"C�"OX,��o�	�}�G�(�)0"O��#@��<i$�IG'֣gH��y"O�9��	C�v�REE|�X�JE"O.�&�_:�PHw��!l��iU"O�}�ACCB/�` �	�!ߞ00"O��k�㟽(k�s��uvH���"OZQ�&(ބB�>;��;?X����"O�x1�N������3`B�H��Y�S"O�ɐ�$�0d��o*H��O���y� ��@��� �h��`�bڰ�y��%v<��-c�~�!n��y��C<z͊���Sܲ�á�ܐ�yrlW�M���Z�����ⱍ���y򏆐k�Z��Aϭ
�fԨA(�1�yr�D�1o�p*Ā�"q�ѵHC��yR�L�>< �8
z�(uMÂ�y�%ø{��Qz጖;z��u ����y���J�&}�g�vH Q�5(��y�g\�@���� "/���	��y��q�X�hC��^�W$���yb�%;2�@c`�Y)1fѪ6�¸�y��ˣ^.���I�ц꟰�ybbߒI�AzR�^$yX՚�#��y��6m4��"�l��d ���y���|n.�AQ@/\N(��e�/�y�{F� ��R�p�u�V��y�+���Txq*�1W�����MJ��yB�.�0QI`Z�d��{�9�y�D��IpX��m��2bL��$OT��y���6���M0-j��mV��y
� ��3���>2dA/� h���"O|�����=�T� ��� !Z�p��"OT�J1kȍ>+ōYt�z1"O,��� s��$O�F�H��"OĹ��`�P��s�\���"O�ųEev+�tq���ǉNmQ�"O��i�_��]���ִ~�����"O�ыa�	d~%Cb)C>w��H�"Oh�������\�ʣHf
*��E"Op%�1�ݏlո��	� [�thE"O�R0��8P� ���إ\�<�"Ohd)c@�.8����DƁ�-�z��"O����ol�X��6�H<i"O���ao�y�`����tX�3"O�\�f��_62���n�$�b��"O�+4
�4l��x�KJ�A� A��"O�H�@%ˌd$ ��T�B\�=��"Or�(�d�>�L+���F��|��"O]�F]8w�D@8!H�3J5LtIU"O,���ƶV�Q���=�<{"O 9�u�4+��O�+3^`��"O�	(�!"�5#Ԡ��H���3"O�Q3�c��Y���Ce^�.�b�2""O<,�� ;Zm:�rf�
_�����"O�US�o do�d����Ar�p6"O�0�/�*<fH�Ip+ٸT\�y
�"O2	�$e��I��
J�w<b�"O�9R�A�}=Bu�2)#%|m("O��x៍?ݺ��C!�s��&"O�	"焋�@Pʧ�
��L��"O(�@����ɩe� ^6�Y��"O6�
$��/"3�YQ#Kl���"O�٫A�T
%XUsv��)�v!��"Ot��3�Z*QS� �Nݹ� |��"OҰ��->=88Y�B����a;�"O�l	G�N~�\��р9��tC!"O0�Z�怑\ι3��A6Xx��1�"OP�����E�(̫0�YrI0MC�"O�d�bL��'�:U��M�	;d�BB"Oh	�eo�0=i�%���M ��Y0"OЁX�+U�Ge�%c��[��IU"O.�;���fj�`��a��м)4"O>�c�B�*8^�u�w!&����@"Ob9��NύQ6�-�3��B����"O2M����0}
���&��/�`�r�"O�9RAE
J;D�h���
*�8�!�"O��&�Ф)�.��w�	1��U
"O�˲�@&0!v�h��V� ��.�y�'�A���е-~xyk�I��y2�S7<�
���K6�����HT��yr�C�pp� xPk:*�@	�
 
�y2��5eL%Ɂ�]�+�~q	*=�y'�(M�^p��/#� �;Q���y��Q��U�&�)3 .u�����yb��7'��d��!��J%j��yBςKC�$�`�׮N��)����yR��4=K�(E?���'�Ʊ�y���o2����G�	R$���y����ڭ�g�^+8@�䲲!�	�y򧐶0[��Q�/Ɏa��������ybA��6d"��B��Q�����"�y�) ~$���w̑�\�~��d
��y"���4B�@�Q�Y#>g��eb·�yAT���1n1��l�/�y
� L�*qO�{��\#�*ءB|}9�"O���Z'G��j6�'��`;�"O����!ف5�x����K�Np@E"O��%GR�R�6䱱��F�0qK"O|��ABD�Y4�A6cx"���"O�<�"�ݳ{"HrsfR�A9<l(�"O��C�eC(G��Y��="1� kb"O�Y�@"�;H�$8��$�5q!B��"O�-"���
n�~dS��"G��	B"O4����7������8{�=�"OZ�Rv����)�Ӫs�1��"O���g��Os||���D�{
���"O10��֦Ϙ�p�ȁ�Ƞ�"Oh8#��ɯ91����EP�V���"O2(�����De��@_V�ؑ��"Or5ʑl��0���Z'�P1n�RD��"O 	�(	5WJ�y�"�[�.�@�"O`ؤ�G�w�i��".Ad40�"O�bE�R�t�@+�"��@�tݩC"O�qӷ�4o�p�x (�7+��b&"O��b	�e�q6MA�_$ S�"O����HךSx\4�+�r�"O~E���ID���K�`Qz�"O��S�i֤1���*M�F��p"O�t�K�j�X ���RX#�"O.Q��	L"h�OגF����F"ON����i}�����ν<ܮ��"O�xrA�d�8��F-Vw1�y�G"O�8��g�=^]�*P�)�貲"O;������W���"O�I���'r'b�C#�
�I�D��#"Op����z�S7Ɔ�A�)GD!�$T�ڼ�쀵M��ёʜ1<!�׮T΂�"���;{����C�L(!�6e+X�@�� �\���u�!���Q�P�Ł�^�Ԅ�dG�B�!�H��ؑB���>���V!�Ď�>��`��x�h)�Oʰ[�!�$U�f�`��&`��9~�����?!�$��wxB�J
�xcv��H��UT!�Ğ00�� #ԃ	����E��UH!�DɸvH@TR$���O���䑊-H!�L?�pL�A���^h�d�=[!���)uk�`�	޼�0�5cخa!�` z�(��C��ނ@^!�DZ�^_�����@4�B�!�D���|���lK[�PՇʯ�!�DP������5����e�ߑx�!��&[�X)X&��Uk�Ф֨L�!�D³/�HTRҡ<W2Ɋ���� �!���"��сB֝X_8=��Ȝ�(�!�$B�l?�-i�'T��	ӇA�Z|!�$�
fg�����*9Y���v��F]!��X�z%�,2U��6_!B��SH!�$��*���V���G/LX!��t%�1���?$����AW�!���.g\�*�"J�|"�X��Ώ �qO,�sE�O s���9�^�6:�Ò|��k}"�cЍ �`�&;��y�+�mPdk#M'�`aat�Ԝ�y��P�!#���}w"�,�����'ʼB�wR��Ig�

	�n���'�Q�&� #$����fb���p+�'BɊu��seRq	Q�Q�k�|��'>�@B�F�^�
�s ������� Y��E��<8���5&X���"Oʨ����0�xY1���	ji����"O&9�`��G�j���A��Z_b�Y�"O`�P�j��)���*�"�)rm6��c"O�� cE ��7��+j����"O������sr)j�N5jeּ{�"O TQ���%ih��3�ZSG̳W"O�Y(aϞ��P��AعE `AS"O��T-�GY)ȥ���F���e"O�� 1������e"X�dP�r"O"��,n����� �"	��"O�4S�^=�|8�ME�,�4��V@#5
`em�"�>�i����5�
�'������"vZ�+4��=��+�O��"$�O�P�QB'C�lQ��¤*I�i�����	4����a�:l���I�K��<�C��'r�*P�	4U�4"=����5L9e�'D�#n���� �����^���6h� �40�a�
I�DB�I%O��0Rs�!LD���Ɍ��͖f*�!��(T�0��fٞ�MG�\c�bex�)M+�J�r��N,;�C
�'0܍�Bi�6E|ɘp�ߵ��,{�ŨM�F6��?9S����鄸%O��&�O0DÃ��p5�<(�jRs%�<���'��\x4�H8P����0>�����a?fxJ@��+F�X
,ᗣQ�+\F��@j ����ğ$v�-��`7 ��$%0�P��g�_2{p\h4�c��iI*Hqy�@�]a�������̈́����C��Q���.+�t�s�GV�wR�oZ�
���g��>=n�����P�3GD�����ν����,�Dlh�(s����I�3�� �a�S�>�4�tͅ0�:�A�)"����`P�.W\� a�
4.���%j�~���I	i�D�	EN@|�a��>_ ���bD�de�S�(}���ƀ.@��dHT��(A9V*��*W���s��?-�LZ��#%��vI%�O���T2���Vj�))��2�8O@T#���>)%����)CIb�� <�	I�My�$��`C����I�na|R���� u�Ԯ�|e���g
_4�)R��ؠ|ԢH(W�*�֡�A�uK��C%��2e�����Ʀ�y%K�0a��i֦E���Q����!J�L�B�$6�����G�d��q�Ck�kQ�1�`��O�t�C2`
79t�	�MI�����8�Fx"��+?:��*AH0^��U�7��79"���+�R���1'M��x���T�� ����[���VU�2�P�$i� 	�H@�!a�/�P4*�'����˗&pp0��9wP�Z�4W�\u�6�.B�F�8�
<����B�ou>�X�`��7.\h��Dn��<�B�7lO�
�G�g؈�H�`јE�q:�ڻK(@��"G;D&�Z`E�C�*����l�r��El�e��qG�$���s��<S�H	�'� X�w�]z \c��`ӏ(V�\i�Deܞ��}� �Ҏl,����Ĉ��r���O��L�.����E�,�y�4$8<�i�O�b"<�CE9=�l�'�K>�@ ��A��Z�T���i�6<���ҦiR��ѿlZ���S�cs�/*��!�Iзg����4�C�#��<���T.R��d��5̉!c�Q�~G�h�R�X2���Črf�sL��n���#�e���L��OZ:�(Գ��D?�b\�CϿ#��5{�CI�a|R�ɳ]�D�G���\ �wJ�Lʊ�!��U�>�|Rs�gt�ˢ�-kZ$��!�UG�"~B�gGc\|���
���I*� P�`v� ��ޮdF��!�C���%?y��d�\��!�*blġ	�厧xo�9B��>®�#�N�0���'_����>��!�9�dxc���$E��7�B6���	+G�!+f�Nޟ���<?���I#�r�����|�Gh�+'�$y�Y��ɸ���
0��p��Q�g
 �Fx�O2���'��]Rr���T�n���Ð,Ӣ�*E�5�iJc��y��`>F�ܴ5Y�0��ϳs$����_y�Fl�<���O.9PFmZ�<�x°����Xƶ�cg\��m�7O�!�ah�>Q�F�O��'zD���ԇ6�z��o�+��ñ'-{�4�͋9��5����\��Д'��M$��Y��А`��n���y�I�!i�I� �(-P�p��8��I䟠X�%00>�2�+)�E�=��Ή#���z5�ǆ.�BE*�d���O���P@ٰu����a�S�T��2�B��Y2~�(�87썜;�Z�(�%�}@�$�C�T>Q:uf�;y�*�ds�� �Y���8���G�����dc�(����H��n"K>vl���%T�8j�䞔j��
��esШ�iU2L@`�׮��gy�HU�g������e�����'�/��C�c�qO�ß'K�䋁�_�6����O�C�ูgI�N6L��E��f��U:P��;X��$<ٴYj����	�G��Og�R��`~�I�̈́6qs�,O���#�O�%��!
��Í}����Qҥ�;=��)�X5E����d���	�*
��������-Kz����Cm̤W�lLZW N��M�G�Br��"<ͧq^x�5aM!x��l�޴P���J�J1S�\�P�FΖK�)!���$��1Q�T>���N(�{�? �5���U��5��
�P�R]B��>i$́5p!����nO�&������O��*tl��R�z-H��ĿlJN��b]���(�S�(;A���e0
��$����
�?g�5��j|����
uοsf��%�p�]���GT��N`;&��7C;��+��)������#"�|1�K�^8��Ғe�!�����]/of��%͓;mن����+���i�|R<�єix��8�F��yô�6;�`<@�H�'f���{G`=D�X�g�f�I	R/*;wG�}�6H9��U!��!����S7�0��c��s^\�dIi��j�,�;
�,)���qDRi��lU�~�2	�<��dE�>2���"�'e�����@-e����L�?M�n����JD�SNS�����@��	,]��������O��X��Ύyz��y�H#_��`!>����{�d��4��̈́}�a蛅�x����4|f�IEJ��٫�����aR��t�f�Yr�51(��C2�?I�b���M�"�%6�ȸQ�H=)�����۟��ȡ1�+�z����3���V_���"Or1bs�ДEnqa��5x��"%v��MX��&�:�[��A����C��� ��P�w�!��h��)��� ���y���hM0��A�/GkXh F��|ى� K;:���s���V��[v��A5��"��Ml-�E�6�O�m``��~B	����-�7��>3o�<�0��y������ل���h���>F
�i�y���^��b�wj� )�*9�$e�0�C�0��'��A2�.$M̅jP�R�T� d0�c�>yL>�;��$���9*�<8� lN"B��m�E��o����$[������~�!]��)��M*,�p��-��yR�"+_���������XtBrjM�Nؔt�GH��X�u�C@
34�`٨Վ�~&���k���h��"0��ne��;HdB䉳P~'�ѾC�܈�7�ʫK�P9��� 0�6M�;Qp1O�'j/.8@�w���i4h	�2O���D h鴸��'��K*�c&h�����@�p�Ҡ�.�$\=���^�!B�3b����' �X�d��!�U��А��=jS�W8�j2�C �MSĒ5�Ʃ"v̘%L��p�1�Me �X@�f�X�R��MKZw� Z1F�#F,`���/�� �Ԩ�W��.Ay�����:���'d�o�n���:�O���7=ܤ���ÄT�����]P�7��$x� |��BB6s���ԥO:Q�8b����fO��"')F��ȃ��v���i��M#�y�O�$�"���H~�-Ȕ=MM0 ��!��:R0_^L����TX���k���l���`"2ŀ�J���>V�d�O����?��4U*���
����Ǿ$�8����ƥG�
e�~8�����"[`³"D�Iz:��҅hӖ�ys�ɧ(.�@QI8��\�'�>6�-Tդ6^�KQ�,���d�E��Ob�I�|Fn��SaO9�2q&јGu�O�4`�\�q�I�����rڴP�b����D~��MW�1���N��.iN7M�=���1�P�7��Hr�-݉.�Q��Y	��y�1Z�n����0���U��+�Ϭ>�4K��Ο�����H�� 4ռ�1 �u��܁E/�*bGA�Uś
�0?��&K&3������[��W�?m�e0'�߯o�\���(� 0������ ��|���O- ���g�c�z�kB*;jjF��ӓ.��4#��զ���:����1tT�F ���ô�Өa8z�xKW�-T �s��L\�O�H�I^����O#�e��"1b�Ĩ3�Xl�S�S%=~xTX� �>I�xhv#L�1U��W�U���ѕ̛�&�µj+A%�Q��r��[>e��YH4��+	��P�qo�
g;��)��IAv�J�[3�9��)�"v��$��Ņ$�(��O� (��#�)7 G_0x����_����"3#��@���"z�5"b�X=d`P(31��-4o�!*��S3��@ 
�s��I1}^3g�"h���&��Kᤄ��	�iCY�!񤁣
 ��@�FTI����A������L=$.�5��D�8�:��f�޾*@4�A�JL3)Z@��G���(���	"d6"�@� &l��9	��<a���$�l��Ar�W���@��^�(P`�6���>�P8%m"+b2@����̡d�_T�DH�����L"@8��$L@�"U@��ǣ�\#.��'��!�D,T*�
$E�j(��y���+�ģ�B�p ��6�B'W��e1ծ�:�������!)�*up�'�>ͳ7i��	�8�8֋R�G�J�"���;&ə�ӫ#=(�xR��Ri�̰1e��i��;ЇJ�g�ʍ#���,[��� ͎b~�ܸ  �;�p=�p�
�$t��Ab�ȭAv��d��1� �ӆ�K�2@a `��%� �-����-�P� ��`���
�Պ�?+\�Ag�O��E��%4��u��I�F�����4Qc��Q*� J�,��b��[ݛ&b�?=�J������(Ӌ�)+9�a���!!��ШCH�r=����+@9&��F��ڨO�-b�.K�
f `�S�o�ڬH���2v�2�٣df�5���Ū4�,a�"S�}��!c�C�/XڭK���h��:��ٙ)�m� B�n&���pc�c�����b�dͩ�O�v&����B<}�Q(�FƼJ$��eo©yH����	�",�̪�C
����S,]��Q)�J�L��dL+
� pqӨQ(6�&ن��0(\4k���i��08&� Zh ����IW������YD�����6b�\h�vAE�>a�i�A^/��h!�ĕ�)�T�����9�`���'���YB�S*�B�i�HZ���mk*O�}A��"I	��K��A�3��և·p$Z)o�75	64��h�"�X�x#(58���%A�k��3���7��P���9�%سb�,czX�>Co�-����,��53�:�&)�@)��|Q��D�Q�0�Ec�"M�����E��<,+�љ��SG����D�"l¬�bwF��a~��¨%�A:�����&"�9FH�q�fO�>��8H��@
)�!d�+g+v����tψ��$&�)"ȱpڴp=�!p�f��$�t��5A���"E�eXў`���|	:\�1IU Fl�I�n�1~� �v�Dɪ�`(ϝ=
NYK�#ףI���B��Bf@r�ڥ쌅t�r<m��U����O�	���p��M�(QF*A#��D�-g �,��`�"d�4���G�)�d�q ��mΆ�$Y~o~�� <��l�dG������ ����d�'��]�$�'g��P�NH#�"\�Av�em
�p��Q�J@2Ca�]�Mn1��'���a!(��pQ�t�$��>+�؅̻}�>HhEI�%d[vlA
� j[�X��I\�l�fiϕO��+�[:*�Ȩb#!��x[B=9�̹�PkAN;Id6-܃S�( �C

�H�c!%��X�I�NG���c�DST�y�kT�S�I',�Ru8fd_/]!��N�#��u�T%M��J�Q�˴�읪�
;Qy��Y�L,e�8Mxw�ƙ* �����unax�c��#�1K�iW������c��7<x�5
�4vtKD ���&�x�g��9cp1J�m_�dD���+~K<�Ӗ� ��jT���So�͠�/H<M)�A��<�x�j��'�=�$���N��e�J`��yTAȃ, 9Ks�|f�y�j��<� ��Tι�;/�N��nFO�L�E�4c�(u��	�7R�̡��ۑS���iX�N|���<�\��"(bӢjօ�6����?¢��e@�n<6����I�R�����\&Xx2yHAg0V�#=�d%K�@�xpje&\Y���1;-�2�"X q�CW�ƱYM��Q�ꐭ�U#Y)Te����
��{��'�<X2!�+�劂�h���#�S2н�%D@�hh���*O?��BLUa�@��e钒p� 9�m�W�<�aX�s�.��`�<�9IB�sy�'�%t��0�,�ONax�D
&�v`I6�Ǘ?b����/��0?�X�d��1;s�q{$��t�ۛZ���PB�ɀs7Bቹ>�p�*��Y�%���Îc
>"?ɀ�F)VN��?��A��vt�+�	j:DDѓ�"D�����J3e6�(��Z&G`���A�<�d�̳���(��i8s$�<%W$�05��\I��J�"O��d΀���\����>gCZ�U"O�qsǣ�
%�"(����@��"O�u)�'S!#vXk��u*��s&"O6�Z���3m�@4
0z�-�&"Olвu�ʹ#�����O�����1"O��ұi�B�|A�IR�J�X�"O��� Q=g�r�%	
�a��t�B"O��@t�ڌ��=�f�J
��\a"O�98 �4[ �0hF����[�"O�|���=@
p('oW�|�6�*D�� d��/�Ҁ�ā��4����H*D�tAW��`�.hۖ���^J5+�7D�t T�v"�Ċ	�� �@��#D�@�CO�O�\�6�S�Tj&�9�.D�43F�4v�̈�T���p�!*D��rs�/a�>���e��~a�y��B5D����)�-KX�1r�	x6�j��1D�1U*L5kB�$�0��	r%���!D�P��䞍^��a�4.�jy� D���� ���2q V+k�4�8�e D�TJb-J|�zԫ#�;m��[��,D����6 &5+��3z,�|(RM5D�t`雿�8��-��kΈ��S�1D�����~P�ړh���:�l?D��d��8X�R���.Ӯwr���F2D��I�aȉP�R�8Qh;�F��J0D��3����F������`y >D�pYS�?����Fe�yC�:D��CB��d�|�ꄐ�ޝ �8D��s�	I�}�le{W�P��a(��$�I8d����S��nZ�Bd/ӫ
�8�O��'���"�F���sc"O��رjG�E��BU�Z?�̙!�"ON|�Hҭ<ܨ���k�`wX�� "O� ��94�o�2� @��s��r�"O�;@'V�:$v���%+�^��F"O��0�_8pY�	�D-G�u����"O�D��(�K��P�ћ#�.��"OhpQaυ(t����Q�<*�j�"O��6�<h�<��'ح'�C"O�%97��'3�dKc�I#`�p���"O�l@b++o�C�B\-Q����"Od���_�I�ڱ��@P<)�*�R�"O�]9u^�{|h2'`�o����"Ox-�eJI2;&s����϶��"OxHkW� mR �Dh9̼@3e"O�@���-���KEG�.|����"O�y(�"Iz�m�I�^���"O���Hϭt��Ȓ��� k���A�"O��铇��.k����C�&���"Of<x��uG��:��ӈ}!��"O4�P���39&�!�h��  bt�"OuJƠ_6[�F�P�ab� 9��"O�u�R	�U����R���Є��"O�yQ��=}1J��
�a�̀��"O���3�ڬ��+N�Ɖ8"Oڥz�șrJ4 Fm��E6��f"O���'įj@��"�#Rv
��"O��#A��=X���`̐�tqT�C�"O"!�ՇJ#\"�i̀P�v�h�"O�i�)!OeR�3b�C*F�B��f"O�Qy�B���.)�ؠw��k�"O����� yѐ"7ټ��"O�$����72���6nK\����"O�͸���Ԣ@��20IR��"O��4�W�MȠ��˙�&`�)K"O��zT�W/�����jU�Ttl��"O�PdmS�Ejei҈�>:Pt�	U"Or-���đb�ʨ2G�q�"OŉW��=���(���q[N��4"O�Ȑp  uY��k�l9$�,8�"O�Jơ�u����+ŕN�6�;"O6��sT��@0xGL՘,�>u�R"O2��p�ߑ��R��8��	4"O�A2��=q�H��`J�.>)�$"OF��/�)K-��Q�$���Ɇ"O�� �c.��ј��F�-�p�3"On	s�b��L���1��t�((�e"O��(O�e���0��
xu�(s�"O"��-E�Z��x{�E�?^;`���"O�Y�%PF����ō��a�"O܄���Õ.<���ʜ�7׬��&"Ol#��GN�tx�c
Z.We�R�"O���è	!}UX;�H��=��m�w"O�4�Ԧ�$�$ ���K9��D8"OZ I��]�[�U9uK�BZVh�"O���R$>2�tQ�穏�A���s"Oj��ፌ�ar�� SIR�46����"O.�Q�Ƀ�)�L�r&�X�d,�"O�(�/<Ad�����\���"O�@���z���[�mֆD�,)�q"O`���yhڢJ�$qa��"O��W� /d��i�cW�W*(y�t"O��;����)��"N�n&�`�D"O�0b�"(�	�bȡ?8�d"O$E��
Q'uʤ:UO��4��"O2�R��	���t�7H�E����@"O6�+�c���,�ӧ��d�����"O� P��c�&y�<�Q���0M"O$�R�dp���6(��� �"O�x��,��p$�B��ҿ� 5K�"O��c� L8���Mw8fI��"O>�!�%&?��Q�BL|��'�8؈R(�$���7B�n���	�'�v��k��A�O�k�6��'�$�*T@�~ղ�`g"�0-6�=Y�'p@��3d	)Pvk�#!X�L��'�aJ�-�)En''���	�'��1I���"�ZDG&��8�
�'�Bb��cl@�R��[�$�`�:
�'HJM�։�4���b��!��h{	�'M�m1q���w�����.#�Pr	�'����kE5yR��!�;�h���'�!Y����vAR����/Fh��'i@P�%��B$�˒$&,�9�'��q3Fķs*PQ��C�#P\r�'p��hw�π/��RC��Fi<	:�'9&��KV�:���!�ΑJWf�
�'���a�aL�a�
�Ġ�"t��]�'�&�!`B��܂a�co��jk�)��'��u�DL<{U�ɫBbX,1؞�K�'�EY�I���3u�Y�q[&���'�J��aǊ�p�����_I	"�';v�R�U��qC$ V�]��j�'��]iFC�;�|�S�X1O	�	�
�'���Q1!�t��SsEӑC�iZ�'x�tsv"�G_lL3s&�%A���'ӎ�{u�Y�J��܃2�ϵ:? �J�'��aG�K
^6�!K�<-Jl��'��,)�C\4@�0�`�єY���*�'ft$S2�G�Hh�8I�1N�f���'njT�А�R1���R���'�$���UFz��B!Ah�
�'.N���i�0W�X#Ǖ;w7�A(�'�|�f��4V��CIk�|��	�'�mÇ��W-��H�f����8	�'w�uxa��5t���b���eJa�'O$�s7�H� 	� �t�
�5�d��'��#�Ɂ�7�D��)[9�v�9�'�>�9AoA�m言�k��er��'����$�՟HIV��Q�]��ta
�'�6y� ���0B!��;XJu�
�'��������� H	�$����	�'qL0����l#r<�@aP�g�x  I<q����X����a��^���3�˯!�d�!H�:q�7>Gv��g��%�!��B��z�N�j1P���%!�Ě7�r\������5�7�#=f!��+fΌ�a�DҚL�����%w`!�d˿]&�L Q�:��w$˶!�!��|��ѩD���:�������C�!�D��t��ha��vx���g�!�B2P���T�3��hJRgV_�!�� Q
L���ѴXR9䀍7:�!�M'��Ps�ؖ?M,��W�C(�!�� .�:AHdƝ	H��U��;}!�D�b��)�5��h���%T!�D����*VI�*�S�3C!��ø`#@\��.$Fh�1K��D!�d� p��Dy�b�)r*�`���Ha!���p^��@3��i���?Y!�D�P�Xj�L�Z�zh1�*�!N!�� |asܼ�t�� �: ��4z�"O0��Õ1�H4�f�{Q�� w"O.my@���+��`E͠p.�1`�"Ol����T�!����	���"O� ���д���3iH�I�(�y$"O<|�h�uD&<�QH�+I�\�"O*�u�ôZ�VD�6�.����p"O�� ��MI��5�^87$��"Ov٠Qb[�V�Hk3LG�TMHa`"O�� Ɋl$@y8��Ь0C���'Cz�3@� j��٪��R8mb�	�'bЌRuŌ�=���E) �U�
�'���)���3�����I&�hH�'M \B�J�x��قMF�C���
�'�h��K�J�j|�R/ �H~� [�'�J�
0���T(��҄V
E�	�'"�xzǎ޴fi~\��O�\�0�		�' E�B�]'e5:��ʮM�̑:�'d̔�3U;n#x��JJZH���'�&l��f�9 �f �TE 5v�Vت�'���K@狹 �R�X�޽kKԼ@
�'0Xّt�?`�^@��ÄQވ
�'=6	�3��_H%��DV�I]J�'���jb
֜�b	�A�Ό7�н��'5�i��](~_��� ��/�",��'8T�rvQ3<�١�@ͭ.t$5��'# `�꜀C�����pb�h�
�'���"c\�A��jF�
$"
�'�~ܰぁ�l%��2�n	a4��'���a��SF�U1!j�7Nr&U��'w�TX�D9 <%���	H�m�
�'�h4FCp~��1!Vc��h�'������i�Jeb�i�-��A�'����C��0��d��JQ5|�h*�'R�% qH�
+�U����t�X|��'�H���.��T	����z��i�
�'O���m�+(�ơZ� X�b:���k.S����$*9W
Մȓ9��P�س Qq@#M�����#�eٸs��98��_3$���ȓ!b��څ�ߦ{K��#�h�깇ȓ/�(�+��Y�(%�[�(		��ȇȓY5�҃�,�||+�d�^�ɆȓV�HY ���7E�h#�#S�7��ȓ^��Ȫ�b�r��Ł�CBLdu���J�4j8Ez�	uE�u;��ȓ���>5�H�"�ϔ���)��=��u:�&�N : �!�O?-�l�ȓ
� �)`mO�)�������͇�Cbdja�lf@sլ7*���ȓ&+�D�Q.J��@1CT�M��ȓ?<n=:���1!8��#�M47Vq��3��@S�ݧy�����C�!��]��T�P����W�}�N�¤!
�,��نȓ`x�ye��#b1V�ڡØ�-��ȓ;,D9�0�Y�y@��:��Y�Q~u�ȓV�N�����Q�z`��M�~��m��aH�y���� �W^nh��BAt����@� ��((V(��>��C#��}~X�[�ƞ"}�*���0��xWJ�/AĊ5+�C�"6u�M�ȓq��1P�K��<l �^p�����s�x��F"I�S��T�@ "~����u>," ,���L�"�K��n��S�? <Q�+Ͳb���1��_G*jx�"OxX��薎����V8>���r�"O�P�	� �4%I��?fut���"OL�	�"�%7�t2�Ɣ:EL|qY�"O@���I^:%��*�Ğ>W�� W"O�
6Ώ�//F��e�x�z���"O����ѠU�"tQ��F�y���5"O�}R2��m�"i��T�Hcq"O6,P&Q,R4nS��כXZ��4"O���b��h=�P���(�"O.tbd�A����
iՖr �D�p"O�9Eǋ�"�t�$�D�2"OX�2G3TZ�P؃��
!P�.�y듃+ ����W�x�1�F߾�y�m��[xz�`��I�$�4��wK��yb�Y�w�x9�0iPgRU'a:�y��_%� Sg�8O3$
(��	�'���c�
Þ��Bф5[F�:	�'B�H���؎ptf��p��*l���'�n\Z*9AZ���ӦK�\I��'<Y��ǘ�B�6�ru���<�\Z
�'hf,�n3c ��!�([7����'� ��p��v�l�!�Ĉ+�'��� �Ю{}��PA�Ұ�*���'<�-ON�cp(�.~�����'�T�3rc�+�84�g,�M�.�:�'"�Ɂ��F\�V��R�4eP�'�|Q@�Q�L�(��ϳ�<���'����e�+gH�@RmɃD����'c�����w#�lb�o�	@��Z�'�r��Е6�tI �X�CST(�'PX�/M�U�4�
Tb�$�@��'�H�	wᙾ{hL�b#B^0$5X-��'W8@DN�Il��wn�k���`�'�����-M
4(ɠ7I,b&�X�'*�XK$��i���fC�-d ��'�HЉ�y��T���s���`�'����Gg��A���]犁��'1va��h�ϼ]�M�L�4Z�'����#I�ۺQ�3�R�zqn��'&Vd���Ҟt� �Zq� ��8T�(�p�ڋlE8qѵ�W�!0�A�"O�](dM#b����eA5h��K�"O�lj��E�]^$���;\�Z4*P"O@�z�����z�m�=���"O�ȓ+Ռn?ԍS�,Y�nj,āB"O���.8��ً��@*{>w"O���⤕90u��򊊜gR�`��"O ,���N�j��I����nO��q"O2qi�C�lM�b��.���p�"O�� "&I����ABQ5$�:1��"O�bWB]g��]��C�b�hİS"O�	�@�!v܂�H��U}��z�"Ov��t)�S%���\V�4I�"O֜�G�s�.�r�W�RG��C�"OVȃD@G`+���WgL:�T�B"OHtR�o�?�������c*R�c�"O��N�l5P�9uo�1k0�C"O&U��ː�=����ӭ-���"O@Ȱ� �L����ךc��	�"O��x�hT�D,���U�{�H�*C"O��*'O�4ZU�v뙵l��v"O����KM^��e�7*�0GD0�"O�a�r'ْ\�̍�AbE�+�B��"O� 
]`6�P#^s��{!�� d�.�94*O���g��)��ى&"ϦY�b"O�|sÂ�@'`!:��G9Y7���6"Of��XM���P�Y0U�p"O� �-ЈM�V$)�j��h�n��"OxA*T���Gp(m�jC09d
�@�"O�Y�%�˭|vT 	�K���Ʌ"O�r��ʅ�\(
#C�8�j�"O��!F�Kzl���*U��Y"OD�1�fe �)t,���p"OԝY4�ƴ��`�͟>�zE��"O�%�ѩ�[��(c�g��Q��3�"O�Pt��V����ߓz",M��"Op��Հp��,�q���O&�r"O��˥D��Xk�M8�uh�r�"OԀ����9�&�0W�XRԄ��"O�m�U��2p(�T	������"OT!j�E@:&����"��Hw0Hs"O���Ԡ�nJ�ǈXv@��F"O~�.eXf�@�%60�Z�˵+	��y��J�mcw(�'Xi���c�v�VB�I(��<��lĽp�,��C�ӄ"�$B�	�h����)Ά���*�nN(��C䉎��#'nX�+v���	��CMPC�I,�v}+3ɕ'6���nD�;G$C�	)v#@u�Q�\���c��L�`&B�ɶ�X`�gH��H�&}��C�ɝ3�A�@3h���ma~B�	0N����"ҁ?���钍�DALB�+o:�x6g����zaKϫ��C�	� ����Enȧ,��tG%:ľC��4²�!"�0שY*o��C�	.k&��'��/g���I�B�a��C�I�N�� ��G�n)��`�$*�C�Y��A���o�$���Q�a�XC䉃
�����%���'�Z�pC�o=�<K�۔Ag4h�p�Z�6C�#�A:q�� N���b͌)u�HB� uh)A�M��i*�aG�tB�`�<P�'����bdV�E�b�|B�I�T�ji���u� $*s� 8?BlB�	�>��IS��1|�yСOLO��C�	6���i�]焉�q�ɏ}5.C�I902���ʇY�xIs��rԼC�	4uzt�bL�,�b]�d�η^�C��5p>��*!۪h#��2c�J�B�)L0��ίS&�0�υ�|B�B䉾u��lp�Nڌs��Т�GO�BC�IZhU��圈Uv0b`ϗw�vB�	�*�٪��_�JT�2AB�2jB䉚q����۠�<�Ya���bR�C�I� d��� �(��7.I�C��/s�Ȩ"�+I��5�e�Ư,�C�I q4��{���ΩX�Ɉ)�>C䉚9����V�	:S�e��C��B䉼֬�K���(�%��C��B�VA���G �&V�~��� �*B�+W�0;�f 	VP\	`s�J#BSB�I�ir���A^�[�8�dC�C��C�ɩg���d�� (ʹ)Ӯ�� U�C�ɧeR�� ����Ѕ�0e�C䉜I=��Jo�lCV�)��B�I&y�f�c�ʹ���P��{��B�	"�`��J��fIZ� e!�� z�a[�W�1�!F�5�&�R�"O���"F�R�؃6�a�\s�"O�|9e�"WYP��!�6�)X4"O�I`������N���E�c"O�k�=6pD` ���#T����"O>���j՛Hlb�4��e�XA[�"Ol�uDؠ#x���'j���1K�"OxR��V� �q����ċ�"OB�a̓�d�D ڀb��d�"Oz}�7� e�|3Q�A�`�"O�t���֑{vV�@RMш^��H��"O���J��Ss�eI7��&Y��)h�"O��4A��/%:4��AZ�x�c!"O���-��g�`9���|�	�4"ON��rd��^��3�ɳ4�&��"O�K�ᇗ 7��+I�J�kD"Ol�����H@�(2L�=z$�#�"O,�I�ĥf��Ix�C enI�"O��p�i]�G��Z�
�'�"��"O�x��&_D⑚��� ���"OD�����2Dc3�řjN�@�"O��"Q��~��p�@*W
4qqG"OXP.���R�a�w�v�1u�]�j�!�dN���hS:W��=�+Ҍ$�!�$S�Cm)�j�)xh�2��t�!��ػ �4l�nN�ULJ�a�K=�!�$W8���:�J��M$�1����d,!�EvA>u�S�r����ѽe!�D��Yr�d[#N8R�*�k��.!�dOU~.��$�d���oV�]!�䟒th�m:ˉ�_�裳��*�!��7L�0��쏞����&J�!�^����RF&�9c��\���O�4�!�$]7 ����Ǆ<E��h���ĉ�!�䂣Bn�1��D�G¬��V	�!��Մ^V�وw�[�HB,	� ��O�!�$�w \d� j�L��Qݨq�!�$�6�fa���;��`[�!�C�!�  V [�*\.;g&�W@�Ex!�DԬ;��$�3���Ac�	9��YQM!��Q�S����=��L���һM!�dK#;�� )� >h�:c�%?!���#/ܽ���!�D	��j� >�!��@X�`��5G�=��{��A�!򄒹(��%#�v,�Q0EL�t�!��6E���FK��Qt%A b�d#!���|Ҥ(�%Q�H�|�����5]=!�'��(�f�!(��=PrһY�!��Y!U����� 8}`��L�2�!�D����W�D,C��m�sEA>�!��sT��qo��-1Z���CW��!��ޜW�J���$
�'�!A�!�DH�}�P�q�Y��X�S@M�"!�dG/J�$I� L�)��\S�nN.o!��SPkb�[c:�@h��N�l�!���T���h��l%�p¤ꝐW�!�D
�R��	��I�1n�����w�!�$�Rid�T$F
\����Z��!��=F�u��R�f�h��ꆆ�!�S��p��j��R�T��!��ĺB���	c!6H�e��,	�!�@��Q�ҁϺE�j]A��Y/)!�D�'+���R�J����ѯ�^a�ȓ{��I��R��*��pE�.n�����S�? �ye�V�*�X��E�@؁4"OQ���1��	#��4B�����"O�-����r����k�.��-3w"O���5��2}�e+��ԷZO�Hʒ"Ob�i�#r�X @��4j3�	��P�d��$!�V�'��T\?+��.ƨ]��яH�d�i�'԰�$�����?��~+��Z�Mƍ��U!���Lɖ�鯟���"oG<�:�pEݒ��5� 鉕v� 蠴aM�yr��"u�Es�T쁟Or�7�>14��sG�����D�9�2��$l���8�O���C1H�����U��=0n%ȳk�OZ�b>�&��s7KK�$d�4���O1`��LPD�*�O~�o�#�MK�4;���Z���,d���p�$�fD����9F����3�?�����i0ö���O�7M� �؝i�HVr�E
�b�d�h�� D&��2�ʇK<��%�2�M T�T���O$k�ܰ\D�=؂O݁aK������Q����(578)CSjM	��`�P�ϥa�Z�R���~�x���~�1^���Hgy-��8ƌ�7��Ml�������O H��ʋ�i�����K��	cq��w2ʌ��'���'%R��;r�� \~�6�qVmZ�=c����	!�M�Ʋi��'S�T��x�I&�aH8�ڇ}�y�d��ޟT���%��ҟ��	Ο��I��u��'-�&�XTa��83��>(F��7@�pT��ƅ4A�ɚ�D��Lf�a"�����1�6#�'Az�'���ݒr�B�E� �i�H����c�ۭ�8 ��@����G����''߸rb�Ign��q��T}�iZ`��%T���2� l�I�KL,��L<���p���>�̐:�6Ƀ&/��l$�p�P�r(<�ߴN+�� "$ױI^N�b"Y�=�D�h��n�U�i>��Xy"��X5�(fK��HjJQ��DFT�ag--d�"�'FB�'z�h+V�'_r�'Ul]�!�>B�^���ϗ(Jh��)��G���`�.Z�+��Y�Wƍ�d���{t��(O��8��ת;�N�� �^
"M�<�M�(`>�`S��8	09!�#��&��<�B�N�(O� ��'�69uC.V����A�96��蒤�Q�L6��Oʓ�?)�*�N��B�Ǫsa�YKs��>�ڠ�"O� �-�5iq:�z%�	v����şlXߴ	���Z��q��ލ�M���?��������޵iK��:w��4��a�BL�!zP��i9oZ��$���:j .�:�B�9C.� `���v���#B %�����K8M�Gv��<��C��: ��H!zQ��zBAOy8�ˡ��(L����e���1�Ņ E�苂c�z;�'�Jh�P�f�?��x���E�(^q�A�$�"Q���)����?�OC�O� ���m�\��>9�5(g�>���4�
�l�2�M;޴>���0�R��tx!�ΈH�n�W�����i��'��Ӑ-sD8�I��`oP����eF�N�����̙:����(Q�oF����J -�$0`�AX��b������`��.rX�J��j��aBt�L
~ϖ6��!t�|A�B�ե�
��	TΦ�H��=hRq�k̏�j%(+�.ة$��l���K��f���?��i{��?YG��4$~��,L\�m�T�'P ,x��?�)O$�=�OY�14���N��5���;ظ���d�ͦ���4�䓺�_w�T���K�7x�d��#�ƵX@���"�� lO���
�  �      Ĵ���	��Z��t�D9,�����@}"�ײK*<ac�ʄ��	ڤ´�xbjR:6�ɈP��}z�$�$�9��K7d���x�H� VM�h� ]��}�F�й�u��� � $q��]�"(�;t.�OiI0Dէ.DN��K@>d��q�R�@^�
+O12�"�Y�Ox�9g��+��R�^�~��=1+b	���
�~��˓H]8lD��+���'�p��$zm�K�O�\�&ϓ�5"�'"�
qY(�Ñ,��xU�)O|�	+Iu$5�D-�$��q��q�t�D�kw&���W
r�Ūf�GJ4�w��<i5H��j���t�I֫��(ìOd���ɯ{��\�5��m�m S�]��x9���r�	;/����.(׈��'��4�I�j
Q�S#Q�=kH���-	�}�⽓[Z5��H��b�`N��[��]��'�(Pt��G� �reiC�ܪ�'�,�9�c)�ay���#{-���N>q�Ky*PЫfAm�,hp ?^]�T;;C�p�C�O ���MށG�'�D9�O���N�J��m���8��(Z��%�pb�x挓O"� e��
x�����<�Rd<Yf���m���;^R��:QM�[3tP[�4"��7/�u٩O�h�'��H�f��<�%J����6bֱZS.+�Έ�O��Q�#�%Z�y�M<!��C�T��N|r$) E����Ӈ�@�֝��DU!.jL�AV[� ���'?B�Y�Fgy��O �҆�އ:��$u_�Ey�n�.Xʅ'�P9�m����0��E�<ɂ�'ܢ��@��B~ ��ԡM;�0$��g�*2�=�=H�$�x�7��O� �'�	�Ҩ�p6$����V:p��b�4`�������9)S��*�'bT�x�*��?��bEl?�By��c'���\�.��Dg�L��8���B��O�]�N��x ���4��J	V��!cqˮ>�F>e^>#<��-��"v�� ��z��C�E[�<y�� # 2  �! =X���ϻ{#Ty!�V�P� ֋�/>p��1N��1��E
o@��Λ/\�n�Q�a�;��F�D$(+�`�A�ݾ�b����P�R��@X�Z�v�	'�''���e.z�xٲ�o�B�����f��wkH�!��Y۵P�/��eic�F�;7���ǎ�� �V`M���'�B<z	��2qB�q���0o"��Od����+D_��x��Ia�=��BV�X�h�@�K�WQ�����oN���捩fJ�`9(�|��t��,��O�ޙh���c�\��I9Y�0E!򏓧�9a1EB	y|���[��ykF&�3V�$��ÏY	90D#����F$�8b7IZ9���7:��ACbߩw�Vy�C�)������Od�Dаg@�W���'j͒r�Q��'M��xD1bV-*QL�9�|pӶ[?��bA�"B�͋㋋�C���%��7O�pD��Kg��QAP)�j�� ۷KOޔ������I������f Q�^�a0��՛k��Qu#�fF�E��&\����0���kb,I�z�H`3��ͫ��'���Agd-�8��m�c5d<{�[=4�f�s�퉃�V�0TGΣg�0�@e`=wY�9��a�(��=��C�o�$(�uJ!�9Ld�ih�~y�H��)L�T��}"������� �:(@����L
"����B9,�B`��
��>̥"&��޺�R�O�j���?i����!l�P�,�W��Q DRq?�����4��)&�������b�/j����aH;�س���*t�~P򦮈N�Ƒ��/�{xJ�C�*
���ed��$�e_)��d*d�<�˅��2\Ą`PҠ@1OąbT ��@ �˩|h��)�AD&���e���� �
 ���D�e���L-N���e@NU�I�/�4�D�lX�X�Q*� I�@ �e.*uL���q���uDW�1&ҡQ�hP�x���I� �tg*:U���Ϧ1���!��°����xB��6:pE�!芆q=y� ��n{r�i�O~B.h�'��uٗ�]�M�%���1��<z���N;�h�ǽiK�h�Vm�rB6��3w ,��ʤ��� �dL='n�Y�1a�%�`�N�F\� !eA�b�Q�IA!O��7̀}�$-�D�C�W
�(+��L�Y�OL����7a_ʼK�
w�Y���x�
�5dn(,7yL����	J�J�W˔��\f�6F�2R� ��W�8��ĉH*���+%) OxqqG�+|O6�3���y���(sl�K萕hto�^�1��g�R��ݱ�A�&7��2���9;��*wd�-K�����$�u�N+$�t�3��oQJ�xOd\ ��
�E�|ӄ�Y���e��I"((�XrM�-�v��,��<�'��}р�A�k_ d��Ah�����K��iť�phd�DJ�nx�h���"0�e�@B��;O��B����0Tl��F�Ũ4扚���� ͢�Se�#U�2 �W0:��O��#�"èD��'@�sd��ړ�D�;3���ؗb�"�2�}�i�*K~�����R�=����e�<���P?v��2%��>\
@2"���j��aÄ@��Ę�2�>�o�E�2�!��)���=7)���ȓzqB�yuJD�5:�D��ƴ8��a�/�'D�X��_t����,�I���!�|K����3|O��ó�(��d��k	���I�R^: ��K
$�!���z�!B���-AV�n����A�I^�OXt� (F(b�H-8��{�H�z�'�(At�Z?by�%kܛ#ۘs�'�4�j�	S+�졲o�6\�<�q�'S�@{��)s&haR�M��|��'�5�Ƀ�ȥ#uf�4J���@�'��!�E�_!`�����IJF����� ��ZfJؼ;�]�fLR-�0�"Op����U�@�5�3cNz�ڹ�"OJ|��̭wA��P�LY�
�,�q�"O������+�4���?a���5"O(�SW�&��t�!`� ����Wu�<a�H$v�!���'E�����Bi�<���T�y�G��#d�t�$��o�<��J��j0�C#5�$����P�<��FQw*�*p�N�Xvx��T'�o�<i`/5A�C�KJJ�����j�<
�t昡GO�A��Xt+c�<AufK��.5NσD�5	b�<����!Iap��A�(~���J{�<	��J�zH@���n}���)t�<���Ŧ���� ж k�V�Y�<q&@��s��2fNŶ`ƚ�B��j�<��#�t�v���	��Vl��Ud�<A��C���8�*]&/�j�����|�<aBZ�;��<��P2%"]s��w�<6ǁ�!ܑ�Uf�~�N�G�BH�<qFE�+i�f�ǆ�<�i�aEY�<���D��;D ">��t�!�L�<�s�ހ|������Q�A�G�<ɧ����քѡ`A����GFK�<	��0^N�S��ӿB}̩FPH�'& �Cr���o�~��dF���ش �BaCЁ!��͒��Nf����8]v<� ����	���;v�p����P}K�HT�nGv}�łN/���ȓ,�x1+��d�P�dOчd��ȓ7��0P �mz^}�s�\�C�HA��l�L��Y�D�rA��H;2�����$6�A�kZ�8�l�Ad4'P��ȓR�"�@�l'���pHW�R���ȓg��p�-�)��|����dH�܇�_,J���U$4Ꜭy&�O�E��4��r7��H�b׵M*�
a��}t1�ȓy��i#��n� �t��A�4�ȓy\�9C��<�"̺��	k-�����8#���lC��ʧi��w�z��ȓ7_���p��U�<�P�����J���y ��È\<\-H����Ώ�ܸ��4�)鵄��q' ��D�6���ȓ
���{r�W23��hkL$��9J|H
ӃH�g�DXP�N	[��	��1��I1r ���Q"S�bфȓ[����s�Rގ�b����X�ȓ<PB��k�g 
�R��%Me�T�ȓb@��C�k�Y\�����mx8�����I��~AP� �t� 0� �=D�H2P��x�XAx����'J�Qg`=D�Dǩ��&���E)J� ����:D� �k�'L` L2�jʥ\��!)��+D�$�U̜4VE�a����O1���Ҁ%D�PRC��>A�X�����'���ʢ�$D�VJSϮ���c�%|��-auQ�y�a#J�N���MF��j9��CT��y�`E"{�0�RUհ�*�k�+�ybm 5l�aΆ'IjT4����yB�Br�92`�IdXu+dҵ�y2$�"�Ԭ�b��nG��Q�T�yr�!.bҐ�6IյO���kR��y"U�cw����c�@�PD�K��yr%�3&F��M�8�z,a6'ѻ�yBhN�!�̂F3+�h�hL���y
� x0z�H�n�yi`2�h4d"O�(�R�E'�L
��F*KQ�!"O�b�?L9��3�ɼMNM(f"O؀YU�F�>Rԝ�PIC;�M�A"O`q@1��:Ɖ�$���&*l@@�"OD<�f�_ l+��*�)p���"O
���B���aH ȕ�g����"OZM��J��:h�m�������"O�Tr�V���m�ʁ��+P"Oصx�I 8�1��Q=���b"O��;L�k�D�����nc��I�"O�X:��L|��Z�ݷ y.�b�"OF1��&��2����(��vB9�"O��& �]@؀S�i�;tD�uؔ"O��
`&��#��f��'��à"O��pc�ګg]&0	���c�H�R"O�LSS)�nT~4[��h�v�83"O�%C �-������8X�"L�"Ond���7����,�f��&"O�R��L"Rp�#gg�5��!�a"Od��$�7)"@�Q�S���%"O@�Ia����gH�3��=�"O ��Z�gQR�O�	nɚ�"O�[vÏ�v��i�"҂��T�!�D�(���KAg��F��T��M�!�P�7��<���!U�NiBS)�$�!��z�l<�Fk(>���K.8�!�L� *�Tp&f����q��#/�!��=N,ja�Β	��u[�M%b|!�dN6i��������Q�Dpu��_!���+$1t J��`ᰓ���V9!�$)'��GU��̥9(�;!��]�Ń���x�8�v�K�u�!�ď7?@��1��1����eQ�d�!�$�&�X�B�&�2�2YiC䘋u�!�$D��~��*Ďa���� j��c�!�d�#�V\(.K�f���	T�O�!򄟆b#Ҩ����)ca d�D��xn!�d��y(,"Q� M��`G���xV!�D�=q65���e�W�`UxLI"O��q �_���`b֊S.œ�"O���Ո���"�#"�G"15���r"O@�K2gF<G���Nޔ6z�`2"OXlx4��/`\5��-9��pC"OuK ʱ$>�5�֒W��	��"O�����|U�b ��{6�Գ�"O�@k���	��8c�Z� \Ҡ"Op� ���7L E��q�"O�9�NM^iq6�4�����"O"����dn<J��C�E�t٨ "O�C�I��d�r����?w%��*"O ���+�O�Ш�$ ��ua#"O��i��1��Aoy&��"O��`�n�Cf��n"u��2�"O�i3�5z;�-��s@�P"O�-s"�IIy��#͐�����6"O:Yy �ͼ N���F�Ӻ:�p��w"O�X���ۖR�\���kP�k �@ذ"Od<A#	^%�6ј���23�V�`�"O�ba�F�V������?{z���"O`�z�hԮxV��Rg�V,A��l!g"Om`!�
p�*�AE�k�H���"OC&��9g�\(�ť��@���hW"O����o����w�"m�0dC"O� �EФ����(�e��-!B���t"OJ�z��RY�H��F� /����"O����Jj�X����B!�i�"O|UQ��E�D�r�i��T�:\"O��t��-
Z�@�I^lQl�4"O��QI)�E��J݋mCd��"O��w�����I	�:{>��U"O�)`���0�̥h�mֺ79D,���'���OP��O����UxQ��my�"O�!Q�Ŷ-n$`b� ��	�0��"O`�8�i�t�`�
v�ۭ3ZD�@�"OB�q4]�%�wO�7>��-
��'�\pG�,O\M�R��"ѐ)��
#��"O �E�E�f�$Xj%gΈ�B�!�iÛ��l���T�8+U�I�A# �{]��#�I3�O ��X�P*��[
Nz�(DN��	*J��k,D��{�Box���'�M�B�0�,6D�X�AQ"J�vQ�`� ȉ6�!D����ܮ5�)�F�ӗ	Q t
�n2D����π�
ߚ1�f'�[�ԒtJ/D���v�Z<)] ,HE��;yJ���-D���@#�E��#��#'0}1��(D��!�f��@�6x����x
�P3+2D����̛;@c$��
��P����:D�� � |�N�J�4�n)��c8D����H�=��a��\�p����4D����X�CqB�{���� �Jf0D�0
�B�-p�$z*�� ��8D���ԶQO�qC0��:� �dc$D�dP�U�L��1b��.]�^
�o6D�Ȣ��N�����)��{4�	KPi6D�,�aK�
�daȿF��1�`-2D��c�ЎB�z�����ʭqGF0D���0I&.6���`B�'��q�'�-D��0p�
9J�8y D��}���9D��A�:S��ex�,�.QXl���D7D���#ڙ)��q��2�:�g"D� z�F�vϠ�B����F|�#H?D���"�C+[H���LO�}`@��,)D��M;uѴ�)���#Cl��BQ�4D�p�O� �ê�o���c3!4D�Pha'T	l��ICeғ��!f!1D�(B�ڜc�1�1#Q�[�Z����:D���C¸
4j%���P)�\(з-9D����2�f����[#%bBP��+=D�`Q�a��u$6,K *v
#%(D���GT�I�1�4��=d�幐M1D��1�R������Ry0 �ɇ�0D��#
1a���+R�	�P1��;D��Gq`�m�򥍘G�}���>D�𸴂�3H��) )x}d#l=D��{"�W�

D�4�M�>f� ��@9D�Ęa&D�?�<�*aI�<m μuI+D��p�mߙ|Y�,r�Ԥ�K�`'D��
�dҴv�"pZ!�G��H4���%D�x��bA�w\�P`�Jظ]��HS��$D�l�G�3%܂,�WE֢����0c-D��D#K_8����&>�YR�*D���v��6FP4 �D�@�v�:D�3�� �L���f�4����5D��r2E�J�X���I.� ���C3D�<�q� "��m��������b��2D� ��P%��l{%�ĢM����-D�@c�Ep�8y{@�A#(	�|P�i.D�� &��A��-'�l�k6��S�x�X�"O�Ŋ�F��T�TI�8h} A��"O 5s���@m���eө_SF"O���u摬d@rt)GŎ�L$��"O�T)6H_g����탕Se��W"O��3B(�?�v���/R���"O �˷�&8��8�K�RPbm��"O���s%W�(ǲ��A#�"����"OX|�`ak��a�↥Y��Y�"Ofe٤��>�4؊WK&�@�I�"Oڸ2sĆnr�����,.�H=[�"O�tR�\�������+�h��"OB�@�Ǚ�����!@�dҴx�d"O �*��,�Xr�V��VyQ�"O(U���ܣ�\�X�h	9� "�"O���ܕH�`��K����z�"OЌq&dDSX�k�Ӣ ����"O��:@,� 7�}��I�/m�#�"O:(�Np8�yC��,C�x�"ORL��͐Q�4��a��S@e "O�	����K��	�>m!`�q#"O���ڭv�����fϠL��B"O"9y�eV,q�(�A�0>��Q"O��:�L&V���%b_�@V��"O� �0�̄'8"Tx��4p����""OX�
��*Ny2ጽ��[e"O��y��"����T�Y~ 8+R"O�Q�唿�p����3
�L�S�"O��;���40{��S��1p'>�x"Ovqy� �
  �      Ĵ���	��Z�wi��:G�����@}"�ײK*<ac�ʄ��	ڤ�N�x��׷��6�'mH��fC)\\�U�bC^%	� ��`�7In����E�֦���W��uwd�'1�����7�.yȕa�O( �Wm�$�j�z$ ���!����~����+O��{�c K��U�O&�����w ��Ʈ�vr�T˄��M�P<��阔��	 ��+�Ó�qJ�I�00$I��(��cľ�Y/�[�%]�>t��G�H��`���I $[�$��C2M ,BГO\%�L�o�~���d�pX�L���J�W	.L1N>AF�[@(%��q�	H .��>�9C��4@S6�ᅢڍa_����23�"h,�Ĉ���\Ӳ�|�ᘷp���!�cؽ$�Ux�lBNp,Eٖ��Y?	3<O|�"MB���ԟ�d��"� n��\:DBԅjg���*�3+���k��x�L�<p ^��O>����Q0l�'>�@�@)6����aIȂT�"y���WhR�
Iz�	8#��s+*�Ē�~�\�q�)حc�4���I�Lr����G��~�(y��q��ǝq��T$>�rk܄4�|�ݩmoji����mi���Һ���Z�v\� �c�I�,	 � >}"
�r<��dIP����z�c�+&���1��L��D�<	1�M8���?��I��,��򈌳1�vp�����#�J���K^}2�ҟH���3J���?�#DY8X��e�9F�P����JS�$�׏L�4h���M�O,4�ȇ��D�����-O��O0�kB�E�*�5k���{kj�01�O�f�B�P�O���O������<3�lx�$f�mC8�5D�J�ؘk��GNf�9𖄁�5w�Ġ��,�f2�� D>�j���`i"i� Qc4H���^�ܳ��
LD��O8L���ǎ@]�'����j�j�ʼ^����1�:֞hN>�P�B�8Ƭy�<���$?��L����;�J�@�j� ]�:	�'�\��@ ��   @�?O�!�  � ��@ ��X�#M�Wሁ��'��ѐ@ ���GN�7��� B"O\X�Tɓ�z8��1G8/�(��G"O*d�R@
����d��5'j*I��"O�j���wn� 3�)��s:���"O �x�F�)#$x+�KӝR�LIg"O򕳵���Y &Ȃr	��.6��A�"Ol�"d��]��йS�R,�"O���OTN�5 畿6�D�#�Q�<E{���R��� 
�Ȉ�o$   �  S  O   ,  g2  �8  ?  �A   Ĵ���	����Zv)̜��Pc�@Xx����W������K;G� �$��=� ����8�҆�
znZ��A�=lM�J0ǌ�4_�1(�͠:h�͆��j�p)��>�8�V!
�!�>��v��17`��pSȉ�e� ��i�e�0��-�䘹�#�5�NL1���3s� �aK��Hl�9��ĆIN�b]'��Dہ���f��+�&�hEȟtt�1��oŲA�N0^�$n	�%u~1ZWA���Z1����1�`D��X�H/nL����"^)x�'��'�"�t݁�I�c:��Dmѽ;�Z���|X �ceE����;�f7Ҽ��BM�����,��A��H�`�`h�$1�6���+�1OL�\�h0A\{J��OH���E
�wmf�0u?OƜ�1�I0q�!�6��>tFp�_��!�'�2�	]?)�"D�(���eC�	W��Ԩ�&QFH<9O0a���R�(D���U����,��|������V�d�A��".*`���F8��T��Bc'��$�O����O"]�O,��'e�%o��<������j���6L��P#,�J�B�N�d����Z���v���(Of��F��^ފd;�;�q����$�p�bGN�
��܁0lL�]b���x��<��˟���bR�G�ZT�6v�LL�Ag��M��i�b]����蟼��sܧ!$�e`@�НG;�UÖO�� {~0��n�'[n@��A$&>P���E�&���޴�?镶i�7-�O�poZ4L�F,B۴�?���?�1or��c�B�%E����E[2�oI6m����4�	"Z�"$��g�?@(�޴H��I�Oox�z�J�+�eE��Zۉ�Ď�o�^8�QN�K����o �z���v,%2�晁AE�+<,С��-D8>n���Ć� ���'��7-�Ol�S�~��e�Q�/�p���M�{206��O㟸E�\c�Tx0�E��f�ۧ��&;�F�zI<A��4�ʔm��M�� ��n%Rҥ�%�6�ăVD*�I��^M��4�?��������U���?鲍�/�QՅ�d�Q���b웆�+\ś��"I7�� ��
F� q�O)1�^�So&c6F)KtA�ac:��%��Oh�S%�i��R��(��#�'�H�浨�%�# �&�Q�ؘ?�ju�rH�O,)��'=��O?E��E��ioB��5�S������C�I
&A���?���K4cP#=�t���Q�eΛR��Ӂ���xtK�4�?a���npr/M�?����?i�?2���Okl�  *	1��UŸ�q�;3cv��ㅝ9��pVlG�mB0T>�<Y��S�:��(�KA.��1rً�U�PM�i�`�aE��L=�O�]s�����	 D��"��Y%pt����eg6ʓee���	�0=9�(��Z��AEщ"�9[�b�D�<�fH(|��1��
�{ć�æ����4���O �Q6C(T�M��]� o��S�%JF�Iۓ�O����O���������?9�O\�ɰR��[���sBK̽+O�ّ��<]�Qje�ި�\���E8�D��X�M�����u�@T��OP6����	ݥ?Hb�9�^��#.N ~���`�A��~2��?/�XPI7�olp�1���PX6 ړ��Oz)�Ffk��|Ҷ�1Aq��(��'�Q�|*0e��r�����5=�t)棭>!��i?�V��!Rh����I�O��-w`��;�L�9�ر�
�5e�6�S�B*����O���N�m���X� �cD��`�P�\E��SUJ�T��M��0��=[5�J�j����o#H�W����,�Z�ƿeH��ɦ��	O�hI����>���a�)�T�ůۼ
:��OZ	��?A��d�B��lz�D��l�m�������3�O�� `�Z�^�pC�p)0�b��x��i>}��O��sF̆.X4�#��[)]8�7U�lY�fٲ�M���?�)��|��*�ON�D�.1+q�V�I
����k!,�nZ@J�AoZ�5��H�gW b�l9#j�5`T� ��tL�k��	0�l�c�Nq�t��6_�2L�1�ƵP���Z�R���_�R�L	�S� c���	�~"$��`l1RA�%(L{'ˀ%�?qAƖ���J>E��⁷ d:R���FnAI�hM�8!�΍��['e
"�4��Y#]Q�O^���k���$�P�{���!�*�!i1�� 
�7��O���#.�K�b�O����OP������{���,&�hh��ڔG��b�nܩq��Y3!N�V��頓 �46�,-�OG��]wg�'����s�ճ~��X[�%��^����n� j���1A��ʑ�i����Td�ãƔ4j���;}�ih�E�K�f��S
�+y~6]�'$��� �az2�KߊM���F s�^��x��҆L&f4�2�7fW�]�0��� i�6-s���$�|��٧E�d���k�0q�"h�e�#�����K�b�'z2�'��]�����|��jܦ��V��PFK
 ����c��Vt��yQ�K5�H����J^	!�7ʓAt�	xQ�C�"��!�o@�h�����T�(��_�1�F��S Շ`�	v��]� �k��xbl^�?�A��Y��n�^h$����#!�ąI&h�� �ݓ? @ �E!E�ay���sx�-HӦ;_��	�"s��I���|��в&7M�ON�D�?Q	n\��)H��dL��xӸ�в��O���O|�� w�V�I�d�?G���i#�P: �z�O��`�[�jH?e8��ç��^��<ї���i"�E�R^�ZtI�j��
� d��D/��`,����^�X� ���M��� .��A���#�ԟ�31/�A��(GiJ,�2:"O@9XB��w����␑%�]�`�xR�i>�z�O>A�WU�2e����Bm�"��Q�@�Gj�!�M���?�-�@��C%�O��R�r��ѹ�f֬2(9�@��n�|nZ� \�UdK�Wt�H3��	}�F=����1m
�T�|�c�à�8�8�#�a�2�!�e���?a���Sl��i݅C7𝁇Ƀ:<��19E�6��!_F�{��,z&lt���-
s���	�U�@�ės�)�y.�XR��R�a9&O�"�U�' �����K��E�b��5 T��(��V�O����A V'P�ִ;UgQ��{��s�~��O(m*Q��MB����O����O�;�?��U��+%-:+bT��C���k�NQ8F"B�g��(��FW�zD0�wJ^��*��uG�x⇑!C{"�cF��'.�\��ɎX��g��%qh�8��j �*ߔ�a�Q?-�Dbm��XEb�ؼ�A�����X1�2��@�Ry�#
�?� �'-�%�Ā�9/p�s�b�+j�x�'���𐯂2*j�;�.�x�T,�v��Gz�Ok�'�FT�"��,]g��p���<[dF��B��a�e�'�b�'v�Jbݵ����ͧy�!�0�Z�Z����1��Z0��p�A&"��p/�.��6�/O�-#6!����a��P�@�˶|�>���O�=��l�n�>Dv��Dn݁�X�� oE�[��'�P��������rת�����D	q|�ca"OE �/�$A���.$X��۷�'�Q�8褭�N��`�2�ɰ,@d���Ƿ>Ir�i��'��m���&�� @�>o=�9�޴ph�E�:
t(��d�Z�J� ��ȓS�j�+��ۅ#���w��?2T������ 
���ZEQ6�T�M�,������N�g���
(T!0\B�;
���q��	�du�p�->B�I�pº���ϴB�\��4�1*�B�	�?z���0o�Qgvi6�P��B�>G�X�cAâ!tN��Â�(i�B�I;���cg�xBg�N.J�lC�	+����)Z=%��x��b%4�B�p�ӈ�:D�h��f�$ZC�I(�:%bW��a��̋�0 ��C�%&p�
�MR���GH&�NB�I&m��Zg��;+
�cȚ�;�&B䉁&�މ�p(LF���� `��J,C䉄�`��1ML�Y�|Aʶ��8QC��<��\k�	&XlzB��7�C�	-_u��d"�,�D�G �oɴC�I�o�rmڒC�9]�^%8Q'�d���*߶y�����]�3��&�6�'p��ɩB��EcB:P�>MB�կV�C�	.1��DCvb�5@"�z��S�6���c�A$Dg��P,��W�i�m9��O 5��L� �pe�AA0I��9w�'��e�CE
 i(�;s@pI$�*&o^�`�V�pS�I;;�ڥY7L��B�f���D�+��$�e��3J�=�U�B9>�'
<=�W�J)8�H�F�]V�M;�t�S�T�%a5�ɝt�AJ� ��nB䉝G�;�n�1Ul��G%�3x~�xFE��j�HW͆�X�k�_��`��I 5t�n�	,���W�)T,B㉞G������	%!�IX�����p{䮔�l��Qʊ�EM,Ш�����O�d�-K3�Е�`f�V9*�'�P��bb�>YV8(a][��s5Đ�
�th�c�M7h`((%�7���74phh�"�6IrT�����0hO qA��f?��nU��Az џ����E�,����M;4B�0ZdYr�H�H���-X��-;��>)��J
pD�a���y���	�R,�CL��Y6\��Uc�'h�@��Y�xٳN��:B��79���lU�ē/�0�ɊJ��#b�>*�	#S�������� �8�"4��YY<Pig�I�
B�$�ۯ ���rŀ�hU�$�Z���#Rp.5�)�:�	4�?wL��t�i e��5��Q��8�(H����0?�1mJ.��fh�c4	3C-�T��삙)�:BK�02���BQ���'!�(���Ѵ	̥j�, r��� 4,�#2�'�.T�a	�3<��d	q?a!jF�EE�6���`��x"F0vbfE[P�P!*c�8r"�bP ��FP�أ�J�0�������8�q���<��#��;��E���?|v��������&r��C�V��\���ۺ{�FYh$K�D�`$���%x]����e�u�'�8 P�	
52�I1�
�1[�9�f�S B���R��T#�1��#��I��L��b>� jY!���8��u��ˀ-�*�����%"*���M-�Tɪ�I�Bw̉�u���)����R���4G�[�'  b�c�9�O~'Eٟ<J��[�
M�E�5�V _I�'��)3�g	
tMlj��J�<��i�7�*�ȅ2I�h:�oY/.|6aze��R\)������M�ǉ7�����Y�2A�9�e��s���
��#x������B�G ��	�T�`l�>��JϲB�nmk��Rh��qwJ�?O�t-(b�Άf��q)���,g������#e�ν���I40�3�L�!:=P"�̻p��	9�Ε�Y>5�.Km���'
�t{@���]p��G�T.q��	�Q�'D�x���3b�5���.
�X� �k��8 �w�H3L� �t�,"y��h���	�>*���#�4�ħU\�@�J�K��(8Bc 22��5�,�����AHP]ʴg�����,4Vިe{� �`If$�<r@`�B�W���p�i���J�Q�8�
���xQPΑ�k�|ѫ��=}���C?����*��2���\	ხ��a��@B9���{Y��!�|(.q�L]0'�i��!��~^�0ʅ�7�HO�X�&H�	�R#BmT���s�>��6-M
 Ĩ�����v��!���fy���Bd��l�&�Xt��7mD�Y840!r!�6�>As&Y >SF՘�K3�i/��a�–o���BI1���)�2�DY/q�T�(���>6�9����m��'�(�b@HɈ4$������aK����'��JG
._~��\���xBl]1r0ZA�]8o��9��jG/+��[���UZ��Tg��	(v��FGΑE[ay���,( ��c���	mɐ��W{�	r�'�d@���?MkM>i�ʶnǔ�A�ھf�8@)�Mڛv��|�)�k�ږ �ҵ�AK%Z'P�o���\��'�(�8u��8����Ӧ&�����ͷhny�f%�Ȓ��F�_8#=���KN���j7���d�bH?����A�=��m�(�<7�L#�����'S�D�[w���ʖ ��q�F:?��c��Z<�DA�c@'9��ݠ�dצ�V�׻h�p� ��[4�-�J~�'ܨ�Rp�BxM�����P>k;�;�)�!7�d!�ӌ޿k
䱲�	Q���%RQ�5
��"=�!1��H�R*�#�Y)֛� rg��F��,�u��T�V���@]�|��k@��b؞�)�5�~W��c��Ex2k��hgdy���Vmy�ٌ~����)ޢ����F�2��8�KޫC`��&_�:m��"�"�!���!�ŁG�0�Z�'B����07$	�G�A�R���A�/E��qG�ć�7���@��:��􏜷L
��l�e��&�|-�i"�ٟUw���@�r��JѺfҞ�[��Y����	���R��	9K��=Y�荒z���MU옑��&γ5�)k�@8�,�tc��2	b-�B\��a;Pl�By� �+1��0��@�E�:��D�����?�DN�S���9f̸o�$�p���*���ɡO�T�؉ĸ����Y�.�j�b@gq��Ĭ	"\��K�$G�,u�1��,�hL���d����X�|F!ɐ�� �\��%����O���c��L�| 	��tG��W/ȫ@���ѡ$7t��(L)�yB)Y�?��@�ʟ�{�"��J���񢐮A�gve[��X�.C�I�F9�ۑ��?�;R�� J���t���e��A43	�E^�h��m���X�N�EQ5!\O�!���9e*Q���X�S�����H�V6��|dTy�!�D5*5(r�_Zw��$Q&&�$	A�̍9���';�Ej�*C���!��]0
(y�'.b 2EԮ;Y������W{VEk�����U[�Kp�����as�C�I�j:ţb���($��i��;D�b�y��[,
�(��Fj� *�BF->���"1r���JTIR?ǨX���
�y�昋7@!RaϋV<"5�gGI'�yB'�#Q�0Pr(�"?AaҍH����@(���"|r
đ�Bx��Z�{�z�� ��]�<Y1�����1#ʪl@��`�ɊR�@��'��Bt �3��y��߸A�`P��k����7}d�쫔�ڃ6���C�
F\p�CN9�$A$.�;m�d2�U+T�9ӏ#�dĤ�f���F��L~�1̥
V`�`��U��-�@�_�<�Ü�P��q㮔9{�t��<	��]1wnJ����Y'���ӧ1���a5"dw౺�&BD$B�ɪ6���o��[5���h�'o�iz7�͊�8�z�P>�<�7�S7C�-2�N_~�	S�@X�����%@r�|���r�f�+
W-���n��;�L�#cb֌r��U���ƚ�&x���/f�7��Z���b��q�LH�6,Y��#=�ЀT�v�k�ǘ#�$]J?ur��:O��/Ш���h( �tv��*+v���4:��� đa��;��'Df��r�_��vtkP�ֲ�X�ߴu�N���ή.�*�X��ڏ�I�.�Vh8��91��AcJ�H)��R1�I�cIn�'�9�&ĉ��R}��Y§ �Y��T���	J����L��e���\��Q�`���^O��"T�)�}2��i�f����S�O+�d�D��U��	�
�?+��M�U4� H�Xt�؜J-t5�ҋP�-�DiKa����̫�F_=��&B��T����#|
U�`�$�0�	��O-8� ㊐`�'B@s	�I��} d�Ck�]�nlʠ�$#���"O�Y}�h��ֆL�z@0޴@���%�_r⓸Ę'Wj}"��nĄQ9Do+
�,��'Qn��BD�t����T�b?-�t����`� dQ� ��P!1�R\s���H���ɏ�A����N� ������*���4b�<P��u�(O�=`6�¨ms@��ӵ����Dܧ ����U �=�T�G4mB� aѠ(�OX5*��Wjĥ���#Tn�zRoY)��"��i��� �8��YRN�D>ȩ��B�K�"|&E���IBf@�	{���%m�J�'zfq1 ��:x"&;�<͠qN�+/>���I��a��P����,ZgĽp��#��G̓B�j��ˋ���x����wnzQ�'�@�!�P�P)6��>�<hxN�gɚy.o�(�Pc�#62��a'�X3X�!A(�!W�6=`'96�3��2 ����Mq!V��g �G�1���2U�f�?[ƀ�y�h�~�j,Rw�EQ�V��c �K�d���:�	%nD�)�J�٤@�7���;�b��y"O t<x®�$&H�����<2��C�K�G,�LCd�\���!G ^�<zĪ�f�������yb���,�� U�&���̞���>�Ȗ�'`vma�kK�Eh�¢�" `���j��{�6�{S�=�)�?,�ȹ�gS�w����\�(��y2fU� ` �"Z&�,����hO�XE4(XH��Џk�@�{&CȸE�T`ٔϊ%9s*�i��Ų_�fr�$�y�Y�7���V_^-�!a>LO}A	D�T���'�P�pqG�d� �@�L͈N��в�+W��|B8
T���+ =kPмswK�7ј�S�*h�*AYq#�2 2��{��'��0�b]�;�H0S��{� �{,�a׬ȡ]�$�+�Í|@v�
��kT��>W�L��[y��z(�aנБ=.v�P��[- ���ޱ):�[B���56`�kC�=��I���"
��6MSP��)�	�y���� ��?,�����H�2��К��J8H��vAK80i��*��,1Or$�$)�'JOxPh��P�&����W�P{��J�D�"5¢όy�p�����5Ip$B�a����+	h�����E+w}�H[ǔ�NYrhc���N�\�pӏ��1�	�ӓ9'�e[�a %�r�����0v �q�W�E\�0P $W<N�g�Y�zdY�i3e ���� ��P���̧7��I�e�l�rA"�❷h}.���Z��LIqC���$��c��:;w����/EwT��TC�_֜��u#S�_��DpEQ?���d��[J�ȑ.�J����L�|(7���8�7�-�bf�lAؔ9�Rj %1�(#'j������.h�sªE�H�!k3ś�]+:��"�g,ZU����vӼ�ر���N���pĦ]���'��q��HYE D�ڟf��YU&A,��W H�� �h�-�5�rq��@9��E� ¯Y2���GX������؁9�����	�p��A"�YH�}�D����L��*�:䬀� ~����*x� �����N
��L��C��O@~%�&爣"&� �׃aیP9�%Y�z�h�#�(��I�����D���cBƄ:���d "����V̽*p� J7Na�G��Z\���UV�ZK"�q��6~��é
Ȧ�(ScI�~����2���m�v�^��2 �c�b���6�#��Y�%Ծ0��9au�Cp�8�ă��M�@������C��R� � BŚ*�<�r�ƃ-q���)�K�T����$�:B��=#A�ذf~�� %˚aW��!���rT�c⟋,�2�p)�*b�=̓����&!ÊA�n-}/���1��,if�ȵ�U:!�D�+-�i�g���4:��I�D�XX2q֮��vxxJ��O����ᘓ6��f���t�X�J�\�x�pԪ��]FXx���K�60<`��#uB����ɷ�az�,j����;OE4�YQ��[��
6� t��QLúU�oگ;�9Z���W@ۊ5��g��ړU$F<�����r bm�;�'e@�"&"�c�v]y��ܸ�4�RW
L�"m2�gυ�MC�ʋ}�v�Pv-о�l���c�
$m<��qc�8���Zߓ�4��BGO18%��g���6H��E�(8�����K==V�)&b��9����NW-�8$��o���y�;hi�;���$��5���QK����?C�@X䮔2)_�+�h�x����%.�(��ɖȦ-� W*]���i��)�d�&a8R���nVŚ�dC�v���Qa�!16����'%��Se�q����kM�.���M g�^T+�ߛaXJ���"?�T���0�#ta�5}"���(�[� ��q+����f�RJ �,��<�VB$@z,�f���h�bԨ Nς0_䕃���y�5�v"O�.K�?�8�x�D�&�LD+A�.i������<1aL����Ȗf�0]��0�l�I#!�d��=m�6��U��	%u\��0� k�'24ݻ���:x��j
#A\~p�	�q,�1��>���䥘��@*r"L��@&UG�<aw�IJ��!�I��dʩ�vgF�'R������98<*#H�3M|��x�ܓ��B�5J�*$A��8F�Fjd��B�	�f
Չ���s��j�G9�B�IIx��� �<Ⱦ�X���?�B�I�
�Y#j�e��Y+�+^>uzvC�	����!��1�zp�7���B{4C�)� �����83+(|��u�mS�"O:�H��@�N�$I��T� ��`��"O�l�1�S+Q��a`$�^�0ƌ�Hg"O�H\
��wb��B���)��yB䌈10phCCB9;<�	qF)��y�B�I�.�9!���9��-)�����yN̈́&�,�kA�4
Xي�kڟ�y�NG�.�0�fB�(<�a�w�I��yB��2
�(5Ň?%IN�[�@Y��yb�E7�,5�2#ַU��XA���y�g
?*���qc��^s�� 3�Y��yb�L�Bê���R���z��B��yr�_#XH�z�ݢvO|i9b ��yb#�D�&8��FI�n�@�`0G�y�KЎ?p6�Bwf��RQp�+Ϻ�y�m�5	V��ȕ�L͆=�eh�&�yb�؈!�� �H�p�b�UE��y��5�|��F�d��e���ٔ�yR�\(l�L�@
��sD�z��� �y�A߼Ec2�Q"X���Z�CT��yr�ȕw���� ��Ҿ�g���y��ǈuޑ���		$li#��	/�yrOM|����?툤c	B'�yr̈́q���'��0\Zy�B���y�`�-N�b��$�\�Q�_��O�q۲��xP�$����J�z0B2�i.&)kei�����a2]5�(�'��H��:+^$F&A@��$�	�'�y ���� �E�C�0��'�N��5O����c�@F����'+����ל}[�@b�B�G ����'$؋���:���.q�����x�<A��R�z�֡s��M�_S$���J�o�<ɵD��ެQ�a�&p�u9! q�<!�'��rH�L aoאW�p�b�m�a�<I@͉"�L9��7 D��q�WW�<��,��c�j�5��4iw�I�c+XU�<��d��n|0�)eD��G�l�<!���T<�P����`�֡xTGt�<��$?f���G ,��r�<���Ӗ
žD�cOŅ1��bVj�<��)V�g��f�)�a$�g�<1#&A�5��)�nL�薀�f�<�4��7���s!��$5��u.b�<ɥȚ4+�>q�� o�0���V�<�IJ�
w�!$ܤI���Ui�<YV���I�x{f��������]�<�f#Yhe�tP�H�Mሽ�1�
X�<�g��9҄��ɕF�بC�-ZY�<	�$�	~�P��b�čQ�J�B�X�<iD	?E��X���
k)�p�K�<�t���p4��ۡ P 9sn�k�<�D��$����BI�����3�7D���H
�|�8�:��O"��0B�.6D�p gBȕI��x��
Ow@�˥�>D� ѶjVu4ҥ0�mL��x��:D�(	��#V:"�hs	�! X���9D��X0� �H�.��U���Ii��7D���f���qKv<QGҘn��Z��3D�4:�ȓ�I��A��O��\pGJ4D��p���^j��-X�lC*O��2�$�23HLR@N?T���"O�͋���"��	#�j���8c0"OLx�P��� ��2iq����Z!�d��8���`��܊r��T���#!�� &xB&�96���E�K�(���"Or���g�D�`i��i�@�z9!S"O"11�Mɶʲс�_i�N��"O�|z��Z"AS@���?pH��g"Of�[�C ,�-���ھ&����"O*!�I�3U��=���6��Kf"O�iBBϟ�	{�%����q���"O��*%��;	.0z���p��(�v"O�IY¨>yIJ�a��'u�22a"O�q�#e�#��Y�w���}�UJ'"O��ȱaV�,%�3��S�AB���"O����	Mm�U��H:���"Or�����'J��U�BJ���h�"O$H����Vn2�Xq�>��0�w"Oz�qn5E6y� ��	��U��"O XG���jjr�yAT�j͚-�u"O�mrPJ\���Ez&.��y�4�3"Ob���5L�~����Q�h�:4�5"OXB�Q��b��m-�B"O���F�ʚR+��Ae�0x'�q�B"O��1L¯tQ�<�$���)#��QU"O<�*!�l��rB��0�"Oޠ�f�B�zC�E#7���/�|!b"O�Z��!~h��B	2 #T��U"O���&�>R���ˋ�,���"O,�x���,��,spƖ+x�a�"O�m�3�ǒ;1��oUr
�p"O� �˟&�xيT�I<s�i�"O�a&�^����Ku�������"O�<AP��+N��H �Z�^\ �"O�� �<42�؟=+ƄQ�"O�T��@�N��D�� �'(@����"O>�0�$1Ƅ��0�w5(58C"O��'㑞6�QR��_"g@�@�6"O^�p��+4�ԡ6�'jOJq��"O�p �a��5-��e�S8�-�Q"OJ5C�� �w(>iT�Z�M��y "OZ��� �3!��B�Kٔzb~��"O���%�
�;���*��{J���"O,���;JS2+Z5N�p;S"OP!BOY$��I�g�@�C% x��"O
� W%f����	ޡ1?�T�%"O�I���;nqh8��bB7Z��M
�"O��*�&��5�aZ1���� l�<y�G�_?\��g']j�)���DO�<���1S�PR4g��Zک��̐U�<����]o��YE�M�y��P�ΚK�<1䡆�?���'�<~����O�<a�J̯t[���RbϷ.?u(b�Q�<�ƏǜSG4����1~�>�C�j�K�<����� 7�B-n-H��S��D�<"�.Hjp;,O+~�^�+��L�<9���	m-��H"ማ�,л��|�<��I� � �cd�)�$E�]�<��LS�^��@�E͜�*yҌAdk��<���	�z��t��gL�Z�z�cDb�F�<)Q�� 	e�(�iV�VD���!/�<Q�׳�h�;�A�n8���g\z�<�g
É@Rf�+"#\�N��,i&�C�	�g�4�z���W�� �E�~�C䉲H��;�䘿�d���,n��C�Ip���!��^2L�V��g���&C�Il}�<��	�)�]��\���C�	)�Ԭ�F�Ю}m�`q�;��C�)� $�J���oŨYA4G��ju��"Oz��i�"�LQ�f�.W�>Y��"O�A��&�?w�<	jbLR�to(!9�"Oꌪ��>1*p���A��ĝ�u"O D�7����UYc�%Q"O�����Lv�.�r���14]�X(`"O<�p ِ>20t�&�G��,�{T"O8�Ⴁ�*�PPi���Kھ�B��'��O��
���*@��ЀlB�N��$�C"Or�93A�3.~�5B�ݴCD"O�r��]M�M��@�e��E�5"O��ca�r������:�v|H��Ҋ}-	R���$ل�x�
ðm���31�̚�Pyr@�6����ҧ� u�$!˵��Mݴl����.g8d���J�R�R}k�j�`��|�*ײ����t�� �Y	�~��#HO�t!��*Y�TP1똨b�tr`&#?�!��Љ(��0f�y��l`UeP7}�!���cP�}�'�J��dy��M�7�!��3������δ`�^!��]�W��#g
�:f��	����yO!�.8����ڹ�SI
!�䌲|������6=�2���ߪ1-!�䜕s�jw��%;���&�6�!򤞹8A ����S9Yt�	����r�!�$Ӻ����@�8W�`�+�!��3ox��[rn���b;�� �!��
��H�,K)>��,�&��!�䋐Nnh	Yp��-58�P���>�!�D.�ҩ�*߫?��ZP@2@�!��Ø%�(x ��O���Ē�%�F�!���"9҂���5`�*CE\�[�!�䝧W#�DH�%ۣt�����d�-!��Z%$jw/�z�
�s7d�E�!�ċ�fzt�
	@p2���#ʓ�f�!��Mv	"�RU�I,�bI��ִ�!��5N�|=�.Ҧ*X`s���r�!�$�)i
�p�PHӄd�&�) !���!�D��g�X�Y�˜*F���ᒀ��!�"z�z���D5+X�#�
�o�!�D�Eʸ�Y1�ŚM#����G�jz!�D�oL����dlp��OV�}f!����tt�E)e%
�WE�QX!��XNXQg�U]�Q�CF�-f!򄉲l~|��"W�����B�2&!�DA[�L4 �i ?��� ��R�!�DG�*ţE�
�F��h��s�!��3w�ɲg�ԊoSBl��K�n�!�_�?�q��.9? �J�䗈v�!�DˬD�Dp����2^3����#�-�!��M�p�͸1bJ(-!�lƟh�!��XA�c%������,�v�!��7]�꩐�,
��y�F��1 Y!�Ė790� �3�K=O�@�� Q�Xk!�$��8��`��!k�=
� �47I!�L�/x��`C��)cL���@ب H!�D�gi����n'^��nP$(!�d�3TC6�z5�Z4hK��!�D�u��Z�A^e��:��˒�!�d �B����6@��*����7�!�$O�I�&�q�L� S�D�è��e�!�D��+kP-k�����ѠT#	�!��O�L���D۝>�h)W
��d�!�ٍw����e�ؘ6��`��fUc�!�� b	 �+ʔJ���qp�@�BS¥��"O�}{�CG�rs����CYa"O@��)էga��jr���|�i�'��k⃞A���I�35�Tz	�'4M�&��3&~����&�.Q	�'����Ճ�U���t��U�FLZ	�'ָ�3�lF�Rx~dг)��\���	�'�bșs�ƘC�~yi��ߙ^p�'�iB�,1�*}�׉�aS�'�����6e�D����Δ>P�J	�'\����`x�ٶ#]<~i�$S�'Z�	KC��	TJȨW���nc�lC�'6Л���z�t�r�##j�J���';��ƈe*V�Y��.xڒx�'O�5����V�"U���n�
�'�䀫���T:�0�����	�'��5R&�D�����C��v���'7V�Z���\<�Z�#��
�'�^,B7F+NS�=+�`�u�n�h
�'�L� 0�[�R2�����l_�{
�'����1HH�z�F�I�#YaLX�	�'ĢPx�b�U~��qe���g�6(�'��Q#�+XZ�Tq��,lA�+�'�,H���F3&W�<�〆�a�\��
�'6�A�ks� �m��a
q'4D��J�*�=ZJ�0� fR� �4(0�2D��Cʚ}�M��*���	�2D�� `���p�v�σQ���F�/D�D�wjT�C�|���țB��Y*##*D��e�    �      Ĵ���	��Z�Zw	�;B�����@}"�ײK*<ac�ʄ��	ڤ�N�xR�˺t�6ٶ d6t��)9$��	��F	@S6{ ��=�XZ���`�����u�o�K.!�eăDN0�"��O�yS��Re+L	1��T�vt���#�[r$ձ/O0p�d�Ϸ"��e�O��f�"ݼ���#��d`VAi��5_D�H����$}2�482b�/f�	�*��,X2d!�T���aSc�
,N���pV�I7���aR[����'����bP����O��%T�G$p�{ab	�D����󆉨{~���L>�2�%ln��%�tb��2dw��ɆUnXr@.m`�2�Yy��	��Bm�!(��	`��- ��|���0;�`	wGQ�/�&�� �1x�P��HP�I�O���*"#+�D­C�b���D���ڶZ�K�48 N�
tŉ'	~1�E޲��:��!�D�t?�r�ϯ	lv�HǝN�`��d8_]��;�T�!L>�$@��f�%�L)�DJ���:Ӥ���
���!�:p�b����<�DT�Z�l� #��e��i�@Ay��ą&���´cԮ%u.���O����L�,A&�X�O�<jqk�U����P�'� 0�RU��J��^� h1A��!Z����xbKsP�����D�U�L���4ԘG��-`��0�>��OZ�����D�䟐�e%��h��	�Q�ts�D�r�X��ı'B�q�a�'?������PyBa�O]� f�'~�H�a�={��ТAfҝ)�2�	�-�!�'��'��'�Ы�'��`�%Y����#��9*��r��Y�}���
�8�*��&�)��,���m��u�ƛ��Y���s��B�g�8����H���:�!*Ԟ|��Ż-�0E�L<qq�Є�~�D`���1ғGP�G�� x��TW��O����b�7�Ig��ᄨ�	t��D���؞X�B��&#�y�<t�Q 2  ���.D�0�s�   �  �A@ �� ��"O��3ȇ1e�>�(эŤh����"O�8x�T�)�~8x1&M��-��"O�	�U�ڙvE~�X�̛�r:3�"O�0�ޤ]9��{0�E�"4��+�"O@%��I�v6��#�&e�Hi�D"OK��i�<�P� Iҥ��.�yr�M23Ͱ��,�3|�n��bS�x"�3���`�O n�ܔQwJ��D���b��6F�ҡ�3E$   !  �  �   �)  0  i6  �<  �<   Ĵ���	����Zv)̜ȀP�@Xx����W������K;G� �$��=� ����8�҆�
zn"\ӇX/nw���gɑ�wn�e�
�����eD���p`�!|熡Pb�J*�T� ��\>
\RG�/���" ˇj[�U�A��(o�p��O �$H�w盵|�eӅ-:AwH� �N��A�p����#m��9����V�����+%tub��٠t x�$ϕ6F�`	2�"V]$8� �_N�H2s��V��`����2�"d 6&Z�ؕ�'@��'s��x��	r=��Z�c�=>��@rt����͙
?EQ��c�C�p��M�(�����05���!�=GM���4�&z���R��5*"�KD�Ne��	�|I�[Ux�Y�Kֺ�y����ud]ٓkM�af!1�f���n?����hO��IAF4���*µ<���0��M{LC�	MY�+ƌ�Wt�F�T�l����ܴ����ПL�'�J	꣭]6kG�Mx��Q*ḵ飠�8�x�ڶ�'�B�'2C�~"���?Y���)����j��8
�v��@�J��ULנ
erي#'MH�X�wn١f���GyNק8B�YQ@}[IrA���Q*^���!�jس��ƚ�Y��1���;�ƹr�� ��'�Ĺ��dk��Y��,�.8'˂�$�;B�ib�7��O���?����?���T��P @�I�O�f&3����<1��ŷ~i��qn�}�Ż���_����'�7��Ħm��9�M�%��Û��'����5�l�;g�ѻ E��,w*dA��0�M/����џ����j� ]1f^6"$���4(M�P��Or�)k�o	=u��#�\�ۀ-x��D�[�ZYjA��*UMD;7�C.Yb�y�j�<F�N(�U,��G�����Ɨ5AJ��dQ�t���'B�7m�Oz�S~�hMა�Q�ީ��D@"7M�O<��F�\c΍H��_�D80w�W��x��N<A��4�\l��M#�D
7h�0̈���N�N� �M�q_�	�ir�\��4�?�����	�&.�D�O`U3&4Aix���
N�1fP�׮�֦!�Ԯ �Wu�u�w�����ꊯZ� 3�#X\�'h7~Ik�����ҴL�w46��ӂI̿�ΈӵR%F]аё��./���+��,�S3=F`�b	����ܑi�~��ɗ/����NZ�)�',~Ą�f!VP���uk�L�"�{�'���0��(��d�ʇ�G�v�!��$�v�O+t��c�(L�V��@g�[F-�D���O���Tƪ�d�O��d�O���;�?��A�PTz� K=b��c�(�ZR�<���Sdȩ�
x���t�a����v��`	C(ī�TsE��>Vx�=!F����hA5��I�< ���ʺ2���I "����v��	��`�Љ�M�ʓ�&��I��0=iS�:.}���Hg�X� UH<���V�';F]�e
�'Z!��9S	�6"���8��|�M>���&:~Mᆊ�
* `J�A�$.�t͙�?����?y��1���OZ�de>��WG�hsf9{pI��
���Ҧ~�h���V�ў �bI�;��xB'J)ov����EZ]�L�$N�|���f�@3l��%dÌ+>��'Ǵm	���S���`1�'��ɕ�*��Ԁ}��B�,j��i��4�hOf�>��ϔ" ��K��ב:���[��OvX� EyR'ؘ?��4K���xD1$�\��D���m�	Gy�Ϛ	4�맽?��O�ޡ�3��<u^}���b�θ��4JR$����?Q��O�|1�R%��'�p� �ˀB�.U�x�����+@��d��Xl�'��`���GYj]@��%��2��ϧT
���Ȕ&	fT2�*ۥ[F�0E	����3S�|2i����	T�'p�l㰄_'��Y&V�;�6��'��~b@ER;�D���1Hi����G����hO�C~�ƈ5H�Q�Ƭ��,,���,����3R-*hl�ݟl�	e�d�ۑv��'� ٢FD�Y�RQ"7�B���C�DbӨT��-zӈ5���ΰ��x��-��=��O�H�')����Fh�	����F�FT:��I�������KJL�n�>:{9��A�*	��eT�q��5L��L�LhS)��J���	�3����Ur�)�ue�.ʪV�Ӆ�>(�R�'!R��'+*lt�ťP�i+(<��}��'��"=ͧ7���xf���1k��A��ҽ������i��'�ZM(�!;R�'��'��םğ֘�QItE{�!�H�t܋��\6�>i���.-h��h
�? �ro�|2s�����H<����r�l�CFME)�<��"k8�}@���4j���)F KM�-���v��Ġ�*59���|�����JVjsF��o��) ¶<�a��ٟ8`ӓ:��a0*�YT���)^3l 浆ēdo�YK���ϰ@I���a��i��"=�'��<�nYJ�N'G��X�Soپ��Ek��o�!򤔩�%���jf�s҃��J���'� B���jx��-S�W��T:�'J������>A@�U?\�D8:�'����1)ٌt��4�7��:Xͪ8��'X����	�4PnP��d�P��s�'ZVm����n�mC�������'��i@�x%�#�J(��y���� ��IsCɃ����Μ!��]�B"OPXi m)$q09-A��4{q"O��* 41��D�C�C.�Q�"O�d��
��1f��1-���t"O� R��V��´a.��w"O�q�W-m�h�
��w����"O<%�����vKɁm�<\��"Ox� aBO�nI�
�2i�P�"O`իv�L���W�5x�U3"Oܱ�#g�I�>�zT��s�"O��E��)�U����tޜ�Ւ|��T��׆�~D�Q{�fU�M'?��@C�*y�3��d�>d�@A&D������.$ナ��l0��틫{�����R��P��iX6}���P�[V�W���zg	B)HEФ�*=4��;uaO���W��3
hd����H�SWv�s��X<��J����;���2?�*���Oߘ<s�h3��0z��y�K׈3h2�	�:F�-���i��՛AM�$RZTC��&-L��*4�Op���k�G����$�ĵ�|� ���D�ÄG�M?6�"vH�M'?�p���)5,]3G�2�^P�D�"D���5�R.|d��@tL�0�nu"Я�~���Cn�-G�
��iDzu���]��s�bW��$�d�ɞ]���Ki64��s��� �<�Ơ�XϨb�A;9z9��*������1`F��������h0�N�T ������%c� ��?�`ĥ|J%�	: FTKs۟B�TE�p� q��6p�A  C�D���b]9�W줱їN�;'�j��� ƵSQ��	]���rp�|���	�t����4��0����@��m��Jr�'��T���։EZj<�'i��C�+G(V2�(��s��I��W)D<r�e-�Ri��3#����O��˓}7��#8F
Lc�ål�=�O���F�Y�4x��6�'҉Rw��Q�f0�-0��L�TR�Pu����Ԃ��"S��H�����uI֊���!�%Č~2��bԧN���d��P����*�8���hR�Ӽb<`:�@U��H�ɑ�y��)B�Vx����@"�`�!ꄅ�x�@�ɬ/xm ��^"NY:e��!jD����'���a���]bA`����)����Ɍ�?�s���J�H���R*%1�O��hRjJ(p(@q��գ,�@i�(��f%�� �J4W�^<�V
���O��_u>Y��a�W��$	4��@��]�'�\���,�4c� `�r�G��>Yc�'֓%~���2�(�d&��<[��,QY@�"灂�@b���"HC����l03 �|YD�K�O{� �0�Z�O�ڷ����_>=�X�'��A��-�!t͂CXr�5�A���>�[c�<1rM٧s��5���#Z���3cW�|8M�K�P<��̕�AM�b>='?�8��|9"VG��)��,qd'��M���z2TM�m��`�J�I��z�R�o��bQ@1@<>>ty�#$� y�P)�"%T������iPy""ӹ'��(h�"��{a���	=D�:4��ʘHrDe8��|�O8�
F�)z�hP	F$;���c��@����ƩשF`E��'L0zF��?	gI�*v�������&ƞI ��ܱ0d��f�[�x�b�$B*��Oab �ऑ����9H� ��K)�hS���HI�Q��� ��>��1~E�.Vjw��Pc&ɳi�]"�G�Qhb4�rO�<U&<���+��y�	�bT��0�*S�~�:0Q��# ��I�H}tt�<�e���0S��`Q� m�I�s �h�@pi]�l �!��I@G�p�H(
d 6�~�R �6P��OMJ�l��5���j���;
)((���>��^����`B
$C���G�_�4�\PK/O�U〤�&8�.�˥C�,zlHPs�ZN�������̠Sɖ$u���g�~�d�K
9�fd� �;|��p���B��yBdV�M������oI��O�:��lX/�vt*�·�T�;r��>0I��{*���P��o�S2u0u�6MS��ϟ"�Y��{��,Q��?�$�5Y�t
HˋJ�ȄAs̋FTE�$���<�`�\8tG��bdLE������q�6�
��!fL�aF��`�(�{A%��N��e�i�'�H0!HN<����KBG}2ņ(��(:7d�{[(��Q��M�l�əa,�%������|��y��2��)�
��p�r�S2�׾E}�(�H�����Q>�,�{*�k�~)LL�����,��B�.LʓJ��y�D\�Ka�c��3?!/F"o�����p���I#g�rpb% �{2B�?�K��*C��p�K?QR�a�{���ڝ'$~Yӡ�5�qO����2���3R?��Ɔ1H��58�lxۑE�((@�·�fӰ��o�-/���`�x��$?�Z���]�Y�,�IQ�ݟtM�ܓA�w-���Ē�T�	-
�ܴ�*O��K�,���F���R =X3"��,?%<�H``��OBс1+B9pN���
�|��ϒS89��m��j'n�3g��z��-;�ON��c�0��?�aU7�� �"<��Z6͗ect�P�D��c��a�#�|
Ԭ�04�! GĐ <z�x�����È��+��3 _�^�^d9H|:n�!a�"��FR�")x��T��3`��'�vC=�t@�������P*��	��㦯KS(��r��*8J4��.z���5�B:k��������?�S��D�O�D��B͌�M�p�V@Վ �<5��MT�TLX�Ӭ�)�T�
4�CsX�4+��%`�R�2��wL�ykG�VSyR>��0���J�1u������?��:���I�R�
���O� X���� �k�ޘ1���Rd��#y�@�!��>hw����
F�=�a�
"N��t���|���O��b�V5���%ݸrp�I��d����A������q�d�T��5A�R��DC�,�:���]�<�!��kt4��*�6T�v�$��B���UF���3�I!W��	�Xrd�?�O$pq'��b�H�{�jV�>���@L����C����w��E�a�G���E���-����1�rҵ<bЍ�&��9�\�z!�[�b�va�eG�Q�����;;�	���$x������B�	�BgX'��i�mъV��Af����0A��H�ִ�C "3�<B7�;ڧYfl (�\�L3�P۵$�f����ȓ�	2`g�;a������CM]�A�ȓ(��8Ǎ�#u���
�D�jp�����.���?�ԣ�:@r�A/�����MP��͆ȓ&�)�'�/~�z�K���&w��'?�4�'Up�S�O�d�:��د35t@觇��C�R�z�'<v\aR�K��<��SM�8:�pyH�x'� �T�t���'�D�#Ď�l�<E�K�i	0���ɔD���� B?<����D��Z��a�&&P6&~f��Wg[I��`�C˞ �l[��3c�0A���&�L�h��J�� ���xJ~
��Y�M�A��K���oD�<��kƙpm٘�d��F���ÀꟜ�N��i϶hp���|�����*q9!��_T����-O0!����ȓP���6�VK�8���A�G״]	Q`�Oj� ����xpE����4+д:�� @�莦fa�\�p)\�ehs/՜bb�Y�Ռ�;p�R�놮:�O8�`�M�L���!�V�0t���؞~J��i�a��]�hdGր(�
�襠��6�F	�'�N�P����	!:!�#U��0�3�œ���"� �E���쁊ȘЧ��Uj�	Q%P!�ц��?��'hK�T ��1����}{����<�LG`34Mꕧ�fu��Ҧ��d��	=�U:��ь.��T@���^�����: ��i����)D���@,�#_�������jhX�@�Up�� 8�bB:ghŉ`FRG[`Y҄��3�r�F�H�$$s��(��ݚ)h��}r�i��k�C
B]�0IF�[3n@���nA��f�&� �9Y���"b_�o�Rp��j�ڝ.�L� jO�//Rq��bq��t�O�v�����j��D��M����0 Rŏ�B"����uLP�5;rPJ���2�����,G�X�+Ŧ�Z�*�5U��R��<�3��4zG\�4�d{0`зi��<�s��ÀH�&���iТzcZH�1��f���Qq��(j0�Kc��_�h�b���;U�z���Ck����u�H�Јui�zu^��U*3}��6$u�bٴ�M��a'd�h�'%2��q���x�o��*��U��.�&����䟼OE�*tn��ذ&�&2�	Eɠ>��hЦuQ4��� _
�H83�[$/�>�Ӧ��#(aȄ��aG�t�PY ��!O@G.�>Ag� +'�4iyÎ��5�"l��OX�(���Ɂ},��[�#ږ<<���H�ݐ�Ê����l��KP��'D�]	F�Rsh�;�!ˇ4������[B�#��<Zj�h��%E*_� �s-��W�l��Ց;��@��N#���yA�ߖ|�Z����p�����F0� ���
��x��_�2�bZ��q�%�7|�~)%��f�� "�ɇ*W�y��O�rj�c ��V-�'Ĝ�L5���Jh�!�q	�0B�d_�iB8���� N�9��3T�vdX�*��inQ㠗#1��1@�hW�5)�8����0u��nĲݻTMث:��m	Rc���}Rg	�-�F��C`M [��Ł��Y�V��ɒ"8iV�W�QhI�{�kU ^,(��nU;UĂ��A�7�1O�����zE@!2N��/.��hgT��*`�QZ�}p3	M+?�}�T��B� �M�'wе0�/��/��E��a
!s����D�0vyS2�M���0�g�(�	ӓ^�<;qE�03Ь����E��9y ��gT7��>��Jw�O g��O�ES#�=~l`��Z��u���2��xÆJ �$�]q�!J.��?�� Z+%�\yuDS�scl�Є�4��S�ڵ�4d;3ʞ�/xH�f��?*]zsHK溳c�[#^��!�GT�
���E?B��D��
ɩs���f��F�'mz�E!Z�uΝg\$s��6�]/ v�	ӇC�����BU�{��d�d�=��` 
8J�T���BXn���
Ջ[-fA"��<q�ث=� H7�%Pr��a�PG}2I�A��	���#ƺ���ݎÐ� ��0HyP�3f���/@^|����-Bކ�huMM; �(0z ��7
m�� �e��WԵb�*LO����O�"�؜��JYNК���)���!�Źy���q��9����G�+b1؝��R+9����π �1�c S+CS�bWl
�WH d�'�X�@a�0+��0�K.��w�W���� Ɲ"��E���]���Ti&ٟj"\)��]>�W��0$?��r�����3BV�(D��J��S*?Lx�H"�	�`�HJc��Z8��A�t>� ��T�������JG���'���
$?�l���a�D��x޴P@ ��/�8�ў��d�3S�LЋB�Ę/f�c2c	
f`81Q��tΌ��f�+F�f��f
�#s��ЈD�ܨk��`0��k+XXL JG���mD���!� �ܰ����4����(]C��T�V(�6�pG��Q5ހ�3(�>+�ꄂ�4^��R1��;p����e�O�@m��"�u�� �c�$��5R�@E�AK0��C+řW����$��e�L����܋�f!���.Ѩ���3^D���C�&��1����Jؼ<�G����tjt�:��ѩ���O���< o�<����EL��|0�Ʀ�a�	�G7|1�®��ApV�pw恘y��1yr��K,��i�8|ɓO�>>�:)aS厝��M�Ǆۧ\9d��E��"V�{"#U� �X`{CBab��˔AH,4�R���W��$���,��A%']�`a��� Q�Te�" ~�7O�mN ��� �V��S�$��xg�$Lƒ��`N�1�@����)�4I�b A�l�`��'��LC�A6�M�d^�q7�A��Ȩ	��I�`$I�Z:ݒ�i�/h��з���N���$ÖP�4��gѣS~ihR�Z�$X�Q4kϹ�L!��D�6nMH��
�yR���ԑjg�δ*Q6oǩ��'��ɰ�c�)�|���a)^#�E�I<!UE�
<F}��k�y��M3�Ǚ2���#�o̧H&��e�@ �q3W���܄��	�5-��3U����%|O$���2�Ђc�}��x��P;;>�#5�X�С��ҽi�$���̦�� 
4���������{�⌃G�I)w�*�O:Y;q�� jl�
�iv�S���s����JX�P��6�ӎ���
;A1���!H}�D��c��-B͌� ��`�0U��:Mt�4H�5�]�J�z��k�$��iC�v�zD����#]�<���v$�{C��_I,	��k�=f�l��<��c�&al�aI�h�l����M�5l��jv/���tK3�<D� ��ͨ@���.�;>Xq�5��!H؍ph8}RcD]���$F?^��P�6(��rC�H�LV!�+^����$G�и���n"\`_ I���6/��ĸw�:Q��mi�@�*И��d[+FT�`C�	��-&sX*���>G|�$��D �(�gS�Q >�"�h^<-R�%�ȓ �Fس�藌SXv�R�M��MϾ��ȓ/>��0j[�Fj�f�۽\g�Ȇȓo~  �� �?6�!hĮb�bE��w7�|x��T�Ȁ� ���A|$��ȓ*S�L9pÁ�axF!�e@��a��P�8U�#�a�;���j��1�ȓ@i<�K�ޡ\�[%�Υ}vфȓwQ҅L����#�����ȓ�z0���ؔ$p%�pj�%@���ȓp��!`L?��H��	�$ƙ��a$��e2R��e�D<c&"��ȓ>Tm8�cۊ{�T�Q��@9>1Ƒ�ȓ(y�)YV�ה�d����ݱI�\��$����I,�<)k�	�	M�T�ȓZ9d�z! ��|�|�MՁT�م�X)ă���H�:�Bv��Z�t1��G�fų�鄘U?�����.8}�h��l�F����/�<�Q�)�4oFI��G9|�[��W� _���"�D�h-�Ԇȓ[5UK�"zT���@ �kԔ�ȓ:�D0�5�Η&�Z� M8�8<�ȓ%R�屷�O�&E�ӉO7rX�ȓ`��C�>�l�´��	t>4��XV����Q�,�BhPd����G&"��U�X�Oo��(�hA�#"fه�9���1�%X4QLux�@ȟ/�R��ȓ��]0pT�K�=�ÏO�y����k�D����d�evǉ~��ф�7!����	~h��LX �Ą���8.�\��D7��zb��gL�������y"��7A(H9��Q�ЈK�)	?�y#ˬ;*)B/Q� dظR��՚�y��2I�Z����yZ|�KE(־�y
� ��C�J_��6��㋗.rZ�;`"OT�����A	zE���s�*Ĺ�"O����(A 2�.�������F"OFm�������1 ��\W���%"O����H
$^!qp��2q����"O�(�c6O��d�����p;�"O�%k��ŮuK�� �a�Qv��6"O@]SDI� 41��*d`�dE���"ON��g���=5`�:�aαIB�0r�"OV"�l
 �X��� �bSNEp"OR���^�'u��z"�$܈�"O�Z"e�N��]���7aj���"O*�RR�]��j��[6�u�s"O�pÅ�X�i�&-��¬�f���"ON� �BI.|2T�xb��0�n�D"O,��F�7���ku#ĺK�,�x�"ODX�F yɞ�k�bD�$y65k�"O�ԣP&�o��$*���/j���r"O��3Ri߃@?*��e!����$A�"O�|�Ј!"���עbfyR�"O�ժp�#n��%+�ړYaH���"O6�j�?b��e	K�xWR���"Op-� `�Jp�$(=(PT�"ONdC��V�/;F�z� F2^T�@�v"O�%�a =$��K�j��5=R�Ф"O�����uC���fTT09�@"O��:���\���"�E����"O���oɕ1Ԇ�(����xp�A"O�|��ʶfd��	�.�b��"O��[�/b����B��8��D�"O�ɳ��O,~�8�e�_?k���"O�͓�)�0
Vh�s`�C�bf"OέYI�'�BI�7��J0��#�"ONY!�/W�l�v Bzx�Q"O|M�g(�s�իa�Ȕ"(P"O�o�?4 �2�D���["O����� +����ԣγ|��"O\��.`���A�ш����#"O*�*0�۲��ap���)�J�a�"O�=�� ��l]��QS�ʎ@�q3�"O���թ��Wxብk�}fh�"O��ȳK��Rꦉ��F6��0r"O��9e�T�l�\s��&E��s�"O��buo�"ue	��i$3,��c"OZ�֫�t�4�q��ȬI��)�"O��A`@d�:����ŋJ�~1��"O5�`/ �zы�"MӢ=�"O��a���XA 1UCq��R�"O*��	�i�D�W�z�a��"O�H�! �}�N��a�:0�>�F"Oށ�ą' $dqA`�&$<e"Of�(f�ީ]��u��e�6`C�"O��:�j��,"@Yq�QV� �Zu"O$c��CT�����%v��鐖"Op��T��me���ü*a<�2"O��Xc
é8�萹�"� W����"O�0�,�^`����-GQ���"O�� �d���X�����S%�z�<��!x�%{���_���S&�w�<�"k��b	�X'L�>�a��HI�<�s��/��h
�-v���tE�<a�gTD'���qI��``�]p֡h�<�2MǮWW��cU`� C����+�`�<Q�S�D��遣*1��9	R�G�<� L�jq�F4�-V�-l4L��"OB�B��"}u�h1\u�#"O2A: C���ѡ�K�K��T�5"O��8G�:)R�h�"
�}7��Z"O����(	-WkB���e �^����"O�Qۧ�� E0u
w+d��e"O Y���4j8AHCi� ] 6� C"OP��R�Кd��ȡȂ�� �H�"Ox�ca�
#Y�� b����vu�li�"Oz�2a��Ƅ�ۆ��m�hk�"O~�E ��q����ᄟ�h>��4"Od�㕈$1 ����iN�\����W"ObD��.�Ĝ	�#�J�4�p�"O�]yF��#<dN���*� �d��"OZ�����yN^PR*Z�G�1i3"O\�2&�M��Sk���"O�z�)��i5X��!e/<�2R"O��`@�N�W�<��4&ը��0��"O�XÒ�D68��Ԥ��#H"���"O�{V�.���9�c�>	21["Ok���mA�ٓ�Ɣ>_
Q��"O&��bK��X]�9�R�O$tL��#"Oĝ���
��a�Z�2반�"O( !,ǔ��3�&J�Q �p�'0��2�A�B`2Pi�AH=g]�Q�'�����͡�X+4��s}:@��'�2�Z�M� @g�ݻ3��	[Ih���'\�Y n9/M�p&��M��D��'
*��g�-�P�Bu#��?St��'UX�R�R 	o���"��<�h*�'�,����׺�`�	ŭ_05m�i��'&��,>�P0���\20H��K�'9�\��gYB�|	(w�'YH9��'�t�2
�e����E��$�� ��'N&قP�Ӄw!�ԡY+}�q�'����G�Ͼ>�&8��(G-����' �Ѧ�!+�(��c!M�Tp��'�H�,oHغ㌋2q�Л�'Rܹ����~���a$�@7�l���'l\�X6�)1�}�ԀS�|X����'�تq�>A����&�r	���';�R���"z��h� �!ھ�X
�'�\����\L��Tj�y�	�'�i�cJ�y��r�T���<��sY�=q�}aoƖj��W. ��y�� �	��p�`$P*)ҍ�#!I�yB�ڛi8v\g�G�	L����S ��'�*7�9�)�i˯D��-�v%����Y���q!��)�bI"'@�-g�H|���%Z�^�Dx��8�g}B��W���rT�5����.=�y�-���@�ֆXd�:P��o���~��4�O���S���6XI�v%-��D�U"O��v��
/q���$ W��"O^a��X��Y�ׂ  D���"O��(�I�Rb ���<1�N-��"O�(�G�WP���Oõ��`��"Ol�4H�QN�� ��V���xv"O��kgc��@mD��d�O?܌���"O�4�FJ�!aB��CB*���I"O>�z�ƇF5Aǂ����"OzA	ge����
�+ߛ���t"O�0�R�]
G��� �H -X�ܩ�"O��x� �(�Иc��.x0yp�"O�!��Aԅ<��3E�H&,k<X�"O� r�g�G0@\� �mڀ9K��b�"O�pS5ƌ�F� A'�,W2���"Op,� [�����4敲'"���"Ol��R��k�2��e �Kܠ��"O����D*?Or͘�	��EJi�"O`��v��*X<�)�WN �" "O*!� @ Hᑃ=a�*��"O��!�8oA�!�H�^��"O,Y�F`�v��e
���<��h2%"O����e�(�2���4� ݪ'"O�$�r"О]L`{e�9<�D��"Ov�h@_�U�H���n��@�*�r "O
 �!�:�>b�(��cʀ(�"O�Q��j�!&ZRԐM�,R%��F"O�Ez�L��~��A���.=��s�"OJ���J�|����jwdZ�"O��F��Nn��H�� H��"OL�(OE(�`����F�@��"O�����\'5(ĥjeT0̊8�F"O�ٚ!�g$.�3���*�汫"O\MPfa��!��Ԣ@��}��8�"O<i�w��"	��%1łI�Y(<�&"OB�XR��6y�qIG�B�.���"O$9C�J��fPd�*VAP""~�)`"Ovq��6XpT��`6R���"O
=)C
B�`l����F�L˾=�@"O:�
�89�MѴ.S��Q"O��A�-�a�@���)�8���"Oʩ���,�P��.V#P���p7"OVm �D�x�x���]w�X�p�"O\������:-�A�O�{�U��"O��hg�ϡ_fU��#ÕO_2�+�"O��:�k®_��Qs��[S���"O؀�3	�s�n�A���6jBЌqQ"On5&L�.�X�xp�DiM6�1#"OZ�Ye#ݏ&C���c��MCʠ2�"O6=��F(1�:�H�	+<0��;T"O~��2l\,XJh�����@�t"O���!���K��):�c�+G�"O�	�B%@�µ��c�5o����d"O�ĀaN�d�ze���Z{HAD"O� HdƇt[p@�� >��*�"O�)"`']�l�t��Ձ�?i0lQ#"O,��a�V%���� ��=h�H�"O�(�e����٨B�<�x�"Ob�+
�
M&:$��M6D�� 5"O�`�ĩV
5`,a��%
�Т"O��۔M�B�y��%R���A"O�� �������
�5�v�Y�"O����O�w/�5pF�f�F|�U"O��0�%X��	ڕ�

�(�"O��v�/%U�Z�"M)�2�"OD})�)	�-���1B
>}X��'"O��	���@S�F҄<xl���"O��!�MN-t��� f4��$"O~I�&��~�<8Ȱ�X�ic�4!�"O��9AD҅o� (J�cБ[�^�	�"O��f��?A{�HI�!~<���"O� �v��Ya�miq��lx�Б$"O�Ш� ���L�����YS'�6I}!�d�2r��1�
�>�v�H�H�&�!�[6U���B�$�BD+�g(z�!��f�=��gD6�<m����;!���F�5A"���;�8|!thF)�!���6I :     	   Ĵ���	��Z�w	;-�����@}"�ײK*<ac�ʄ��	ڤ�N�x�V�!�6�?1c��C��[!t�\�Ê}��cs��uORTc�OT֦EYa�uwBܹ!&���ʖ)4&@�3�`�OJ�Jwɉ�|Y�*ăV�_Ve`��W�s��*.O���e��: w�>���%���2uCb̨ m;S�bd��.H����9�
�(�!�&��'������C�i6pz�O��p�;j�x0��Ź93��Fk�~��k�|ҹ�5�O9�����7��> 
�;Q��@�'C�TZ
�O:�9��NXC�'���������D�&]���w�C)k�&Ī����~����~gj=;O>�J�6RwXY'��A�b�"~�����	Ze���dY�3@,��r�|��^4�!J>0�N$>�ٔ$6���C��X�|Tz0Yr�Iu�~i(dA;�$��I��)��P�h��)>���pd
B�wՐș�L�O�A{�F�K��'�0���DV��%��@��Z=@����,�iXh���|u��Ol}�pOښpl�'�t��J��M��ȚP�b(��*?�z|�QǦQ˘'�ΰ��[Iy�OT��G0��	���(�dO�ms�EyU���( ¶O�}�ʄ�N<�`胐9��)M|�cH["�@�ҧ0*�qeNL�M�q`�X�XZe�'�R���Jny��OZ���MD,
����3y��H	�<֠!p#�'rڼP	����+ ��<�v�'߾ ��I	������m��rs���@�	�im:
�Y7a8��'��'�8hFy�J~XP%��M��y����u+E���7E�5T�"8��Μ�}�f$�T;�|y{ub��Y��_���.�$JZ���-��T�r�a����I�<��dK�!%��A)o�$��x��-�8@��^{�p����9!���ч�����䭒A�9*�%r�j�&	A��H���Q�.�8+�4�yB��.3 d  �����'����@ ���+@ d  �@ ��C�@! 2  �?���'���e��6p�B0ȃ%�%�tZ��˺a@��A��^�8Oh�5l�'$���[���r��-�3�W��mZ���z�OI0qq�`��8\�S6C�2Y��l*��t�'�4��@Η���~�F�B�jK�p� $�S���R
6k�8`��$��H4�YE�*�nQ�V�·kI�dڠd3E��D�M�y��8��G��?$B���rmV�5���O��
҄F�G��h1E �@[(�{�"�r�Z	���-I���q'zա��њӓ *%��F3��Ӡ酤BJ��O�C�ᓊK��4aDD"A��\:�F��p ��$��D\ Z��W>��x�B)�v���t�E5��89��S�ꔧh1P�1�(p�&���돺1�XIҶ�q٤���:=���s����R�)筚�s��N]��֨2��	�cB52%'gv!������Jw���/��!��aI��Y�H�t���/"=�����gk��
���=���?�%�Ce�eP���O\2����+(�Nj�U��,<to�tr��V�$�@��$&����)�Cf�-X��`(��F�Oe��!�O۰=o^����pjh���>�t��D`gx}��[�H�@ʓ8�Ƞe��h�6�C&C�F=�e��͍\���ƈS�m(�q�*�74�.1öA�-W�Z�hQa��:�FB��O�B�S���5)���`G!C�"���4.��X�L�2��u(p1�`��H�Z��O5(���H7!�'��]%�4��R%AO��k���<W��������i#���R����h�&#��4�=�`NEJI���13i�=	�a� �B��� �ē{>�I�&L�z߲�˴eX� ���D�ڱV��Q����d�,�ӣ�p� |�
Zx��E,]�6���"����	�V+]Z6����nX�(j���v49���9	��b`�<� DXn�0pk���y���k�O��@W�:F����*x&b)���c����C*�7W,ژ�wOflbp =
Ơy4�0�nh�#(�$ h����'Һ�kG�>�vL"���?	��ɀ_?��A�w�����ͫ/>����#gz�#�'����S�]�
�v�� ��.Yb��ިPa�a�P�f�ѡ`���%�\��f��`HN��O�c��� c+:�%�=�T1��'G{���r��Y
��ƺ󦙡t��)��(!5���	�0l�bGi��p-���Ɉ ⬃�V�%�XKF�Ur"��'J8��,*(�L�	��tm�WV΅l�q,�E"�m��L@3#Ǣ���S�"O�� Qb�2.�j	�G�X��Mk�'$�'�	��fJ8&Hb����w�X%��$�̑pc,H�H�i�'�\-7焙sǞ����2(Ҿ�T���?rL�)W��z����F��5v;(�*���5a��-������8�ӫ*��a�M�*��1n��M��х�?�q0�O����Q�*����9�e�4LO�>�P�c�_�<����C�"�`�tC<E3��[�i|�ԇȓ`�4���� �#��'��"�^��y2�Z!��:���r���_��i�ȓ!�Z�C��!?BԪ�Q;<��ȓ!���r%�:M�-�A��
h�~q�ȓ a�O�<<�u�ֈn��L�ȓK���)�	d�l��څ�6݄��^z��D+�=�0oS�OBن�I�p�$�&��*�d�--��؆ȓ/�Y�eϮ���Ń*[��Ն����Z�h��f5���
R->D�<�# s ��M�/J�<Y�l=D��sf��[r )Hc�ǏO���0�8D���ՓVz�b@`���̵�@2D�0z��,|��#��ã8�|�C�>D�8�f-OXȻ��^�X�<0V�<D��h�bÐ:�j}XΟ,��<JĊ9D�h�FF�6�fzFzx��˧�3D���V!>t���Ui�0D�����3D�����+y��x��ݥM��+�o-D�hJ��Do�~�Y��Ǹw�\��L)D�t�6�
BL�B*E�[�T9�r�*D���Ϟ�'n���@�p�6=���6D�x2`��wt�A�	Rk�"�$2D���F8of�҇@Z��ҵ�2D�t�To!8P�i_�(�ij��1D��0��I�c~�`'b	I����S)D�� @���	?#K�RAI"�2�C�"O��p���}݀4�f��LK�"OF����d@���/�>a�:��F"OT����S��Q��'�Ȑ�b"O�&j  ����r���/9�3�"O �R�B�%�&��2�A��,��"O�|CfN\�m요�Q�W�r93"Oz%������	sc��h��A��"O<!�営 �d��.,G�*�s�"O�= G�p�d��be��#V"O�1�Ǆ*4R���픦~c�I�#"O���FE׽E������"���"On�vA��a
-���Xs"OPL3�	ǈ y@�@T,�Z�dP�"O� qO�\�޽ڕ�����"O�q ��!O�U��ψ��p�"O>�1�ʘ�Ը#�l_������"OR� w&(XB���r���M�8���"O4$���@��aR��"O�K���)��i�� �;a�
"O	p`�M�^����%?̨��q"ObYɥ�7�%���'��1 C"O����+��z<B$j�1��Y(u�'�p:�h�l�	�]��E ��Td�(�q��00-B�:bX0 [
�>��(ԎQ�)ɪ�|��a�ݣ?Q�ӧ�����b��T��|�5X'LiR�&"OxTY �Q�r!�BH3Bk�������I!� ��F�Z�3��b�4�hs�� oN2��������D�,�q
b�E��vt����tU
��'#�VLQ`Ǘ�=�DdT�(��*�Kـ7�
0��֯C�^E�ïީb��h�`��2ԭ�4:��:��3��s
�.B���&��2�ĥt������t���E~B� *"$)8���T�S�.0r�d���Bi9�[1>��(�2C� Jf����iՔW�1ˣI�"��D��~�De)Ѕ1?��杊��}["Ϟ�u�~���KW�~���x����K\�^����\������E�f�
�"��Hsl-KXP���$�"DJvd!SP
��(�,��1�@+G�dEzb�+��0�wM����Ire��~�l�Nv�����Ft����*�=��Q���ǯk�D�X4�_8�:���G�%3�X�ń.0@�AX��ݨz0fB�Ћ$\N"<q��K	\a�6-�t����qL��[rT��&ݔ���N߁}ȄX����Kh�U��O��[��=���Zp@ј�Ɯ����U��}ʌ@�e*7{�~u��K�) ؐ���N���S�-��)]<�N��/�,	h�ju��2x���'=��l��ϑs�M#�B{m����i�X�m@�L��2�<��'��/>��h۵/��w�eC�l�yj�䮱$��5y�e��@VH07��6t�,�S��5^p!�u��!�2>��1�Oȁӆǌ�'��l�G�̖,(��b�N��xӦ�_%T���B0+]�� �6n"�}�坢/ � �� {�'^D�aFZ�R��;4��|� �@Qf�lF�1�MмA@���j�J5%۞���H�#Lлu�G�2Y
h#MɪYѺ�2r�62����'K�J��Eȵ�ʯ'͔�"���>I|��'M�95Ff��Η�����\�P��¥�3���(�ز� ����-X���M\qF��`�:~�P��e�3���`���1����j��(�t3�`_�b@ÆcrBu�*OB��Q�	V�%@UEK( �5�G�D)ڤɐ@e��R_���p��T�P�Q�6Mڗ�K�,X<H�愪O	asum��y¢ � �jB��T ѴU� y�G�ʁ(VpF�)I���@4)4dmH( R8�S�ʿ&P�R#��g�<�a�C*0a������Te�T�E1X�>t�F)K*Q���w.
��8���n���Jūʈp�*���J�0\�*X��i
(U��	�`�jua�ŎH'.es�I�a���9"���P�ؔ�Ӵ��c��DB�� ��AQ��H�"��I�Dx\�DzE�Ȁd�l���BA�$|Ĩ�e�&R�8F·-�L�8<1�݌B���C���D.�2�Z�GX�a/�|�3�;��D0�L���gK q>�i���_%Y@����Iy�c�'Z+)7�޹@��ĸ5�Q#L���k�]�4�BֶC�*M��FO��'�С*:tydH��z�a�S ;*��a�ÊO�����!l�]�P��$��Dʛ��?�$6*���
�	I���:�c�$g�i��C�h�lV��P�J\����?��!�ʹb�i!uh��kD�3��k�h�SѸ'f�I�'Jf�L�e��H-^��0d$B~��96H�5\���Eabd�`�P�M�҄hN�T�(���,j��md��M;^�YA%5����^j$�`!}r/�,k��y@�!ρJ7L��eQ�v��8e(��(���h�JI;p�.�IQG΍P���oˌg��'�	���J!�N]'7!���Q����bl��'ӌ�,H���!2xn���'�n��!�|�ɣkv:�X��I�g�T� ?��H`&C83�U� �nP�p%�Y~�E��-̄�Q���6ǼMX_~�}��@�	f\�h&�?e�W�H(d`صc�kz�`c�$xގ�RV�@\;�١&G-?�l�G-)gg���@nt�J�#
�|ր��A��g�HzP�������ze�բO� �p������j��
4�]�;{~ �ņV�y*���cG�e���3��3h|-y �C8-8pHz�a�
8$�%��W�q:��R���^Qr ���\��؈Ф�`�@����F!;�:��u���ڑ�Ǚ�th}�Q�9L�fZ��C�	z�ݯ1_U��QG�ph��(�U554h���+sl����L�6�b<�2
ۙ��	W��� Ԥ�b���GA���";5��P�L�.�JD�ځJ�=�#	��ʀӢ��"AN�=H�D�#:4���/�I8b�D��Q���ŋ�>�v��;#"��k�;LX�s �:l?�3��C>��)��H�f�'�&E��l�؂}�tu��F)s�HH
$�JU��5��i�<b�EΓF�!��A��;)�|�SB�%�Ҙ9��Y Y�m��B�%>.��8b�̚G�O$��x/�ۼ[TfS |"�9���7��q8P�ҽFa42�B20Y �\�<�SD&�`�'� =b�+�+W��pWk�5�����#������Js�fea�*
j�j-R�+�_�ɜ��.��Hs��_��@�G�-[ɐ%����7@��� �pJ��C,V,gΜ�B2K�	
&����<B��c�Bή z�hط�#:,0�c�84&�8.�
�Ӥ[:@"��2��F��MʒYd<��PM��-n��/��/h��U�8ٮ8���;
о죑�֠��)	 K���F�N�~�D�I3��Y��ۺk��,��,�0۠u����e��|C�.�x*>x�dN\6�Hf��5�$����C�L��i��!�A�O1>��G�`0�#�?,b$%C0q0d�1�OƟTX�c� B[&,C��g���(RR�����-����K�#��*5�.~~���a��y�Ph)b�0���,A 	B�j�1ќيtk ZP��ي�61[c�,I��~���T։ͤ@���%�V8ňO�i�	�4�-U����NLc	�+�L�$���D��*"O��fdZ�q`,�@�+H��{0�O8���Y!�VQ�vo�<E�S�W'�-Cs�2~�t8u�A�!��dX25��$�'�	S�x"O���8�$4�|�R/b�X�3��H6��**}rH]�:�j�+5�x�K�v�	�֩�!2�tP�&�3��SuG~�8�#dZ���xr�F>���r�ӹCd��$�Љ7��M��*��
G�`ѩ�*e��Y�D�I�!�^�A�.#>q@�l���-j�*�S΂��qK�1`��3l�e��� ��;��a!6\O�hSFǎ:�|��cf��#��i�^�����0DB qwď�uU�	����H6z�)sdD�wE��aW%�:L|`���WYZ�Pk����iE�)�'ʹ�P�͒]��ɀ"d���Ra���������7� "�H{�4�3�a�$����N {�Mּs��c"|��
&|��� ҈���4 �p�b,�&d�h`�5gI"-��|�"oA�'˖dZ�)�^q��2L�.�`P�l�`�ft�e�� +��'o���"Ǘ���T�F��'���I��DO�,tl}���lͮd�!Oߞbc򠔯n�r	�@�[k΅BAVfD�ڦ"��M�f �5�yZlzI(�L̟#��+w�Ʌ8���ea� �:EC8t�q�@�f�0���Γv���kTD���Db�+�k�Ρ��W�H�6�8�m�b���Ɠ4����w&K�T��5��_��U�H��zb�sE�܃N��\٥(3�������U��!�H�Y��e̻b���p�$���h��� CH��I� �1�D�vu&��i
�Q���F�D�J�[7�R�����O�iAB���=p~21ɡ	��S��O 䨣==^�CE�w��i���	;��C�ԸQ���A�߆Zl$츃֑A����l�FZT�p�O�t.d1�@K�	����\]�ė|�(��&'�Y�O6�sD�\�.��y{��]�0{4y�F�O�}�U/ۙ���#)7���x���H�MHԠq�N�\2��V��ك�Q= Lщ��N���	�{��#���0|*�`��	���_0k9���G	X9A��0�'��I��O���Mkd`��������ㄬ��l�q$@�H�#��B���݌B�,ON Yr�Юv6D%>���w5L���޵h\l�	v	%0��`�>��Y��Fc�FX
�'��h'��l�AX妉Q(O���6MՒ"uL� ��Y<���A�;+,^5"'��P�ڸ��y2gD�R�Ь��#��S���,H!��'V����L�R�V6-�,j���4,p�*3��>Q�bFiB8�Q��
�^���e`0 �n���[�
y���1*
�Ç����ӧ2�/i�^����æ}r$	Er0T�8 �؜s�ԕbv!'F��d� 4��Ag��aiR)e>�(��p�ډR&�q��pg!�m{��� �g���C�v Ӧg��	�n�h�/�;&X��`w�|��'�t��Ü�L�5�v��K�l��d�3��`�"��0j�����Hu$ C���4,	�)�6�����iZ�{�
�}@���\�V��`G/pA�ц�L���	��Or�w��
�I0�U�Y�Z��4�'詐�����aF,�{��	��G�*�. �p��4d̬Ţ��x�Ծjψy��!��?e�����Fy[P�W=fs�K�C�n=���\Ժ% ��^�:��)��5�rq.�?��4:��5I�͋�1�?��>Sd��
�݂��t�%���~bnW�R� 8%��.]�|8꧋_�1�~#�.B̧��'OT9 "h�Ч�J��8�1��a�'熜��^�-�| b0��DH1\�D`�>tg��c2�ѲD���̉+D6���K�#��'S�t���t@"1zFωH�V���"�2=��Bmɬ13b��tk��i��>\��ѕG��|�Hu�v�d�<(�Bqj��3?0<�B���9���� ���`S�(3�m��	��j�9�jA2?6���Z�8�굸����X���� H�1HӔfm�Z]�I�h�`*�&�<EaN��*G TH4E���U�P^���b���8H� E�D�	"�����=z~
��d�	Q�\L P@C��̻��'��� %D�2ܱ�+N=��to�	>��U��g� �ZdxXH�'jl���X�3��`A#��E�0�T��_o�e@K~�a�� A����	�)�p!G��RJ�ɠ)�e��ڂ}~D�A�d>��P-�1 �GG弃�%�9-�8�qiG�)6��2��V.}�s"ˠ�h����B�,�*���,�W%�yYxE"q�J&H������x8�C �|���0�oyZx�'����Hks�t�Ò|�H�it�P�`�19s�ሕ��H���ãJW�l4�C�ݏ�e�'W���i��B_5������:(�}b��O(��ѐ@������]�P1EOY�d8@�� ����!x�͚�J�)y���� h	�_5A��썊>O�q�U��tkƩ���P�Y�ظ���Y�Xp��P�&*�?���ON�y�u'�L�$� zAӇ�?������
S�8�"SY����. $�Z��iH��͓U�l� D�@����U:1V��#��!����څCR�s��8c�2R�kA0
I�I����ܳG�.$�|���#	�AI�@ZSBܼz���z��ƛ[1��#��M%7 Γ�����M$4'�����'!�b嫴L�1oL�!�ρ�	��m*�Ζ?I��l�MG��:#E�N�����ׅ3`�u�t�@2�V�D
˽�vA s&&O5�	cmēJ����*�5m�y�d� �|�w�^�. (�UF�
y;0��O~X�DX��,�vd t�_~�$�5eͳG�U(�k� |�t�ADߏkP�4S4����%��FBL�ՀVe3G>�q�����02�Q�T�X�_�@�ў�;�#�"%.��sV�I�v(��4�Z~���v�<�� �`��I��Ug˯hL����n�w,��da߸''�*���=�����ףw���~��
�S�I�=��)�d��H��~�ک �(ͺZ����(@���Q��,��^h�˵��l��q��ˀ��d\�q���!�݋d�,�g�\#*����I�enX8DP�K��\�6�+1��]뀍S4���r��������<�|t�A��}�z͠�/\h<��N)����#���l��C�P6?)� �R.*;�n誁N�?�Y�sO�*�����'�j��#/������MJ��\���0p�d*V��r<��͍�ȐY��s4�pkCl����L�dkz�Y��s��`Ad�(�ذ�F�q$� ��xr�ּJ�Aa%G˛��9�@����O(�#Ve��)e.HKg�C�do^=���ӣ1h���E�R�OQ:�S��A>�P!*�F��X:i���;��˓I( ���H�M�0]I�!�s�*��'�0����	����p�R���=*��ӿMR\@�pO]?�2�80N�� xpP"v�IP��)!��i��a��(����a(R���NҠ`H�����>N�*1���x�,9ba�.� �c�T�R����ҢeR�ͻx�j��/�(>:�#�Z)R:Q���y�d��%lX6sjJe�T�
��ެ��JʻXƈu3�F�JH����	�����̙�uf^E����'�B%+`B�	4��1�	�6(z�-����@�K ��"fŤ9а�ɇ�N�Q���uN���*�傯\n�Ⳮ�:Z�>�1@m�dS:�j�E���<Q&��-2������	)�<mB�I�Ty�擢|/��ti̥IZ���b۟�q%�%Ib.A�"�D�Y��bvc��z0�X���]�A�����i($�$�5D�/����Ð� -+���[Kzu� �O<9���1e�X��D֗,
���G��1+E2�,���*�<vDŉ��JA��j�O(����R�*��V�������N�'f�$���!��}Y�o]?i�*R�.�$�6O˻��Y�лÃ��I�D�)��eX�4O
�킧ipzP�MC"�~RJW�t0�+Ƥ`��	Y&kD��?y�/�l�hX"6��0=	����|Ê)��b5��\�sbNC��E�k2n͑TG��|�n��Ci	�M��O�y�6`Za���^i�؈�b
�_��C�I?dK�����$A�䠃\&n��[���[�$��M5����,�_�6��Ν ������	o��H1BΗ<�!�d�m��US��7vt���(��D�FO��p?���	R�ti���K���jBi�<�r�R/-�Y�f
�O��YePX�<QG��'"�ei��AX���`2(�C�<	!�g�JSIP7!qʄx7m�t�<A1� ^�~QI���\����b�r�<��I�6K��%�"?%�Q�5h�l�<�P�b�N��b�אvkM!�b�<Џ
�7��m�t�ډ
w̰1�Y�<���\��E�\�$_�����T�<��T/�����f�T�8d��P�<	� �8}��`�"+A>[�);��MR�<�v@Ȏ�J�T��5^M� �ǍTk�<�ǅ�.9/6����8b�@�ѳ�HL�<AV���Blă��H���r}�\�ȓpu���f��o2|C�㘡V�Z]�ȓ1oN�c��=$B��c�M��ɇ�}S��K J?Z��*�'��e����Z�0t��L�r �O�C�H}��E�汛H�ex�� �F:d�ȓN@8���mL"���:4�69�ȓ��9@�AZ:cMDY`�P�U��ȓ�4�qDO�]*����I�D\�ȓb7��b�(K8R���ч̗6e-���ȓf�j�`�J�1<��1AA�Y ^��ȓ).I�֥ $.*�8��0*��Q�OBhʁ��)f[�����Nݤ(�����&N<�Hwf�.t�Ȥ�3�:lZ����M�@�Ů�v�e�3����Gŕ/�����g�P�B��٪�M�"��=���[��V�Y)����S� �ܣ�G�U�akA�)(�dT
S���J`��Oo~ĺ�cW�Nr 5���\D�2pN>���A���O ��+�gWil����M��6��,O�%���)�'$C~�� 잴S8Ui���D�����c�F��'f�0��L�V&4��AC�-��1# �Ί�O���I��Z���8">(�6bO��%�W�lŜ�ْ�i;F�:'�I�(j�n�r��)� �&a�73����o?i`'��t��ODp�*V�y@�Ks�6�A�^�"!_���d���|z��I�9Y�q�u�>g��ǀ������e[gyO\�fp��X� pvKE�\,ZfG��A`�m�)Op� 8O�yO?7]?	
�O焴(!�T� �%Q'犪8�B��/O��Upʁ�O�i�U�ӮpH� e��1ÑM����t�8�����)�'}d8�J6m��c�\Ah# Q�4l��d��2��>çA��07�RB�R��w[�t̍�*�S>mJPJM1U��pB�2K��0A�`�H�!�'�%�$ˎ���܈SClea��W��Q`���5���I�u1f�2��B���Y�D��ȣb��ؐ/V��<
`�iӠqD,ט�y���"�!��5%��s"��'FQX��D����IY�'��	��n	;��?��0���V�2BAS�]L�Ac�	�	�,��O�����������[�/����#�vu�dAx~2+�=����)�'��A��.+��Ȇ�T�[�~	��Y�^��M\ l9H���p�a���R�E��C ��Q�/2E�*ARAy��d�a�Ď ����d�T	o���۴�.�y2$��r+T������d4b	�t�T%�y2ǝ%c��]�f��^ei�7��:�y�+��Z�FP���M�\{�tKp�ؑ�y�g̈́)�|���Qf����M���y2�	u�ҹ��/P$�0BI�yi�2`���VL��Ɋ��y2[ ��'�� a��0�#��yR�?������\��dpS�J.�y�!V�6�x`#Ela�pY9cDX3�y���<�jQ�s��#�I���Ι�y⧂� %��Ү-�b< �+Z6�y2D�>-�x�A�����V8�y�cI�xq@`е�?��oL��yBm z���-R�W���H��y�&:���O��[�T��y�LX�9�Tix҈��]0�Y%�L�y���TQ�K4��%�T�Z��y��΍y��Yra�N�:��id���yb[�+�M��'V�Ae�m�2�߈�yr��,k�ؘ��.A�:lPز+���y�Ł?Pch ��ȃ7���g�.�y��̑^� -ɒDƮ	V*��j�%�y���c��i�"2k�܋��¬�y��2\,��tz|� ��y��0d������! ���0@��y��"6}�	Bw⁌)�ʥ��#�yRBܪ!+��q��$�X���yI�?��Y3�
�n$ �4���yB	�� ��z�IV2wt@id!%�y�R��i5�
����Ѳ�yB��u32��FZx�lYQsK̖�y���1��UY�eW�Y�V�೤��y��[�&RhqZ��+����R)���y�AN���c�kD��,�����y��J��`a�����S�HQ.�y�lQ�,��ͱq�F���S�����yr≘l�B(�Po����H�S8�y2f��.s� �h�O���d*��y�O0��(�sI	3g�r健��d9�S�O�F}���&<3�x@Ҷ>�
���'�2`�1�Au8-#!�]1���
��� ��#4 �,-[Xd���	~2�]�!"OV�B5��tW����!I6-)H���"O�I���8Jx};D�_/$���F"Or�C��"z�i�"��m
���"O<�0� 2�|3H70�2�"O�DA$N��]i:WN��\��J�<A#aJ�<���T�"ؽ���D�<q��1	��C���W�H8a�L�<�1̏@_ZY�AӷМq�q̗]�<a @>np١�N
��h�Y%�n�<1�iI�lqHm	��_�TCB� 櫋l�<V�iU�} ':J���k�<1���.:t��̅�
0J��"�Og�<�0�3�\�(��0c�&����`�<9�D�\}t�C�+o�� A���E�<q��P�������Qg�z�<A&��)%�0���L�(nԼ*V��u�<�ˈ�Q�V1
�@��(�3ԇDI�<�OÆ<�`pի 
Q�8�Ӑ��E�<)�Z9$~�C%䋬ws��[ ��@�<)�%P
4 +��)�\�qf�+m�!�T�A�y�H�/���ㅅ,rv!�dޡ��h)Q��[oz5�Oݗ!���$ ��W�)0>��Cn!�d�&zd�Ix�N�i����&6!�ā=rT��@�@
�:sޡ�M˱0>!�[��6|�	Y�$k]�����!�D1����bE#hE:��B(�Zv!�d�P2ru��� w)�L��&Y!�DYҜʁ ѮGs� ���ڤ�!��1f���!�ڲaoz�3�cT5�!�DX���L�&�˻Df�%��W�w�!�d�>)8�p隟mK�W�� R�!���8[�lP�d�ԥ?�yR���!�ơY/.�5*��s*R�Cbp�!��/?���WV<V�!�=�!�DA�oɌ���N�3D@�H�"!�d�	K�)���H��J�k�9L�!�*GŲ�RD]��Pj�gF�o!�d_�,�d�J��r�\+�&]3�!� "LQ)�eB$-T&\{���F�!�d�X��`eT%\&�1T�֋P�!��[�K<�c b�"E���C"O�!A�ϭ]�hT��`)i�  yB"O �:��9j�K� U�����#"OZty�G�x~��U��C^2���"O�|�4 �Ji.�A��2F��#�"Od}���$�m�B��u�)��"OQp��V!k�:�w*�'V��+&"O����jL�+t�L �f_1ju���"O��+㧋 ��`䤜0e�`G"O�Ia���)l�ա�h�Sb��2"O����ٺ7�n�-K=D����"O�P�rh��d)ݗD����"O�]�uoX�ZUr}��a�E��+�"O�\�3�

�,p&��jݠ1�5"O�lW#RP��H�v�_�\Є@!q"Ox\�.�� 5rU	�2~a�P�D"O�00 ��R�J��tE��oH�XC"O�-�a��Y���#b"��E��p"O�5c��
7b�kơEi-6]	�"OҜ𥅚�o0�R���/U.����"O$m��iQ� >��g�U����c"OR��g
.1�TI��,��D�`���"O� ``h g�-��`X M�g,���"O\��S�B�#�Z�c��ɦQ�@�t"Oƹ8�˔9-$�e��ؓ	�Pq)�"OL�be�&&�3�-D>6�ٙ�"O,��ER�s
���0��-MD����"O�������	@܉t8 xy�"OP1�f��k�ᗌ�D#�,��"O8 FOrS�d�L8ynР"O�@�1)��u&�R��=���`�"OJ�ɦ�2٫ ��ZkNܒ"O �`/U5�6T��)�h1�SD"Oh�c�eF�DZr}PIX�[y:X�"OČ���L@ i��
Z;���#"O�U��)ڻY����=�m��"O~�k0H�i��-�N�X2v��ȓR���Ӏ=� �Ҳm&l~� ��y�d�R#��!<�"Cf= Z����_�����N�K"�"�E~�ꩄ��jX�r��	��l:����za��Uu����c�֬���P����ȓX�v�T!ZըIwZ���z�<��F��#���7B�dCP8/�r�<�&bļI��=�c�L��@��ew�<�$�=� ��4M�:������q�<�5�sP����E	Lı���Q�<�����H��h�%�9��M�1�t�<��o���fi�5[Қ 9�r�<���d��A�S<>[�hӱL�Y�<�"��R4l�"�):|zY�Ũ�T�<�%�N�X��Q��8:�D��)Lx�<� Ė�-!ִ+wLP�K'��Z��Rv�<��Ƥ "��GF�<	t	���g�<Y1� 2��f���p!$�d�<9�(ϩN(��؁��Np����i`�<��F�@���1ȔU ب2Jg�<�3 ��Ƥ��IL����E�a�<AVl�7�&�#�/טB�4�XB�G�<��F�p����aǽaX����B�<11A��F�"�� �Ҽy��i���\s�<9����&axcHG6Valq�!��o�<1���| �l�O�l�V���ɝk�<)dM�RJ�B�Bq�Sプ{>C�	;-�L����2�qr���=|D�B��y ]Pdʓ���i�g���{rpB��Pv�	:$a�bbPMV$N~�C�	)E��[0�
�_?Z�&CV�s�BC��@ӓ� �9��#u��4>C䉚Q�^�!gч	~�aks�U�B��B�	�5��%9��Ҍ(�rb�ȭ)��B䉳�j))u��~p@9��C<L�B�I6��J6b��=����BB�ɉ.�i	�H
��tC��Z�B��22� H���)vx�hK��I�T%�C�I:3��-�-^�5�t��-+�C�wlRʱ��-R��� �Z�B�ɛX6�X /
 ����C/�:g�BB�v�`�2��;A��`"m"%��C䉻}J^�@�O�Ъ�iee�!"�C�I�y�������
N'�E���F	`C��&¶��e�M�q9�9�fLf[BC�I�7��y����O�����-�B�	74I��{dj����>B�I??��)eG#z8IC�2f�C�	w(� N���$�˕o�+/0B�)� ��k�CԘ�t�j1H��\ɸ�6"O�It-�3m�(��m�W�F!�g"O:!�sȝ�4.�ST*C5g���ض"OXt{��1wc�1��Eq��4ʅ"O����5�ZI��	��)�J�I0"O��(/]�a�,L�)8r�l(�"O��p�i��z(����ǋ� Z&͑T"Ot�2�	��YP�
q��>����"O,	�V/@xr�	���M�(=�В"O�����!���u,�?G!%�f"O�ap��?�� C�+J�w���1"O��Q+��z!Rx����7\ 	��"O
�� ��H�/>=i��"O8���C#E���A�@�G!4W"O����&U�=��BD��&"Oh���>7~`��E�T)��Ex�"O~����Old�RF�@�	"O4)�EA?�~�f�K�3�J�d"O�u{#f�H�.|�E�B�e/L��"ON�	2��"o��}T��q��@+B"O"x�����W_���*	�8�0L�"O ��P��*�\95
� �2mj�"OXQ�,�*�����#D�I���b$"O�i��&�}��B�0y6�՚Q"O4M��j#.���Y�o۰Hv���"O����l �,TnTz��b4l�J"O���M�,%`L�UmTx��y���O�Q�B�MӍ�	5�,Ԙ��N��(�s�b� /��?A�k˱50��
� �ަ����00�Ye���/J�,��ejK"&���pSN�W�N$�C�Հ0����K����H\���§ɖ@�Wˎ0y���U�B� ������D??,"*~�̉&>��O��	�У�'��v���_h����)�gy�eU$�P�9��T$E�p�ŕ*�~�F/�,
�֨w�N�/Ўȃ��D!��,4�1�����/6.����e�R���<�'������4;�����H��˔%��x/b� ��D
X.�h�'��v1<a���G����㟰ĳ�w?b�Z%��! %T)㰌N'%�,��X�E���"���<� �+a�Ұ#P��Z(�:�ħ[.�.@$[�`�砓V Hp������	8�M���>�1,�n��?�ݜs�<xK��U�(�Z4I��YΎ�a���>�"�5N2Thb�*��?��=j��t�.��<��i,�7m2�$�����{�`=�ae�Ib<Z�M0H<�C��ON�Q�#����æMr�G��؊�T� $��a��93�����Ţ,�e+C��)XLz��сu����?���C�T4<���-*��`�Mɞ+�Td��GC�Y}tm�!h��Dx��&|�������'(�-XU�0{�@�֜B�4���4�
M�I��Mőx"�'��xrb[�cB��֯�q.�f�R�1'£=E���v4��˙0hr5 ���qQn�t���a�	7�M��'��I��4|��m���h��֭[�n�TꟌN;�A���*Ol����FW�=!�-˴<���桙�8 b� @@�.Gd�Gg]�$wFE�C�5�M��$Ko��aY&�E�2.�)�ځ���M�e8<Q�g5M��([�P�O훖�ĜޱO��8�';�7��%���
����~��ÈJ�(����_�d�O��d:�!��������A�W^޽��
�x��B�I�9�P(��δj��fk��i���8Ұi�7�<!�I�5���'��Ou�nЧI)<�O�쒨B�iZ�0z��?Y�!���8󧯈`�(��ć]�a'�M���B�?řq��$�j;eKH7J �#�K+�	r��y���	Z���
6!���1�'=3���!"C��	b�hma�-��'@S��H}���0�I�~�bb�5@uS"���<���Eڳ.m�O$��<I���:+]n�P��|�:�!���J?�����Ms��i��	Q����,���Ka��uF:�'�Lk4���'j�i>!�SV�q途���O�i�"	q�-
�>kfQ��L*�԰�*� N�|��3�Ҧq�R(�ȟ��I;�y׋�.pV�H��O7]���)�>$+$��X`X�$��(h�*���,@5IV"��M|��3ﶥ����l��#rhݲ!��9�c�ş��ߴ_R��(��"|���2E�&*B	1v ��H"���"S(SΟ4$�T�� d����c�GYP(Dʏ�|9���ڴ ;���	��x6�=Z5Ь�]z�Ye�4@_���'j�'>d9*@ ���   F  0  �  c   ",  �7  �B  mM  �U  ?b  rm  �s  %z  {�  ��  ��  >�  ��  ğ  �  L�  ��  Ը  �  W�  ��  ��  ��  U�  ��  ��  P   	 : �" l, �3 : X@ �B  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d&�@ƹi�l�ç
��v�F�7P�-���Z ���o#x�0qC�i=zA-�Jj�����d�����~&��;�Lӆj�0iIq��
,:9r',9D�`�� w.�ʎ�PZ֭Ŏ68�0��I��)��їzW�TB�Лb\2��Dg��!�ɈK�^��V&x�d��"O`UI��l�����cӯp�B��@�|�_����S�y�6Ń����X��R��"0 B䉓X�Ĭc%넯e@q� G�/*�	b؟��n�{�8��
 	=v�q�FM/D�<%蟗\�aA��\�;fy��D,D��C���?��<q��۷=�Va!E7D��7�U�|a�AT����uj4D�T93%��|CN%���ߘ&Ez=�`�1���'[1�0�pm�&k��!Z�- �Q��aB"OzY�ē�Qxdy0d��f� 4ZV"O�ɉAKU�?&ԂA�5y��@�'51O�uP����U�͘ր�V:�)4�>�H��ቭ(0�B��çu�eYDث�����ܫ��$������<�������, �ҮCA�R�Zq`�����K��N�y���t����#�Q����hBY�2"^�|�!�@]����jM\BCo�,h}r�'���YDx"�>�V+�#�QP R�EY���q� rN<!ҡ�,����K,D�x�&H0"�!�8|:�l�	-���R�GF�M���Ȍy��� j ���ܤ-FuJs �j�u���'Nў"~Z��	p3��z��S���5I���v*�#J�xI���M�!�<�b�^����FƐ"J|�ɜzda}r�X]m\��j��z������.��t��D{�'�d�i�V�3�n��;}��� �НyO
ԅȓ&����-�4���*�������<����=����OPNI�i��0����f�UΪI�	�ua��'� �y�!�'!13��	Z�Fلȓc{VQ�T�L�$�s/�eY���l��И���i�0�j��ڇ>�ꠄ�Y��AB�b��ƩݮX�x%�i�ў"~nڪC�j�gc�(t��lA�_�|� C�I+%����2�F&ވ[w�ǲg��B�ɳT��P�-�=��� Ԯ�A� C�I8E��b��rU��� eؙK��C�	�AΜ�`�*?�2@�C͓�m�B䉄lH���P-�$�"���A��C䉝�n��U�6 ���ƂV�X{pC�	��Hԑ�b��U�C@�	k&C䉲t`�@�!��OF�a��N�4�
C�	,L8D�G��l༹�RQ�x=�B�ɜ�H	�Dϝ�u���3�/$g�B䉣5-����+ cLp�1ҫ�3h�B�I/=��`)Y7&�n9�!΋8v~B�	�	j4Q&��C�buc�$�	5�C�^x$���
�xIqޯ�jC�I6%F0}q '
�E���d6�hC�	�B������BL`� Q
�<o�L���<�`H�$3P�y�p��p���JNn�<I���`�q�&��`tQ�Pf�'M�?j�-ؓuj�d�0�O���(AJ4D����&ĿL�F���*�fT�5�2D��i��Ǉ	 H��O? �Hd��1�Ol�p�d�+d�G`6�`�]�N�����s���Ī���Z���G��"�a.D��v��-�~�� ��^�
H��'-D��8בU�B�; �1r�%�Ы8D������t�@��a��I��	;T�C�$S�ws0�hAR���a�k@TH2Iz�'��@�@ꅆ[��x"�a��'%PD{ߓ#�Ya�O�i��^8���8�E=|<x8jd��.ړ��Gf2��6+�&� q9J��� Gyrh����D��ap�z<�P��s�ЩV�NqC�I'B�)2�՜WUt�1O2w���D ��?i���B8�f�R��"8�f,��J�!� R�hZ2bT�d ���!�qXa{��$U�*��Qc�d�-��!B��	fga}�JyBj� 8j`=l��a���'uў��@AҶo�8&Ҹk���+]jd�剮�HO�S"[����R�Q%BI�ҧ�*���F{��9O:!��M� �����)�̉�'��P)�pUM����	�> �Vn�h�p�'R�s�'�]��P��7wH������8�Á:	�T�{փ��L��`E|��/Z�8��N�9�&�!#�X�~�x�q�)�i�89�6�e�(tb�@5k�MR�)�it�)	恇�%V�s��Cw"�)O���dהfNL�C���G,��MM.w!�K�E�vT��D�*�	*f�Ja!���l��9g�Ĕ>�ȨbD�{&�zRgG_̓b1�)��}��Յ( �ȓg��AA���]B�-���?Mx}�>q����$���QY �F�7z`�CT�7�y���O>@�1S�ѢE��0 �.��y
� ���	�H���0a�I/��8��"O�M�ƉW%=ĔyU�ܒ6i��i]8y���5:v�)��.~>ehS��cBB�I�"&v���n�h�� �ܫ�"">������V��@a��'k;���@-�0!�\!f>�����]�/)�� -ɸu�!��]�/�r4��ȏ5F1�U�=^u!�ՠc���ƉI
c���ū�H�ay��|��'%.a����),KX��eO�*B�XA�a/9D�\��
��!��R� PY��5�%�?�VAu�n�	:�-�}�"N6W�x�KpC��*.��jP�k�'a�d`�0W���g���]�����y27�2��?�'�T�Y�*E�xg�}�m�Em��1�')0�	��^�OaH�D ��4��	�'��zR'3 �����
>MhY��O�EX�
پL3@5�`��Nz*U�"OX52*W�\��}Ȅ��VcDh��|��>y���ۺutE���f��@��"W!�DS�6�pi6�X�!t�	�fٷ]'铇?Ɏ�����R�����i�Y�#!�ˁ:�>��)�vxP�Ҥb�-w!�SgjT�q��-f6� �/,�!�xD�4gח*6��«ļm��؇�UI����
��u��)p���l_z]���(O�=9`�\S���!W�M�|w�䫳"O�e�bo
�s����� "`��ё)�O��;�S�'Ҹт$x�.��Ag�T�݆��?)ƀQ�1ZX�Z�,��r[�yC�� s�<�Al�0f��` '��f=3�[k�<�ЇD�7����JDm��r����xҥ��r%B����Ę�B%ɖ�y��U'�tՀb��"�ؔaG����y�E�t�4$�t����l������y�⑎�L��L�5Z� �@�@��Py�Cȋf�!Gm՝k��cug�f�<�Ƌ�L������� m�<�O����A�J.C��l��Ms�<�&�H,�bp�����C�Mx�<��˾r :�[�dT�@L�uQi�<�%��3���("�\��#h�j�<�!�T�Q�d�C�"� MD�y�u�	d�<�C"<P����Z�[ 0�����b�<�@ÐB4,@�t���@�yӈ�c�<Y���A��ґ@�{s�EQ#,�f�<y���c�)"�A�x���x�o�{�<����#d/`�Z�/�(�Rc�a
t�<1��ҙ}�a��熁^	�I��W�<Y/V"z$�wN3����Ag�{�<A��3}���걉�H��x����S�<�eeN]�&��ǩӟ,Pt��#h�<�ဿ���p�M
�z���k�J�<��S��u���
t�����ZI�<�6J��BX����$��+�C�<�᧛i�2���
SD�ҫ�~�<���r����@	O�fK`�h��Ex�<6�o�t���B�[C(H	ƍJ|�<��j]%P��!F���6>���URQ�<�ciȊrB؝�uFS9d��/�e�<�q
�{�Vű���?�J��í�b�<Q� 
s:}�׃>]��9ȂLA[�<�'אt�p�q�NY���*�W�<a�a��.Q�bH8h��}���Q�<1���=B�(�Ѥ-@gE+�AJ�<q���8Cd �P�+r��
r�M|�<� :�P!c����蓪
3J��l�1"O�t3���Bm�H��ER#�C"O��#D[�(b��I��(�f��"O��AbK^)����)��(�RH �"O��TکgV���O��6�: "��'��'�B�'���'1��'���'��k�)�$j�}�$A��L6N䪔�'�b�'R�'n�'`�'&��'�F�"G��??ԕ�DO�8�BL8c�'�R�'�R�'qr�'�"�'���'���	��y���oѵR�֔P��'cR�'��'���'V��'"�'0�UC�t��9c���<���'���'m�'�2�'���'2�'���vj^41���Q@�a�ԉ�'�2�'R�'���'�B�'B�'���Q��]�VQY4�^�s��u���'�'�2�'"��'I��'5B�'��$D�f�p!��b�LZ��'��'w"�'B�'��'T��'�����J	M���〄�vy��'���'�r�'��'X��'���'oT�[U�x�t|x7#
�3�r	��'E��'Lb�'��'��'���'�ph�(Z�qN��ò"ƴ ��9A��'�"�'Y��'A�' ��'n��'�U�W��1�i����`P�'�2�'�R�'��'r�':��'�tH!��ɼod��3�FǟM�tk �'v��'��'�2�'�RmgӾ�$�OhE�&h��&�I�LU=*؀�jcMDy��'��)�3?-t��(=/9H��i݄SR�����(5�2���O`�o�~��|�<�6L����Z��@������b67�O��"-kӌ�EU�  �� p.�O�6� �M^t� �
���U��y2�'���l�O$���V��;n���g�*
Lb=���j��t�5�$�ӫ�M�;������w2�T#�J�n(�(aƻi��7m�@ԧ�O���� �iv�N�Ui����
�\Ԑ�ϒ�q���ߙh�p�@�
ŌA�.�=ͧ�?	���JbsnQ'B@�󡦃�<�)ON�O@|l�s�2c���R���d?5�Cj��PI���\��x���4�Mkp�i�D�>�bτs���e�ua�����g~R�ڍ1O�M˖�1јO7�e���De�	+�<�)W�.P#������4v��'���͟"~�2��%aې/����D�͝��ΓV	��&����㦱�?ͧ,�1Br&���0R�K�M|@�Df�6n|�~��T� ip66?��KD+Eh��"�#CL�VC[�U��Q���/	�)�ScJ�YGV�#v�.UX��R���2!�D���P0x�21�D��;!��I�`M?Vvp�Q�#�l(��M�������+1x�!�ǝx��A8��
b�P���8a l�f�P��`8�#�Fn�;��!?ʕ�$�ŇP��- D�]3%��Y���ފA�t蕬�Hp��3#ɝ� �]�����D����ŅZ�rڮ��Pl���6mA�'���dj� 1` Bf�>����K�F�ˆ�t�p�A�
�}#����&Z(O��3Э̃T� ��ǂcXp���,8�:ؙv�-��i��jg��D�Ol�����'<�mV����#�)-��B p�$�D�O��8��)�S4b���*F��ȓJ"H�6m�=T(�n֟����������|�S�f;�`$ʽ9��\�EK��G՛V�&m��8���?c���I�%����ۥ}�@�l�W�̪�4�?����?a֬ː-V�����'YR���\������(X+�-ԮN���?���(�`��<����?��E�$9#c%�8��!f��&g�z] 2�ig�ؑ9,*O���O\��<)c�@�)��%�EWQx���Ҭ� 8��&�'��qa�y��'���'V�ɽ3�����+6���Ҭ�ci��@qAM����?����?q-O"���O�uRq蔌Dv4Q��H�j�\h �#��q�1O
���O&�d�<Yd�U�h%���FI�;g�B��̈�׻;�	�����ܟؕ'��'E�0���@�����N�0��G�
�<�Y���	͟���oy��(����`�!Z���ہO�>*���a�I��L�'&��'��Î�/	x҄;�-Жĸ�_>��l�ܟl��Vy2�>�n�����k�:;^����B#􉋱M�-�vW��	̟��â=�'�nڱ_Ґ��Fɜ:WM��,W
6��<�v/Y������~r���j����c GՖ|6��{s��'
�&�V�j�����O8�j�&�<�O��L<!H߇����ulܕ^i��+����\��M���?i���
�x�O�>�X�/�[v���!�k�z��#�rӪ�A�@�<����?��g��?Q��Q3-΅*C�
0|�	��듯}��&�'dR�'v�TZ5�4�4�n�$�O&��._I�Jq#�-	fY�`}B�'X�����'rb�'T����#J����̂q�r�#�*jW�6�O(e
`O�N�i>Q�IP��g��i����.�1f��&��O5[���O����O���Z��̈(jF��Do ,~����(c�'"�'*U�����@����;?v�irG�o�hq��C��c���Iϟ��	_y*Z��
�S%P�p��=��TE�R����?���?I.O��O"p@�\?���m��J� D;΋8$^L�x�ˬ>���?1*O����f���'�?�6���@8��<8�����O=Db�f�'�O���@�_�-���x��%LtKwKE<M��E�� �Mk�����O��6#�|���?q�'PK&�ؐ˂�6���B3�+sx�EH����Ot�ò���t�1O�3� <���M z������;H���Y����8V;���	�$����X��KyZw��i���"�L����#�F�p�O��#L�2����I�Ɖ:�!��Zu�����/w��.�[���'��'V��X��Sß܀dc��B�,�p�6A�0A��MӀO:䐨�<E�d�'�6��FRZ�`�B�Ͱp2��c&hӒ�$�O`��Ny����|����?��'H�=Kgeȱn�~�0�B�[l*%�v� �{-�O
��'��ę�:����p@�$O�E�#غ-���'\H=q�U���	ݟ��IRܓ@��P��b��(ۗ&�6z%�̫A�2?���?�.Ox��=|Y$}��>M�p��a�3�p+�d�<���?����'#�%�*���X4j���#��}ÛV�������Ox��<��.�l��OT:= D��! �Hp��Q�z���4�?q���?A�"W�Xj�Jl�ĕ��`��&ː��c�ɔG$�P����؟��'�0[z�S�\C�+�0���xV��vϺ�OL��M����'���,	0DO�p�� ����p��o#:) �i��R�|���yL�ؖO+��'N�tJ�A���U쟽�j����5�"b���I>G���B�`(�~��iGP��]�A�܆'��&kI}��'G�e���',"�'���O��i��
��4]p��6�CqJ1����>���V�p�e�C�S�%H� ��l�9Zh�Ţպ�m�5>�A�	ɟ���ן�Spy�O\R&!sj�u�wa.�>�"P8��k��U�����1O>Y�əZ7N��f[1l�n����>I�%qߴ�?a��?��@>��4�j���O��I8B��P�'��3,.��*�?9Xvy؋y����1��� ���O:�ɓj���*�f�%{bF��7�[�u�v6��O�i�4n�<���?�����'{9��O6�8��.�4�\�!�O���e�W�v�	���~y��'�.E(�f�2j9;R���cI�Qm�1� P���	͟0�	D���?�g/
�h�l� B?q��|�!I4m��s�y~2�'��V���I]T�m��9'�5����"���愽F�T�o���P�	���?i�~RLe����Ys"c��r���զ\ &�Ӵͽ>a��?A+Of��Q�z�'�?�1��0q�|���W�6����c��'��O�$^}$��!әx$P�?X�Ĳ�(�e���V��M����D�O(e:B��|j���?A��V����ډԂHJf�N1R��9�����O�b䡈��1O��B��ݩG
;;�4Mʡ�R�?�n��?����?���?���_w��iݑ�S��d0e1 �LF ެ���>)��p,�@��Ra�S�'&��������T�
��ܕv2FlZ*4Ϫ!��ܟ����t�SVy�O���+z*����p.(%{��[�g��6ͅ*v5d�����S쟄����c��T�� �9N�D��tg��M���?q��hv�8�/O���O`�$���J�@ߌ6K��y�ƛ8
ƨ�A�O���'����p�<���O~�$�O�f.	�5�F���F3Y�j��2�����	�0!s�4�?I��?1�l���M?��[+#�p��R�߫	
|�oɼ6턔\-�=8a0On��O����O��Ħ|�!%� *��<i���1����Q�RY\b�il��'�B�'��맊��O�I�q��9�|<�	C�4�����.�1����O4���OV�D�|���z����i�ȡ�Ɲ+X����SO�2P����|�>�$�O(��O���<��brL��'2�8��� a(\���7�2r�i���'`��'CB�'.��Kd����O����/X>t�V]�V��g��q�M�ئ�������cy�'�Ȥ�O���O��A�`�8K�:ă�Is�I$�i�2�'���'^��Da�.�$�ON�D��p%��������P'ҿ������¦���y��'�јO�2�'s2� ��MSѩF�eĸ��1d�;T�59������I���U"�M#���?�������?Q��Ԯms6M�CԮ:�=�b�/o��I����՟`�Ivy�OV����	(k��`�1�b��m�I%Puݴ�?����?�������?���m��#��e��@QS�J@g�&�i�6�!��'kX��r�S��p�r+�+E��puߗ��t+PN���MK��?���,��}�G�i���'^��'�Zw?��x�J��Vl��z�"SSͶ<��4�?�.O�)YC0O����	Z�c#Ԣ*	����N͋S����,ۦ���>+�Ibٴ�?9��?��A,�^?q`KP�+[P�Awi�F=���dDZ}��Z,�y�'!��'/B�'p�'f$���Ɏ*���ů�B|-����u�6m�O���O��$_S�T_�(���u��B�&�1J�pL�DAB�Vݔ���g��'D��'��'��Iʶ/��6m	+@02��C(V�8t�`%+3�T4m���X�Iߟd��ʟ��'|rdF�����\13@�C�"�!�Wq87m�O����OF�� g��8ʈ7�O�D�����ᇤ�u[	�4JO����i���'�RX�����"s"����)�P����v���R���

��o՟���ӟ���)L^���4�?!��?Q��<T��XU!U O��	B4���i�V���I� ](�X�i>7��|���������xb&ǒV�'���9��6��O��d�O��)���Ā.[tt<� ��hw�I	�LE�j��'��+�O+��';�i>���&\J��!��
*R�_$�ױit<M�)b�j���O�����H�'�I�0B�a��ݼ�t��-�	%z�i �44���?1)O��?����� ��BbEO�訜j����so�tj��ir�'�2RD����D�O�	"5���O�kM>��@���7��O��C�XI�S�D�'��ڟ�u��X<Q��;(�||�P�t�i0�ϕ4x?7-�O��$�O:���`���OP�&�VF�6(� �4 r��i/�$1�f5�yb�'���Or�'��'4ڈ�R��#��!�EJ�u.ه�	%-Z6��OT�d�OR��GK�TU����,14N}��+ }~��a$ևl�X�v����ٟ��	⟸&?��ƍ�M�4�ĸ4�B��I("�l���� =���'�2�'���'`�ԟTC��c>7���I��ň6Ɛ;2$"��3GW�y��'�B�'@"�'��#Ǣ}�N6M�O��d��J�j�b�bS�h6�9��ڗ���o��,��󟠔'��옣����'P�D٣r�t��3�(�P��ݘw+���'�r�'��#�1Mf7��O���Oj��,J�NA	b��D�Г0*ܘ3E�8l�韄�'�r�&��4�'P�i>7-�; �.![�N݈=`�K��[e��'j�JJv�6-�O�$�OB��������'g0�$(4�Qn�ܩ�0OCY����'��H.E��'D�i>m���3J����'� vޢ��w��Px�X7�O����Ox���b�D�O����$�\��CQ�v����
�r�:�o\.�,��֟D������D�'8�˅d�!=ؠ��KSQ�݃ +~����O���Z�x��o����I؟���֟�]�W��%���Ԉlr���!%Q�0��7M�O���/A���k�2O���?������2�eF�.DJ e۪M\�z�`��M���nx�8���xB�'�2�|ZcP�q�'�6�;�bפX��q;�Ou�E�>�$�O4�d�O$�$_����"��1MŪ�ȝ�h9"��[�E*�O��D3�d�O��� .l�0A���� 4�h�aS.�:8
Fm��:O"��?���?�(O�hR�a	�|���\�re%_c����s�m}��'���|��'����ymC�OG����9Ps��ؗ��9+P듂?1��?�+OX|�WkSX�S.L.�@7%T���q�j��M�M`�4�?�L>����?����<�L�h��kH�6�JEr��9w_r$�b����O��d�������'t��j�F<^Ě�e̳�.���J^듭?���?ٔH���?�J>��OXvlX�)_�t�2(b`�؅BC�u��4��dT&ьn�;����O���Ga~���%p��ag��25Rrc;�M���?��5�?YO>�~��H͡l��4Cr(H�f�\�Y��¦�7̔,�MC���?����RҜx�'n�������n^�tʴ��b�k�$��e �OޓO>M�	o���fo�MD����h����	�4�?���?��'�?C"�'3��'��N� /%�D��U�ⱨ4ȑ�*�f�|b��{T��Z�D�O����7�\=:�eU�Q�	��e�1��oZ럼�����ē�?q����k�P>p~��oީ���:1�|}����y"_�����&?�B�.r�u "1G�(U`���g�x�:O<����?�M>���?1��
�p)x�*J�8f�0b"�A�6ɦ=I>Q���?�����8 d
)ϧ9� �{����Rի��>1b��'^��'��'_��'� ��'������{6���d(�PJ�>���?�����+aڶ�&>��G��."�0���L�[S�����M����䓵?��u��m�����7�1�5���w�h��U�p��7-�O���<q�J�o�O�"��5���&G����h�M�9�T���'��MߓE�b�|����F��X!�qyf�,�R9�c�i��I�I��$�4*������S����k4�������c��E�	�T�+E⟼��K�O�d���c�j,`%� �Daڴa6	�V�i9�'���O8�O�	�U,�4ɒd�;"�dыY��l�T�&��Ity"�&ҧ�?�Ӥ��k~��H�n��l���I�̴(���'H��'u6�1o%�4�h�'��yJQC���V9ے%�)1���ٴ����O�(�V'�H�����	ޟ|J�Y4�����`�& ��Y�tğ�M��];68J���?��P?m�If�	4�
@�@�;鈽�ǔ�I��yq�O���'
�GY��۟��Iҟ��'��06CUUf,�	����ȭ9��ڄi�RO��D�O���,���1r��fY��J1"�푏Z$L��N?��ߟ\��ݟp�I��#c�}"E���J�3aV�S���qw�U���	ȟH�Iw�IȟL��4MY�AQ�ec�d�H%d�-l%��0c�0[4�2%[�`�	џ���iy�f]0�f�T	��1O�X\ɶ�F�i|@�@O馵�	O��⟰�Ɉ]�2b��2F֡u�Y ���&~4�c�s� �D�O:�QSxM�6��D�'v�D�5�p�9�|�%��$ �azJO����OpX���~�$��1.C�P���Ӈ0-h�k�Ŧ=�'i���@aӬ]�OV��O��6:Ĩ��I
V���pJצB:�n�؟��	<+$#<�~J "�f�֬��@�"C̖d�p�^禵�CmY(�M���?����ʲ�xb�'XxQ�B�$x���� 8��0qӢd���)§�?A F¿j�<!�@�[�:T�4K6aZ7jӛ��'b�'�)C�:��O�������2NŪl=~aZҍG60&q˴�9��&iBc�t�I����8鬌��^�\]:Tzq�BbD����4�?�t��6,�'bB�'}ɧ5��'`�(�6W�zi��Cɬ��$f�1O����O��d�Od�w�? ��b�a 4�1f+��P 	B��/���Ol�$�OZ�On��O����+�;"��a�@�`Av1�a��1O����O��O����*�Ի.��sA@�g��a���~J,Ql֟�Iǟ�$��	ǟ `jg?V��!h~)[��T+'T���a+�D}��'���'���'��C@Z>�ɳ)*l�2
[zp�.*�XQC����IJ�Iܟ �	3q��mA�e(�$-��ݻ#�ѿ���K�As���'@�Q���P/��ħ�?��'w�D5�S X?`��RP�Ӏ!��v�i�O.�ڄ�sӆ���N�Ph���<d�( øi7�',�A+��'W"�'��O��i�9���$�RyB�2[*<#d�o���O��	Q��:{1O���x�BL��v
0�@A]�]��q�i�����n�@�D�Ol����%����b�<�z��� J��P�a�7m��Py�4s�HYDx����O =J��؋A��L�G��EK: ��	�����ݟ��I2c���L<Y��?��'�����G�����wm�+����x�ZĈ!�<!��?��q�h��r���d��]+�c/p�����i^��F>a]xO����O��Ok��{�\��� h5�e���ߟD���2�hb���I�����Ly"�G�gjx�!�Q�6�"��k�OT��6�&�d�O<�d>�D�O>�d��w�|��c��t>&��Dx>�a���Ov���O��H��I��6�Pp
��^(X��b�cU~e`eX���I۟X'���	۟|�Т�>��eϊ#���Q	�.�\D1g�_}2�'~B�'���-& ��I|³��^�4p�
�2p��0���W����'>�'���'�����}�ڭpݔa1��(.�r��T�M���?y.Or�:Q�x�Sꟴ�өpo�]��X�ZU��ѫ�i�J<���?�%�Vn����W�#���УLD2e- Y��O��@�fT���h���M+ T?����?���Op�z��}8$���C^%�Ӽi���'\�X���)O�0�v�96��ؤe�P�V��1 7�O4���O��i�`�ş��v�k�8�ьL5	Cxx�@��MC!�@���B����$]p@I��PL��+�g'bxl���	ܟ<��ş��@���'�D��^K���iL�*~�AAg��H��5Gx�&!�)�O����Ox-�冟!��a���g�i�������	Lt�X��O���O�R�'����%����6(��1�e�M�7E~��'���ᵜ|��'���'m��'������*Q��	F�*g��]����'�	`y��'�'���Of�C�����8�	����m�(�(Q�i7h�H�O|�J�ˬc���M��6��7�W�~T��ΧDN���B��ޤVkR��8�*$�����p�h`�>�4�=A#M�k��9�a�=0���"�
�|�Q6 ۚY��"�K�4�������9:tR�8��$��#��
 =��À�ؑ߲�cM�.8�F a��'�My1�><�\퀥	�O��<tIԮgn��$�U��p	t�̷H���q�b3:Đ��M��}�>�jO��!
�h���MڟLIslC&
f�BV풵�$��f�ןd�	�M���Z�F�9hIL�8`j�c�1cU͞(7lH �OK4���j!od}q4K$h�
�N������;~�@���H=g��mi�d��/��?Y��L�2_��r�E�`CC }b��?���i��#}�'Q��p`@@p�2s��-B��8�O�x�nK�y�J$Ȇ$�^:p����'��"=�� �#*���A�h��+Z���DZ,*��V�'��'{�V'��AE��'7���yG�F�pe֌a�%�47H\1C���bE�� & �z��
�z��2U�|��
:e`��aA�-�\|!�$K_wd ;B L[oȬ��AhT��a�J"2��'?0�����s�%�う��T ��Ԫ7iz�8DO��'h�����|����$n�e�%Iժ&=@�hd!�s!��	0Z̰�����b�NI��@�33���On�Dz�O�2S�;����X,�' �� ]Hѧ�V^�0g,�����ҟ �ɰ�u��'c�2����2ʕ�r��R�iA�B\�a�ʂ����&��PXw��5�p<�t!��x\D�Dݹ7����P�j��k�E� ���#*�>u����>!��F� ��"�v��4o|����P_PuIA��?a��hO�⟼K�N��N�$Q����G���CG"�O��Od��%B,�A�`B�]�� @���צi��JyBj��맾?�RiԒv��ܻ�i݋-�@T����?�����P���?��O�6��K� � t3҄��6Ά�U�,�dCͼ��y@�9�p<@�ݗ�~��X�`�J4�"�X��j��ß$�z1��O͜vwd��ɩ�d���O�ʓLb�ݘ�需E~bza���\�4%�<a	�@[�Y(�GF�m߶@#C��,?�=���?��&�!�h�e&�1�!)�E�w��^�l����M���?	*�(�J&��Ox�P#a�' �ԓ�%��k���-�O��$ì];�X۰C�$d�b1�����'��)C:��i{ e� qj�5!����)��b�dJA"E�	'�e�T�Q-TjQ>ᢤg����qjR-L)Tʼp��'5}��Z�?��i�����Pe�Zf�H�"� ���u��O
��d�d��`c�F$!�re��n�}axg;�S�? �=y �}Np��IJ/C�p#��S}��'x���)/Y ��q�'s"�'�R�w�H�o�;H��$P'`

0R���N�d�t�wO�Of���6�1��'�D��Pk	dΤ�Q������0���/�T0	��O�\��������� ���.W��r��V�	��B�����n3�O�ў,kr��*Pj���CJ$Rj�Y�s�;D�(��! Lh�ir�d0��kר-?I$�i>%�	}y�̖�g-�u�R!_�����m��p�b��V�*�'���'%��ş��I�|Z��ۍI��Rc�;W��q%�I�[�xa�g3�L���#E�|sv���	�R���ZD�ɋ�p,�jЊLY�pR��Ѵs�F$�a���(�F����$O��#�&��N��qQ� )e�.m� N�0i�~��lo�u��v���A�6���Bq��Q"O���b�\���yA��DX��d��L}2[��٣&K�MK���?rT�h���iK ��P�h��?	�� u����?A�O�f( q���-��S*O�qԆ\��RX`�Ǝ|j��:�'ѠcB��(/R8�)O�h�����p�Ŏ������'�R�"�_���Ȩ>)T�U�@( ��D�S�*<�I��<i���?����I�,I4�C6Lտn��L`�,{�!�\ӦEA�JC(F��3G�NbdF8bDs���'˒5؃�uӠ�D�O��'7x\\���:W������_#���Ӭ�<7�������?q�Q����°�c�T>��O4*���ܣv����b�È/�`I��X��`�X���Ɯo&fz��Z�*;��BeG�DKb��|���Z�Z�&5��X=��$�̦i�ڴ�?	�����Y � ��
F�),y}�4�<����<��B,tY �˵��e�Z}+C�T|�\0��2=E�C�+�GM�M��I�.�$oZß`���x9�C%��I��d��ӟ ��������D���x�}��-�+�y�����IڐH�V��M�M�|굇y�l牊:@�)�κ,��"#�kz90����Sa��=3�=!r�4.�v���<Of�8#m��b���[�o�"��T��ɦkڴ�?���۩�?�}�'?�D�6Ky)�E(O�
�5!pIՁ2g��K�Ts��ŗa�p1��,\�	4�HOb|��'�剕V.�Y�"�%8�.����� �p����	Z[�h������	ڟ�Q^w���'����
6j�k1�G-m�]�������%ۥ<�TRB`ןBRb��E����bc qF�y�C��Y��Z��!������s7Ozd�$ b�ce �$,>rlJ��'���2�ST=���� g�r����P/@|�B�3BZ��cd"m���z�	ϘX'"b���O�ʓ4ϬS�ii��'mTl�ahO�|���y� _���s0�'��,}M��Ꟍ�'0�z���t�#��L�'h�T�
I�3!TY�ab�-40T���y�Ш�,�!!�쉆�u�"
KE����=^D�}��ʯ~.����?��,sӬ���O��ˤ�K�]F�}Ȥ��-2j�1� �O��d�O����Oʒ���Ox���gI˖B�24ɢO�qn�"�<X�E�+]� ���B�a��	gy�ή���?/�RpRu��OF���^ �(��L5�-����!�?���:�
L)���
^��\3��ZH*��˧Gp���"̵A��`
:kN��Oʩi�Fd���q.(%����5j�(l�O����3�%
AmI�l��3L��S��O��D%ڧ�?��͹tc�p������=#��ϛ��x��Q-�>�� i
28lf��0<	 �IY<���D�6Kߦ���.�h���Pݴ�?A���?�"dʘX��dS��?��?鱺�5�Ao�і���D�,03raP�	p��[`G9�3�V�?��*��B�WYN��G w>��'����Q_q��'�P����Y.���8�܊1*���eu�T0�'�R�	�S������x`�H��[�Pi��jE�&����tHKh<!U�e.¹��J�pV�IA�S~2�<ғ���<���
o�K�k��Z[��T�oJn��`P��?���?y�n��O8���O�!���$-��Q��M4N���Y���5'����'��XP��/^:�zψ�����䙰w�|�ƅI����ir�B��0<)���?I{6�F'ѭx�؄J��$RT�����t�O<a���?i���*ap�0�NƂ+/֥1TID3ɸ'�ў��5ˑ�V#u���ڀ
<�c0�Ǧ99�4��.3*Zu�'��Ė�~�̼�u��m�r�d$m��'{����'[�0�l  &᜗{���Z�C�c�7��a��5�ꔺo� �C �je�x��5g�bQ���Pyp1,�����T�z�@P�W+|�����
\`J넩7ғO�V���򟬖'�N�I�	��C�j���̸��j�y��'��r��O����@Dсr'\���'�6m�Hd���CB�dc�E��ׅZ�D�<���	[��˟h�O����� �U�ץm�Vl��5+�D�z���O��d���ґ�Y�g�,�x ���ʧ��X%tR�h��ѭdG���d�ӹ|�r�j�R�^�@X���I��H��d�ՌG Uf�c���eQɢ�>�����	l�Om��ӱL���
���(	�ЈiQjׁF���� B����@}�,�!��y�ax"(���+t��/e�*U��ꕄ/���p@�i�"�'�B�Ō(����'���'dB�b�	�N�z�< ��ɞ*
+<1��� [�@��tMK����	9I��|��>G�T�*�ES�l�9(j�Pz��N5p�
���ש'�TI�q�=R�$��}.��I�s,.�u�U�Wc���Q�]@D���W~��;�?�}��ğ����{��8Nҏ:���[�	��BK��7�r���]�X�T!�,��r��'N�#=ͧ�?-O&Yb��>d�[��o��8�@ ���0��OL���O��D�������?y�OC��+U���n����Խ>��X*��߻j�}�#�қ�HmJ���>U�џ�c'�ߪ��03�Ӏ�f��.Ui�rKB*m��Y�꘸���Eb,ȭ{J�вw#<�����)7����W5�f&q�~���<����'��0���M�����؍1U>���'!,LP��:M�ES��=A��y2N�7A��Z������u��'��#%�P��)� ʰI���#=]��'�H�bb�'%�3��уwM���!0���+R8�S�
�2?ݚ��-ҍl�����ʁ��p<��@��{l%����;�v c�ˏ�z��Ń�P eZA*#��
۲<8T�ݠ��Q @`9������7�M����?�Uo֤D���@�-���B�O��?1���?��?�M~
I>� Ð J�HV��,*=�W�R�'�ў�Ӻ�M���K=$A8I�D(_�R�ђ��I�?َy��(��I�,�EAa*٪=���T�E�>B��,>��Ec����a��H� Z�&B�I�5yt�Ad�_!W�n����(!B䉉�(�g�Qq���� c�$U�B�ɨ5�h���#K�Uf�����4(B䉜S�I�&�P�%p�z����C��:4qPzc��9��� p�RC䉻4����̎-Ngp)�T�]�3�B�� c�~�{%тI]X��v��
E�C�	
����@�m��*a' �	�jB�	�y���ؒ#Шv�4��! �,B�	T�H��NC)"s|��`�\�>�DC䉴�e��	��gz4�gM�:�4C�I%ـ,��j]
I��8�gH�K�fC�I#G/&e3sN�v��H�����2�B�I5ЬT�6�ս ��0�1(C�
�B�I�=����1�	�x�ĀcA�Ն*a�B�	�[��Рg-K�?p�`�Lҏ	�^C�I?_�A�QGM!��Pu-��PC�	�`<�Y�k �[eF@Z�l���nC�I���A7@L�]_bth1Iͷ3�ZC�I;���E�7{�:���%0bB䉆8��l[UG'A�0HhÏ�$z4bB�	�0$°��	N,��r0�RfjB�� @��U�՞�L![R�R7FC䉤w�'���T��cD��C�ɢz�&!�*�+�Rm��lӇM��C�	�p��8ӵ��aV آ�K�:(��C��8.Z��J�I�t�4qA� �@U�C�I�#�e��B�05���$/GnC�	�2��t���2[P�������.HC�	$^W���R֦��HPha"O�u2�˶���P #�9�L���"O��@�n�9&���A��&��a�"O�������aqO�����pl=�O��tdM�~["�*-:nD��=K��Rr�.�ڿc��ћ��ܽ#�d�C�M�-A�OFx���,��%�!� sڬ���I���X�c6%!m�B�-V�Ek2�s�8�x��|}��vJ]�
jk�@�.���;3�˽.'Ԅ�ԩ&\O�ճ��6l,L��a�x`p�i�u�ӎ��iv�M;���@�.��c%R7�~�i�q�$�7v�Kǖ)H���a��#X�4i�$"O��I�EG�4T�K�+��ڈ�� [��t�KD]��?�"�%�$���|��MH+1��=� �%i��G8N6Fܓu�.bT9x��'�D�q���d4�$&�2{Xv����Ʒ}��m�vnP�	�/{HL����dԅ���O�{Gn�Z���"dp�r��1ғ}M�`1��Pq3p !r�Z��� �2ۺ�j�A�6��|�$�׮l���ԥˉf�ĸ#��u?������	�.��h�cGV��
�C�
�j�=k��|B��B'+o�vd@13�(0����@*y�`��5�2ь1;V0'��d��j�D #f�"o+���s�˹�^���O�-��?y�����*u�<�G�#E,( ��/��@�eh�:X�T<P�Ȃ2�Zq�p�t�2r~�JK��'�tl�ҡP���BHX�nPT�(rf�4j�
��d#���O:@RS�ѫA8tI��ĵCF~�z���=&d�T���5�z�pa^|{�䆨Cyh�0a½��`\�W�$E�*_�.W ��ʩ�HOδB6"̙/Z��I�O�o�h�	e�D;DcR��GM�.3e�|��;�v�0�ժG��M"W� ��n���^������V�=1;��S�c~����J_� �z�m�0�)q��^1�M���08�:�xjaf��)R�X>� ��˞W�6O|-å�S A�l�S2��e����~b�Ÿ:���ґ'5C��N�� ��<a7�O����a�G%��J��2���8uF0�Tò�V���^`�$��`3�^
c��smZ5���h����5H&���Y.{W�T�#>�n�V!����
y|y�#�	$dy;��-6
:�� �?�{�(�i�'��X��$ߜv-p��Yl�TH֥ޣ\����`�cV�v�8���r�:%�V�AN"3�O�J#HqIf"��8/�T�'!��<鴂�`.qOJtXłZWI��{���I�̑ᯄ��t1�X�A�nh��n��~�7͉ �6$�=	^�l�WɟS���S�)n�Ot���@�82��D" �Q�]:�~���g S���
4d�py�T<�(OJeB,Y�qc�
��QZ��E@�P��i^:W��8��y�'&�d�a�Jd ���8�*(��BW�F�dD���ڇ)Sx��4��0>�t�k��Ć*+��M�°	��}���܈t���3X4��p�݅/B��Y@:�~z�"ܤ�����#�����Ҫa�.�	.�}�TaRP�߯�HO~�Fa� ���**0(���?�ŉ�� P+c�κ����t�hK ĳ6N��KA�Q2�~�KK2@���3VoM(6���r� �PH��Q)�5���'v��s��i��<(�����0���N�2�ԡ:���qO��`Y���G-$xD|ه)�6	��lC5O$�@�OԷ=�L�#� ��	��O"�(H�\���G�F�đ`6*�����ߵ�~��>����D�Ɉ�F�̓{����)�0:�&x�D�K�������-�G`�'�0<��� ,,�q�T�Ʌ0>�0D�?r��1�:����O���ɭ)]�8��?�i>��R�x��ʐ$V-#����1��H���8H�05Δ*|��! %��/��Pc��"cL���0O`����D$���m
#Z��4�'[y<rs�?���A�`��t�ቻs�`��$*D�p\:"���|�|�D^3Ɩ0xe�Xa8���v��O�T2g�'���	*'}�\>c�|Y�X�A����j\�^m�l���#?�5�Ř\=�����ۧo��i1 �ԟ�g}�f�pV���
MhƔh03.�,4��c-�{(�Ň�I�0J�еbZ;��p�["�	�L.�������O�$@tf�1O��'�вScG�0̰Z+��UJhu
�O�ѰW+A��h�צ��%4���A_E��%�6?�
	�UJS���4RǓR�b�F�)9�z�D \>��� �F�$��g��0�����?c������?�0P��+y4 ��df$�3#\)Ðx�E�h�L��QlJk$4L0��Or�;�~�i�9'�*C��?)2-��~��t�͘��â�q
��j����1�O8-�Q�݇GfM��)P/Y�����6A�X�2�2*���	o`Lb�O�扌Lp�4Kݦ��禅���ǖ}2n�W���yznIx7i8�Io&	U	ïm{d��5����9O����ʆ=�0�sFg�'R�:�����?�w'�\�t*����3�{��� �
�B ��")A������J"�Q)P	��a�2����ԟ�'t�d!�Jmu�ӥaF�T)H���+�fو�PG�'�Z�	�d˚HBH��f�.��9�ƥջ�y� �Ld&��4#)�i��đּS&SOp��x	8y�d�*�V��I"Dc,�	�!�9.f�GT�rI�l"gθ?7������O�1�ua��ve�-�2L޼��ܴ<�M3�� :PJ&��uTHEx���!i�'MA�wH�$�p͓|��L1�Hߐ,�٩%	A�Peȅ��-C������'@h�g�'7��#�?_�b]�	����!��3b|�% ;MP���'�n��ӟ�I ���<��c�.�Ļ3�����Lt�׭�w��u��$�ot�����b���#?a�����?O:QiƉ: �Q�)
�/����Op����ygnC1&�a��^-2�"|y��ۅ�M+���p<	��#V\.2��X�����<_�|��sć�(��Aș�]������M#U�\���1��i>7-P<�|��ϝo�ଃ�/\�l��i��]�L�x���a �W���)�����NKỶz�APIԓ<�0Ik��ҍSDR��"��?D��?��'"��ӂAj�}Pv(��C�xl����=,Nda���'%�8`��-w
��fL���)��L���	/u0Zu�1��1	�0���$S6�l�fG$��'�l��V�n��<AƆ�9]s20Q t��3���% �h���0��s �)v>!a��,��8w��|�;@m�8Q`��_h��c�BP��&��Θ3Ev1���:�V���b�sb� 9��AH�p�&�{9�1�����}&(�Q�O���U�хt���1E�����|2E�B"I3NLQ��a�|)��F^�O���G��f��&d�?}J����O��*W�Q8��b��&bĘ�O
\,r�!��</ֺh`L>��<7(֌?�P��;Z&��*Ҏ*6<��EM}G͠�i�90."�f˃�T���s,�l?%?�O-X�ʓ'ܹ.#�����ɐ@�z��'g����'��"����Ey��IJ��c���N����͔N��ţ�'ed	rf�_��u�O�O���,ub�2��Ϙdg��B���TN�Pc)����K����i�ʘJ�8�(|CfO�Z2�$Hb-�Gl����$v��~���`�p�����S2�G�n����K)+��%SC
c�'*b8f �*�%���bh#a��~�'O)�5)U  ؠ8z�G��X!2�쁢��'\X �)��0(���w>��#!@ǜ[�A�)�������R�tͻq� �1b89uh�-�~����'�h�+@(p0P�Ȓ�
��0
у�<[�$�� ��
 �� pӘ�!�Н#%D�9�O�|qb 3���+%�ݩ`�"�4�ɒC��q�s��g�!5�v����R��0f�a�VP�fW:~Q��)�i�-#6.�t�ֹ��&V�]�B�!4f�	x�$�ϓ
�b$�q d��-2g�4h�q-���S�F�H5��=�%#�
^�h����K�'_su���`ꄤy��	�"�f#! Z&�b4z������@H	�ɓ���D?�J2�����̏)"���fLi�Qa�:=Q���V)B9�H�S��yB㕓㞔x� 4 �!Y�.���^�Ƀv� �e�5�|��;g��<+����51�1: 'Z2V�,R�ă*��$
�C�$�e�ٲa�L�ʧG�@���+�s��IyU钊.���	�� 4�Q9G��.��V�I0@��D+nޥc0�	i�jA�q��*����@"HZ���t",�q�LI�S�7�T�S���(\��|B)E3S4�;KP��O`�V��8����("�S�%j��܆&�X02ƤO<V��X�����lj�#���aA�)�'�~A7u����u'M�_7@��é�M�uQ�I	��%�q[�"~�*z<c�gY9�Ezv�:1�@٠�����ē�K�'g�����?�>�.ŋ��@V��#LEKV���<�4�� �=��lA���Ox�I�JX�IEZ�o��YY�ҔC�0x�TY�,A��p<��BC.Y���ϻI� �U��	Q5"�����O �jT8T�X2��4D>�ڤ�'*�N?1���Hcof	Ò�B�䴂AH8�a��۱`F�����Z7#�JLS��]`w��� P�t1� �d@44b,O�c>��r��	C��d1���<x��I����Q��@�c	�,��cF�<E�3�n\Q�G�+��R�B�6�R$���'�T�04 �
E�,uk�$U"\�n]S���ΪO|���De��.E^�Q�͚���M�Ԧ)�V�=^�����O�`����i�R1��:�XpՁ�;&;6�T 1����I'Vn���4C`�}��V�\��i��n8����W?9��?�rˀ�h֮� �I~J|Rq�� T���͉3~n��6k�Q�'^f�;���D��
r��V.}���b�P�Ј�di��~Đӣ�d����ZI|�����5��	�WJV<m�
Dˇ.�,BDx[�C��<%d���PTy*��I4�d$:�Bش�N�F](�i�I�h��'Ԡ���(P�S�b� %����p<�F�99<���  H���Ǚ�<���Гon�I>'���C�?aR��xF<a��4o��84�R�O<ܓw)׽w�&���h:\O�\�q�͐I�WJ��Lp�t��Q��İ���'k��� o[ Xd(dfQ��rd�y�M������g�����s����D�j�f����a��q'䅏sf$��׏�p�禵��$�+*�l*�.ɗOR��z�C	F��r����~r�Ǜ �ZYr����6a�����	"om��s'�xoz}b#�ݥ<� !�Ү�|�bh��'}����;n.�#����֏Ԕ�ހu���`T&M3��O*)}Xl�U�
��yBm��p<��O�-�x<�sI�U82u�3g�l≖u*pe�o޴V��Y�m�'�.6M����۶Ë�p@rƭ�Dc��S�EN�z�L���Px���4'H4�(@�ŏu��03O�ZxHq�LӭB�X�Zӈ;��?�27G��y�c�/X&xu���h�"9��͑��x���;���U�-�$��T�G�P������=n�v�с��1p�H š$}�N�kr���fW���RF.����<��nG�E���PB&��=l$x���˅�=�FL'�a:e�ζsj�]Zԇ�)D$1rF����m��I&3O`A�v!�ESo ;O���PM"�����g2�{�� F<���5i�Ţg��&� �B�'�hL)F��S>����L� C��{"o�8_��!AkZzt �����AQ��a��[Xj�f(E�\�!�d�p�I�EDN�xbB�j�ދ3�!��H�u����6J�mF^ "D�F�<�!��sˮ3��� 9`ٳ.��)�!����ʕ!%�܌f� ���^�6s!��4߾��f r�j�(ej�$Jq!�DƴLT `t�܏dҠ�j��ȋ4_!�� \�@��Tb�(@���)�v�X1"O&���%�H�4 �"��`o��Ip"Of)x�-³��%[b��e���8b"O�|A�h
24��`Ӵ3���:A"O\V���s�
1���Q�A��)�"O@Y �����ș�iH�y;�P�t"O�)�ub�>iش���!D�f��c"O �գ����!C��]����"O$��C�Վ(Q�M
B�zy�A�S"O�Yx����^��I�1�F� ^�8��"O<�RJ��ep�G��kR���"Ol%Q6Q��b}��BU)?�p��v"O��	$ϔ=ʆ�2a�'}�X	CW"O^��q��)DS��(#��-i��d	$"O�PK�lQ�c�c�$'i�dy�"O��cn��
eK�cZ�~�0�[�"OJ�r��;|nl�f	&A1�1*�"O�2׋ٹm��{7b��E��"O�ؔ�T;r�*� ��"�zY�T"O������V؁��L(�\3"O<i�V����	�B�ɉ-�=1�"O^Ue.N*&Q=���K(	r([�"Oh�4m� 5J�M���W<�����"O���2(�n�p��ή�% "O���%�#��P!pB@��R	KF"O|�cA��0A�h��*z�!��"OP�AP �.N,3��|�v�9�"O�QBe̪qie��, �`xJ�"O���"�7TM �C�@$	����"O�*�b=;�0�+g��G��`"O�`���Y?/��k��u2j��"Oh)�%��,�
	Xw$ʆ#��w"O&y��`+a��ӢT�/��t"OµR��'G��Y@�H�v�� !"O\�c�0r�1�/�&Qı��"O�R��#|9L�ȇ�
:�ic"O����*ٚ��ރA�.��"O<�@U�U�@[�X�ǌ:R�D�
g"OxMb�%!V��^?��\�C"O��x�dBfŐ�O��K�x���"O��	܍K��e:�� �q�"O�9P�'��9M#vNכJѴ��"ON4h��%D�p� ��ͤKʎx��"Ozl���U;ԑp�A�6H"\��"O u�elíj��|R�"8RxF8��"O��I��L�S<
l0� ^(I�q�"O��ӥ�+��P���8DѴ�	�"O2U��GP1Rb:M;$/�?%\^e�"O�A!��H�d�;�
{����"Oz5!W��>r�I� ٔj��I��"O^}��J:ak[���5V��z�"O�!��I	�Щ�lН�~��"O�;$�ܛ 9�)j3+�)^����"O����P-��d��*H�*c��"�"OJ�9�Ä�Lj P�a�l�V�[&"Oڸ(w��?΄u
�#W5WG��y"Oh�"A'�G.F��"ٹ0ƴ�"O
���e�1TM� �X#��`�"O"<H6$�7O��1���ڜHv�`�"O09�m՘:GpĢրό`Uh=��"OzHqCAҠ߂d�Į[:S���"O@,�����
�@�5��:&"O��h�&P�E�dq�kήx6ȓ�"Oޑ2Lͫ(1�|��F a!�K�"O� *0:Ti��0�Ʊؖ��$`�� �2"O��9b�&̆��F'��;�I���$$�S�S
�N1j!a� 4 ` s��X�rB䉆��pѐ��'6[�Ђ����B�Ic�j�p�oQ6C����HI�C�I9��)�X)7��eAu��gC�C�I5W�����BT�mr��,DglC�	5Ig��a��P�qQO�`�dC�	�_�	�Bcِ88���1΀�HT~C�ɕ��u����"��c+��cVC��1/.,q�B�;HT�c"�B�I�&,� ��&-
h����6��C�3+0�rSl>�����T���C�I�==���gLذ�`5,�=7��C�	< YȔ���N�l!e�2	}�C䉻! |T⠠K��pL�bJ-���D{J~����20贐��v`B���f�<	ě!xn��WmU�S�q	�'�W�<�%��U��D�`�Cy�&�����T�<	'��$8Jq�[�)������ �<�S��E�g�	A�X��#�/(^�M��)�t%�'�}�t+Я�7"��Tn�s~�)��8׀�"քI��h� CK�*C�&#>����մU�A�S���S��yH��O�k~!�d��U�ȸE/��o���B�hZ�}G!�Ԏ3��{D��*{$�Rt��8A!�D)-2���pO^&-J��)G
f�!�$�ź� �-�kC�yz��ڞoz!�$��L�X5
E�wFd�A� ��U\!�߮sHԢ�)��hE���5�]'h�O&�=���d3�Ē�0�65jS�ޘ���j!"O���3�>@$�G��v��� �"OB�)E�� oV�� �c.h%����D����v�T��"F�#ܝ�1*���F{��9Ot��Dl�5�L����'k��`"O�}��!�8� �M��(�C"O���&��.Cn �n�#<�P�9�"Od��jλ��y�$LקG{��:O�=E�$NU,SA~Lk�í]�F����yr%ׄ8�8I!J��?�����O��yb�RU304 c4������H�y���_��iɧi 4j���SdZ��yB
�F�D���1:"~L�#���y��+�ʴ󅨞E�n�fR��y�i�(B�^�P��.���c��y�#�5���pC*A�[[�=��MX�y"G�j���/E�DxFc���y�i�%/�x����<X6ؠD&��y�ǜ�E��-Ǎ.DL��A"�y2��&_���k�"���c/�)�yBAɘC�6q�c�Q�F�.%p��
�y�MT�Q9"[`�L2�����y��[Y�@�QA�T>(�(˵l�y���)��`"G�)&��ѣ�?�y�O��F��w���)"d���y�"�o�<� ` ��y��Jb�ց�ybgLZ�h���u�XA�Ӂ�y�O=z�|����E�,�Af�ƿݨO"
�eA�%X�@���
hhr�r�H�g�<��dԥ��A�iz�\��Pd�'�?�@��۸9��Y��a_&U'��9�g-D�tIG�0;#�(��h�G�� CL?D��ش	�4'6x�SD��^4���2�=D�hkF��-:��:v���c�*���;D�� �ya�Qr}�I��	5:�|�U"OHa+T�E�InL��/s����e"O
�Yt��#*�e[��H�85�Ųb"O��g&�2:T�Q7�W80'�� �"O����Ӡkܸbw��1p�⥈�"O@���j�o��X�&�۝(4���"O,��%ꉳ	���A�:�f�$�	Z�O3��HĊ�x�C3/�BD䈺�'6:8���H�P��E�R(<���'����>B� y��О=�I
�'h��'�[�TDÔ���h�x
�'��U���g� ��ccT-~XX�I�ą���K6ru+�R�?9��b A^��B�I�{��c�� r��P�1 �+��B�I�P�պ��N���G�,VC䉻J]���eU�n���s�:�<C�I.n��[�d4�vx�&���RB䉧���#�AåR�p�*�@׺0F$B䉢Te�����E�uj��U��a��C�	  <���@T�Y��L@Gg QU�C�	�i�^d(vKެ�t�fGֺ��C�I5EŔ��F�H�#����v�@�~C�	�p���f��r�%^nLFC�	,V��L#�� � �,E9'J݌]�|C��3!CP*�U�q� =��HΣ�^C���(Y�e��$�<x����x����6|O�b�$W�Q10�t�ϑr�\��H4D�b����X5Y��W�}�`}*u�1D�@R�ӂwP>�BV�W�m[(mYd+/D�p �)��A;�Y�V�)���f�+D� �₞�Vf�	CSL�%&+� ʅa+D��M�6w��ڢ�ӄ,�� �DL$D�(�u��6 ��R	�/?��dr� "D�x2���|�>�)��
�1N��P�>D����̪{������!R� b��<D����.��W�.�+C�ǳ)v��Yeo>D����X�μ����$"j8S`o!�	̦��˓!-`M���4Py�d���ՆtB�`�Ɠ7��Y@V��]�$�hԂ���2�'���/Ԥ �\i��E!y2\�
�'_sr�J�L��i��s?���	�'EZ��v�yX�=)�"@ k���{�'��ph�(�?0�Bd
V��s1����'��|!`���9���u�N*fq"��'�^%{�"��oI�q:�뚍\�����'�0L����,%5����қDp�|R�'�>ij��Xh���\>9ȕ�'��� �A/���a�;b�B�'�j�1N�8ᐹ1���4D��a�'���㏃� %� hR		4an��'G���JGx�ݘ��å!(�	i�'���r�,R}L�����&�x��'�-��ɍy��]��gX�~���q�'��a�D�T�s�[#sR����'�c���6$yt�]	|�x���'Ѽ�qC��+����"�8E�na��'u���f�."�b�q��@�v����taA��2��UĕY�Ʉ�O�J�S��0�Љ˕�@l4��5�|���˽��Ts��|�8�ȓ5��<*��xlb;ҫ�)���ȓ<*N���$R <�Jv&Q$>uJ�ȓ�)��ıf���B1��!y`�y��]oX��mM� Tޥ��)�3!����S�? ��[������7"�o���e"O�X��(L�Mc��<��Q�"OE�Uԫ!2��	�+˵6�-�5"O>���JɼJǹ jH,-F �"O��B4�ļ1��}*r�T�N��"O��@­ߝ5�u���Q~��80"O��@ǌ-z�=��Nby*h@1"O��6IY#=p����b]|�a"O��8gB��5�`�i���B$p���"O�����
/kr1 ��#z4��0"O��w\�s⊠��X�r��{"O�y�bƟ0���2��I�^�ʕ"O�����R�Bȭj�*Uv8��"O�P�p�@�<��sU�^�lXa"O ��Q(].M[ah�2��0�"O�;��&;� ���G+"V��YD"O&���Нf�
e��&M/��@��"O��÷���_���)F��G���"O6(H.Ȏw�l �$ٵ/ε* "O�[�^�X����=�,�1�"OBup������Z�a i�č�P"O�D���d?�) ��;�Z�$"O���^�p��0�GHV�B���X�"OVT���+/*��	㇃�Q�����"O��3ԨӨ���5��K����"O9�w�P�8ƸE��EʎT���P""O��K���Ig��S�U�P=��"O�PT��=ٶeK��UnO����"O�	�U�}�(�sᜏvF�5�G"O Tc�/n����ox�����U!�$N�^��!U�/R�k44%!�$ɱ0Xna;�eAL�ၵ��>�!��M�T�`��wcթ,�sDѲ �!��^W]������sqC�k�!���p�� ���Ĵ=���2<�!�D�+1�n�%�ԕK�	`b��,(z!��-M�n|�E�"G�h�T�~^!�$���`��L�������޽z5!�$�|*�e�cS:;~�٢�-ظ<#!�S�8��F�Rp0�ZO����ȓ`����������/�n�����``�MR�G��S?Va� ZM(�Ԇ�:�]����7 �R�vĖNIxB�ɯ=�$1��ѓ9uڜ��bT:ykC�I�iD2!��!�a����g��B�I�~�52#'�X��M4�O(��B�I5|x�e0�$��{�L�b�<3(�C��	PrX��J.y�D  &R�C�-O�6HQàB?T�P!c�C�I/#�i[p��8u������be���D�M/��Ig��g��ؐp���U!��! ��� ���.1���N�A	!��Âՠ�W~�X�
 	e�!�Đ�rT�*7.[g"9і���!�$у#�zw�	`O�`Va�x�!�d��#��Cd8��`Qd!;k�!�V �4d�@�&-w�CGF2e	!�Ĉ��(z Ė	�"x��O��1�!�
O�>�XWJ1�R�RDβ_�!��u�l��3�.e��̓P��?�!���n���K�S~��b���)�!�I�S0~�	�!_-+R���#L�*�!�ĉRf���
[T�QK5`ݙ:!�9%��p��oώY@d�BeI!�� ʍz�	бL����b�P����"O<�*şj(F`���ӎ�Āx�"O��聀�9j8lhKb�I�^*pi#"O`��)��a�����1ғ"O<]#�G�8�>���Bm�Jԓf"OL�bU-ɏ%>���C��%2��I�"O���6���aY���b���l��A"O��A$LX6a��񏜻O�
��"OB]I��B� C"���9F����D"O�y�%,	�e�R���)��`^\ۧ"O"`��/�`t(B��9hD&�!�"Or�Y�A��v!�|�e�?O5���"O��0�̎P����%�]<n+�"O�8q���=2`Q�R�'ʝ�$"O^-� ��`�xb��^rq��"O��[��I7Q�����f[�] �k�"O�Ca�
I6����oޑ'���0�"Oޠ(AL�'�Y+B�]���r"Of��'����R��O� ���q"O:��bdF�/���P�Êt��y �"O��;ԁ�%M������86�8Qڡ"O-�IY
H~�ن��$.�zH��"O�D�9i,�i$g��By��
&"OD��ǂ� MԱ9�+F�Z��y�"O�DK��&�P�y�
�KX��r"O��1��#B�I3�ٛpN��R�"OX,[�n�1 �R�ר&]�Ѣ�"O6(�Ǟ�Hz�%�dM��u"O.����N�F�#Ρo�"q�"O�����F�\��+D���0��`yf"O0ъrT�\��ɉ�-��LR'"O�9�I�<	v���IH>	#�=
a"O�I�%�
�t+(Yf��B�L���"OF�1��ˣjFM���g�b�"O��[C��<1�0d�3�/���* "OR�pՉ�N�{B�S�v2���"O�ա�������w���,v�E+�"O�����Q2M���b��_=�mٓ"O���(_>J��E/F)h�xc�"O<���Ɨ�8�jĐS�M$|��U"O��'A	c�iTIP�45�"OX�a�������!1�ڴ��c�<A'�8U��8p��.P����Oa�<�6nF�|�Ɲ��b�'U$�m�V��D�<9�i�+�($kG���+�����-u�<�����vБh�D_! �4�y#eNu�<�f��~A��Y�Q)aIے�u�<Q0KP��x�y��V��Yɢo�<�`o)w�I2��`hA�K�g�<�&)T�kB ���E]�{�n-y�Lk�<1g�͔O��kqD�_S��0JOf�<��@զ��z�銤S��i���H�<)��/L�4K�O�	���C`E�<�n3rm��zd��[��3w�:D�x�DF��
��I���@�bI<]8P�:D��x�U�|����@J'^��}��4D�8��۽d �ib�*9��A8��3D�������Co�ݓ4��m���Bc�,D�x��̆(dlR���T���F/D�hI7�6<41%�[[wR)Cѯ,D�ܱ �՛Uzu2'aZ?y�<I�Ҡ+D��#��50�P��Xr��XQ�c+D�HjAO���鋗� �0��*O��2+ӻ'{����{{(�s�,,D�� T����A"k� ����=c�m��"O���o�n�>�;ǩS&r��
"OlT{�D�)'& ���R�Xd��S"O�tA�+����42R���4IҸBa"O�<�Y�<ub���(ń<:<=y�"Ofq8e牋zO�⡥��-!x�6"O�1�4��-.@dd�*�ܝ�w"OlY��L�'�|�tMFC谡r"O���A�-WK���q#ęP� XE"O�Y���<m���C4��,LѴ�+4"O���p눙j�ߥ%���J�"O�0����a.XE�Cϕ�5�>�1"O�����D;l.�p��Ĝ/F��"O�08@e�+sڦ� nX�JAhU�ȓ4GTu�<�lu;�	]t�<=�ȓR^�cCǴ	;���E�&�n�� �p��C`ɮ$�p�߇X��̆ȓAd��6�ʦjQ�a����yrh!�ȓ^=�Ң?"ک�Ꮌ$�0�ȓV���ysā�G�0]Ѳ׏�"1�ȓ\����B�>�y� /�	Qc�}�ȓu?��p� �~Pj���B�i=��ȓ0���A�$.Q13kߋY^hq��%�=b�cW�!N�\r@O
@�&����D���	���(5�v�X�ȓnl���J_�{�d5p拚���ȓO��p#$���5yʉ{�	�	s��\��s�(VB*�谙���Vd̈́ȓ|-�"3�
�D�/�#� %D�8{$�S�7T:����Ġ`G(-D��JfL�hR�����ep�{2�/D�4x`O�l� 1�����r����FN)D���D@ ��@$|g ��+D�dÇ��XA�8&fL����3D���iЂ\]
�Ye��,�Y0?D�hyr'�/�<�q��*Dbj�p�L;D� a��C��J^�p&NȉsH:D��y@ʫ3�pR��1�.D{�+D�� �&�h:^ +���/G���%�<D����P�it�]���:{R�]O>D��J��̆	"\HK��9J��CV�=D�$xG3s&��c�KA?O�I�v`0D�4��;FJD���� *{RQ:�$$D��a�ͽx?�DІ_ 3��c� D��ʅ!ݭ�P�Kq�[�kԼ��;D�\�F�(Y��ġ�o�� �fE²�.D�P�#k�@��`�)�RL(��.D����y��;���#�ڬ"��*D���C)~�Le�!_��[*O�A�')d؈��I�n2:ə�"O"њ'�A�P���Q��X��Z���"O�$z��Z+�̍ѣ�Q����`�"O���.�-��Q��#�3a���7"O�����637c���"�"O�8�	Jr�L(�򢂌4�l��"Of$�� Ĝ����]�$���f"O�u�T��hޜh���Wh�`�g"O~�ҥ�Q(n�J4��/3�T��V"O<����Q�,���ˉ#���"O���El�+����U�(��	�"Oh��ѬE�s�>�Ң%Fiof��"O"�!�Ҍv�D�G+z�]�u"O�IY0��2%0�m!Q*B0l�V��"Ol�a�Fb�4�E���J���"$"O� \ɰO�,Uq؍"`��)#�l8T"Oj�x�n�Rx�qq���2"O(����8&r�Q������x�#"O04a�C��zzx�ec�����`�"O��i��g8��"F-dl�j!"O&E#HJ	�~�!4'��U�"OJ�zC�H^L�����>W�l)2"O|t����lNA���Zf�y˂"O�hڃ�ܡg�1O���I�5"Od��'\*G�Y1-
f�
�3"O���$�P�nX����>����%"O�y���5jt��T�-�}c�"O��ɳ�N%zöřa�nLd�"O�D��	Q�u5p� ��"OP�h2"O@�0b���qnb9)���2d�B�"O��A�7Jp�� �J�V���"O��U�Bt��@i��R&o���"O$,Y�Ǔ� Itpa�ʹ6��"O����@�!�JU��-E�'H���"ONQ '&!稭 FF��!?8Q!�"O2�k'�X	ao  �Qz�"O,p���L�:� !���F�U��"�"O"]�MR¸m��+M�&U�M@�"O��u��4Qo�YIT�%=�P��"O
ɱ����J��J�.ӟ�6 D"O��Z�dǮ��!Z���3Sψl#�"O.�(6*�.k˘�� k�
R��q��"Ot�3ri��T�T��?��ܚD"O�!Ȱ,�%i�9�tC
�iF��"O��x�Ζ�,X�Pu`��a9�H��"O�]�¯�@�P4 	��SD"O�E� ��E��0�VHW��8R�"O�������C��}���{>4 &"O2XzSOxm�`ZQa��Kn��"O��)e�ϲL3g\�C"O0]����.��|vL��BV �2�"O:���P�� h�@�|>^MJ�"O�����n*���a���
���"O~-K��{�z����l��\��"O1d*c;(�9�.�!*��x�"OF9a�3Ȭ��� !4���"O1q�K[� t���\�֩+�"O�@�[�;Ĭ�!�퀄3�L���"O���C��h���a��@���"O��RlJ7�yPCOS �z�6"O�EqqD.&&�q��\��s�"O �ӃIʂ;��,R#�Mm���Q"O���b�5-�Y�OÐ*���""O��atO�N�MA��O�`l��Bd"OP}�F�?tM�/âCر:�"O�!pA:_�&x��M]2.,<U�"O�	�j�]X.�A�ƏZ�l� �"O�Q��*��s&��x���"O���A��4k����#A�	�s"O��ASB�b�L�v)�s�"Oja!�A@�HP��2/b	c"OjQb��QS���1D+�ݓ�"O�hA��&R��('�W�"�3"Oؔ r��-P�l2a��(�9"O
��wO�3#b�"��|�@�!a"O���e�G�����A�~;r��"O�z���N\�X2M��yi�"Oµ�AYz��z��	^���"O��K�^��0����%,���f"O� ı����4\��!�ޔq+\l�$"O
�����V��qQg
%+~�B�"ODA����-h0ꐪ A҆D���2"Oȗ��[;~(u�ɗ(���"O>��3O渹A��g�2�'"O���腿	6q���ȤF�ЅA "On���a�5�����£	��0�"OL٪V,Q�q�-��? �d��"Ob�b��nS4��ɢYN �"OX�t�Ŕ
���2N[�-B�H��"O
	��C~�E��N�n.hz"O@	b3�^<����8���*O>��A�Q+J���V(N3h��$�
�'M��⤊E�$� ��b��[,�x�'�
TA$��;;� �(�đ�@�H�'�
ٻIȜ.8n�@���Q�'E�аC�_?G���oR�_]IKT"OƬKBd�!yîy��&�a=��` "O�Q���F�W��(�eh�= ��"O����]; ����u䙷o/�t;&"O"�f�\|�� �W�w�j���"O(�:��ߋ{X\L�P�ţd<�a"O��R�S ��V���r|F�bq"O�}�p�߁3�I����.yPu[�"O�=*A�ͮ�Iz�F�tj��Q"Ob=Ҷ�$���EO�q���ٺ�y��J
�ʤ8�a���P�R��D$�y�+ޏ-d,i�Ԉ
�Bx�w�7�y���8d�2�,>Ni)p���y"�ٻ�|�G���z��o���yR�9*j��y2Gϛ{Ά=XG�I�y�b7�����*"r�w���y2�I�Fc$�*�N�"~�`{&oG9�y�hL�|�.u���{(�@v(H��y��^�!	Е��J�	S��6���yr�ָ7�0j��ɦ M�9	&a��ybdE�O��I��
ݣw�rp��J�5�yB�¸/���["'Η�B%��J.�y̅
F���Dn�;x�6y���H�yB�Q3g��B6LH%w�|���i��yҢ_�J𸌘C�'v=hػ�e�yB+�$#�K�<`\�:� �yr�
t�i	D���h�L3�V��y�
%	~Q��b�OL@	��+M��y2J�(*�d c�ѬK߮}��%���yrƀuh���hwb%Y�̜��y�/M6((�p�!�m�6=��[�yr��!'�z�s���i\R�"(�'�y���x�h�RFf(Z��E!2�_��y�Wx��$.��#}�0R�>�y�Z�" tA`mEuNt�pǟ>�y�,�@�s!(�*.~^��QK���y�d��_@ٛ�͛�n���1� I�y	�6�x](5�L�a<B`g��y�cV�+{F�S��4qV�]x�	�yR�^.'t�в�nD@FP��g�=�y��R�y���S&ܵ:�� �ٙ�y�DC.)-n�S�*�;6����5R�yB��']@�@GT�5��Qkd�T:�y�nX��2��T˰*"�e�ph�yr�E�j�2��'�4�[5�\?�ybl���0V	�+4d�Y�K��y��Oۆو� "�}��æ�y��
('c���kҬ��& �y
� ���ӊ#��u���ùX\��@V"O`	8a�=�QW���ZS<��V"O�eiv%��G�Nr	�?HW�P�"O��*�m�zu��G�lM�1K�"O�x �
LjŰW�P;+I
=�"OH-P�T�s�0��5��?5���W"O~�s�A�1k�TtC��տG m��"O腉gHՊw�����;)	��#"O���QH1z�#��m�f��"OV����цfKXQ ��A�RDq�"O̜�Ч�<G�B�����;���""O�(�dͺSҖ�t�C ��ˤ"O���#J�C	B�0aX-_y��""O~�ˑdV�^��ir`�8�l�s"O�%��c)'늽ʲ.�>Բ0��"O$�j�ڃFޞь���P��"O��B�'�W�=񃌟�OF���"O��j��	��-u��s2�5{�"O�S�?]�����+��*���&"O��BҮn䴜S��ǽ'u��7"Ot��%�#S|tp��)�_�V`�$"O~�{Q&W�4x�I"� 2s��Z�"OH����N$���ц�?iZL"OV��姘�My<�9Pe� B��w"OȌ�%���Vf�0� �G�N��t��"O��;Uf3<sbq��CX.����B"O���FX�7���mF5|�8�"Of){e.M4J�B�AŬ^�;\z�w"O�H�NM�H����li�"�7"Oֈ)�F�p���Ð���^y|<T"OR��#��c=R`C���Tf��a6"Of���nJ���[�C	���p�B"OJ�P�H4X`����cɽ{��dc"O� 0A-f���
R�E�.�DtZ�"O~l�w&4mԄ��B�D%�X5�"O<H$�Ѓ���쌓��}1�"O �!R~@yqK>[�N�%"O(py#aɞ0M^ �p�9sZ@1�"O�)P�@3I�P�5�B�O����"O�t�Ca��J�J Y��K�,�xe"O�\�Љ�W _�[�&
'Ů�yb� �[�R\�k�!P#@a���7�y���oL��Htǝ }�R��r̋�y��286�z�-�̽�r�ފ�y+�^���dg�%qi��1��M	�y�`�,y��0�̂c�������y��ͅP-��P�+^�UEDa�TNY��yR�@,�*�)WH3�f,4����y���4�hRR��:�(Y��N�+�y�J��* �BGj��aX8�H�'I0�y���t�(j�(U�K��	3���y2��$�ٺ0��sG����R��y��Б:�B�O��j�!�gk˽�y�K�W`8y����- <릭��yRj��kp̄�c�^�*�(� �ý�y��F�Q���Ps.�$��"
�)�yRLF�HunDA&ǔ�S�1�&-�9�y��F J
J��E<%;,m�6gO��y��L�Z�)Wf՝:$U�%�<�y�nJ��a&�[�\ٛ����y��\�ln`8�K�,��3/��yrE�/WԐ�B���T(rSK���y�̰:��3D_�h�5,���yB�[�p��P2"��\�fqJ��"�y
� �Y+�D��@�~�a�E�^���"O ��G'^f�qX�(F56�4*"O�ya'��B<�3q"´b��z�"OhҢǾ1�$� �&"l�1��"O�9	pkҩr�����,�bik�"OJHUC�FB)���m]8Ś�"O|(���[�:��XSdy��"O��Ђ�%(9����q<Ly�$"O 1��)B M�7@��U'���"Ol�:`H�l�8h�aW�P"O"e�
�9���pǍ�x̭a�"O~����@2W:"��@!A���b�"O������#vXh�s?��"O �cC)ӆK�fI1���?%.��u"O�(!���#'�0�%�w:�ht"OP�Cc�?#�lkqC��S[v�ۓ"O�}���U;j���@Hz-��"Ov%�s�����g �lD����"OF1�� ΈI}��E��.B�$��"O. a��T҆� ���S��1(g"O̥���
�z�*#��h�a��"O\�sT$�?r|����Ȕ�@f(!�"O$ c��8 �&͚����	;��y�"O͂�k�7��Px���U�҉��"O�t��\�U2(�p���9@�!��&.�f��@���t��9"&V��!�d�{�2T@�A	Em� S�fw!�O��v�hu&¢�\�s�"� �!�C�o�@����)I� �qQ �`!�$<L�4�+�i/���s���#!�D�.{1�蓔KW�H�b n�}x!���%�̊��Ŗi*x�cW̝�0q!�$�Sr�0��]�vzDa�
�+uR!�d�@>���.�Hƚ��HFi*!��%����-�@��GL D!�$���"T��3 �=!T&�!�dJl�
����H��� x�E\�D�!������ၣu̠q�����!�$�D��uBqMMUz��䣖�VQ!�D0�Q�Q�He�ؑ��4jH!�ĉ�B0^���ED��P �\%l<!�$\$~j�q�T'1I'��H�"��4!�	$r���I
�o#���U!�5B!��U5�R�!c�J#�	@O�D�!�9L}��-�r$pD5�!�
U�iq@k�+M�l�b$Ȟ{�!�]�fhq0� ^��q�S��!�K� x�i�k�4�p���9[!�$�;���'j�+��t�Xr�!�dԅ Z �g�J�ZǈQ�E�ÑgB!��$u����+�<y#X���g*!�׊�^�¢��5>d���ޤ<!�d�z���A�t��33$I�U�!�d

`rt`��J	:��w��?�!�DҗP0�Q���q�y�7��)7�!��J�;ꊔ��!p����i�!�D�0)F�	���.M���/ܥ{}!��H($�~|j��oy���QEP:�!�U6SO��� �!o�1��D�:W!�D�:g�DP��\z͈��Gc ]A!��C�TU6��qg܈9���q�9r;!�$��1��M�&� w���.�=0!���f�
H
���q��[�&H�%�!�$��%ت�C����n��fIR�!�� T��V�)�d�vʎ5A���"O x���T�l�����N"8&�ŀ�"O��C�">Nq(�a�	��6"OFA�����a;r�C�S��'"O����ʥuvv9��K{�:��P"O2؉CK����*R�U"9��v"O� XvNճ2�^�ka�9H�X�P"O�"2�΢^Ҽqt$�g�<T��"O��g�(Z5tq�ቁ�s�����"OX-�tj��Ǻ�']��z���"O�0x��S�`J�XS柏.����6"Ox��d��N#�n��+4Dĺ�"O���,�&'��ڤm�}1�9�"O2pk�퐭Ww���j�8��J"OzT���W�U����@	��).J䪥"O�� �̊1V�Гh!. 3"O��!W�N�?�
�9��I�F8l;�"O^��&�v!JA����i7�C"O�M)��Uli�|���'�]��"O,����r#�3�ȏ?mX�KD"O��85ٝ�"$��
��{����"OXJ3�M�.���x��.z�L��R"O6�"1&�Q��(��+��#"O���J�Eb���X�Z�B�[�"O��7i��V�`'nCؔy�"OP�2��O�Ȝ�6��s���bd"O�L���VC���#�*#��1g"O�jSKƖ@�Ny�2D�`6��Z""O�C�i� ���S�ҷF��\�"OܠcC�>���$A�;uT �� "Oޑ��I�V4^8�� "X",J�"O�MB�
[�~�zc@،xLҼ`�"OPm�0�Ȅ,@�"�	�KH.��"OP���L� |�ax���0C�P��"O~�i)��T(�@!H�H?�,Ҷ"OX�"��˖K�� �)��H'HВ�"O�8x�!��L�[���f�! "O����kH�3��1�@]� �"Oڈ��K�Uc���G�R�ea�}��"O�4p���%�Aa@�}A��C "O���o�G3�!f�ݥ</�r�"O�L��d����tm��T,p��"O��yGhR-`��L 0tQ"O\��ɀS%.�H��߫#sDtH�"O���fcS]�d�r._"�4p� "O�WOR7�h�o�'�p�R�"O�� lH� {xeXE�ޖI�B��e"O2ZWϜ<v5�<J�$ճKƪ�P@"OB���;��}�w#R"
�!�G"O� �D�t��h��:j�^��"O2��T"�$bv���ŭ"���"O@��E��!8��󎐥 jPpU"OnHPdA9
Z���pm�<�V�"S"O���w��.� �H@gܢ]����"OV@�v%�4:�2� ��bq����"O�cՀ �,�jM�eIZ�Cd��Q�"OfYS�)E5n��lH5
+���"Ox�q�e�0�a�ҩ�tD�%Z"O��P!D؋
�p�S��J�!��IY�"O���R,�T��m�F��#�&�"O��5�gdx=�M)l�lʑ"O�YA��"=� E��
�d��"O����*�j�ґ	��#;�Z"O��	�;Eb��d�K�T3� �4"O� \U�a��&5�w�ƴy�y��"O�(B��B�(��񖪚�kZ�B "O6A`�GL�z^Tx&�5K �Z�"O<L�	P�y$Uj6";AH�=[5"O\T���A�c�l-:��]�vKe�*D��I�Ȟ|bp�	�']�I�t(ƍ3D��2mPt�f�q�M�1h�*5D�z� `E4%k�!C>Y5����N1D���� Y�:	)g!�^z�J20D�,��%�b)Bv�#T�b�J��,D�4�4��2k:�q����=R4qS�')D���T�ƃH7�h�C����$��¡!D������7u�ԅ�F]�.�H��B,D�h��&9��P�"��(�8<k�*D��$'@��7�7)���-D�t�aBĝ3v�t�� ��V��|��,D�lڤҚ�h��#MO,��,�b.D�t $Ѧ	��%��)64�ӡa.D�؂���_uؠ[4�N�^���A` -D�ԓ��P7�����k�1M�1r� D����dT1n��2v��>�x�Jh>D�4��fߦeM�HX5�L�y�\(q�(D��cp���<��x"񧊺)����8D�TY�	�&N�
�Rc�(8����-7D�T;D�-t���G�%%ԍ�.2D�,��0���p���VB�h�QN.D���SP3%s����jȲ᪉�-D�hI����aTL�)g�ډ�,�Z��&D����H�5t�[�L@�͛�n%D�$`$�ŤAk�l�e�df��KӦ6D��q&k͇C9��r�T���Q��&D�dZ��,�氈!�_��)8g�2D��cS�U�mMP�"1f�2*&y0�=D�\���+,G��ad!��V �LZS.8D��"mD"�c��N�/���ꆅ6D��������ܨ�E�-��eY�!(D��� �ۄP:��[� L�;n��� 9D�b�hIUIL[�I�# ���5D�����p�Y����=�1D�,�Dď "�ް�&� 3}�lMش�9D�(:�F
$� H���	$0Q�1D�,�P��
[+X�(B�ԓ<�<,f�/D���&#ǦPa2���EU�|�P���	.D��Sƴmv�Y� �3K�) &�!D����������0ä�1U$D�l��%��P�@�a�G��v
j��%K%D���0a�] ��!�&�8 ,A�UI#D����L��`��1��\�W��LQpb!D� C)Ϥym�x*��$8�ms��:D����	3����FNՙ_��5Rv�-D���j�=}6Q%�Q	���AI-D��J׏ƽ)Є�hE����Ѥ)D����ܦ-�8�i�ɛ�S[���;D���3�	�b�|���l�ynj��m7D��T.T7!^���F�8Q㖆2D��2��D�*�9�#Nb����1D�D�U*ԙ�vezT�M�"]$8)e�0D�\�&��Y�zX ��K+ �ʇ�-D�0i��7D���GI��]��n,D������4!%�e�Եw�>	BV�7D���a�\R��#��,Zdd|�6�*D�X*!��2u�Ve$퍽Z�Nl�#D�Բ�߿X���	�$3�0,Y�l7D��@�"{��@eǋ2n{�cBB*D�� ԬJ�*��{-
��#
h�A"O��
�h�;n�|���a��1��#g"O2�[H�MԴ����f+��8�"OjU�%)Ʉ��$N�wf�0�"O��z쌄m΍���!;��Q�"Ofx	���l~�Ĳ��N𘍢�"Oh(� 쀥+n�e�Q���P�\��"O���C�ɲF��}��Z�*�b���"O��� ��tj��#�ԈT�,A��"OZ�X���V�� ���ʽM��z�"O R&� uGhxid�]�1���"O����H�}��9�"%�*�l��"O&�h@#@����E��*�fI��"O����W�}ۢ�9e M	��-�"Ov[��ӛR�D��n�'�ʐ�"O4����B�fI�^���(t/�2�yR�ǍO��hBE2b˜�0m���yrIX�%+Fp2�R���a���ȓ%���A%�3[=��'��E�ȓxDt�3�"���1��	ܢlИ�ȓ`Ӕ$�ej��l��$C�&�>̅�;d��4�с�V�2Ƃ�O�ȅ�; 4 9�"��O�X���(�c�
	�ȓQ(�����T14r��a�C�`���ȓ5���`eN�9ۋ�^*['�ȓ`��M8�d�J�P`�ҋ�?
�ȓBΈ�""/EK��cE�#m�I�ȓM��и㣃(&ژ�כyq���ȓL8���i��7��l+��<艄�r��8��^'u�H�*gd��$�l��ȓQ 4�� 琋~��=8�g�6Hf��ȓw�0�y��[�a���+D1d�2��ȓ0����E�]�����.Hȅȓ�Ĝ���2��3BEN�tQ�d�ȓ-+����&@!JB�<���b�nd��;���� ��A��C�(G#eDt���r�PZ!��!A��x��7�1��f,x�J��	c�~y0C���ujĆ�`�HaL��\�L@v ���\e��CAL=��,@N� ����=P� \�ȓ'��Zφ�Y+�\r�ʼp�$}��Ho�!���ӯJH�����I-	����ȓj$,�+P��>�H��a�תyw�I�ȓS�����Ȣ(U$��p,@*9�F`����}�e�P�c�:1��.��:5�X��t\�{'Ձyr��� �XG�y��|�հ��m��E�����2�`�ȓo0�l��(����`L�"
��ȓu�B'�ia`̛qa5<�|X�ȓr�Z�)�U7��C6��fɇ��R�����:+�ؠV��=x��ȓ-�
���{m�0H� ����9�ȓTC�[Ip�RYct�7r�8��ȓM�VPc�.g�|�ʐ�4'R�(��u+X{OQ��@3*/
����F�ؐ��9[�V�p�#��%#l�ȓqg�K��5��uP�o�!�F���;�,�h&i.&Ah}*B*�1��9��u��4)��._:�M�!�-zV��ȓ.VɊ�%O���і�*(���ȓU�2\��
M�䴉U`E?'�F@���ԡ@$�ȅ��ࡔ$�6ho��ȓq5��aֻa�\Z���2Rzq��i&ܱ�q
���D*�,��#^�-��S�? ��*ЌѺ53�P!�fک-�:�P�"O�pHH�>h�}�`'ɭ<�`�Re"OP��Ǡp@����U	s�R-@�"O�8i���-~(,�5�;m��5�c"OL�g%P 7#?u(�̨�"O���R� ����ψ�.!jԙ�"O��p�=WEY���h(�R"O8)0���" 4L��e4H��&"OpĨ�AÌƍ`�O�SK��Q$"O ��g��y�/�3��� �"O�%�T�ƢE!���w�νkƮX3�"Ox�q��Z�vyfa��F�&e�6�*�"O�"H�?*f�Q�T�k�Hq��"O��i��,��h���jl:�"O�|�e	��|�"��H�oE蝻P"O� ��X<=
�����g(ҝ�"O���J#V��,�%&5c�ݚ�"O���]1L,d�I#p$I�`c!򤀯Ox������&2��z#�܇�!��W�~������i�0QzI�$�!�dTLV����|�Ƞ�Qh��U�!������g �%I�8�w	T�6�!򄎲y����/K��C��9s!�$U����`�X�����Pa��)]!�$֏h�4����>��e��/���!�ę%"U��jÍ�l�tg����!�d��h��a�j��*צ�����9BP!����>�Б���!�Gɴm?!�D�8xN|:�똖j�V5��春Z#!�D^.lٶ1��Y�~LT���:!�$��_&��#է�:-`2��ń��!�����y�ᣒ /�>��f/F�!��O��
Ê�;����E�
�!�$F=`܄q���$r_�����SH�!��4a~��CtGF�,ջUɀ&@o!��	^6�T"��S����(H�!�dF�B<^�!���qm� ��핛=�!�$E*����B��}j24���w�@��C��"�-�	w�T�	A(O�u��>"���@ɝ�8!6��W�ݫ�R$��0���b�̪)�>iŪd)��)D�p1$ˁ�t�P��	��G�(D��p�E�*�6lya@͎Nb�a��(D���#C��V����	9Vǜ$��&D�x��阰bz��ڃ�XӒDi�n)D��	�	 �K�}�4%�<V0tPa&D����M�kUd�b#���K�ƐR�F D�|�R
�"��Т���9_0v����<D�|"2���� ��G�����@<D���$T�x��c��WoD��я�s�<a��K���"#�>�J�2�Jp�<���G:[Xy���W��B���A�<�t)٪<�^�1a�[�6���q����<A3HC�ѣ���,|����p�<�0+Pj#,���A6��$�0� H�<9 ��~m%���~݈Q��@�<�\i�(\���ԍd����W�!��^�03�U�� Ł�l4�ʚ"�!�$@خ�H�`�w��8:��M�=!�d��2V�A�HF;�P��J<e�!�
�C���3/�p0�p�
C�E�!��ʝf�x�9���!��İÈL.�!�ިmͬ�@q�U�<��dI�L�!�D�W���	�}!l�נ��&�!�� �d�ud
6D��ccմp��ա7"O��J�$��Ot��䉩<�|,��"O���� VQ���D#jTF��"OjT���]<��	���O�@�"O8ݐ��7Z��uR"
T:HbZ��U"O*13O��=#�)�$*��`"ON��'��$m��$�F����DzA"O젪b�C'a@���jY�F�Ɉ"O����
]^��4I5\A{T"O�=���F>y���v犪o�r� "O�����1uд��/�o�``T"O�L30 ̿8��c��OU�� "O̘WA$y�@@	�0pF �"O�ӗ��%7�훇�V�|z�"O>�2F,̲W&�%Ё^E���Z5"O��%���F����`�0@��"O�a����J�r�Yr	U!>����1"O�!p�*]����[#Έ&	��t�"OTqG)"�����Ȯzx�@�"O"`�C8{b%���|a�2�'j��d��K	��F*,����'E�4��� �L�xu��' iB@z�'�S�$E�oO�X�%���  k�'�rL����d� ������'qj؉%L�=l�(E�����p��'��!�HW�,���a�ǵj�-�
�'n�o !�ܚ�ǋ����L�<q`�Y\x՚���<[�ZW�G�<a�Cg$�K���JI�����y�T�3� �yBD�4nau���y�ЋT��Y�D.�(��#$+���y�%]"=�<��I�#}n=sa��yҩ��~ٛ��͵l�~�#M%�y"H�b��1�铫����IV��ybC^�u�r���Z��k���?�y��#d��8x�h��'��C6	��y�dM
I�$��f�N��f�ٛ�yR!�#K2ڥ1�e��7@�Q��*�y�ę�g� jT瀷"�X����y�@E2m+BI:FO��dʧNǑ�y�C0;�(�b��2)�p%�D��y�I�fdI�G�߅$�B��ƋC&�y�� %4Q�-�D�X�l	"A�Kנ�y��U= �^�s�&�4i����"'Y�yB,��NV�a����a�rL8m	�y��G9�rفE��	��J�@�yRH7{u�E������	��KQ��y�f�5m-F���cѴ>{h4��m�y���|��T�燙6���bc�P�y���kdY���ķ^��YX3/L��y��4oz�b�(��(ۈ�q�ύ=�yR`ݾ?z�`�lC�'����R�'�$�0�OݞQ�z�2Ba�=��'2݂g�
	f�XTZ��Q�
�n9��' ��Ġ�_���@S���j���'E�@Cb��-p�*e��	Mte��'y�xYѦ�:]�~��T�
V�d��'�qQ��N#Q����$�7b�<��'��Ր*�U� �@�b�2���'Az(�3�lFP�C/R�V�Q	�'s<x07%�"jeH��O�X��ٹ�'�
���T�pS�{��H<b%�=�'୛vi�AO�e�$Ņ�а	�'�ha;g
���U�T뒟VV��8	��� �aW�T Hx5��FQax���D"O`�rR-�6
��<�҆�	ez]�"O��Q���?����LRb*��1�"ONQ�u�޹_(�pkN d�@M�@"O����FX}�����L} �Q"Or�k�˃����eӲD�*��%"O-R��""��X0�W l8�"O�d[T�Ðy�T\��M\�i.!""O�\���C�E6��y��+Vd�x�%"O�uK1K;ʐDk�;BJL��"Ol8�TB�!��Dr���?TA~��"O�z��
��������ub�0�"O!P dP,/�����&��R3"O���fY�CX=�V�XZ�,�"ONTs���7T�.���ȏ<H��A�"O�z��S�`��`�.��l>R�AP"Ob����ϸ0����M�m*M��"O�h$K�����Ћ#N�ȕ�"O�-2 I &Z�X�
06�nTa"OEqA�Ӵi������!(LY"O֥a��%+�@�u�L�[��"OP�fݽfJ��SF�?d����g"Oحs�*߹S1��`�=,����"O*t!
;��t@ ��L(
U"O��z&��k��l���ؿ\}���"O"0S�KVwR��%	H4Gf�d�""O�L��#�
1X��kC/QO0�{�"O,��P�I-��(�Щh��l��"O@ea$�N�62���$IrP|0�"O�T*#䑪7��xG	L3
�t��"O4m��(�8|T�q�ߑ(L�m�&"O��1��F�s�e3a. zb�tX"Oı�d�K,P�I�3���Q��L�"O��gH�w�������aC�"O��&#��R��@ⲅ_�*�"�i�"O���f%P�Y��3��Y8Ę8�!"O�#0"�]7��	!-�W���(B"O,x"�"�(X�s��(#{ �Xg"O�Rʇ�\z�l11�.m�K�"O���%��Q#B�:���?mlFT#�'�6�	sˑ�we����I�3]F�-��'UL� ���VĈa�#X���+	�'�vI��S�Y�z�R6��)|�d@	�'尐�Å�
�b�+#�%u� �9	�'$��{����}	��/E�$Y���~�<q���`_Y��`�+9�d�8u��n�<��o	�K�l�SgJ�~�Ct)Vt�<�AHF�i0�l+�)Ҥ���7p�<i��R�\��Бp!J�y�j��c�k�<)0�����4c��ӆi
f�<����J ����H���K�<T�_�=ْ&Ȏ?�"=��L�]�<�v�JQ���k�1�B�ʠ*�N�<� eL+c}�Dc�`&[\�e��	H`�<ف��>j$(�iv�a�.eJ#��\�<"
G7<�U��E�6���]�<�e�
:X]J�{�Q@z���m\V�<�7�9�TL"��Ep���6E�j�<�p�U J)�?f:� GA�Z�<a��ƪ%߼�� Y���@���V�<)cG�)Z�ĊG/�2�(��MO�<�5FܮF<�05`�}�i�C͇F�<)�, A�$d�)�0�{��n�<��(��p�������>Y�>�;p$�p�<� r|�i��������F�hx��*O����Y9u�y���#(X]�	�'�ă�� ��������� �'�F�P3_f�s�	I�e��Z�'��i����^,`�T��Yt@Z�'t1�t�RYL���t���X��)�':��RrC
$D⨺��D�RZ�'M��q�ߢ��⦄C6�
�
�'��:4�L�f�����%.d�(�' $�fG�:�iX$���"t ��'ozD�w���z���KA����'��!�g��#�hZcO�_�����'z48����C~�i��ODXq	�' .����$���CcբEe����'o�łǩ `f�Y[c�0B�PĚ�',��(��H�f>���wa3c\l��'���fj�I��\�g/_(%�t�
�'�u���L�����'���	�'$8��w�Э)���?M͒���'b�p�Q�	?A����EC�L���
�'����G�a��6�͈I����'�����4�V�k��̭F}Z	�'Y>a�I��4�	х�3Bc��'�4@�T�PO��A)�4E��
�'i�˖��/NsT���-^0�B�j	�'�a��oC�R~������8K㓇�#Y4��DJL3Lh;$��xx0��	�1Oƴs��@7Y��9lN�ظ�0"O�<8$��J��%ˆ��� �R�p"O�!;%�͞߲u l[�H�.�B�"O�q���s?t1@�ȵUeu��K9�&��>1�'�ܨ���ڊ|���0� +2^��'Y�e��@�3�p	U*'���;N��%��D��d0D���GI�u)�[#
Д�0>�H>�� �n<��2���6c"01�LB�<	�q����`�2S��%��@�<��D��a��a�L�܌a���a?�0��_�'"F�!&DǥG�v� bE˿#K�#���O|�$�c����g�a�L͜5+�KQ���H��$LO�O.,�c��O�]�'�]�Y�O̢=Q���:{������r �2j��{��$���;d��<�^����ɳvq!��!e��Y�6��&�l\� ([i��hO�j��&K,jn��H(n���rǳi���'k
��� 73�@��O�z=�ղ�'��e����	-DX��^�k��'C��+E�Q��C&���Ó�hOm��$�^E�7�_�A f��'*F�"�c"R_��!�d�,{�4�k�{a=ғ����)h��T�q�����oI�j�����\���&Hӿik����̏q��P��I&D��c7��l�J�����ZX�dXgy��'��~��)�	F�D�c� ]5��Ӥ�B
	�NC䉝hV���кW��3��+ �"<��	�f��QN��f�6�
tIX�@Y��D"�P3�����~�B�E͐&�� �'$�'�ў�+�T}QF�Ŷ̂��DMJ�B&C�ɫ}U U!�#@�w4e�r� ^C䉊Wd��a�ϯ);�]S��D8��$ІL*��8e��0C�T$3�&�%$]��
O�(T*
��4�0V�Rn���"O��{OQ�gӖ�+$l\�R"O��[���xT LY(��y�"O8�
�"A���Z�!˄ExI�_�@F{J|Rq�O� �!�#�½��ѩ2
X��8�"O*<��h�y1��+��T�e"O�|p��J��^���&B=�6�pE"Oµ�aO�2��9��D�P��"O�Q�B�V�h����1g\6R��'�Q��ۦ'�x��0�TA�g��e�!�>D�(j7ݣzp��Є)|�aвh=��s�	Y�'����5d  �a\2?�TL�!��	y�!�i�Q(բ��'ĄaXr�$��p��	7 }����#  ��R4��C��,J�\�Am��M�*xKFJ�<`�|�	C}R�'�򙘁%U.,��}�����'0!H"�Z��0�Q��UL�d��{1�����'x�#Ҵ"����4N�:�y���B�u�}i���7kv����[�a!��F�$W>���:i4����Q�a�O�*�RJ0l���c�(�)-�^G�p��f��4��5����6�LVچi���8�ab,�X���,�T��%'Z�X�l�ӓ��'��qC�č&u�h�D��%�c�	y�<qpA��T�Ԅ:�.�	ypi	"�9��'���	1���n"|λOC$a�sc�z�cqeۓ0�| )7d=�S��M���km<�K���s�����L�<A�	O��Nз$��G�������R�<��	v%�$�ٻߘT��d�j� ����k�� �i��-��a#��<r�n�ȓ?T��`�`
@���Ɗ�D�T@�ȓa��d·;o��b �17n����?q�B5k��J��|��dn�c�<Y���(
4�S�)����vgh�<�@�ld�XrfBSa y��I�<i4�� i1�}��w�TH�CǊJ��By�~*��A�8�A{��$���GM�<�'�H�	܊}��ᘁX���{C.�I�<)�K%�,�A�3�̙��G�<q�#K�R���:U@��S�UW�<YA*��z�^YFh�9n(X�$�W�<�Ď%McT�'�	S�Q*' �O�<	�C��>�J ���$R�"�BQfX�4�Oޑb�I)b� �ҳ�YU�0�;q"O��Ǌ�<.���P��� s�p0"O�q�$F�0��	#M_�f��"O��0�ݐj�v(��F�4����is��J�[��\��MP�}/�ı'���~f!�G�W��Z5FZ3gw�}��ʐ�+�a|��|rD��@28,Ѕ��;<�-�m��0=q��ϙI��aI���\� ��Ą����OP#~R����l�bxڧ%]�A���@�u�<�7�+�=�!	�m�n�PS��u�Iw���O�؉�s���D�dc�Qԕ:�'i��2B`�	E��� ��q�8	�'�^30�0� ��ҁH�l��5��'�>��O*X�	 ��ښu�����(O��j��K�0��r��1*r8��"OD��N�S6*�W��d�V8����pE{��)�������D��0+�6o��hO�^���Nu�P���1c�[�c+�佟���I��2�����aH��V�vY<C����M�%G�%���ÎV�c����cPm�<)�=�Ε��aL�xN"��ĎP�<��B�<Q��@a[8{�u�W�JI�<�U&Ħ"�,h��^5I^TEZ�G�^{xFy���'�P�!%�.!�|�R��<��2�'yx��D<W�n��ր(Z�H�aTh����x
� �EH�+RXx|ph͡N��jP����G�$�\�H�:��j�n�r��V�E��yҤ�?�NB�F�g�v,�7�Y����4�S�O�Ѕz��\�
_�t��
 ����'���&�1v�y1G��u�~��'�^!hgAB%�teX�b�k��"	�'0dY��e� �`���MԨq�B�@�'-�UJ2A!j4@����1:j�|��'�����R)����S`�3%�m��'J�,b��4i��9K�$�1��}��'3ў�D{�&�b��	��	7۬,;�Eğ�y+�-����E��r��I���D'�OT����(+�6�3fNz�n%`""OM�7�4b`-�6��t0��%"O\���ʏ�d��8���ϭ_in,h�"O����r=&�1��E>q_"%2�"O�m�ai7[���g�?,�z�8�"OR$Hb�B!l|�0'���V���"O�Ikr��#og��B3#ko�$8�"O������%.ܚ$IF�H�$�Q"O���f����I�PH#YJ���"OJ ����r��D�
�lY�"O̥��c�z�qI2l������"Ov��fJ�g��D��I�F� trT"O�(���^�<Z��Ǡ��,�"O�)�,�,h)��B'�{W�|�"O� �1@ح���a�&��mH"0Q�"O�0�6Jh\X`߷t�n��"O�u��fH,�p���
T�A�G"O�8!�jZ> B qfe�)D7�<��"O���e	�uR`؀��K�$�A�"O�MS dȀ8��DK�[\�;7"O�X`uHP>d�l٢�ʝ�AY4��"OP ��o����kN�Yz�	�"O��wf��zNz!C�a�|G
lPv"O��g�'mz`:Ņ	0!���Q"O�,���P0 	YB��6�Q2�"O� ��$X�N��P�;{|�}�"O��ᗢ���<c���<�6,3�"O�a2�l��4�����gd���"Obm9�� ��x�@�Aw`��Y�"O�� g�\*�1+��'_��b�"O�M�� 
=z���M�UEp9	�"O.�k$iO0T2^	��N?=&Ir"O�;��&oLȚ��U�(��"O|4x�-s��E�7'�9�"O*��ը��	���./+J��"O��k���26�`H��������r"O�
��	*I�VT���Ԩ`����u"O� h��Âl�$�p�<E���"O蘂��N�!�f�Z&g��~u�
��`,h�jO�/��hcB�G,b}1O�Ts�'�)uج���
"3��$�t"O���F�ρF�I�e�/yT��"O��F�}��$�5���KT��"O���@˹f��z�&w�� +F"O� �
k'�HP��NƸs�"OT	�BX���S!�J�o[-	s"O��-*��i3�dg�HBC"O�)�"B@�@(p�/�4Cҥ"O��Z��L&(�BӤA8ohZ�#2"Ob��P���,�WŚTf��"O�P�	��0n�9��J84I�I�"O�(�i�YW�I:3)1-� ��`"O.@��+5��=�7G�;#�^ ��"O� ������ �*U$A]� HQ"Op|օ	�i8ZUۣO�NQ�e"O�l2� B�L[���Vw�4ѣ"O��0�kJ&#�Љ9cx��Qb"O:$C��RJ���V�v�!r"O��0LH ^jq1����U��"O4�R�oN�W�	@�;l���Cu"O:HR�G�=���N��)4�H�"O$�W+�5W�P]U̒�Q&I�"OV�R��ǭd�f�f�Z"`* J�"O���S��32��m�C*�=Q�9�"O��1��;�v���S>AH���1"O�%	D�
�Q�V��)6Q4� U��w�<�WF�2�:YU��&|�f8� ,�V�<IWh0V�^\qQ�յ ^�� �RR�<�􇛚1�n]� �Ӭ\V�ɲ��Tt�'7ڐ���74bz�nZ�O�vQ7�?�������ؑX'��t���9D�`BD`�#r�tXbw��>��!Ko��E�4:W(%w������2U�biJ��9�P���㖼z2f��dZ�2Hx
#"O�8uJ��D	����dڵO>0qӓ�� Q��cԀK>M�Q��c�?��)���(Of�W�M&%�P  <0�r-"t�>A�� ya���F�yV�!�0��('U�=�u/Ƈ��:"�_3
�ԐB�Z�џ�C�H��.rWm,xa��_7�ZE���v�b9�B�W� ��1y�'�<�;X�D�ŭ&{E�T*e�>N@�I��aZ��i���5z:����!^����ʟ�/����kZ���u�ȟ��
WBO�I�̠x⍝.	�0���/Z.q&�X���$����0��[���*wb�Ψh��]��4���?���ru�r��@eҪl
4�s�-V$mؐ��R(��֠�?2��b?-����49�V�h�JںX��
�ګAh�%0���fh�KX�A��@[h��q��H�t���D��%%��� C�n�jI�!n�!��qb�+��/<X��^Zr��#	+s���b ��R�����G;{7��
w�	.[��9�@��C^0�EF�M��,��N� -bQXADų ]f"<q���2BhL Z��%��O,(h��v�-Q"j�ri��8���F�kΨ�*E"��"�vA����.-l���J�V/r�Z�V��8��b�˽6�� �`�;��B�CL�XJ-���Ɣ7V��a�E�����E@�y`�SN�>EKE�1�����`&;�d�����6QZ\H�mݯJ^u�3�G�M�2Qc�52����4@�8�n�BM
9Z�S�p8Fl����OE��D��Pf*�c7#ŅfP�$N
@N=�O&�	��?'y��D�/��a gҲ=+�t�D�C�;LN4�2���qz<��	�Il(|��š,��IX�S09#�'XZs��"�� A�l6�l�P���6�0�12��"�ء֣�4�P8Co��'�����o1�p�P�D�7�L�)���!Ǌ����R�4��-Q�+�6�H�Q��8y�<YcCl�R��s�BY�F��< �n��s&��mN�գs+a���hF��l�$���'58�R&O�cnY� �H�hE��ۣ��(a���8�AW�g����]�!���'U�W�q��I>�a�O�5(��P�*7�TXSb�2
耪���$D]�RÉ3.@���Qtp�
�,VX$jF�[;~��=�����@�Ѓ��D!`�����X�\@ PD�=*[B:�)��K&H[��D�:d�B�dXª���);E+G�8Yi��!��kA��N�2��B�ʓh�@ �u%WU��[�E�'5��3#�V]Wj�x����*+��H+��ԙ��ח_2DY�b�=̎��'�bh����0z!��ۥ*�:��E{#�M/�	�G�8Y�b��[�I�OL(ig�T�w���&f�;,�L��
�.z�`�	
�E��j�	�p���a↉0��̚��-��I�d,U���\".��f�w��V]�i����E^�_�v�aM>�e�� [�`�!勁�g/�6l�9_��	����R��kƀ�?{y��c���(U�H��ň�����&5����ϡMGz@Q�L9��0I�C��~H���He)�F��0���U�[�P���EVv�۟,r��%YbHPTѕ���d����%�[�FD<�D�����i�!��i����Ā1N����a��0���BB0��'�1OR9� ��5GS�%k�
s� ���`�IKd�=^��� �4"U�J�0m��,����Q���G��4:'Vb�THs"[3|Ϩ��mΣ3rx�H�n�6#z�!��l;}�̝
hM�t;VO5<���!d�B5q](`�W퀅f��H�H�/�"@3�B�x� DXf��e��'���̟��A3A�׆l�I���&�� �p[��:�Ĕ;A���M�����lW�!��-��e �i��u�t`R8-�n�j2*]�UPX2 ߭WZ&P$A��$[�I;�Ф@��) 	��"���DjuJ�J�f��YPZw�r�֪�9JSЀ8��%+P"�m�l�l���	2�|T�"ՠ�t�֊ǸHUޜ �n�/Zb�;i�<0���ζ����Si��� H!��1C�@#Q��;;��t�!���2$��T>Q
S��>V<��l7"!��Q����pX��C/)�Hd+2l�0�۬m<~��l�7 '��1��J��0�%jC 2�C��k~�)c��6IRhh��R�=ْ9�Vg[10�52���&"����Y�lq���Q�r�^)��D�O�d���G�z���B�Qc����ץc��"c��;x���	tQ�\����'F�ܨ�c��/45��8�卧�Jqr�L͛<���bc��p]�X�!�%B�ָ�s>��E�*���u�T�X^T9�1o?�	 Y[X�^u�t��0��T�\5�Ee����A�S1˦\�D�̟&�p��*-%���	�
5Ov��Y�-v�R�KH(i`�(�~Z��zޅi ��6<~�Ps $N�"�Pf	��r	�;S��0@]��jCa���AG`�r��d���0D8�P���H����$�>i��-T@C�u�K��^FV��&���: �p�	�Oc,��p��0B ބ�RǍ��`񪄦B
<�(c��L�/}���N`$���-�dЮX��`8Q!�����sGɀ#�"\���Z�L�{ K��u�"=�d�\�|�'M� �� j<)`�6?��Rъ1��+�.��Q�pã��:*ĉ'�D��sY�
��s�����������W�𡃄^(SбO�(�WjT�h@�&�f6Ti��'�{�N��%V���Ӑe��J�#h�%_���,؂����GP:��Gҫը�"Վ�6>��ٱ(F-_nx�h��Q��a+���f����F'.�&E�8�| 8a��bv��G�׹D�=��� `� ��zvv�s�_�jr���' Z8���P1�\�ς�y$�Ń<[���`�(li!�
����}�h@
���L�P��zd��|�n�pfN�j�8%+�`X��j��RG�̹���͟nv�Y{�k*��KGE���>5y��)Fͽ~�ƞy4�Qv�L*@�!i�n�<I��'t*���ۓez�1�Fo~"d�%:��S��_(�?�����{�y�6bIe�8d��-mL,�ɗn!��@q�3@�������%z��?�;B�T����5s�Np�s�X��~�:�x��ޱS��L<7h3vz���+F�0(lYg@� 9k��i�v�8&f��)�5�@(P�g�:����b`TOܹ�F�n��(x��٢���0��;Qn���䟝�� s$��Db0RG*ͣ{K,=��JR�;��ey3�_���Ё�$R�[� ��c�5���p�'��ܮ2��H��L#T<D`B�-}�YD+�d��D`hj�PĦlT��P��
Jf��FVF�6س�Æ G:�4(��R�o�:xydI#�P"cC�YR���خD�(���!:8̸��ZG��:$��S4�lڄ�����+i�-rp��(���!O
�	!�F]�J8�6@��M�!�$��#JJ�	b�	S��5���\=R&X�!��&D�(��Xl?��S�A��D�A�A�W��!���?T)���;��D�B�+g�Z�[��:Ժ����`�H�d��0ȉ��VMl��S(��7�RY�D��	x��ue��>�\J�K��@XVax�)�R�d�t����=��D�L�@����O�,"��C�5������=��ȷ��2"tQ[��¨��GX6ҾA��W4$r!�D�1R���+�*O`z	�,��d/ڥ[�#��(��t������:>H��Q˂�Nb~��c���wU�ej ���s���'��~��	�'W�qR�C�$N���0 Cm�pA��'�5J}�Mψ 7܉F(��x}xa�H��`��A�l�xU��On  d��F?�`�G̫EN��f�'nF!�qH��:nH�`�"��
6�WH�64��W
+����!*A�y�paSsA�t��"i�:�X�O>�2):��ORiyW���Z`��I�KY����'�Đ�nְ/
�q�BI+,���u���hah�FBuY1�R[��!��.*��,��(�O\�I�E�$-*#�a� �
aP��WH��z��we���\�PfEk?9_4�M�Fg�0uH�"�>Ch�d�i2	�#\y� �A�y��@s%嗖%�$��̡r�_X�
�Hמ0���~�V:���<k����b@�x�R�I�#�=O~ɫ�]�/V�	��mʃ�^4u��7�Qy"O�VN咂��sФ�CB�33p�A����*���7�|�*���9g���6$��8�'��jf�
����f��`����'��\ 5����M�p&޼9��IQEV`[�K5��ՙ��i�1�Q�?�t�5f� 3�.y�K>�&P�2�(u�3�<�� 2��fG@�#$*p:�I�(;c��b�g�5W�xa¡HB�1�0�Γz�Ek�nV��:P������'5U�t}�ш��)�tAWg�Q�W���D��ո���3Jr�qfY|g�LK4�]y
�-�T���	q� ���T��d��&��d��e!q�L�k�AZ���>f�Axf�O�h�6MP�P��D���e��OlY�
K<,S�D��?����Dq����B%����3�	ZIJ\G���.P�@`!��;�����՟���FI')��4���<(=�(�ţĹ;k�T���
���컂c
R�I�a7ꉙ�� �t� G�H]@=��g�*�0$�
�
�*�!<�`��AՎ~�%h	$�0=�*A��l��5Y�ԦG���.Ӻ�#��a �@�i�����&T��R]N��Zp�pa�@L��8�O
�r�m��68 �D�X�a�NA`���Tڰ�F"hS`��S�!tޅ�ׯ5���A�>��=ѴBO}��q`��?�e����H#�b>E��KؑI#䐰W�Y>u�2�K�+ח|����IV�l��c��C85�p7M�O2�"փ̚z�`QX7�/-��'��՚��Ǡg֬��K�8����̋+d(V��N��4��M3]î��B���`  ���=���e�
ɟ$6*̍ejAQlY�+0�Ŋ��N3������0Ȇi�Bl�D�/g�%��eG7^���Y���ϖ���Q'{�8H��
T�r��ٚ�جz�a��*<�TyJGj߯-H�����z�6`�
U�v��Ū�dX�c���)�,�
1@�%_Nv��ATS~2��H���
�#Ǫ#��a{��&X,@�k	.��IH2.<A�W���9R����+��Eޖd������*R\p��@��iD��i�)j>ɁR��4Z��w�J�R�HUҌJ�eK�CN*�˅�5v&i����+#S�xI�P#�O^�P	d�#f�B)�-������㮅r��P�'%�2�N,�p��i�0=2V$#&R,,��%��#$Wʡ������k����tT0)��\�v�0��i�;%!~t���đg3ā�P�#��kb"zD AF��
v
��W�ߕ<�L4���!��yA"(~b�Q��ē^*qO��Y4I-e�htm��T�sSN=�`�s��{��DAä�
���#a�ƹVS����6Iu��N���`�{%e�z��LQӄ�~bW˜�Jb��q� �B���[B����A,�����6�b�K�i�8>
�9Ԣ�(����#��-��ޝ_���a��:"�6(
@��J���(
؀��~���wm�*��9�T��]-fM8�� [f��QC�1 ���Lɦ��O�n=��C�8�u@U�O���cf���I��G�#BD��D��Va���W��d��d��E1B��"u��4l&,��,�T;d�-SUlpc���2n������0@��b��53`<zcF�.�V�C�S	��$��/B(
@J5BQD_A����0ʂR�P�g�N�M zu�t�S���H��H���p�Nd�0���N��t�I���hI�M�S�>� �u��E������G�)��pYT���,X� �@�$w>�OS��%�X�����A���a�97��iR�Śh!�pThZ�
�L�$�^��6�1�ەB��r2��F��I9����Y��ɱ^�f1�b���O�E!��N"[��uy��[�(7h�H_�<�B����D�"����G3W��]�3���9�J<�	�;x����5<��Lб&4�%�<ّFr�F.�9|�Ku���:��d�f�6�9����j�Q�D!���b��T7�R��P��\<�B��x'l� �D�^��C�&\-
��'b�!��m*t��: �i��B��|/|�@h��?��s@^�k�Y!-���h�I�06D�'�Xh<9�+ٟu�(5ӗ$R�Z?@��߂#���Iw�3|K8���#@d��	x«Yv�8���-X8dQ[���)��0T�����yP,Y�r�3,Ob�JS+�� ��p�pH&5$�AP�܈ /~|c���%ET�5z��Y� �ޑ8�BG6R��q2�e�N�	����n'Z��6�z����A��K��'��c����r�*U�@-*r����6���4& !�i��Z\�!�Vx�\�"�[1iN�a���'�h���I�a�R��� �n/�Q�gd�4	s��D�O.u˦bO�7|I`��R�d�H��@4m*�Q�Q�g� �ݎ7�h�P��P�is�<ʳ�['v�B�I�y`5�j�;O0jH��E@/�0@���9�ب�CF�*V��bn�4.|n���L�I<~h��%��.��I�.��D`[ӢAˇl�g���� �4��m�F���<��I�d�E!������p�jK��WL��Ex���.��H7�׳B�j�-���O:��U���7���	��Αs�6!(��xʓ� ��E�h�%U��K�֟�� F.��ՠ
�T��$�:,�yK�.P=	�� �k%�O"�9��F�x�$Tʀg��G%��PӞ5|�����%�?qt��.�yq�G�|�(DҠ�ODd�w���� ��?���C���&�B�'�eʡ(�^�-[1 ���a�����i�z����@��t��(�V�1kq@M��4�V���ɎH�.`�FT+��E�牎I�&t���� (��IPs�i֪TZ'�Y�ef$�b�� ��OP�0s���	�(8G�8O�� @̀*��@��*V'.��	�!�֧/���q����ڥ�#���M���n����)̨%�j)��  �a~!���,5� AE���B3� ��W�O&��JÊ�U���H����U%��O�$]��]�&���@Ǆ�^���Ɠ]ÂLJ&�:P� Q��,G� 	�lH$d`�(2�O��ه���vX�2b��,��B"�'j�`E�Z�.Sq�`�����lV(�ZC�
2�C��!>��b����Е� B䉽H���p�ڰJ��	��J�f�PB�I��hq��A���"��ȑe6B��dL$��U#�,]�Y��E*ee�C�ɢFȹ ��~	��
�Gp�"O�s�胏ug��DHSM�t��"OX�凰ڂ2��B)\�H�k"O�`CI�?5K���PO2{�Xљ�"O����n,j��M	y���"O��a�X�%h����]�R��	"Of*�ץb���zP[&'Q��s�"O�`G��:+r]����9bz=�"O���D#ɖL�J���H\�؃"O`(���1'^ȉ�#��bM(p�T"OPa��-�9x�X=����Ĩd"O�xٵŔ�b���6�N	��ɱ`"OR9����T��(�h��%��-[v"Ov�8�n�i����Y �"O�	�·�@E��!rEE�;��!�P"O^�ASmB�!P|�b��.=St � "O��Q�]I昳"��cu�T�"O4Z�Z$8�&G��mfj�[�"Oia.W,cf�#���	,v]9"O�H���3 *Hc�A);�"O�p��c҂US�نG��}q�"O�]����+����g/ZD칊f"Or�	�&��1+��½1�`�"O`����C�R^dS�Ú�(�r�"OH�4��?"�"LA(ơf���"O�����g�U��	��}h4{�"O��·i<<�f(_8d Yt"O~��f�Z�V�xr�W�b`��"O� d��0 �::ھ�E�*yT 3"OB���M��f��s��>���Y�"Ov�acC
���p�'�"%��]��"O<��B+� �w�T��z��W"O�axDf�?DF=���e��1"OD�j2D.;@�'�2^�b(�"Oy�!��`R"a�E6�%�"O������q�x1���E�bF\�G"Ot �`�8P4�p� _�:̝�"ON`����	�vL�� Bp-���"Ol`��¨t}�W�1v���'"OdPX儗�C�^�j���.���2"O�����I$��{#��"���y�"O�q���Zy�2s'�5��Ȳ�"O�y`􊝵^.���	�;yV�"O��Y�#�%H���p�d�2OV�q�"O
T;�o�f:���^��fD@�"O&�:��s(p$*��<E|�3�"Ot����5G�XQ�k\��V"Oq a�a�4$Q�@��0�v��'H�< ��~��"k\��l؂`8�����y�@�D�r���#אD ��&��ՔH	0�S&S�"V��fPTjs�H��1 d XC�<Qt���
���5��T6p�{��l�trl �+Or�c�(L|�g���p�ÚW��yi�gZ Y��C�Idw��y�
M�4K�� �l�,7-f�a��ٟ4�ޘ{��Z3�a{�fէbЌ�b7ִ�P�B�lQ u:&��.w�bE;`/U�<�Er�M+��]8Z��Ek	#V�I��OC��(p��V��+C�8r�^I��nJR�%0�v�+�O(�9�E�"�d�`7��.��k���[r�9�*�u�"P�R��B�&��e��f�p��/��	c�:�f�
7��7�,2���&��H�d��PI4��N%Ѝ�R��L�'wf�Pd�9�Ș$Od���E�h@��3��L�P��Q�;[-V@�����<����E��O���(+H�
mbC^���(j@L�;L�&�x�v�*� �1�6���R*@���,�z�r(�22�6��i�4P	�\˓b�" ������p}kE J�8.��0"�)�G@8�5Bw�6\�Ǘ�[��X�B;,r���i���T�����E4��@��^�j���J��Y��H�A�9	!l��iG(�\��5-�6���9c�]p�8�H &`qORi`ɓ1*"�Q7>��ز@CE�8	�Ow|��E
5sQ:a�W��;�"�ǖ/Z�&}S7�S�y�@��iC�)r���S5pU4A��M?�,ʚw[�q�	�4n�j�zW�_36b�(���\���D��ƭr9��F�^�}�Y>���,M< 2@iw͆x��L9C*Zg�E ���	Z,���3�$ȕ��Q�Ƽ(a��|��lq�J�_m�e$���MՑ � ����0R�eI�eE�R	��1\�� CaE�0Tj8T�T%�0�5��1\�qq�ED�V��@�
ʌ8��b�=OBA!g;�0 �ɡ~"U���Ts�B�L���&"�TC׏��޽�'&�j��p��#�"u�,p���۟����2v1:�Gρpʑ�'�D�l��H� c� ~� 0��|�p
s�0<��d)W��=�XX�.7?�r.�rڙ@*\,BdF��S/�8� ����W]�N>dx(�K!}� �0d�!\zݩDGv��ڧ
 "K@!q��H3|\XwKM"x�
,���ԓ$Tt���P*�*�����4E�̊@D�P ��(,�0AK�ѥʲ�� D
� ���g�Ɉ��S���8�� ;�|ћ葬2�$T�\�X�"�I������z�9�W��� "�5����kT�E;zr|�+�0s�B����ʝy�J��''׻w ()GK4�I�p- =K��,Y1�؉w�E8~�H�����+�]�$8R�ܱ���M-�t�"�&{A2�E�=?���8I��PB�
�9R�4���E �nd0ԇİj�p��j^���'�t�e*��2��	�~= (���7y;�*�/��tN�8�G�)F.���ʉr Pt�D�9rW���
����Q1u��a�h[>H%��nA	h�	{7NJS�Z� ���@,T�XׯύL����E�Ԉe����r���$�'�N�`��F"F�0�N�H�����ƌ�j�#�4�lI��MC���Ec��S1���W��8P�p�ٖ6�0y85#N�6�n�i�T̓]O�]CbMZ-F3�0���Xh̠��D]5&Ӫ�:��]]����
_H�u#��.@9�,�M���� �,<�HxFH�<%�!#��Y��%���`������]� 霹�O��g�ĸfN�Ǡ�� P��bܳ3��Q���ܘ5���h�a��,t�-������A�	-�ѵ0�{f��&$��X�M�!GL"P��LZWP-vP�5�[4s��һ�~�S�K�ܸ�ȃF�qm&��QV�9��:�͜����x�fT't`�a��ƖO��'a�m�s���J��ՉA뛉beVQ�&ߔ;xzt�t��ߺ�Q�L�*��zj��Ք@sGϥ�x�2kI��Δ�Qm��4v�p�a�̥*�� J`�L�М`#����Q��lS5IZt�"���B��	�@��I� a�4��.�^�j��ݣ
ڐę�̓5���9s�:H3���2L�L�ؗ�@�q�&g�3��0Veԏ|�)QDNضnv0!3(��`RJ���D��p;G��"ި�z�ʏ�Xe�9�"G�t="�HrM�)1��T��%lt;'&а�
c�Τ]n�(A1�F7p780 �����y�Mnd�z@/dGz0��,^��HO>���&��
?~	��"A1&7`h���ܱQm�c�&�&Xb�7�:�!SU東tl��qF?szP�#�ݳWo�5gF%]j��O �ID��n�b�� �a���Ғ��ևc���" ]&D�T��)W�
[v]@���/
��)�0�
([V����h б��8^J4;q� �d� ���� �����S���O�|!�{�? R��<HV��y�'��J��E�d`d����XS�@9"��,\ #�&'�� ��A	J�.��NZ��u�u�A-6����k��a�A�6_�
�
��O�,���dS�lJ�L�.�8e��d�g��)!�&���
�9�b��-L~qp�R"o�3mN�P���x�$�'d҈��E�z��H�`W���2�dI�^_>Y��U	���Z�+�sz�H�D��,�&L��k��u��Q�Z 7f,|в�%z���i'���D�'�ve�Sہ.�t[`&�X��	�Z��[�·2�sU%Y%

�O^]Q)%�`�3́�zN܀lUe�*�LE���!��8׶$��+H�9���<�q�&eZJ>�qE/�&���:�dK]�:�~Lq�EY�v�~H�R�I�ҹ����fY�p�G$(�>�D�D?�>0���O�>F�:T
M��2�0����,"�C�� B�ى��'��Ј4�\(�}��$j)�ɭ�>5 M+���@��'�Z
nsd�3�i��a)V��� ��?Q���-@(/�BA!�˝�����I�Īs�%&�DY�+C�`�V�?Q0�θ��T+q�A.��'-�ı��܅:�cgL���@"O�MJ�-����ps�lǦK7�aq՝������O�d����y�O�� U
����;-3aPRϋ.[�t��'�n��c�$��좥/�!W�&>�4�Ѳ�A�6���5�j�2e����-j��^i��g+�3�DCTՆ�{�S������1o�:YuM���q� ��R����[�!���Lԧ1
6pSI<	�bDy#Q�S!c((��p�O�L-��@p`4�o&,m4�E����	ő�а�S�:� �S�۠S ��k��ˌ):���7��5@�xX��cDG�A�X�"��M��Eٕb1}RB�-�桳��#yO��X�ȑ�Z.T�����:*�\0������8��6-��>�D� ���t �Q!�3�` �c �(z��P��v�tQ�P�
v5���@�&���V�)�|l�FY�����qݹ��K�^�nCDB�H�A(� )�`�I@(˨&W!�D�FG��
�����E$��X Ҥ#�Mk�NL�uܐ�H@�SN�d��1T���gM� L4���D(?�L2�-!��\0�)����F����	+d:Z�ځnȭV;<��&OU\�4�@D�9TV0��d��0ň�	�P`���āz���hƎ!O� �n��l�6 �a�D�>H)���d�#��c&f(�� �c7��4m]%5|�@��F�,��Y�]7%�r��7���������i{2l'��G�J�N=�-YQ-8jЂu
ժ^3z��DфC���<��&$W��!��*�H7�1qam��kՌUZ
�ze�xPf�� O�n��Q��+�bB�ɀ[O���@	�4`��c�:Yi� �5dJj�tٱc��>�p��ņȂ^D�<� 1f��3M'?���R�1Ov����rTRЁ��I��a���9Ն��2�>/�N�Ywi0Z+	 ��Hd6$��(ҕq�l��"�T�y��悰-�2E1w�&��°,�6A9�O`m;�G�R���R6Z�Lx��ࠒ����ڵ(����QA�-o���OҤu��g^ tI{���[���f �Kj"$�GE6iK��e�>A��J�mѐ8���خ.�n�sH�yRjR��7��ͪ�)��V���P�Rp��H�i�~�Ke��~"�׿�D+�.+4(��]+f������A�,��@�@i�I>8՚��J��g?���8`\4��@#qJ�Di���/���;�%�k�8:�D��7.��\1-@#@��%m���<� "A�8�h�3u,��#����D�! 4�skF�P��	#"/�	�Q��r�O;coH@�=�&���̗�h=Y��"�����8Å�5YN�XJ.��'^,@���f���x)����*D�L�@�kgf�(#�`:��?�D��) �l"�_/͘O"�hn?^�D�hE�R�i�޼ ���<c�:9aG�3UA&	�f=O,��Ӑq}�+��k���<b�2-Qw�N2ֿ����A�H�K�9F�\Lb�-��:�� D�98d�s��E�Wވ\��˚�@�J˧�yRe�/i�9�ԅ�8�J�ɠ�ɍw�`��^H^����h��?q��V�5X��T�ܞ;�L��H<9��
�F<D�L#BxPa�k�Z��U@4!��c7ƴ)ć�g����e�D6Hc�'Jh|9��O�Z�A�fB��8?Ft��$ٓ���C�f�_����s�&.M�'������HT�8K�ߵr-ָ�e!�
1
:���Q�
�����2Yz� ����l*���a��x�z4���O>6m��=6 cu�V�M��B�?P�)�O&+b�����3B���MR΄�g�ԁb�j�h�g@�<b���4�L�x�'m� �RT/��N�Ό�1�O�^��VѫG�F�?)��:�l]X�<� h��l� B� ���t��0J��C��X)�F
   $�!�Ʈ��O��$ׄU�̈́�@���@šؗ}�v� ���I�@�84�Ϗ�M����:����ڊ��ٹ�*�����54�V+
�s8��
�k߬ �i�s,j���Q7��/C���BR�<�5����v;��Z+,!�U���'��l�ao��zN@`.�SӸs6Nۗ�ּ� �E��!)%�>i���h�e;�ʛe��I�RCߙ>��	2��ı^8�k������3��"�N��	�gđ�����9����1_<�+A��	�����C��'#Ȕ�R+���}�䙟�1EV
v�8��&�5�j � �E^z��o":d��7r���!Įz����� GI<[C�O@���o�>E�4
D�A�6�	D�x���S!���{�-ػNR���`D*S�yC��_�Ж��D%JN�R���C��|:�6@�b���Me6� d��.�͛��R�m�6|d	�%�
 ���>1���Im&�``����Io.��B.eCGL�?�ZDk�N��9���qD"P�w�j؃q7p��Y����F'
QKgLF<�H|G�O�Ӓ��&�*p��ܝ�N)㑊ð-Ax�����4A%!u��,��Y�W�E (�'w���bn87����	�9ؔT:��M +�@�[��*�j����%�?�r�O����7)�y���bd���H�e`(�%��ɑ�>�`T��5�4�J�C��t=i��D����a���C"ژyb��,hq����9% fQ���0���⋶'8e�7�6!�l(St��F-�|k@�Sx��IS��3G & I���		I��"- � ��R��6dh�x@	H�@����	,&�q�1f������E6ġ+�$K�D+r!���Zx?��QD#�:sK�[��W#O�������E1ȱs'$J�@!j�$<��AT#�i-pa��J�M(�R3%EJ��DK��P��l�S�W�W���R�|�b��Q��2��9+�
�$P�.�7׌��x�n��D�T*����`�!���&� ����^<^`����IL�~94��5<��OPHr��Q�+���0t'�Zaq��'`���ΏA����z�ѐ*����M0�DRa>m���݄�15�ʶ:I�ɽb/�+s���O��)�
68N��@��T*�%8b-F�Eh4D�LҊ�R���P�%�zla��%\�"��� ���k��I��옥�P'����<���P����(2��"���L�\�]b�(��#���E�j�`y0C	 	ǄA���H�"RPt��o�0ǒ+Z&�R�g^������v&����+p�e��!��h�$[��S*Y"����;h9:�`�DЌ_�*����!��=�Ɠ�6-S�eR��r�A�q�z��O2TT&Q��ƜB�0(Y��F�>5k5eS��|�id���t��I�[�����NҎ�4�� �GE���8pI*��,�,,� ����S�ǌ�9v�!�&!��v�f5
�͑>F{�����ޠl�(ʖ#��Oz�"�<��}����
J)4�x	:5 �P��-X]�h��g�=,�<�{�C�%������0z+(!5��
�P)�k܈��-���b�� JD�����s�d\^�,{�m�"B9*t	��;5I��ɥ�L�Լ!��B�ԅK��^�8C-{�-��� V�T�S��6u4� !t�5$��#�.ԝi�h`��	�^��1OYE�J��6h�=a�쀅��1�@��ԟl�r\�Æ]� �_�$���Ʀ;� )!b�շCњf�:,O�z2�)j��S��Q4F�8Ԁ�	�>!&��IG�Ԧ��)�CȂ�I�r�R�Ȟp\A�'i�9�&�����3���b!ę%�`(20d� ��'J�`�@I��)�Âw]�)"F�(X 菱��B��?C �	��9)>$�X���-"������td�a�K��0�0�B��h����e����*�}�f�N�pl
�!拎+1����5�yG'\�����l��Sz�M�HC�	",�,8��֥GTB�j��z^d:��̓uVta�4s$B�;�'(�0x7�קCSN�!Z>��I�#S�8bf��$�$����!��yrAP�&�(� �-� ���mڜ� 8�q�%�u�e����O�T�d��Z��8;��,OEB�X,R�Թ��
�?L���$�(>F���!P�!v��0���m�!�M�S	����	�+��%H�E@��
�>�!�d��E���m:4~P�V"@~(��A�����,�Tl�CP��OK8��Y�SB�3z�� �����yR °~]�4�F(?+�tt�'���?����3k� �������!��#7��jC�u�!�O' &P�PK�yg����
�#�!���$� 5���
ER�4c�!�ă"r�pSv��x9Fe���[��!�\*-�$ '�#0��@ʝ8!�h)���-.��:��@�-�t �'�P�!0X䬭ke�L$�V�b�'��PB��c��|I�M> u�a��'��}�rf� e�	
��}��	�'4h� !�'Q��k��1r��b�'�V�Xa&Gf9,�pP��2_�`TP�'�8Q�W�Yy ܃2%;I�T���'d&�0�.DiC��! G+L|P�8�'#F�)��ڱ_9ڭ�+!>ʄɱ�'W��jw�X;<O0�@$!Q1��X��'s 	p�ϠD� �,{'�S
�'�Z�1���F�rh�WT v��[
�'ݒTi��7ޮ}�r@��J����	�'t&��ICbe��ӁfNK�tQ��'6��b%���~� �'�EO0)�
�'��y���L���d�8V�A��'y�u�Q�Աc	�9�.Rs7��'l̸Bf/k��q��N��4�r�'E���K'����#˓mζ���'F�8:�!V�~g� ��Ƀ6n�ʔ�y)B�i�Ԩ���K |�����ۘ'�B���"ɰ-�l\�ċ	_�~}�6	I*��r�f�z�*�K�//�a�D���C~݈"�\,=��p�D[E(2��q����'�cl��r�xZwj.�b�+u���ӏ�/ ɐ��"�a��k���������BL�I81��	��'L:���$�&p/DE	���<;`�a������ēywGx��� b�fg5TVU��?=bpI�w�i����"꘧���V)��:�Z�h� �(�X�����!�M@'K��ȟ��9r��|�L�*e�ډ������<�ךxb�o�1b�p�N�"u�:���bM���D��)���F��O����)�'G=T��3n���0A{�cu��	�g��z<�����'��O���f�t�N�#hM��v���+Qj���H7^�L�Af:�j� �-�>.)�����Z!x^`E����2�`ʓk��}�S���9�.�]�z����5���b��!7��'j�I�!6�zY�O��HA�#�6o�$�j�'֠\@���' ���>��O�>� ��ìU^�`����)���EleӜ扝L�~=J�"���$�.a��b�{0��yr̅ȟH�`�)�؅@0��XV���?����FX�R��J?��-M�bYB��	W�b��$�ɄY��Y��3�p�"��O$Ȫ7�(�"���O^eQb��)�z, Vۼ T�1���O�I�CA0�yB���}���<Jɲ���$�%�.�DFZ��Bɫ�K�<Y�O��iq�`R��$h[!t�v��)6��hr]��7m� Z �gkt����uq�(�$0�=`O܋~ٸ���G�p�2.��aK/�����DߢZ[j���N6��x��MM�)���֮n���hc*�7pia����*��@j��,��)��n��A�AՀQ~"1q��>�'{p��j����%o�
q����ȓj
�<��X���X��B �vp��\��������K�8���(� x�������]�w�L�!Ђ�0�"@��H�N�H���P^��얚aSЬ��l,2@i�fÜk��M ���mRZԄȓ��9�!ٚv����E	�e1�ȓ)��T'�ٗ ��#�V5W�4��wI��S���p��ĊIc��ȓ4�2U�,#r`����8M�&1��Z ��	�i�g����T�1>�V�ȓv��yj���<�R�do�>y�I�ȓ��1W���_(�S��چrҊx��}�i�س3yd#��M4Ɇ�Z^�:��H�" {Sƻ}v��������f�1�"ΒBa͆�i����-�<'����Ug੆�H�2@գ�j��N�\�~�ȓ;X8;ᨘ���2(E�B����ȓ"c&�Ñ��)Yh�%)qm=c�Ȝ�ȓO��Q�
V�33�,��w�7D�X��G�W_�QQQE��q���I7c2D�0�u䈎s��8�Oɀ\�-q 1D�t��ƽ��9E≤ Ȝ�!ק-D��Z��'qv����F4|��u+2 ,D�8��)#��L���?&��W�%D�|���ĊY�}[��^�~b��M6D��Qv+�\��YJ!fY�j6���� D�(ƥ˙M��A�ѺbF�fI>D�R��/���CG�܃5*�{P�8D�ີ�[����A�.��;e)+D�P�$�lӰ��O1����+.D������6�d)�`M���S�F+D��㪈�>5,���'�	z9`�6D��q7�4 �a�W�I-	8J1�"&6D�؀g@�5l��,�;Y�����3D���C$�SR|�ɴO�mS܈Z�1D�dj`��6����l���S�1D����ˉ&1ߘ���EO)���[�0D�����*n�8�@��E�(Ay6�-D�\	�)Z(J���zqI6N����g/D��p��J0u �q��`@�V�����2D������M)b�A�f��A�ͱ`=D�� �k��Qzv�		�~��f+9D�8p���8��hSnʒcY&%�1-D�� z�����)�3�揆8�|�Д"O�X���S#V��ɥ'I�Ia�iu"Ol��`C1g�l��� GF��e"OL\��ި"����)�`+*9�c"OnXA�)��=����aȒ4g3�"O2��A��"�'��Ll�"O���V�A�O'��ELXAAE"O*�C�\<t��=��ϛv�M�1"O$A`R`o�e�0�ht��"OB�ⴃ�\*�AA �֔q#"O�m�fO�,��� �M-t���!�"O�1��C�"h�P����	�]��Z�"O��an�^��x1N�*&�U�"O�@QF܃>��щ`��+�h���"OdT�䑱"��q�e�i�"O���a"+10��ц��5p�Iۓ"O�U��.0��i%)��1`�"O � $l�&y�5q���;mXt�6"Od�:ǌŠwGDH�튠GQN��"O|!S��g��!p���  U�q�v"O�\��i��"EzD�űgg���!"ON����W�Jc8�_�++<�I�"O2�Ps#�}��� JΊZ"�
�"O���fo�?,����fY�g��Da�"OT�yE	;o�ڵ���V���i�"O�B�H.i84Ԉ���B��eJ�F$D�0�s.�:1,�!aw�:�tq7�4D����U3���;�*�R�&Q;�	6D��	t]J龱*�ʐ�vj�T:1�/D�����I�"��CZ��s$
.D����A�3@$��R�\=J7Vd���9D�Lj҅ �7�"|��$��tԣ'$#D���A̦,�*1Hi��g����,=D�Hʒ�շ!�T�{��φ+P�Y{e�&D��-D���Z����B�Q �&D����BU��έ�G�ưJo:5A1b2D��0���Y����A�Q�vpE#5D�Xa�E�4^l|��-Q�UM ���	3D�P3�MM�MH�ɶ;7��yK� 2D�X���& AJ��'
Nj���BR*O �Gl� c���f��8��<�"O.���#���-^��(E� n!D��r�IX��h����]h��A7/;D�#���:s),�"�]b?4��Eb$D�P���Ѧx�b3Tg�h8���#D�p�e�Y�v��e�L-/��E>D����'W��D�祉:�z� si D����Y#�HaS��>bjL\���<D�|���b�h���#��]�4l��=D�Ty��D�3�@��b� z��X0�:D��%�j�*uf^&`g����h:D� �T��[^��#s��M@��"D�4`�$1_�f0� k�<��%"D������;<xdY�Wcˋc�d-�u�!D��:����D��k�3HE���<D��)�㍥pk`i�n��hW"E�B:D�\Q���f�L���;F9�1ѱ:D��r�Q+0(ޙ�c�R9MJ���8D�L�d"ӝa��#�B,�c ,D���E��(6�"�� �
6�X���k6D�`�����y0������"c �P�C5D�$��/�}���#���tg}Q�3D�`�ƌ�hDީt�/f���Th.D�LH�L ��8u���Ǖ;����s�?D�� t8:�S`x�rQlU4e&,�sa"OD1�Q�9� Kl#��"O6�#q�ݿ�Mز��F�i""O6�zR%\Xy ��բˋS<��'"O�lZ�� I�U#��8��xf"O<��'�Q�-à-�e���/�|�0"O0���K>�MP O� cc�M*U"O���FOؚ��Y��NЂ~4ޤ�R"OɊFC�(���'.�:E�|�A�"O>� �Ȅ�'�6��ϵ.��iG"O�۠�VW	�Q����\)#�/D�p�!O�]Ns� :Φ�sի.D�p��C��pU�ĊMn$zrB+D��)�ix�I�HD��T���--D��zU�G�Nb.���!�"
\��G*D���o�	k��g,�r��w*D�IE�٭�R�;�F_b���;AJ&D��`%��i�6!���+)VY#s�%D��z��ʃY4�$�qi� ��� D���UeY�4Ī�)lS�<�`:D�q�O.��h{�D�?+�����7D��4"�"��H�f�
=�\��;D�4��+�����KS�2�����3D��ڲ�F�|<�,��L���I�'F1D��3���1;�H���b��u[��.D�c`���rˊ�Cy�a��-D����LC'`˲��ӂ4iz�z��8D�ؑS�]�O��be�O).k�Q�r,D�@���û6�A����4@%&ɸ��>D��$��F3r���b�a �Kw
<D�X�� �1 (�5���=@���� &D��2#�B�s3X��"�2�x@A�"D��2���;yZ!��*�o��t��i?D���υ}n|A5�jc���a?D����=~(y ���喀e� D��	���M��P��.�!$�=D�|�vl���� ����A��=D�����Ed����-S�����<D�4����(/���ak�;y��$�p�;D���e��l�<(��S�a(���Ǯ:D�l��ɛ�-x\�20���|�[W�+D� (w��B��A���	E��mCB%(D���e23G����,7P�ե$D�`ۀ�1��F+�{����-D�$*PJ"yI�DQ�Ä�ܼ�4O,D��5i�l8x)��.[�5B**D����5A���G^.�}AR�&D�x�7�H�\�p���P�?̸�h�d#D��*�`���ڄ:�.Mo�`����!D�4+�a��`J2�S���
�$i���=D�s([.sa��vfߝxE(ɳ�<D����˒�G��a���B�E�5�'(D�4�f��0��B���?[�9�u�0D�ȐD�P8���rd�9(48[�a-D����l(J��ƴ/�j��j)D�*sB3`pQ���]�j�Ti'D��"�TT�:	�U��6؆�G�9D������Qz"�	E�X�	H�c��,D�x����4𑲑f(w�Ԣ��+D�d��JF���)�À�Q~����&D�L�5�8f7(M��N���Nl	�G$D����K�����x�ʏs�hq9�+"D��C���)7�1�CD���N�zVk?D�4��ĩn�b�˘]����d�"D�� D�����AസVM��|�X��"O�1�H@�A��D��L���1��"O���ÌI>4�����5�"O�q�w�<xJ��b܁�l�"OՈ���jW�����I�u���"O`4���4�,��ҩّ��a�d"O��+�a��
�pq����$�f�"O���e��A�*l�ԍ�`]z���"O-�eF��z&���c�7h�0%��"O�����=n�@�'�з��H(�"O8�*�ŀ�`�����#;;`��p"O.��*J:�}���K�z� }0�"OT��� ��b��sA�ТsbJ�;4"O�����4I!��������"O��ش�ƪ.@�2�F
j�8B�"O���T@	Pꬪ�D$H�H��"O�m�"��!�C��pO��j`"O�� Gf�T�h�L	
G�	�"O�hP!�[�s���0�`�"O6� �Z1�t�FG_�N��|Q"O��Y-�+|~����=��h�"O�isD��(Y�=�vo��N�Z� �"OF՚g�q�PQ2�MX� t���"O&@8g�4��(�`웝WD�T��"OF}i�   ��     �  f  $   X+  h7  �B  �M  V  #b  �l  �r  Yy  �  �  ,�  p�  ��  �  4�  w�  ��  ��  ?�  ��  ��  �  ��  ��  2�  $�  � 
 \ �% �/ N6 �< �B XD  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r��R�( �gVlɦ�M,H�IT<�7�)D]���%��IM~���Bb؞p�4)9�$�\���`�	X�����|o!���7��3���n)R�,�.W^!��b����]�:;p�櫔�'�!���a� ����Y�4!BP���-6@!��L1KF�1Q����Z�9�%�-'!��3��4��ɞ�Z�,��&���1j�͆���0&@њn�8��ߏ	>��ȓt��  �C�m|h��po\�-@i��5�� �d�b�%��.�_�`�ȓzN܌��E��Z�E�ic����5>��J��ۮ3\r](pE9)���
$ �z�f�0'��J��̳vO���ȓV��8�l���%g"��y�R�8D�������>vxx��лX
�-`8D��2�A^�b"}3.�S}�e���1�O�.�?K�~`Z	� PVd:q��6~���2<Ox=� ��[���xD�0Fq���a�|r󤃾�Ms��t�l^���B�Kyl�`�ɋ�1�����S��\������Rx����m^��O�~�] /dD5KE�B;efL����<�a�нl�X��4�F�pl �Zg
d�<���V
o�N|�qc��n�@��Wc�<1Gd�%8�1iܨ:��`��S�<aw$�q�*���&�D{cMi�<� �U˶`�E[�\�I՝�m��"OR��'M��j�HI=A����"O��#�T f���%��4$*A"O
�G	OV�T�h�"�dŸ��ĕ,�(O�q�p��v�;+3����#���ʸ���:���*��f=�q�@��`,�2�;�S��y������r��Q|P��T����3�S�O�y�3���]����%k�u�@2�'���7�O�M"0m�9t��׼$���Ɵx�J��0<��'t�J����ޝ!�&;F�l��'�ŲƅP�i�TY�#f�u"	
�G8�_g1OB˧FIz �&g�8z�T���H�-���c�'�^�YR���	'
�(�#��=��O
�=E�D��hج�R⤚����Z��Q��y� �H�v` 5E1$$ �o��y��)n+`�R"H��S�Z�N$�p?��O �Ũ�uR��Ca�YT�`sO�1�%F�tm��+ *ZJ|��AZ�<�4��5��卅�Ej���r+RX���?���J�]9�x8�J����]�(�S�<�q�A����/ƀ�|a�v��f�I�S{�d*�)�S(?2m�g�
c	�=P���OgF7�/�S��M�J\:6�뢊��MdZ��k@�'�ay͎1d:�9H�@ T$~ )�oF�y"���
]y�@\�X������d&�O�p�s���1�0��*J�&���p�'��'
H�C
�Np�C��q��Q��'�ȵ;���>��do��8�L	�'UP��5�E�%�BFz��)$���U���s��<s͓���pc�<D���+V2%y��b�ݣtf��i:D����G� Ć����7��1���$�ר��9	�F�@<�az���?*z����"O4H�$�-P��r3���fW(d
2_��E{��iӷ^�V�	����p���b�;���9O�̲@�߲ �l�ض�K�8IP��>��m�����,J�.ݻ�a��~�����V����&�!
��@���P'�y��`>�0Ɔ��g�T�5� �cDDx2�)�Qˌ;Tx~Uv��7y��%*��r�<i�#��O��)��1$�|��C��HO��}��@� (�(*H(녩�0� ��	|}r��`Ĵ�ׂ�p+px!d˴�y�jяU��32�H�i�X�` o�y2(�x�캵���*AgY#�yBOʨ��i�0k1���ԃ��yrAQ%e�h��I��i�����ybğ�mNRB�!RЦ�
Z���:�S�O�pH��K\�Hn�tJ�;*z��ȓn�iZ剌5UN�TM*s��e��_�>`�2��� �)2l�%f��ЇȓJ�*E�/�c��L��,�K��X��K��9��2b�0xx�k��GJ���uڒ�X� $�d��Я�DŞQ��X���5�o�&p��ю8�)�ȓC�>��Ч���m"d���j����JP����a�
�	.؅j�@��{���t' +�<A%N�a��Ň�rDP@��k��3���`���?���ȓb�VⰈ�C��p�B����h��S��M�2�]6>j`�d$�f^��ȓJ��Aô �w�NaH��Q^ꈡ��s�$9���<H5I��_�T���}1�=;��Fo�&����.�����?� ��*bm�3�F�Hec�=3ĭ�"OJ$BDe�/%��up��^�A?�U�p"OT��ʅ
$<E�d�عHTMb�"OY��EH<;�Б�g�ČJ?����"O�82�dШdŔ�8�a		�
XR��IE���IM��(����-t��c�\�\B1O�=�|
�-�m! �KW�O<�x:��	A�<d�^K�Ԑ*��ْZ:�Y���{�	�?A�}�����QB�
����2J�$��*l�!�$�%}���f"[�x:H�u��#j͊⟼�)�g~�E_�&e*�{�?D�<�0���x�&��3�2I3��m�i�d�P�!�� �l�@$�据~o)餢P�;�a|��>ѳ΁P�Z8b"�Q��lzСDB�!�DO>�����Ɨ��NL��� (����?�S���	�aUVA���?Ϫx��L1Z�C䉱(Fvy����'%�nl���'қ��'B��r�LY� ��k��P&��
��q��I��M�.Oe��f55W EJ��H���y+�I_���� �T8�pCs���k�2z���ē��
8�Ġ̄!��<� F����U�r����	���ZХ�=ܴ,h&�\�{�.����<#��/����cE�t���K���u�<��+A�8,���/3�$��0�Y�'Y�?�1��� j٠��ҍ��d���(D�8c��!B�
��`���t�;�N'�.�SܧrF0��M��n K5vLFyb�i��?�!'�  b����
�@�j�N�`��B�	�I0P$)��/2}��`��(2��d,�	0e�݈�c�$+"89���6�&C�	�JA[͓V�$�x���D�FC䉏6A���l$R�� ���+vU�C�0P4>+�'�>�#��@�xC�I�B�ZX���Ǟ/�$=��� ��C䉷UV65;��9J�A���B>Jx�C䉃mc$]��#{t	�T  �&�B�	�6���mK�=#N�hDd��>�hC��'rLa��\���d��̢B� o3�FJ�O#�Y%���+'�B�I�]\��R9�U%��3C�ɺQ;0D� �/9̬�)���C�	)3��-kqnѭX;�5�K��"QnC�ɡ=z�ʑ�O�1�����\�\�C��>g�򹈑#�t�"�M�1yפB�	�N�+�@!sc~�k`n"�B�	,3
D�J3�Ș8أ��
�8B�	D�̕ڀ��e��FȔ:>5�C�?@wʴ��J�{2ƹrЧ�M��B��
���
k��D��}� A�A�DC�	�&��(��&Jz�8�aJ8n�C�I�o�0@��}\�i*�'I X�HC䉞X��E㶠�M�����G�9$C�I�>��h�� ���&c��j�>B�	7:L���T�����A�'{NB��D�LL�"ϒ:�񉗧>r�B�ɬ��u(�E�,;�p��.��B䉜�����>A��P3D'U^`B�	�js�)�U�_���1q&G0,B�	(2�62�)W�M��ђs�
���C�/8r|rg�\3���&c��D\�C�	fZ��C8r����2֞C�4K�ޙb�I�a�D c�(,C�I��I�6Jq��1 E�2)�dB�I)9�,E��KK�$�|�aN�7HB�)� �I�W�ـOa$yҠ�V�?E�)ZW"O�L����2: x�� �;�T	3v"O��R��80FW�v��2F"O��*��Z�&SX��毄dq��*S"O( 3�M��[Nb5J4A�5~�5���'�rT�@�	埨��̟�����|�	*��`�5�7#rE8��f톹��ԟ|�	Ɵ����@�Iӟ��ڟl�Ir,2�z��1|�༨c��^����	����Iҟ���������	џ���(Z���VE� 5�:�,�}f�������I��`�	���Ɵ��Iӟ �	8+���I�.Eż x�F_P�1�	����I̟�I������Iӟ��03Ǫy��N�c���H�e�'��}������	ϟ���ş ������	��`��/ 6X3��Í.ڲ��㛎^fI����(�����I̟0�Iʟ��	˟���8}Vb��`I�5�Hm��BY%O1���ݟ�	� �I̟L����	ʟp�	-���v��	5��Q�g&E�B�d ���� ���p�	˟H�I�H��ǟ$��<
�����~Z(��¢:O$N|�Iݟl�	ꟴ�	֟��	ğ�����T�ɞ�>��P�d 36�)�P��㟴�������ğ(��ɟ��	�x�I�D]N�C��_�n��At�̒M@����@���8�i>������IП0�	����@�f�6%�
�#R
s����Iџ��	����	ߟ �Iٟ�ش�?���C;N�8���f��a�O�>�؉��S���I~y���_�d�ܴ3v>��VĂ�~`�q��[#6o.9�q�]Z~b�o����&�V}r�n�ԡ��*V@7��q�2v(��@Eꦑ�I MU��I�N-?q�^Ȉ��7���
�$ɰ)\��X�#IX��'�2Y�XD���Q�z��gU�|�����*Cx|7��E1O\�?-����St�G+'킅��&�|v�āu�I:%���}�L�	]}��T"_�:l9�'o���X�6�z�y�j*Ȃ�Þ'���S��k�j����i>���OxA;@* Ԕ!���	�4^r�Ity��|2�f�� (����b�0�e��QL�X��� y�2㟀a�O5lڈ�M+�'.���,
^�p!�͛e�dq�~B,�"˴�%CY�&�|B�Z�����GQ�y��K\9#�>�:s,Or��?E��'�P�Y��|� �����v�B�'�6�Ě8��#�M��O)�0��֖F*P@��,����'�l7M]ʦ��I B{X�Z��6?�FP*_j4y���(D�s��}�N$	FNb����'������II	U�,��V��uf�A� *�%P��D��Lv�� ;��/b�
%�)[��U�P%�#h&Q��&��z$�Hӆ	T�A*��B�VxJ�ˆ �?w�(5��'�7@v�D%�0x��,k�!F[�(h����)j�&ő��ͳCv� ���2��B�-s��[��BH�d��r��#~�v%Q��=�H��"��%'�^��U-ǰ[	��&��qiX�V�Z|+p��5#՘�J���3��u��/ºs@�S��6�d)�4�'h\#�֣
�,�����ui&`���2��0n�џ��ş�Ӥ����2N���;6�����uI���'��n��y!�~�����O?�
�-��X{�ԪE��x ^��	c�Z�k��O����O>�$���ʓ��	Q�s ������
{(�;r�\-8�qm��S�l,;��0�)�'�?�6�ښv� �	���ՀSb���%��'$�'6����'�R>���B?A��ڜ	.�g�6H�	ʹ�1O�R��F��<���P��o3>b��Vh��k�	p�������'�������O��O��ak��h�����J�iZ� �}�G�ez�f=?����?9���?���G�|�F�؍w͒Xq+ל��-
$�N+�?q���?A��?N>I���?��3-9 N*t������Vw��K��m~��'�B�'&��'�Z�I��'��=`�S>�`=�H��F/�D@�jq�H��?�I>����?YP"L�)t�Mn� �D�� �,$���p�*�0"2듫?q��?���?!�ϑ�?y��?�'b4z/J)�3&&��L���(t�V�'j�'QB�'6*%�5K$�ē.���ZǪ�1��r��U�m��\�	yyR��g%t��$�kLҁ:��4��[|̞-j�c�"*�FW���	���{� �'�nZ&�����JQ�B��AfA	q	"6m�<�R��1h��"�~j���!�����m�E3���4���t�i�E�bӼ�D�O�����<�'�?��g�	+^Z���c�.�B�p��Ӻn�Ҥֈ]�6�O~���O��)�P�i>�h1B�> F�yUE�I�,m1��M� �M��D�O���1ON�$�@(��1"z��qK��b:�nϟ���ߟرE��9���|���?����@���EO�v��"��t����,��=�`b���Iʟ`�ɇB���2��&��9aY#l]ZA��4�?�Pm�8So�����'��X���M�'}IR\!�*�x�X�C�]+�M��b	��<���?Q����D��j�!*ٗ?p��Ho��PqA�͹n��'���'��W�p��۟S '�F=z�3"�K.���e�	p��b�4��۟x�	xy"%Ź=���S�ȥ��Y�<uKP�E�X�>��R\���	ҟ��	Wyr�'IB�Q���ФN�`]zA(��x=E�V�1������	柈�'Y8 ��M=�)S:$2.����a@u�'!U'^0�m����Ihy��'�r)?��O�X���
�5yf�!��&[FUYH��l���D�O�ʓ	���
2��d�''�\c}�� 
%88��.�2�F�8�4����O����[�>��s�� Fq�e���rpSI�nK�e���i��I����Aڴ(���͟����DL:K�(�Ȃ�-B|����兰p��v�'XR�C��)2�g�	�G|9����
t������%:P7��g�N]o���8��ǟ������|j�K[*'���Ё�D�l�Lxpf�(Zěh�8;�����	�?c�|�	HI"xQ���J����UA���/��Q�Iß�����.]i�i>i����TPR�<K���C�]m,�*1 �=��D�O�=���?���x:��gg��*d��4�޴6?$�j5�i�����M<�'�?����d�)��QVb]V�x�'����n�c�'�R�'��X��'!�� 'ح����<"/|=�$���P�l�H<q��?�K>y*O�n��5G|0B*�1��M��Hס. �Ov���OJ�d�<)Ga�Z��I�9t�u�+!�L�5�^�AZ���\����'�b�IX� $�����:J�,�#�fġ(K��ğ����@�'LL�"��=�I	(|.a"���'�X��э`��l���|�	`y�'�Q?�3�Cܑj9�d��F%f�Y��g�����O�ʓc�l������'��\c*RecQI�"<����
���4����Ov�d/"�1�r����� �8dU���!LY�i�y�*C���d�O\l{�f�O~�d�<��'��p�#LT<�梁�*�1uQ�d��U{���G1�)���-�<��%E�?��Q�Ȟ)	�,6m
:���$�O
���O����<�'�?q�E	-��fJ5n�6{r�@v��vh�&e�&�R�y��)�O�������	:7 �d����6�䦹������I� �=�����'���O�=�d �5t���@�A�� N�4'L�z�Bp���T�'���OLe{&��
���c�=�� �i����2vj��8�I���=q���"�;���ym6т��X@}���
0��O���O�˓�?a�IX<jb@�Plɠ�aY�?)�0�+.Ot�d�Of��:��̟�
��<�b�ƁQŨAɆ��d�|$&/,?���?	/O���;9I���$|'���I��e�65aW$�Ev\7��O ���O�����WD%���`Ӓi�⛉8S"�����*��Z�x��ן��',R�׵8�Ɵ�XA��%��
q�*$�`���[��M���'���T3.Un�yN<	���a괜�p��3l�l�(w*F�Q�	\yr�'.���\>�'�����v��$ϙH[�x[�ŅO�*c�p�I(z{��!v,�~� �?;T��g��\g�� ��Bd}��'���A��'<B�'���O�i݁p��R�ű�89qHPϰ>��� �p��]e�S�Mk�IµnDk8U� ɹ&��m>~ȁ�	� ��ޟ��S\y�O|RL5��TԪ���8p��ڌl��6m����(����S�G�%	t(A��	L�Hzq�S��M����?!�#��Db*O���ON���������Y�hk��X�̹IUL��'������:���O��D����KL�Y�L�	uDu8E�x����/X��˓�?����?I�{��Ed�Fa���[t�L���vI�'�y��"����O���<����(\z�(3"��� c������&����O���O��t�	%r6:,��F��!����PS�����P^���?1���$�O�]JD�?!q�c��ek�8\�F��!/�,a���'���'(�O���բS�z\��iy� �O�m_���l>~�a�O����O�˓�?!W#�����O�(�M�A-�����2.�<�U�H�5�	E��?1���e5F�'�0��!+x�C��>A$,ҳ�c�x�$�<��$*��X+�:�D�OJ�I���6+�3�&	�:Z���>��2�N����S�S���ş%0�$��-_. �}�#��1���O6�9b�O����O�������Ӻ#CD]�P�jJ3�ҋ �F�hD�_h}B�'���%��Ř��O�*��W� �Z��� F	
%��i�4$��%��?i��?!�'��4����Ƚ8�.�XR:8d��X�{ ��m�e!nݹ�H<�)�'�?aB�=xǪ��A�C�Zq�L��l��b����'5��'�LjB]��ퟨ�	q?!e"A�6 ��.Bj^�P�
�-�1O�)ؔ��f����II?���_��pA �u���CoY榽��6d�E�'�b�'������<
�gN�`I~:f.��f}�I�J����/?���?(O��$��r�I��1v�+��,q�,�uHD���d�OZ���O�P�I�%�=@�J3e ��5����fo�[����?)����OXu�Ǽ?��0��}*�i��!��W9�<1Ht���$�O��$%�	ߟ0�3c��.O�7Vb�e���1OF�ա�@n�I��X�	RyR�'j�@�Y>%�fZ��l �2\�#�ܐb��mZϟL�?��Vb8���Q≏��ٰ!���J'�|�@�ţ��6m�O�ʓ�?I��	����O����%S��� �^���$h{���"K��?A%�C|�<�O{n��bWL��ٰ�!.*��?�V�]��?����?i���+O��Z.7��5�A3m�j��DiO6���$��B��5�lc�b?�Qbg��ҬQ	�k�;%�ܣPs��5��c�O���O��$�$��|��,�������ad���S�u�$Z�i�@,���\�ݘ���OAb�'G�C=� �}d�7�D1�$��u�Խv�i�rQ��B�ty�O�b�'��$�`Ybq22�]G�JS (\�<p�<���Ҫ#o�O���'�䄦Q3$$6�5�e��	E����w'�d�'���'{��U�P`�RC`$�Q�۪p���"qv���>?q���?,O���B$�l`e��x؂�K�'�� *�!v*�<A��?�����'���8F����f�^_�X��%�"&��8� �����O���<��w���O���.r�������}����ڴ�?���?����'�,<sr��;�MkD&4cV*�dw�u�gOI}��'�X���IkQRĔO3B�T�(V�̙(66�է�6=|7��Oj��͓=��$#Gl)�d�:T�������s�	��L���'��I� �׋\j���'�B�O�^�����<��� �٫����k ���Z�	ۄ{-c��'^�I3��غ)����M�4�N��'�2��8h��'�"�'��DP�֝�6��q#b�N�NRY�c��`J���?�5��|�P��<�~*��Y�D��10��h:����&Kͦ��4�P���I՟D�	�?������'�R!���B�i6�ei�k5M�N%��lh�>���*�	S�1O>����	 qA�£��ِ�5QE�4Y�4�?1��?�E����4�n�d�O���,F�ă�J�.�􋃾i0	�y�E�b���l�D�OJ�ɨ+�0���?��I�0��;kOt6M�O���1��<1���?����''���f�C��dⱆ�O]��Op`b���0J������Oy�')n�	� E�$ `� �Z{ �����(w�	T�I�� �?a�}��h¾�'�܁JÜ� �E H�X�5A�C~��'��^��Ѧ��B�Qd��kªn��d�0���2�jY1`AQ�i�	џ��Ii���?��(J�:z@mZ�HP�*�K�>i$������h[ ��?���?����?y��D7}���'R���?�%�0|8N����H�9-��׹i ��'u�X��ɉ+���c��i{:%�1!Q�3�p��A"[7ba���'b�';����9:�6M�O��d�O:�I�K�, ��h����H�6�j�.�d�<���}^���'�?�)O�i

�k�,ϳ�NT�q� ���۴�?q�<D� �4�iR�'���On���'ڵ9qMC�����D:ɰ���Ĩ>Y�&��HA��?�.O�	9�t���(���%N�R�P<+!Ɍ��Mv�(��6�'��'���Ob�'{Rf��^���+�Bb�8���-v6P8^1|�D�O���|�M~��� ��R&���"�����8"D�i��i���'v�?=�07m�Ov���OB���O�N	X*�!˼a���̆(0��[���� Ӑ,���)B�'�?���X��(�G
?*^�1��Q<JU�� �iM��˜7�T7��O����O��đj���OV�����E&
���i L&�qr�_��JJr�x�'���'���'�r�W;]O����ϪP!*5����B�ըu�{�`���O ���ONu�O+�ݟ��JF	��K��X;�tc�`�Of��I��0�Ɇ)����ϟ��O�L���s��0�7�
<v���	�-�d<ɱ�����쟰��ȟ���Oy��'o���O:T�qEd����;�h�
|�*�S�nӌ���Oz�$�O~���O����֦��͟<Y�d��@KX0ɢ˄�&*:x����M���?9������Ov��2�N�'����� 3	 ���!4O���4�?����?)��E�51 �i��'���O���Lv�����Oʶ0�XI�o�>���<	�� ��ͧ�?�/O�i1J�
��ǃ~y�Y"�I��� ش�?q��y��ir�'��O�$�'A©�u��8C���ç��yB�[��>��[,p���?)+O��#�D�5eB�����с���z#�:�MC�KS�g��'�2�'��t�O0��'��N�,Y�ԙ�M��4LB#% t��7��x(���6�4�����D� #��=*��I�uH�gܩM���nZ��4�	��\�v�&�M����?���?Q�ӺK����0x;�!��s	���B�ަI��FyD�#�yʟ����O���r��i��ܑ@���$%�C��m���@�����M���?����?a�R?���J$� �g��A��QD F���'	���'���'b��'��^>=�edZ(1�� Z"���;�Z�1�m�)^��e	۴�?A��?1��$a��myr�'(���Α�;ijD �A$W����􁛫�y��'��'8��'m�S��.��޴p��9��_#;��a���=[_���s�iD��'Mb�'~�[�0�I_���/pѸ,G ���f��a�&+��0+�4�?y��?���f���-Yx�ܴ�?)��!���!-w8<�h�f<�9���iB��'�2S��I?!|�S̟@�f�B����˄�����Rr��mZ�����X��=|%�4�?y��?��X!��r�E�<!�a둱)*�sQ�iXBW�H�ɈQݾ�ܟȔ���4[Ls6��-z�P�RE���lep m���\�I!lv6 �۴�?Y���?��'�"��>���1�Y�yiQU�q���S�����Cg����씧�4�~:��-B���B�"=�e�e!YǦ%	Ʈ�(�M����?	�������?i��?�F�ɃuMT`��Ă�b��PZ�nD
:�&�W��'I�i>U$?5�	�&?ܡ*fB]�/�T��L6 ��h���lZß��	�Ԉش�?����?i��?��*LD�k1�M7�<��� \�
Pl�Jyf��P�
��������H���OF���Mw��csm�;"(A$��æ���D���h�4�?����?�����Sa?��
�iKB%Ak�~��BVeg}2cX���$�Or���O����O����Y�? .=b�@ʺ��Ÿa�G�?�D[�f	 z���'�b�'*Bn�~�)OV����ȠI��f;��!��O��n��<Od���O6��O��d�|���޲/śV��\�8��� Q�8���D�r7-�O��$�O^�$�O���?P�M�|��F� ��8ˤTs��rH��.��6�'�2�'a��'B��-6��O��DI*�R�I���2]��3c�ß��Mlҟx�	џ��'I�↊���>�e�]�¼�Z&���A˦���ן��ğ\��&_�M��?�����a�,?6.P��'�3v�H�ĥI�x(���'��	�D���v>	��By��MF�_�3���1�dЕm��9QѦ������q@]��M;��?���j�'�?Ѓ��\�S�C�#�>M����74���� +ϐݟ��ILy�Ov�(T
�)H\�[�Y��#7jjxm�YqPߴ�?	���?��'�����?���^ze�`B@O�P�B���Q��@�V�iJ����'U"Z��S`���$H��
�@��Ac�P�Ay2�c3���M���?)��
�l㥶i���'�B�'�Zw�"��E�����M�C*5�bA�ڴ�?�)O�X�:O��şp���������Mr6MG�97������M���o��C�x��'���|Zcθ%(2�ړ1R*�I�h<f�vA��O`d`�/�O�˓�?����r�: )�n��1���.Lǒ=x��ؑ^�'���'��Iϟp��۟�&�ޟ"��!6����	M��Z�	Qy��'y��'E��Rp&��|BW�7R�>`�'I�F��m}��'(��|��')ҮD=�y"��h�8A� �b�(�`>(��?9���?�)O��x���Lⓛ3��+0�>;Ӓi;"	Q)�"5��4�?AO>a���?9�j��<M�@�tM�+}���a�:�&@��H�(�d�O<�3	U������'��t�C�:�#�E�0��9Pg�'R�O���O���4:O��O0�Ӻz'�q!����H�ځS�@���6ͤ<Q�hG�}�F(�~��� ��t��h�o�f�93��w���SRk��$�O�)����O��S�O�*R$O�%mǤLc���$�*D(ڴ'�RtZ��i���'2�O��O �D�"V�l��j*��b�F�q
�ymV�©��q�)§�?�#�7y�ʤ3�m�v��eT A���'G��'�h��K(��O����ș��}U��� ���b�h��O��ZF$P��d�	�8����?D�S*Ȁvʬ��e��,�M���8��x��'m��|Zc�p��aʋ=�2�zA��[c(��OV �5I�Opʓ�?���?�)Ot�pE��o� �P�Ӄ.x jF��aX4%%���	ӟ(&���Iӟ�!%���֠k(�t��(�l���zy��'8��'��	*n��۞O��x��O���V�+=S
I�O����Ox�O����OfHZ�O:��uj�=B� Q�b�Z�OQ�S�Vx}b�'�R�'��	y�R�0M|�f��&r0���re�~�R����|̛V�	iy��'��ߟ<�K��Y!"gD���
��c�i���'�B�'vT���'E�[� �S�g}�� r`N�8Ƅ���.	�|�n��L<������/|���]�M
BH��dͶKxF}Rb�� 3:7m�<Y'�I	C𛦢�~r����3���p�?dMV�cG�|�����5�N@���3�� f�k�+�]�$�⇏D���>p�"�'���'�$�'�2\>��0��P$�q���~�di�Gդ���RQ�b>M�	Z��u�#y�q�M8�~��޴�?y���?a��,(҉']��'@��_4$�Pi(��.�4d 7A��±O�q���O����O���*�Cع��&z��-�榩�	�3��p�J<A���?aJ>��7h`��KGm�E�y�r��'��9�yB�'LB�'��	�(G��2�F[?yY<�����7]è`0Љ^����?������?���"%� dY"K̔�s�S�-�9�"m�N̓�?i��?�,ON���V�|z����t� \ke %=���:׉t}"�'b��|2�'c�D{y��dZ�y�G@4Yn���e�����O����O:���Ot�y�C�O
��O�$St��g��%���=7+�}��t�	�x�'�xE�H<�ϗ[��YY�"�	Z,�Aq�/��q������'B�4�g%"��O�ɕW6�l� ,ɣS	xɹ�J��n��oV���aD���L$������
W�LQ�e״s� 6��O���#LE����O@�D�O�I�OZ���r����s9��(4n� Q�0�r�iTb^�$suh.�S��Wn��S (Ŀ8����bD���7MZ3��l���	�8�����?yA̓�:Mi���X����0,dٛ��y����$J�B9��B!Ͼ�c'Xd�,�m�ʟ��	��pA"�;���?���~��ݵ*��k����cXfm�����'�Ԑ�yb�')��'֪���͂'q��3w��P�z ��mӾ��~m$�t�I���&���\�b��B�;"n��&�����<�6�<Q��?Y�����
.G{���m�'mn
�3EX�i��=�B'�o�	���IH�I����f�4 ��U�k�D�PfE��J���-�IПd�	ʟ`�'�<4QQ-l>���\<s0���`/qB$tp�#�>����?�J>���?�ʝX}aG�._�ՙ�>`��2�"�0����O����O�˓D:�(�P����+� � �#.+Y�����A�S2:��@�i"�|2�'"HW+��'�R}�i+{l�B��p=��4�?Y����dF�(�n�&>����?=�5��4f�qbf���*-@�Ó�ē�?Q�x�8�Dx�����+����U�$���jR�i��� f�>��޴2��ß|�����^@�-�I�9��e�q*�?��'AR�ڤ�O��T� 5�݌`�Q�T�U�:��U�3�i���Qll�j���O����z�%���I�q�a�@��e��@[����D�.L��4fDXGx��)�O>A�vD�bs�![q��$��9���Ц�	��@��C�
X�'������<����clH=b�aK#��
-���>��g_p��?����?r&�\�\zSé7��0�Gm��
\�P�����0�'JҖ|��o�
a#�	� ��uxlWt+�O�h����	����Ipy�B��$s��	V38����Ք0�+�>���?���?���)[|}�=x4�ߙDР-�ՆU�zz6-.���Or�D�OD�$�O����O�H��� R�z$�fHùzo޴Z3��	�	Ο���_�IΟ�'�~���4s�l�i4IZ=
�@�H�燐+�N��'�"�'nb�'7b�7D"��'#"Í���� W�S�p�N��"7��O8�O�į<	q�s�ɡѦ�{��9���c  �:����ME�[Y�P��OzaF��O��@ EϽ@fP�3�G�r��(�"O"�q�Oр-�,�4bD�g�4�jdA�%�-��a�1I-XT��/��L��B.�#ά� @8u�z�+�C�1І�[�@�c}r��V:f�l�R���؃$n��N
!�vI��M�W��(#],J��Q��쐩-88��݃+�\��@&s�UP�ϯ`�2�!���!�����B�S��	r���O����O�d�ﺃthY/V���Kؙ#Z�cs'��t�=KV�ӫ�y�ɤR艌�L>�ߤo��cg�ۿkl�y��D",���Ӆ�M#�y"+S� �}&�tHEf�UK�S�&��49\��`�¼�M���i��ij��,O ����^�~@�4���ԋt�
1�B�ɀ:l����CD�]2�P1�_�^@�D����ȟ8�'��Xy����>,ir�R�~��s�jL;Hp����'AR�'�B�~�y�Iԟ�Χ��m�+0���y"�j�@�m��݈��'=��TA\t�,��kL�OR�Tٗ�'F�TT� H�8��'GŌm��猈��N��<9��x��e�(Y������W:n���'iR�m�"l ����X��p��Q:�^]�ȓj���.�ф`0B�T4}P���<ɵ�i��\��*%�E�����OP�t�H%!�����Ѯcg�y��.�O����O'<�D�Ob�S�����w ^�s/.��D�ˬL����o	�/�X�+!.l]�����'�`�+�iY_��U8u ��t�s�Ǚ�`�$�7�z(I� [<��P8��J(2!P1а�|��J(�?A����҄4=q��7��p���� ,1O���R�V:@J��E
\n�݈7��G{�Oo�7MI-66��	�@۲m�2��n�)��Ľ<�P�M:w����'��\>]0��џ�x�N�E 37%P�75��K�̟���5W2�ux�'��$	y�
Ȗrd�.���';���Kd��� ����ȉ��8�O��J���-_�XE��-E�RG�DAv܌���o;!fX�˲L���	�|C2�$��YJ|BK~ҧ̕�	��mdj�:߄���e��?�ϓy���#�D����0��'(8ռ͆�ɶ�HO�aƨ�E.� À��w�\8�ISۦ��I�|���Y�
Y��+PΟ �	ٟ��i޹��5gJ��t�Դ$8
��k �]���9 ��t�N�S��k�F��|Ұ�>���)5�
G#)Q#@Drgc�==��{�L�FFz�:!ƸP*,�3������	ΐq����w�,LH�Ǯ�2bDw)��9ãcӰ��'$ԸC��|��'��'��p�w+c��R�$\}��z
�'�<Y�#$G���+T�ӣ�m��'B7ғE�F�'��I�M��\J!�]$DG�g�ˇ�:���6+��q�Iğd��ݟBYw���'9�)�$+�1�vG@�.�f�A �£,VҬ��f{ȔH��K<m���	������ʜ�j^6pB&��^�.�T`+M���DF��Vr��H�4��ƯQ"(���O>!���)��TK���1JuXu叆G� T�I�M[�i
�O���~� d�q�j4p�	U4>R4 5�B��%�4��՝\�|�)&
�\�U���1�ɡ�M����dхP.�OhR���E��4/��#�֝,�����?�%��?����̧;�xi�Qƍ�r�H3�O��3��H�X=�F��qt��d�'��e6�I��hTc�-0���h� �d�t��߂ah���_�kџd����O��m���-&-�)����o�ȉr� �-21O��D9<O"L�\�?�8(S��\%]6QOܱn�<�r�)B�P�ac�#?J���EyR�J7��6�Oj���|�s���?!�d�e��X���L��&mI��?Q�A�LH�(�}�D(	���b���,��˧Tsʰ&�R�>@����L`�O�����<
=����"�*1�B�ܚq]�d!��;� �}���$��fF֭�(�/!\�%J��>Q�i�쟸�Iퟀ��x�g�? �TА��7�H�r�=:0���p�D�O���$D�e�BɪA�߅66<l[ ��N�=�'/M����&g۫,p�p���P�0�J��ۿ��$�O*���U�\0�`m�OR���OX�D���I� ��$*|����V�X0؅�W�89����eR�+/`u��eQT��c>�OT��"*Y�<��i���԰Ad�X���x���Ӯ>^H�c��O��=����V��ˋj��;b���bL��M�\-t�	 ���$�i�7-�OYb@��Oq�����G�|XT��ϊ�:�3!�Kh<�2(�o��A�1I�\�=���K�<���cl����DiH�'v�]��j�� 7�Kщן|�%`&G><Ea��'���'b2J�~����@B"�xh�M��y�U �K��̒r"�`�V��'��ib�yR�ߜVD�9b��e���X@*�>j*IFTP� qE�2��yfTFBpa(�퇐 2M!��+Ƞ��ݛv"d���<Y����'���y���t�������i�p��'��A���ОI&fk�g��`�qˋy҉�`�|B�!�	�p~�̈�mX�4Aʤ��JΉ=!�$�<��"�W�&���qG�F1&�!�ĜN��Bd˜ sy���h�	�!��Y�N�Z�3��.Ko�����۳B�!�$Vg�JZt	@�c虻&Ĝ,VF!��)~���î�m�����^!��,��-�4�Ȼ m����`/8!�ُp�eJ�#��=O��RE.R�CV!�$�KI���M�9@dR�ΑBC!�$&_��5ꖏ�.g�r��B&!�dһ˖��d`����)!����̋�cN#u�=��,�n#!�V�xaB�"&G�IjaH�X	!�D�;S��(��A�rv:m���œ�!��B1n�����y9 �@g]"A�!�T_RV	#�Z����F3G0<�ȓ�iZv'��S� �]�#��i�����f�Xr�Sw�]�j�ȅȓ�H�D�l��d��kۚ(����'J�]� >�nxXF�O=8ꑰ�'�����W,놱{�c�y�� �'�LH�$��� Kt����'XL2QI�7z �� Ej�L�i�'zT �A�>?N����_� �'��a���Á3t�����^���
�'��ݣ��ˀ�uQ�O��xؐ�'��D���έb��HJ�.
���b�'�$��T��S�����NI[�'T$l�pm�&!ld@�b�U�C� �
�'���DI�}+H1gYE�ڍS�'��kU�Mi� �D�XA%L�a�'i,`;C蛚/; H(6.����'d���Vl�!zU����%')���'��u�L6i��PX�ɘ�o L��'�x�@G�>��{Gطm��0:�'Қ(���B<���:��״w�LL��SSbHi���;L��U ��9r<���f�]�1p0�� EN%P>��!�J; ܒ	�P1K���5o�E|Baע��Y6�
&i�=�⅒A�QHFo��A����2V�&��d�<�1/St>��g̝4cl��h�bH�<�D>F�H1��ɮf����5'#��h�$�#и�G�_0�@\��}#��X�;Ӏ� �'�
@� ��3�_�%a��C5+2�R� �h���䕾!5�p� I�`�t���(��l�a~�['�,�D��!I� ��E�xA�'Ֆ5�D�X�� O��}��I+C�P@�䋬	��c�"S.,�����5�0��bJ���S&"TiT�� Y8�h���!�B䉄#�Z`"�,��[50`��'BH:�"K�8��4z@1꧘O��9�8�����M�n��4� OCͨ���OxuZ��Q�6���7�V�R'�bצ!A�O�q6ҵx�H�*P3&,K��^;�Q��c�G9(Z�ɐ�Y�R�j�P�O�p����,�?)��>A����<�䤵|
C l�? �t�������x4�	b͜<A��X5}�p:�J��p=1RE��U����V�=��A�3G��[���+.Qn����O�88C�n>Q����R�0,H����]�OX��A���N�L)c�F��0<�'h�dt``B	w: �c��ć�N��wEӓ94�����saҡ�<���>��皆g��ij[wΙ	�ͩ��9�C��(�F�p�ɬC��D3�=?	$鐳�̋b Rgp	�M�hܓ�Mc�L߻��ݙ�D�aG^XӇF�Tyro�7PA�{eE:i�0����(OЕZ2F@;��q��� ��HH�L�a���'#�<G��䍆P2ДX6NPY�'x�!V��d$��#��D?��3�� �~A�ENRH��杶zPPMQ�AەhӇ �o�bH��!�]�����KJl rI
w���Z�^<Jg��~�����'����q�@|{���B6]9$���"ͰB`D)���qG�����(��O� '*X|���9�m���@�X��i�:�k�AF!U���Q�	�`~fXz�O �J4,I���p�K'26�*H?��e�}�ȡ5j���-걎@*
j5��<#�؃���Bx��[�ML����b*?����OK�!U$��Z
!�F1���	�q��Y�E�>�O,�wP�l����@�F�zt�I��%:���oS.E�r�b��Y��x#wH�&���'�/�|���
,1۱l���|��׌*缐%?�Hl�*�8�)�L�� ����3�S��l[a�'wM����"T~�y0�'f��(ۣeǦ䐬�V�C\���c���}�vm8E�
.�>u�ѡ�Y��,���l.��3�ŸA8n��Č3��I8p�Z��놬hZ�zD��,���G�ܴ9�B=*�,_�x]h)�{I���� ăbM��2��ǥ6"���0j��<Bb!�g
�}�Sg�=d��(�2�d���x��ʧ|���ʟ,�m��=#�ʆC�W�
z.$��K�bM�P�軔�'1&it�Ӑv12�i ���<����V��m�̠Y�+��Bx(�WaO�(%h�����U9"�)����8�R������mJ���7�\$S��]�w��">��)ǀ�� ����$j�i���<�b�U-��`§N� ^�f%&�6�Z���<jD	��� b���i�$�]?Y7 0�$m��*F��"1�IG��	R&x�dHRRC�Ur��R� 1E�4"�d�LY�L�b����%��ɺ��a�cޏ�~"�9`�Q�8X��I�-�69Y�GV���h�N����چ`��u��c�G�Vit�'���.oZ��پso�����P|wH�ǹXX��aϙ7���qu ��p<�`��]�^A�i��A������x � �H(��{k��s�d�' �0q��$R����ԟ�u1�!�{��5�Շ��u���I�nf���e#̇F9�Q�l�2�S�v�2ЙE�6J�Q`AӶ.�\Dj� �� =b�L%6�4�Sܧ-�H��;$��9:�&��>D�%��ϗ�?��dΓS���E@<5l���GTDe88����(�p����k?�(��Ɣ���3K�����@H[�b�i%��c4�<9U^,^�S����DI�[m��ԁ�7'��0+�1`	Q"��d
Fw�4�P&Lۋpb����,s4�L8�
0fW�s�����d�Z�&I	�SALx�1�#\�\[G���Y v��0L ��C�؇1���g�%`��`IG=|�\Z�O�?�Y̓p� ��6+�l QQ%όM��PP� QZ�">�bm�=@�*��7%�$nj4�&FS8���Uv���ږ�͝O�������51Nt"���)A���(O��xI| f�(6}��.L�nq���^��`#��D.O&��	7N�\a�[0A`'�]/�>���w�'B��n��>�2쀵,��q���<�Q��oKy��#�;w���f��\�.�<to�;��u����\HH�AW�!7F���dN�ii�̝��t�tg�_�6�9bFK�(�r,��4l�.|e@hN���7@�xg��r�ҧ`�����>�OT̑B�ΞT߸9��D��<)�4O��K�[�C�N�B@�ݱ�D��ƅ�|≹g�	��*�D#�ɉ3>(IgJ�f�!��T�i�:�Qc�Ԗ�t��A' LLt�"��8uF�'��Jl{EA�[�b ��8����l�-Hz��a��A:�"hB��'�4 J����%��p��A��:�6�%�N�$���c���T)�'c�	��uI��]8��Y�3~�p(d#ҖH�Hm���E���2���"l����&8�Z�S�O@<T7G�0�u�G��?����Su��92��!e���N��d8����Y�\(]�f	��$��˓3!u�F��0|�/Ey�n�8A_�i}�t���z�'�PuQ3�O�frd�u
��`S�����|jV��/�R����ӝG@�0SgX���'����g[-S@�AI�ǟ�,M<I�h���]�W�TxD\�#���4�����5?�J��C�"��A�韑�8���8J��Y���L��
yhxӺ� C�&�O��As-�5o�����@Q�bD8�#�?tW" �Z�'^Q�|KA���v�I`"�	y �aK�I×T�8���@n�$� �Z>�Ӂ�Ĩ2��&�R�`FjH�>)�i�I�/��ZR��x�FE��$�b-�)l�����C�-C��Dx�mP
��"�K�X$pCc��?��$e ����sfМ�3aV�L��aY�{2#M���-(�D`�1����O	P��(UP��0�hγe8� ��A�n���-g�=Y҉�0 ��'���2N<�]�H�l�S�lONԠH)3��#C�4��ĖEI���@��r���;6�^C�'��A�A�f��B��W��	ʡ�	!73@,I��(}�Ib�'60bW������a�i��`k��3b+6�y�a�� 뺍q�#!�� Fd �m�r��e�4/�\�	bD&00@A�""W��S�!_м}q�.@��udI}�	� ;���Q�)�M�'�4Ļ5��Z�� l@�ؔ���?7M��\+v��q���|� ��*Q����|��� �$ �T�� �J�U;�����`� A����5>�1@�V���R �q���Z��=C�h��3�����9�!S�����Ӏ���΍[����%H�OΌY���y�g�	�K@�sE��������82�l� NЦ�#�Y��;aӟ\��uŨ�q5�O�ښ90bգ �I&�@Ƞ�l�:����+F�p?YrI��F"��(�КG$�h��A�e�d(h �߭2� �d���uY�������	�Q�`�q�e�	�����K�9�������qyqk2��O<�D '���Cm�ANdc"��n?aL8*�	��:E�9�t*3��dR j3�Dx��A/Nm���G�OD(Cd偤	����E6F=p9s(�2K�d$�}���j�d�X�-ĵG�B*Ηm��0�"B��5ZB]y A�3��O\E;��v������)p�L@�E�S����}A���޴)���s���xbV�ʧDmA�]�)ZI�tʖ�/�:�%H�6$������譑!-V f,�̃s�lG�mJ���:YRb`��'�>����<9&fC�Mt��� e��h7L���`��ڀ��<��f�i����X��?Ahqt	i%n�;�����Yc�&�Q�A��R�&�х7O�p�l91�tk!6�����H 'O�d�91��<6ޒ���@�t݉'�$#��סzi�@��'�Bt�+O��raf�1KX�G�H"B$IUk�m��f��4:��f̂S��Φ_�v�R��E�1)���4�(�	�'�*;z�Y3T��"h�HQԄBz~��<�"��p����G�7o���S�R�L�Ys�F3�~��㨍3F>�*��ԸuGl��4�FŹ%I(lR�� 7!�"_���OB`��'	Y��o�h���R$5�i�,#��CfF	� �qa�վ/�`YC7�׺�0<Y 	�+k.�|��
�q?ּ!7��@�ε���ةD�v)��X'��I��]_t��
dcG�<1��ߙ@7δ���ȉ�*��H8c����zn: ��(��Oi���0B�%�'�p�/�!]IR�]' �DQL��9O�(��댺 �A	�//?��Q�� ,�ވ9��8p���+9eY�	�&�=�Pr�]@\PI�5O��3�>�@a��S����<y��	�r�i��Фk�����
dA2y���4s��)��j��oC,��ШH1�ӼK�
ڼl�F��O	DL\�����P���&c�<������F��V��SZ�LQX�̒-�T����Q(�y�'�-O`iá�E�i�a�q�J)�fH��oB�H.b����S�n�⑩!��W�6��d"�>J�.4�B0OQ8ekB��b���4�␫%��6&�$�/#����S�O�pjVQ%�ҕE1�ɿvaԍX&B��orűal8=�J��~��itpq���?��-�&*��kQ���@#1~ݑDgˀ.*Rɹ-��dQ3�=<�dA#(�H�d�1䗦i����GAG2prM�0�xӆ����G�|
��i�0,beƒ����q�qsW�H"}�R@�K�&��#�7u�%��Ӽ���8K�֭�m�&9"BM�;9�4,N�m՛6M֦f�T�+�����?;.�l�
DΎ/5Hl%QQl��4&���@�'�|�Cf#��"���3��&Z�P ���� 1yW��Nl�#��O 89t �7U���L�����ڠO�m��[����'J00�B5�#�+��$^� �,�h�W��nx�R����y�n�|�88)��( �w����'����ݩ��9�f˖5���1����'\�n<s�c�/Av���-Q�{i�|�!��g��`G� 
\Ĺ�>��}�'Mz���$��
��Ё�B�aV(�� ����b���Ӽ��C	<�(!� ЭK�@�����	�Đi�ry��Wt�.���ؗ���3�~�{��5��1�0�'��5��ݎ?VX�Ӽi�����+�<�u�@�<`���ٛt��`d�S��A�W��>y�Bŝ�wi�F�n(*ņ��v8 ��F./�!�D�9�B���ތW.�q��U w�!��T��4�%��g�
@y�"�2eh!��#*:��jV}��$�3GG�K�!�D�3;a^AS�/��
��bu�߆x�!��-r�p1�T�*���È� �!��R�S}�+�%H�zV���ș3�!�$Σ[F
���Ūvh@�A����!�DJ�^�@ �gXrˎl�@���h�!�d�C��)b#�+�|Lqf/J�z�!�¤k|�\@c� �\s$�x!���(z�����ׯM�t�S'�W�t!�D�b҈1�g����X c7�Վ=�!�dA-t~X�d,úJ�J$Z�@
�|�!���G��m`,־B�6�Y �%H!�*5��h0�,�ܞ��`�f:!�x
.�q���\�I'��'2�!�D
d���	Q�O�f�zX	�	�J�!��ܤ��h �´S�Dmvi��5!�� @�� a*h<��F:{\�3�"O�A�%]�a�0r友.�P��"Oh| 1��<7E�l@�O�+hy��xF"O~�q�A�&yniH�ώ%g�g"Od�v$�L# cō��
�<D�Q"O�3U�;V~�P)���b�L!9�"O^ ���M�b��P$��O��)Q�"O0���H�I����ÿ=x�ӆ"O�)��kA�r�zPQ��ڝw�e�"O8� ��0&-�ȃ�p���`�"O0�Qc�ܒ\b��q�'�+(ǢXf"O�yP-A�mf�ZR�>[�x�ɰ"O�� +�R��k'��r���#"O�0��H͘@��ZŌ�K�'�H�e�\&(�\�������:���'r�@Q'gM%�MʐM�Ф��'c��B��.�F��/��4�<ES�'����s�[�мJr��Wn�<�
�'欹�(��T�;�NɧHO �A�' :x�ăY��%�ߍ9�ll��'�z���c
9Z(!T ��I�2�P�'�{����}�H�C�M:Ө9�'z8��`-��P�R�F�_�R���'OZ�WO.J���R)B�@9��'��aZ`I�!����#�*:\�=��'7�q�gc�w�n80�* 7h��'�6���f��eY�k.��+B��;
�'ƴ��AK?gj
|�g����	�'�]�#��;v$�h���iy�-	�'�@!^]��BDU6]@X�:�'p���ǈ�9�F` ��� !���p
�'dD1�FLW&O�(��'�Ïc���
�'4f�:⅕$b���p�
��S��h)	�'� ��b��w}f�ɳOV� ��m��'y����]�u��<�C��<x�zi#�'�&�`2�׻F�q���oLA�'��҅L�%D�*���/i�D�	�'SҘ�w@�`�Cc��5c�h0��'��iY�gX=s>���n�X��1��'�a1 �>��]�''��J3f���'�R� a�ګ[���1�-�⺸z�'m.dH �ۮh�9FB͓[<�}��'Q��a��&l�ȉի@�Q�N��']�0ŉ)o�E��,4K�*���'f&ذ�׿.�F8$�4��5z
�'��* G�!j�:)ҳ)N�1ݨH��'I4�����R�B�%��%]j�b�'{��bA�=	��dC�ɳI�����'�.qsE��Y����ͮEgR1��'�`�1@I�|o��$��6��u:�'����w�����C�<��'���I�K�C@��旻7�FP��'R6�;�� ;Ԍ�C �V,��Ĩ�'�\�{��K& ���ƫH5YJ��
�'iB�+QH
y>�Ë�d��3�'.���� ���]ɱBn��9�'����R_�f! �Q�|͒���'���@��!w����`��w#|�'!��˵�Q�Z���i�'�i
��Q
�'��l�a�V)�8���(�l����(!�S��?�@&
� �"äݚT�6T�"@\q�<���ؘ���[�Z?l�dQs��]r�<��łK�\՛'f�X��"�I o�<)��r{.�3�&��+o�� ��j�<� ���,^� ]��L� :��p!�"ON}z�JQ,4������
D-
��"O�����_U�(�4L-|������rx��cG��E�T:�ʕ�Z<�u�9D�d�Q-�,���[2n@�� =���6D�x�0�9M���X�cĠ �5D�����ǧgm�u2?c�,7o D�PK���5+(�����;e�f<*��?D���,J�#������ӗ]��̑��;D�<k�+�70 ��3Q�oӐ��=D��1嘼�a�
ra��&D��1��_�h��TA�
�P��&1D�d!���$<Q����['�F��c	4D�l�b탽(��h��ؐ$��i�C0D�,*7�۞l��d�c��,}<)�ǀ.D�HS���k{���A�C�9
�x��-D�� j�^rd|���A.p@\�i&D�h�t.ښSr�ܓVN��t$�q����hO?���,N�1z���L�@Ir�/U�l!�$�-j��Q�	7� @���΢lq!�$�{ʪy�/�6XҰ2��a}>I��	\�ޤ�T_�]�\��7@�k�<���/�(��H� �x\��K�j�<�7��&s�|�r�D�E0E��P�<QD]8l8���6Z81S���E�<�	��,@E(��G�w
x����@�<Y��L'QO|	�p���`��s�<�f�ٖ,���e��4	��r�<�5K�	b$� ���ȫ5e���oE�<��HX�<�nK�╪I��7hU�<a�X4�^}�RFW%���(�BO�<�7��4*&B�!����fq���V�<�$o��<�E`J�.�����l�<����
Q��a(T�xejwO�|�<��@H0���&-�����Mr�<�`��NO~upW��`e4��c�<`�fpe�	*"��צ�Y�<y�M�'g�T�2DG|~@����A�<	�ᙊf��X���P�5}ukD��}�<y)�M,��k��s�`D�1�Uy�<i���6���"��T�@��#tJ]�<A""!2
�^�a��D]�<����9K@��
%� �}}�\�f�[�<�T��l��x@SCE� I���k�L�<�@h�&Pi�&��
��`�c�J�<yF�E�u�41A⡘��8erH�B�<1qĝ T�BѤ�-���C�H�<��� ����
O���*s��C�<ِ�NW���@勻z(Ly����e�<�A�gv�USb`82̖ij���F�<�"���P	1�Ɖu������A�<�R�lTI���K�@U���o�z�<�#�?�8t#*�rX�����x؟��N�D*�j�1"��	E,O�� �ȓr�$Q¤�[>o����R�O�<�Fy��|*ǄF9���Ra��&f�V�O�'JQ?�م���w��y0b͚q��dS��1D�� �@+���q�Xd��t/D�� # �A�X�3Aɏ?dm�F�-D�T�5���H���AnA?G�D��r�?D���>:��X+�c@lrF���+3D�|� `�(PU���Ѭߜ��U�0,5D��N׾e��"�^�g�Q�5D���J�6(�X)b��W$[���	�>D�� ��Q!���l8� �+K�z�R9H�"O��a�Lł�p;��"(}��["O�-� ��G�j�[d��=�� ��"O�;b	�:P���Ӄ�>��Ļw"O���0���q�0�DQ/�Ҵ� "O\��F�қQ��j�Ȕ�BZ({"Oj�9��>P���g6<�Q"O6I�S�-��)A�F�.N,�1�"O���@C�z�n-������>�"P"O�8����]u� �ǒ)�$�&"O>�IP"b���R�A�9Z���["O��# _79+�� ��Am�ԝ"O���K��sU"-��Bʢ���R�"O��2�*0R���� "�7y�r��"O��p��*��PQ𠑮��`ȡ"Oh<r�g	03��	,�  
�"O�l�ņ��xQ\́�ܰ; �iJ�"O��hd2voU�6�b)Q�"O�L�ӦF��@�j�D�XA�QaQ�P����0���9�d�Z�*9��?�B�5|�z9�bL�_��1q�Y�C䉄`�4	�W��>�Ԕ�5a[�J[�C�I�.���I�*�8;�����W8W�hC�	�e ��	�%Q���!���+N�*C䉾�`p�J�9�t(�Td��^��B�ɸ�4E�#��4�P����4YHB�(d��Z�*t<�(�.�Z�PB�	'^���m��M�*��5��g
V�D:�
��#�F��s�_
S�4X 0M!D�t��&B�WKza��ңL ��K>D��rQB�$$L�a'R�u ���=D��S�� &4lH ς_���)>D�@�DCܓl����%M9F�	+t�:D�d�g��.k��Պ �^��q�.D����ѩ/?���g��<Q�U2dM.D����('Rn-xp�]C&��3�,D���	͗l��EJ��	
��0�E+D��c6!�%q�t�+`�*hP��k�N)D�$����i���r\�\�%N�_�!�$^*4���g��,P���ʘ�!�A(a�@��Y�C�2���hܕ2�!�K�[�Ļ"�_�m�x+և��Ww!�D,Ș���P�d4�E�	tX!�ą�^!6U;D&�Q �-@ ,c���>��/ɲ�|x�%�8�"���T�<Ɇϖ9'p�! ��1Q�IR�<A�$�q�l�s[P��P�,�X�<��@ Y� ���85��E����W�<A�F��K3�ՑCf2�8���Q�<y�n�3����NC+0)�`j�Y�<�c�4)���s%�C |c�w�Y�<�"b�-zY��c��1M\�i��Q�<VAE�-������XŌ�=�"B��${��B!Kʣwu�u�e%X�'NDC�	?���H�v���1�NW�o�BC�I Q?�T#�W��.P{vk�x�,C�/%R`�/BE���#"܈g�C�I ���c����A��:��C�I�ql~�Q1dٝsX
�X�H#�B�	>$����'��:a��a�'[ie\B�I���<0S��

�,�i�J�h*�B�ɇU�-ґ�D�y� ƈ�/'�B�3\���Jga�(:H�gh	q߼B��0�v����$;�>A[���J�B�)� �l���қ7�b�	���}��"O^-�$�ۗB8��Y��� d��X��"O����k3?��e1��B(*��Yi"O*�
�I�7:3Z�K��\��Իf"O�X���hkgF��b��"O��9tA��R^z�2�����h�"O�̱�%�.%�ԭIP�%2�*d�"Ov��֊2�١��K�Gj�H�"O�q��@�7���k⣊�=��Y�"Ox����8ò�Y��-,9,��"O(�����S��h��K�T����"O�D�r��<p��ً'GT��"O���C�����p�_����"O�P6�ˑ=����n[�2��$# "O��������,��Lt�y"O�@�B�'4.��+H
5��V"O��O��<Lt��bi�da�p"O~H��$ �e�0K׵6�\A��"O�@�O�$�����!� af"O�]
�D�'�mI��,a)���%"O ��	�L��a�JO%?� {�"O�{  �
I� �J;�Y��"O0�B�0ke&qi *ƻ"��Q�"O�t	_�^�����J_�����"Oj�0�#>x�w�ɡ=�܌h%"O���(C$W�^Q����^���Q"O6�X@?7LR�����&��u�f"Odݨ"���v����3zF8�&"On\�o|Eڵҗ��t<�*�"O! ��Q�E[�ț3��fV���"O��e*U��B"��J�$��"O�ႃ�f��MР9<0�X%"Ol��%��9f]� �<R [!"O����!'Sڨ�� ��%�4�"OR�r��3c��zHʍR�T��w"O6��C#�;Lh0�&R7t��i��"OB��浲�$�G��,v:0j�#C�<�c��
<�@��D$(�x�	u�e�<)�kCm��!`g`�
m=`sS#�|�<a��˫Q�<4�͍,��@��x�<�D*��s� ���&Mm��а Dy�<���,?��t��A�E8pb�z�<�h͠[�T�ҕM�i*�� A�<�wG�6w����R�X��Ex�<�eD�}$��� ĂJb����m�<	��HrJbF�=+�J�0�'j�<91�ݱ+;&� ��1\ˀ��3�Nf�<�Ɠ!����V��A_.�ɠ��k�<Q��]L���'l�./���2�He�<��Ç940�( �?f, ��
�d�<9v��*	��Ԑ�NH�,�6�)�D]a�<!bgN
G��ۢ%�\
^����JD�<9���KT�؈"`X�T�v��TC�<yGB���}�E.R�09�f�
V�<�N&OFN�i2�J�������T�<A#λ.1�y�e�� �M��˙N�<�H�m�^=U_�3[ A3Ӏ�G�<�#!ÿ)x8�Uip��"��|�<A�J �f�1�a�,��Ɋf%	Q�<)�b�*��d��O
*��A�fS�<y���frar�hߋ~�l��	�c�<�ˁ�4����$�ÂK�^�Y%k�^�<�e��N RBf�I���O[�<���p�8�;Ť�bB��3ǍT�<� �m��i������ML*W��-Ӧ"O�(���ݝH*8S
!�X8�"Ob�IW	V�#Bb�Vy�+w"O����7~�����
^ܭk'"OtL@�� F��ӠU�Oޝh�"O,�ॡ@�D1�Ds���0.��V"Ox�z� �4`;��� z��"O�di� 8�p���ي�"OD���8��ܫ�	��۠"O��A0�ΣTz P�m�+�L� "O��2�j��⤈�ι2�TL�"O�!���3@~��*��i#����"O�)R�kA�w������3�")��"O<a�(֜Zٜ��r#��A���!Q"O�x��ϋ6t[��Р٨q�\jB"O@ŲW����04b����"OvŸ��F�s���b��԰Z��,
�"Ot����L�h����AJ���"OP����J*Xn�uk��9�Y�"O `�0�����ձ�@K��L�R"OnU��S�|�'��?+Ȓ�[�"O�bpL���1�腊B�@�"OL�c	�uX���F<�Bt�w"O���#ꕔ=��(���@w�Q�"O.uI��_,D9�H�쟛PV�;�"O���C��FH�y��K�z�z��"O�`���ķD�����IJ�%�$�+�"O��fnD�}�rݺv꓃o�JЃ"O�	Bbe�0�x�p���p��%P"O�-AfE�(0��bB)yl��"O�d��69D��he�Q�x@�Y��"O$eA4�K��DXe�$?�2}�6"O�U��%�|��ciY5t��+"Oy��d(R5�8�קN�!�*X�"O&���$]�kߨY)i�6�`5kp"O$d�mV�o5���J�>�F���"O���p֢E�(h��� IJ�dq�"O�(�H�.а�4�D�DH1x0"O�Xɢ$�+=�l�U*�AD	AE"O �q��ia%�&^�D% F�n!�$&��8ycj�!{�@�z��VC!�dH�X�~�Y���)�b��3��;H!��a=���d� ����0�^�!�^������B�%�,�ƥO�9q!򤀊Oтa��%̆����8�!�D�4&��j�e��Ce�	P�!�B�\��!��t����	���!��K�#C*ճ$Lߕ���cSi�/^�!��'KWDI��A��0�j$C��!�Ċ'C�D��H��D� }+��ϛZ�!�dL3W�hᨳ�Vk����Wņ��!�D'ε�!n�8�J����	�!��_$��0���ŚrA.0� #�	t�!��=|6�ʚ-i@�j���x�!�d��V'��!����c�>HJG�R>=�!�D��W$�\Q�ʓ�wP��C�I��!�˻1���Y��
�<Ȱ{�)��R�!�Z��u:MF�İ"�咥(�!�d��Gޮy�NLNhn �t�«,�!�d��[/$}�vJ��xBB��dGÕ�!�䂙;�D�)�C4b� �~�!��K�0��ၳJ�6eNa��dV��!�Qܠ=��	Jcv��'ZD!�L�ơ����+�č*6'�6v^!�� \��F@�CL�T�۟]k2} 7"O۠K�4�zIǧh����u"O�;��=6�� ��K�'��<�W"ODi�O}�|[ԍMe�TL�'"O���ǃ�S(�$��"\B}�u�7"O�4�í�>E�����K7`?� {�"O��+V$̃1BڕB�(��hr"OD
��������!_;Y��<��"O Q�)ޡ����B'˂1�u"O��Дj�GFl���B��h�a'"O@#@Ē[���1"ĵ�&���"O�p9�Ϻ/��i:L�e{�\��"Od����6w�&�:ъL @��"Ob-��K�3pA�$:Ì�k�"OX���ѩ+��cd-@#���e"O�`��B?xv�;��ޯ�2-
�"O��0�C�1'�m9�����誖"O6��3�z/|��#W]�Ԡ��"OL�;���zc$�"2�ي�&��p"O�a3j@��(I�v @f�Hi*""O�B��L�h�~���A �4D2�"O�	�7�ҸP�`�Zv�x�"O^|��D�"�jb���Wf��Sf"O�ܐb$�Il[A���"SFSa"O\���U�c.�8Iv��-�U��"On]k߮Pݜt+ݯB�dh�"O�q$�7j���h�4;�Ᵽ�"O�y��Mެ=ǀ!j���aa�}p"O�i�cf�2b��BDyJ `"O�����Q`��C�>�12�"O�ucnٳC�`�Q�у�6�%"O2��1�L�#E$���G�S�Ll��"Op�GJ;A.���A �~� '"O��R�HK3'"�b,Ǟe�Y�"O�p��%~8��r�j��"��ɢ"O0 �Q�¾&�@Z���>�(m�E"OD���.ˮ)�h���5v��q�"O*QՀ�.[�pg L���Q"OBu*���Q>�9��&����$"OZ ا��z!�Y�#��?"���� "O�!��@���xA�3?��h�"OB�;��
0 i�KE�[/Vv>���"O{���hj8�
���7]�"O ��'H�*�R�!TJH�=R��{�"O(] �兠m3���&'�M>,�P"OZ��5��v��y#bۓj_��"OP�k4ۥ`H>�(q�ӟ>Uz\c�"Obx#@��G "�b�H��vL�<(7"OfqS��+6��`�H�4����"O��`���FMXr�ƀdbli�"O��?W���KF	&Z~���"O(!�q+�0;�<�)�e]�x�"q�"O ��gcG���t��ܶdֶj5"O�X�!�R�l���5c� �"O����(Yd:���Nѱ`-ء�5"O(��BC�)J��` [�K�T�"O8C7(��d��e3W%R�V�S�"O��I훔tK�T���]{�z"Ohx@үX�=�.1��[�^Xf(CG"O�qRE��|Ό��b�4+���"O�P��#�	W�f�1�/��az�u�q"O!��T7K�B���@��|��P��"Of���g��d�ۣ��2-{"O(����݌4
�.wy��"t"O� ��+1�U��И��K�a�P�s%"O2��!�;0/`��'H���"O�ģ��;���� �u.|��D"OrhC��	j����텟v�k�"O��Q'I�'䨼bW�h ��aS"O�f,��Yޖ��B���d�X7"O�Y)�)Ñ�����w�\K""O�(����^�s!̴�����"OJ�t 
� Ap�%�,va6�yq"O� �a�7���������lK�"O�8���\�N=M 1C�"��q"O��"���!xp�K���?����t"Of�r�KW
2�2�h�k�8����"O�u�6�Ѝ:R(���N�}��Ȉ�"O0�F� �+Ҏ,��)[�{�,��"O���^<E��݂5�P���"O `�0k��W�~��i�1bj͠�"O>��fEM����Ă6_d�qS"Ov�$@K���M�d"�8y�I�"O�m��ޑvp03K�9&���"O����L��KdI�2:��"�"O:��eDx<���d-�>4=4��"O�D+�d��+K�e"$��7e6��X�"O��I��)�D�4�A|L��i�"O*D���TG�<%yeG]�2In��V"O��J6*&oR
���G��]K�"ODչ+3:�<R�f����"O
�rCV;-d�ydk�cJ�!"OnKw�.�4I"���!y\�4�"O��BP`\���1�ϑQ>H��S"O�$��9�<�BoPh/fܡQ"O|u�s,������~�"��t"Of5�1A��C~Pц͂YP��f"O$abQ���B���PF�
L��"O�0���ʢf���vD�:Y��8S"O\�0JY�Q�XIyP� /�$1`�"O6Ł�F�.Q%���!!�.�iu"O~Ire�V:�`[g��4x�����"O‫�-ô[���q���U
�"O��*�fW#�B9����n���"OK��LhֽӐ�H�n�"0y�aR��y
\ "�yz����dW�,3ց��y�.،<�H�`7ś%l��욲�y��\��i�1��iRń���y�U�3b�5$�,u��$�\��yr��R)S6cO�#�ac�В�y�HO�[<���ee�� Պ]H�A
��y�`�M����wʗP�*�/R��yBijˈ)�F��D������y�!��4CjE*.�!4D����^�yB@�5���������t���@��y�GO�����N,�F�qj\(�yRb�5&���!�AH6 ��c�ĕ�y�"֢o�1!��_�����/�y	��S0�x���F1�Xf�۹�yB��*(�}鳫M9S������yrk )H�HǞE�6�%�� �y��[�H����'c]���`p���yҢ�6�a�3�	:X !�)N�yң�<t�ʕ�9EZ�|I�	��y�}3��ɳ&���c!�*NJ�ͺ�':�5���Ӆ�ʑ�m�4��ݫ�'Kphq��R6��];a
�Z����	�'W��h�r������c���`	��� ~a��9|IׁC�pI��v"O.A1,f�4	�N�>~��RU"O�p�sN[�(��da�*�1��|��"Om�G^�3��٨�
�-o���"ON��*[�J�ސ(�Ț4�A��"O����:g˦�R��9?Ɔ�)"O�ȕ��muf��1lZ�L"O����&�`if���I�  8� "O��#��ΙUx���E��(iXK3"OV<E��(Fέ���B/dP��R"O*h��B?�^�S�,T�P0C�"O�a�����^��Y5���4\<��"O|"tbܴb�n�(��.��"O�}� aI�S�vx8���<3�(�"O�e�0��V���w�h �4C"O�=�U��(��Y-)�eKg�3�y���l�H�!�S+/LyF/И�y�٩� d�R��=5��$9� 2�y��/�b��"ؿ%���"E%�y2�<#�l�c������)�lĂ�y���!�$Ĺb�D��`�'��"�y�,R/�FM�Q�U" >H�6͞��y�`�o�r�S�սsH��6ʲ�ybU8_��LiC�o���UM3�y"�J�}@~`c%�ޢ���B�٨�y"@� 2����&\���ǣ�yB�9zњ�Х���챒aH��y�M�"��	 L��dH��Z$J˕�yrL�.�jr�OԞ.X��K$����yb�VZ2v��G�̅""�E9�f�yb�],6�D�c �2U<��$0�yb�=E�J*�A�'���j�)K��y����ؠ8x@e�&4��IY�(���y�(��{�����9sD��7h��y�f��aO� 	7���`�������y���>ILf};g��Q��D8v��>�y2���Z����M�6����p���ȓ���q�,�f[PY�b�,^#fŇ�R�*�m�.1v�؈��*Z�}��>�2�,��0}V%�w��%0�C�	��=	�d1�*"� �6;BC��1�9`��<T-P�t-�4*�
C�#"\҉8f��|�J��1C�	/{����C1�y�d�ş[��B�ɐ[~JYj�'��x���#
�	��B�	-UW��x5��8t�x�����B�	<T#�q�0ڼ�P�K�X'o��B�	�-j�lh��l���a7�H�!"O�@���.Z���pR.$ORH�2"O�đC�f�$���@!PO�+�"O$��Q%ٍ0�V�˰��9Rp�x�"ON�����a�H��06��J"O�x�1'Ӓ=CY�"�=�U�0"O��I�s��2w��h)c+�=�C�I"H���
t�B	O��4s�d0E�B��z��&��4��x��D�{��C�	-e?"I�F+��z��<���@=D�����^7��ƫ�'�\���?D��S)�`)V���)��CK���S`8D�v�_�l� (�®���u��6D�����R(Y��&:@/����6D�z��������*]���{v%?D��;��U!O[0��ʃ�Nݜ �6�)D���d�O�ܔ9$E�;A2P�Gd<D�� ��C��߇bq�e� ښ`PĚ�"O�(��F�1N5��9SE�P�j�"O�,3����"8�4M�(tq�4�B"O��xe���|��L�Lև$k�ɉr"O�i`�Z�>Ry;D�]�)b $X�"O�=���W=F4�!UE�M�U"OV����Mk�6��Ά
^(��j�"O���g�ǥDE��ClI�J(�"�"O���hQ�U�����4%
�Y��"Op��V`\�!^ �� ����x�"O��Z�e@�/�hx���[+vv�R�"OV��D�0洲 aA^*���"O�������Vm��`3����"O�*vh͌NI41A�*5FN4��1"O�HY� �mi����9R�<�"O<՘b�G�Q����ZjG� ;�*O��#��L�*��s��R:��=�
�'��\�#hN�+@��Rd�L�AT

�'%В�ڌB�9r4H����*	�'y��;��_.�PP�&f�$wY.���'~�U1A�H�H0n��5i�m5�l��'� �a��ߚB�a��k@�]���'����"�*qΪ�ɰ��j`�e0�'���*"K�NG�HI ��P�rK
�'��U����T�R9��B��Y%���	�'�.i`І�;��kG�g���'n`�qF&�*���:rf�`��AR	�']L�a���?I�d���Tј��	�'i�x��.Arغ֬�G�v5�'��D��'�d�!F ��
�<d"�'�PyRWl��L�\��#|� -�'�V�@P�C�x<��ܜD4D̩�'OD��QA\=.�� �K�.4!i�'8��l ���ǭ��l��'F<��%Ιp5Z�P��*JjP�']���Y�74e2�õ�D��'n�P�@�D���UK��y
�'�����^�u���K����Y(����'����^F@D ���1&]��)�'��9�vB��"�T��H�i�24	�'\�� ���64��k�kƙZ^��H
�'Q��9�!O3�4�Zb�ϧ�A�	�'�@{&�\�r��@���QM~��'��z0�$�Z|Q6�W�Fh(�!�'8]"q�����kB C�24��'�Ș�ď]Ղ�(���5�6���'��LȓBQ*E�r���לV* �b�''\�Y C~t���n��dI��'j�92���&c:ά	ף��f�hXA�'J~�b�� H�B!.VYu.y�
�';D�B���:5 �[PPVt�XI�'0|<�gÉR��+�&�G�ޑ��'�̱Z�h�O����>A�j���'�jPy΀ f����߱Bz�
�'��0�d`�qD�� ��?L	*@�	�'*ʍ�ЋO�	|}� ��00wfy	�'(���b�^�&�p���Ԯ$��D0	�'�NI@]�ޜӇŀ" Jx���'������*1���h/�<��'	��� �s����ن!�ȁ	�'l��h�=V(Ih4ϓ�g��H	�'@�EbU� ��i�6b'9����)i���9.�9 CuCU�ȓu䒽X���	X3���A�F�5%����S�? ��jP� _vm���MV�l"D"O0�w ��Ṟ�m�&� ��"O�9:�ІBCD��cA�_�H`P"O�%�%l�c��E���=|�ĩ8`"OX��P�8sN������"hu84"O���4�C�[x�q4��oi8��"O�!���ʭ1��Yْ�T@U��1"O\e�-<.X�P�cBö�R)J@"O�II�,qO�Ѫ5l\&t��@s�"O�q� R)FP�0S
�"IL���"Oh�0�
�-bB���ɏ����"O�xqID�C��00W$��T$�s�"O�q��i�?(�2�Ү$I�"O��y��Q�y~ԕ��U�W�p�"O���@f�5,,H�P��"̹"O���b��%]/b��1"�Z� �C�"OJAI"��H���1�;���"O5cƬ��$4�x��O��Sm�b6"O�J�_�։*��Qw<�	6"O$i�%��F��EP%�_z��9b"O���G�ES����Q⇴��p��"O>�i�-p��B%!�&�\,!B"O���	C+T.4�B�B���"O��{���-���	�4�4"O6e�A��/)��� i�)v��i"O,�"�X)Q�"�j�@�V`�}ف"O���U"�?xn�"CЪ@M��"Oz��$�p�{�A��ELTj"O����^_l|���A+�D��"OfB ÑY4(����2�L�*"O�D�2(N������V�c$�D"OźG$*���cŢU�
Ɂ�"O�P���.��r���#����R"O�T��F�[��eo�
�*�i�"O����o�����,Y�GiR�R"O.�Sꅨ\��:2&,� y�"O~	�k���`g
�=I���$"O@��#�(Z�1�oOI/h�[�"O���O��ߦ��!̂"O ����%}����)�xZ��"OJ��a�5!���S�ڒ3��*�"O�aҋʌ&2�|)��\81��DP"O `S'�ON�ց�#��{\,�%"O"P���z��B���(6G���5"O�4�DJ]5F��I�
mE�� �"O|���]O�D��&e�;1�H	A"O,eA�N�n�V` �c���t#�"O�E L�G��]�UD�+�n��w"O&$�Z�k��q����=����"O��1&/��#�p��6�u�t�"O����hQ>$����L����*O�����N9S&Y��L�^S����'��%qs�Q!����
���P��'tZ
&(�`�ܒ�K��lX%�'�|H: S(u�b�I�ƀ2x1�'?8@���������^p�Aj�'�$�J�М�Qh^-$F�-��'�0�� ��@�1��L!G�e�
�'v�\xV���� aS
͎bS.�	�'B��%��xQ�gΈ1c�<�'f(�'�ļaeT@���+,��'� (rP_��n��Q�Y�$Ҕ{�'�@��@��KHP�s��I�%�u �'�e1�
B�_B�8�*�R@.B��� Ta�2K�'RR�D�v�%8��ͨ"Ov9Q��Y��I���ןU�0�7"O6�J����HyU��&f�~!kT"O�%s���%C���󤗎��m1�"O\4j@c��h��47DJ7qlA�"ORt�4<X�D8w�]C�]��"O"\���T�'��3� \(kB����"O�x���ߕQn��O2�$�0"O8p	FQ'y���Nϳ�4��"O"��©=x&���r�	��B��C"Oj�3�&���)AÆ�7m�$�!�}Кz��UHaH���
_3�!�D}�vt�vÇ�e�j\����,�!��L�b�c�T�A�A	�"Hw!�V���k��gd^L�6�V&T!�$�%�m��K�cr�3���K<!���>UP�AN1c~�z!̅�9!��tN���o�K�bA�v�W�1�!�$_1(��i4����� �AM�!�D��p}jVǒ�US
�5]�3}!�dUK�>�sE��yMXuڗ%�5W!�$��D[�Ԛ�%vA��b�Î�<�!��	9VH�5�Ì�N6h��p)3`~!�D�%f��!\%q+:	�f���b�!���	�,�i�jݑ=0���$�%Sw!���&(��Pm]3� �C�a>ʜ�ȓD� �$�\�BZ$�v/�TS�t��3u8��tDR1F�������#5U� �ȓ(�d"D��bQjY�V(BPrm�ȓf{�(����]�`�K���(&\�ȓ䰘"#DB.�"��0F����!h�,G�8-��bT):SV%�ȓr+`)*�|�	�&��(d����ȓ$̃�b�5y�>�0�U�z�݅�Pl��8� ��*H���B� <f@��XF4e�F�S�h�(��"�/z��͆ȓ87�Z�hmpp60}ʌ��F�k�<�PQ�@1�P/�@��f�<��J%�����J�i������G�<�
�w[�kր1z�D��RG�<�*�<JR4˥$�/�!�&��~�<Ⴌ�!0��F ��)�"�ѯ�a�<A�'�9j#"A�H��BDu�<�#�����dK]Rt�MRǊ�p�<a����𔛓�L�$$E�e�
m�<A�LD;
q��b�� sld�ZU*Kg�<�w���#����"�
 Fd0�c�Z�<)��F��y�1�U?�.�M�<IC��'�$m� �;q�<�@G�<q�*B��aa�a�.<��l#`oOz�<��$(��&@�!#
�����q�<y�"�R,qG.�%��g�<Q&J@����ӯȺo.0���`�<�GB���	2ā 7�f�b�M�X�<���!c��G� X�f<��O�<a�G�6R h� +�+�^e��LM�<qL� 7��ʑG]8`�e���J�<�`jN�\њ���4oRV���}�<�b���lt{�-�6�@D0��{�<�Vʽ7���ɼ<�����
p�<Hı;_�Q���X)�L��Ag@v�<a�œ9N;(4:�Xv�|���G�<1"�A������/�!��-����<����rf
��	)����3�l���S�? X99p%�y8j�80\��b�"O��C�Jep\H��%���F�J�"O��p#��E<TJ���F�L��"O�Т�Ͱpj���viO�~b��"O8;�+����k��+8j,I��'90�Bgw��s��&xn
�'��8Ć"F�Ҕ���Jk��,�	�'얕A,^�& ���p*\���
�'U�X!�)(d���?��]�	�'� �J����6�hy�����	�'YVj!!��O�ZسG�ؗ]j`I�'�) �@�"N�#7&߂��M��'��5��gӲ@�>���8�����'����u�׮T�2LpV��1*x�Q�'X����K��ot<(�Ղה'�`p��'��E��)d�����*��o����'c\M(cN�&���xV&P�PP�<��' ����� /6���r&kRD��}��'[>���J�V�R$��;�!B	�'�aH�	ȁ)�f*%��!�D�X�<��	�XG���f�&)O|� ��v�<�e�PIA����9n��B��o�<�q�ʡtw�m�� Y�]��H��*B�<!�
O#]*�s��߁-�r�y�<��澄bR�H=K����� @�<���@c�	�Dյv����S��~�<�ԭ��G��UHw/�Xt����{�<Y&b��Ix�A�c��oR��� g�z�<	f�F?M�����ED�X����.t�<��b��~�A �^�(3��Bq�<�ะX2�A%VX��C*�+P`�ȓ~��� Km�tXk�"��9�ȓE$��8�M��<�����!S'���/�2aJRǜ�g�vܲ����e�����N 4�I��ߊ��:���1�^���5�	�n�78�:�.�x�[F�R�<�s�-kl������ Z&�����F�<��KՆR:�"�̡A��͙p�A�<��͂�o��i�r�4\�
u)�	�V�<7a8`~��Y�!�YBvYt��R�<���`�杀&l��/T�j�N�<���C<k��x��	RNh� "�N�<y�C��N��d���C#vh��"Uo�<��AD;�
H�F�VAX�d�F�j�<�a*и-^A`u�Bu�<0���Dg�<���0~1E(˅�)(�`@�ΜW�<�������s'i��Xq�Q 0f�V�<�"dZ�$ `!*�ER���'j�<�ca[�Y,⬐Qg�#��36N^O�<٧$��
5�z��ڑl�Ak��J�<��愫b̸���~�j��F�}�<��ŕ�)	t�2�I�H�d!��Dz�<I��]23���b!�I �����L�<!b 7=Й�2�=ٌ��#�XE�<�dc�0l��C����)�D$K�<�V�O"@@��s�-p +�,�o�<a��O�)M��!�� O���sGHG�<*�2;��1p���X��Հ�m�D�<E��0�t�c�h͓J�FM��}�<��&]�VH�3¬��0iQ�x�<�%�@P%���&`�@cRw�<���>a�|Ȃ��t��t��OI~�<!��C�A8p�"��X�8!fh�R�<�2E#^�iX�&�	�r�����c�<� X�x��WdL��P��k�Pْ�"O�	��^�Viq%��1@����v"O�UWL�9o<H�P����T궅�b"OX8�b�>��8C�]�-���"O:���:�bx���((���U"OD���l��G����� h��R"O~XREꏋ]�(�� �|���"O49�!��TN������e��;$"O��BUͰ1ޘ���(#>���&"OH��p�;6���4&S�K����"O��R4�&����D�,�ʴ�r"OF�I'��G~W̳MA`� ��r�<�$�Z�0.<	� ���X�"�g�p�<!�)�	n��J0a	 Z��#�B�t�<K@�oJp�;!^8t�ޭ;�&J{�<y ��S����8V�DHT@�<I��2j�ⱚQ��9q��3�Gy�<��B�$�p-���ʩce�JL�<1Ѯ�j�H�j3hں*Y�q�M�c�<Q�&�\��( �H3
�|D���b�<���o!����-9K�b�EB�<!g�:R�
�� )�G�9b�PA�<�͜E�8`b�	�u��� @I�<qTE��B��s�tUv��,LC�<�W`E�7�\=�F�'r+<<�3e�{�<��զ5e:E�K e����5��y�<iP��=�q����[Z�]y3iO�<�g�֎lsb��� �_��m3aJa�<CKxQ�d��I��R���e�h�<y�D��PiRp�N?d�Px�� d�<�s�� %8E��䐎}�� զGe�<ٵ�� C����� g� ��AF�<yQ'̤,���^1$T��1gϕx�<�F	�Z�N��H�-[�d;��Y�<)#��$;4L�"Z�d�����W�<�fW�fz؁�喝�> ab��R�<����8PwF8���0-cTBAOGO�<�v,�e*�pE�% ��Q�J�<r�'��P�e��I|j��*�A�<�u%?�hX�#)�$.��倴��c�<��d��=6����=}��'l\�<)3��*J�H9
`�.>��)�#��<)�#Dx~�0�	���cC��|�<�udT"~��Mt�O$tp���Dx�<�q���p�<!�A,��]����P��r�<�BO�>;������!7�X�1ы�S�<	#�Q�{kR}�!�I�ή����G�<��f�1��I����1'BU���DG�<1aȠ\���3M�c����o�B�<irhҳ*�DJ� �m�b%��"�B�<�w�8X�8a�
�w���A{�<�c���mSZ��ci�T=�l��M�<Q6mزY4p�C�	�
5& �s �O�<�q⍠�	��M� K�� b��M�<��M��ru��A�-嬬P�%�A�<���NF��@�х(�|�K��b�<!B-'Y�X�"㗬X�T��r�<A����PK���+q�@��C�s�<)�c3(14h��YG;��� y�<�1�fJ=��fĎaF<}� l�r�<q$gN:*��(�FN
t��;�nQV�<�C'ΓD&�A*�S�Jy�Ư�N�<i�/;Rl��s+��w�V���K�J�<ak�tǚus(�->S�h�uNQ�<� ��EC@�A�lQ�w�����{�"O��k�+	�
[�`�vH�4[�����"O�ԫ��6p�T�0g�"���"O��C���h�.����<��y3"O��Ia�9��ƅ�k����"O��8��7	�p���2��D07"O �Y���;]��0�Ҁ%q���q"O���#�J0��uJ!]\��JQ"O�y �IR�p� 9AD/B=>d���e"O$h㵤]�P�2��ؐM��g"Oh�;�D<J�����1:/��g"O�`���=ԈF͚+,� (�"O����\���%�`#@u�"Op=�GKp���R`�5>(� a"Ol���7���0*��.�x�"O���*�)C&���	�"OnH��D�2�1I�"�*^`�i2"O��DfYz$�e�ЦqI�K�"O�r��M=��]k"��1c:�@��"O �k�&�m�c���@44�y�"O�k'×�F,*8�&�C�J2�A"O��Q�#V�@�Ƙ��.@6q�i�"O͐�)fnR�+4�E�S�Z��#"O2�k�c�J>٘��<6h���"O�[�lC�٨as�k�+����"O��Zf�"rQ�ř0*KX*LI�"OB����0�p�g�\<�F"O�0;���?}���#�5��X#�"O�b��� z���x����F�����"O\���[�b�x�:X��-@�"O,��WWD��"��� \���"O�d@�NE2=��x���6�䅓�"O���#h�R�d��U�޵τi�q"O6�T��C�$�h�	ͮ~�@LH�"O�Q�u���bT`� �"��F�4"O�d��T)��]���25�´zw"O����	+n����`�.�:0�B"O"�� �غ+�`E���[�XZ
 �"OX���MX��`�S�A�%o�})1"O���L�'' e	�o^R� �"O��vE�%H�ԡ��+���r�@"OF���㝣A'h쩵��%'��G��y�A�}I���I?p��,�y���*HO�H��
9sy�@k�"&�yb���$���(Ֆqx꥓"��!�y�(�x�0�֋i|�R�=�y����9jD���GYm^,%9��J.�y�G��7�$�s����f�= ���y�"M9y�)C��"c�T�Y2��yK/?�\r#L�-N�|��NH��yJW���pfB ����A ��y���K�bXZ���K�@ѯC��yҪG�?���81��#ZxL��ɱ�yR퀜7O��@6`��|�Е�׮ܦ�yrd�.ƅ��GD�y]�������y� Y k��!cD��+u@Ȝ[�c	��y"�I�3&x�AFAT4rG�i#$��
�yBE�
M�4�7 ��iR~�pgD��y�!�K�,y9�߷gא���l֥�y2��~��հ��6Y0(�pȘ��y2Ħ26X��4
�P,�8 �ߖ�y�߈s��p�g�]�Bz��ʪ�y⣜�d��T��`
�q��D��yB�!RM��yDM
�,��lK�!�$�y
� 8�����=�j�b�H�BF��"O6��`��l�
��F
=����"O0����=�P���1VƐj�"O�`�֯9�rT�J��Ria�"O�#�����Ip�Y�G��ě�"O ��nT�C?4�1�L���1k�"O�T�PG )vp�őc�L$x�"H��"Od�������� Ű�ڵ d"O¡��/�zl��B�4��"O���FS�T�&��ǍA�
��s�"O�i��,!xE�FF�]�6I�D"Odh1�?.�BlgCϿyb!K�"O��TB�zϲ� P��hk`$Cc"O����E�q�x�R��.�D4�U"O<EY!bZ�!��Q6��6p�djC"O>Ђ��E�3�μS��x؅"O,,���U!2X���k@9$͢��%"O�E;^) l�*���X��(K6(�{�<�sc ET��G-ơ>�r���j�{�<�NS,lĘ�k0�V�2�����y�<��c��M|<���	܃N�I�A��n�<IuL_�{��Ă�K\Ԑ�4��f�<A֫�>3��\�/� ʤCA�c�<�Ł��r�Z5�>*��A+Ë�t�<Q�K��Hx�=RX��ڸ[eg�x�<In��TU�r��~Xj��t�<��ߊ\��Q`�ߠt�&��"�U�<��0��I:�`Β<��
��[K�<YԩV'Y��1 ��G� ]���E�<qF�{�b��'T\LMB��UE�<��+[5��t[��g��"g�f�<9R&ٌQ[�Q�Q��'��ls��_�<)&�*vF�qDʄjJ���5E�X�<���!�fbG"ռP����ύ]�<1 �H?�bh���wr��/�V�<���M9Mf�����W�s)�)!eh�O�<QU�C�)II�P+L�_!�y�jP�<aq�,E�M��IX�<�4�O�<a�L�+E�0�	#FҬ^4&Q�g��G�<A�Hś8��	9'��>9^�P���FB�<��� '4	Y$I��\i���O�s�<���:2��-j#����1
��g�<y�H$
 %�5*�| %���j�<	��%|�=�B̀�]L(� H�^�<�TcP�Tq0B�$W�$�4��N�C�<Y�������Э:Z��B3�SG�<�4,ӧMb�k��D�V���"�MHC�<)fôK��y�2��)�X�dK�@�<)���46��{q�LV�5Ȣ��<	4��<�Bp�<#�R��$G�|�<� O�0q�8d��!l�f(��Fu�<��L�6s�&��@�:b�h��X{�<��6\6��UlZ4�����Ct�<�B3@N��asM	�Lꕻ�Hm�<����/܊�a�dG?=�B��c�<����U�Ey���~����C�I�i�p��,K�9�=ؐa�${�C�I�-	�^Z�p݋�F�[��B�	�}�AK��$A�\UI�ā��jC�	'$���+���,��4��lΩ#�!�D�?����k6@5pP����C�<��AV��G�]#�J3��LE�<	)�p�h0�,>�0���_�+	!�Ȇ`@`�(�j:L�$���0�!�� �����½WԸ��ʖ- �0UB�"O��!vOFp��� b*á<��T��"O�Ȓ��r�����nQ��Q�"O�P�!C�+*<YD`ˌ	�ШAT"O�=)�.z6��q𯈍W�r ��"O�2ȧ|���ɖR��k'"O�`�m�� ��`ٻ&x��14"Otl���B-/J�3�O�2 Y���"O|y⦊2T�֬�0�ƹ*RN�"O(�c&!ʅYX��c�G>pY&"O$1��Bt�0!Өύ. faW"O��Г�PSԖ��5):�*�"O�(;S�*Fd|�wg-d .)!p"O��8�Dǵ"x@ԩD�ŹX�� #"OR�XV�0�^���H�FWRU�<1��ѩM�$�k�KK�I�z�Q�<I�H1�t�����2+�P�<qP

q܌�@�
K�@�5��O�<��	ێs+����ކ"s�)�g�R�<��1N�lB���->t���@K�<Q�╻&@3�l�- ��z�@QG�<Y�ff$9�c,+/8\�G KX�<C�	*D�(8�H�@8�U��V�<Y��T�<�f�VHʲ! �6|����u���f"<8�R�P2KPTh�ȓCKNZuf�75n,a��Ckة�ȓ��T�����2���Igc�XUP��?r��+��	,_��L�T�*�*��ȓ+�N�֧݄6b1ɵˋ�vo4���צQ��C9L�1e�"o8 ���)H���@�N�)	�����9JM�ȓ&����'+�f1���_0*t�E�ȓw4�����X�6�{s��6<��\��j:B+G�_&K��)S1NŞMxl��s$%��jC�J��@��
�/Q�2��P������K��L�H��<�ȓqt���树 �\/:���ȓ:��Eq��[��T��0 O�j��,��D�Pz��	X
����
$I?�C�	�v�(��3F"R�e�l�rB�Ʉ/6��A%F�2=�t�$�]�
ZB�:7�X U�B�@
��cmOJ:B�Ƀ(�ZT�l�0���p�Q2+�ZB�	�D��YbЋ@�(��%cM�0w�C�I�l�����B�tCޠ �!�Yn>C�I< _�aҴj�>셚`�ōY��B�I�54�%� ��ָ� i��C��7j}�ͺ�-L�� ��U�=��C�	�BeQ�W�"ͼ��g(�<r�xC�	�8	y���K���
D��o�vC䉛B,,9!E��~�T�hA"��+6B�I�'�^��G'a�"�8P�o��C�I2s�]s3�¨e��ii(�E��C�Uj��rA����ZO�/i��B�	-V�I�" N
h��(�0�@	��B�ɘR9���Y�b!��Q�^4Ly>C�	]|�h� �>HfXQ� Ά�NZC���^3�^2JN�xz6�ڃ*C�	�V�"��#���:�(YO�B�P�
��b�
T��T(�G*?q�B�#R��l�����ty����x�B�I>s+���TiѢ"�X�B6�Ǧ!�2C䉵B��p��H�z�@�0jǡ�.C�	���Yb��"�*!#�k�#(t�B�)� ���
�� �R&!2zE�#"O�\����P+F�Ή8�x%"O��@�$F3:GZ�Ѣ�*c.�uI"O��Z���&wι��-G�}5@%�A"O��Ҷ�F�j��퉰1ƞe�"O���&���b�82ވ��W"OH�8���7'E�p+�4*@�CQ"O\���j��qJ�)]�l'8���"Ot�I�AEjS1�ŇI�
@�&"O�lH�/�)=���5�	T�D�y&"O��q��}�^)�t�_�e�j�S"O���QH�7�z Gģ(��D��"OL5���>Y���x�K�z�>�a"O��IE�V�q��dQ�H�LHs"O�i�k�6i.�h�B���^�:��1"O���DCQ�'tƭ2f$	�A���h�"O򅈖ٸ=� `�7�&c�f=I7"O�]�a�*�B���������"OLe�6�ì�n��e�X�P8��'�v�Gx��R�GP�N�J��3
��H�<�ȓZE\�Q�.F�0�A�	����Ul�Q��M�T�s�J�"5�c�T��V�O9�̉��"O̬3�拋{��8#E�/?ҒDx2��X���<ap�y���a�d�b��OzX�\Dy���g���22,Bd`�6�E��?��'�nD��H�}5Z�ؠK��f�`��'��Yc��v�F���υ^6L���'�$��A�єg��8�!M؍EE��S�'�`ݒ$��t�v�p���?���'�B�9G�\�1��;ġ��:��	��O��D��F�DA�N֜*x�i{�BO`�'-ўb?�	U��m�B|t�I'��)2Q�(D�D�pH6m�p�PņM"|�Q(E�D#>�M��O>�C�ᇏdm�e)g�M(?�~A��"OF%#�k�	|uRa�U�O.K6 L�"ONEr�
ø>��`2eL�i��t�����#+�t��0�H��۲Z����ੂ;>y0�3�"O�ըUc�_�*�'D�5\&�"�	f?A��Ē��1n�V_Fe�#:�!�䎒;��P��'L&7W�����.����j|�~"�\����i����+���1vdX��y"E��&k��[2�N]RРL&�y��£_> �z�ڣ���'	��(O"�=�O�H��5�^�e��4Jpf�_�XY��'ϸȂ�b�lJ*ѣ�aG�n��'MqO`�|B��/}R�,?pV`YV"��9�J`
G��
�y��@��t�Ɏ�0���6g�4��D;�O|`�r��+M��b&�1:@U"���W�O�R�EJ�h9��	�T�l�9��$6<Od�`�`��	@m.#A"O����D�1G� 0,���m8�"O�h�"�@75L��Ŋ�%�}���'�X)'��XĀ�l>��IӬ�z��E���5��nZ���!��^`Py'�D@C�	�-wp��(�'BH���S�4 ���5?��Ūx�NQJg��~��h�\�<	V���L�6=s��;,��P�ȖY�'U�ڥ�ޓ� �V�4R��հa��p�<AI�('�
$�t��X=f�(d�K�D{����`���L�L�b� �:YF�C©fӨ�<�O����ǒ2�! h^ _^�YxC#�>y��6W桂cHO�#���ЃW�6��G|b��aI,L���� �L�#��o�c���IU����Ńm��Z��A�u�LC�c	+�!�� 9Bшܕi| tIB'ȧ98���]���ɇ
���*��)c�<K��Hƴ���%�I�:����)��N��ee�����O���$I�8�hx���Y��!�.˳N��O��=%>�(�j@�R��!t��L��(9�0D�Sv�&oּ�0��F�<��>)M>�B�>9�������D%$fNt�WlX�<�ET�s��a�۷-���jSmDצ]��-��}�.�2q�Nɻ�B�c&���!B��0?�*OT�ʐ����'��jzP	Y6O$���� V�)ʭU�l�h1��0|b�'5Wr�*s(�	ݚ-3e�bX�T���$�L�����iC�P>��!mň0{���C8��'�џ U��F�Yp��U�o�r)���.�DT`���O� �ѧeۺPl���CI�T̼�
�'q���$J'�|�"T�Pۖ�'�	ɟ�Ґ~�'��b��͓�KK�,��	�,+q��H��'���AN��B�� HN֤r�"~  I��D�?�����"+K�#�ݻӪJ=VԨh����(O��Fz*���@��Y���bh�]���a�z�L��TX�Ȩ0�ۛ	�UQ�N��@���鄌d��"~��,R�E��(ՏV�������=J�B�I��n�B�˦��`���A:f��C�ɛX����C�ֆo�({�K�2�B�I�A�b�B���1�`Xp@��X��KL�,���^�pk~�`�Ը��̄�	z}�"�:= H���	()�$�Z��A
�y��&W��(8B�D�M�,������(�S�O���Yǉ�:��	Q�Ɨ0 >Y�	�'�b����.1ݠ����"iR���'a�P�V�܍lv�$�Я��	#�]!ش�Pxl�zEP�h��@������-�-��d�<)�-��m*%��C ��WER(O�� ��PB����oX��u��AY����_Iܓ�?E��'�B���Їl,����ҰZ�v���'}0u��)
1�u�G��*<ͼt�'��]�d׶E �1��_�����4\9ꓽy��O����w�SJ��R\����'����%���芸v/�:��ÄFp��ծ&�	a�����I�ON�3&��qP6��),O��<Q,H#}G\Y�	�F��qb�LL?�J<���?Q��ǆ(�$t�PᛳG~�US�"D���@BŊ�r!�2s5l�#4L�]_B��&?����ʜ�Ny��PfV:S��"<!��?�g��3@�d�!UՋl����%�� �y�H ���WI�3uR����(�y"�O90"}�������"����=ѨO����@��@�ƌ.';��7�׫
��4m�E(<a��5&���GnN8���(1jQ8��&����\� ����:6�q�F%D��c���?��E���?4(���4�&D���A��E��$Qs��m��tC�)D�РG�لc�,�1��vE����hӬC�I�<f�*��-a)�_m�8���q�86m��r��u�(3`�)���6):!�$X�)�B�*��	aM���p���H�!���,<�x]3����b+����Z.(!�$*P�9��Ǐ+h���j�+%!����l��gԡZ�z�b߫<^���ȓ"���%o�,.@#�+Z����ȓ��%Ze��X@Q8S��P����!�Đs �>}��- �ܞFJ�͓��';a����C����rꕮ*�
13`F	��y2��#`�T��Ā-�L$��N��y
� �1�7�L�z9D����]Z��z��/��$�lEBh����3gJ8�%��
/�>���:w`���	v
���$��h��>��}�BF��uW��L^�C����.�9m���ȔN�B�	:'f",���;U��Ԡ4K�Z�xB��f�c�ɪB�홒!Ŕ)�C��Z�>�9�
�"QZ���%�.Z�vC��+9�a c��5d>n�
ŧC�6�"B�	|���㡮L?}eb����@�C�bO~`�V*Ӈ2�BPCO�0uc�B䉥.�	C"׆Y�0P"�`�%Q��B�	4g'�" Aɵ|=���I�;erB�I=}f1�%@�a�U���L�+P6B䉑=?8��I]+�b5¤�/��C�	/\�2|!"�<IrT�:�)�9m
B�	�1�� qN�:%�B��C�d��C�I0�>��vĚ P �*���h��C�	!��I��D�9i�P���<�zC�Z��$�#V���a6��Og�C�	�=�,]�c*��	���ЯV�+�B�	6	���2NO:���p���_�zC�	7� �0'�`�L������.#�B��Jf))��Қ+�,5�4�Z�&�RB�	; �.m��i�;>Fb�XW���BB�I#���D!�.�6\�$�M?�C��:����\�kL�J2�f�C�	�t>�m�oǤ��WDU�ne�ȓC >E�C.zELaX���8W��ȓ'~D�"�G�͒��Ƴ3���ȓ?H����Ǐ�/���Ճ�[�� �ȓ �*��ѣ{���[�V�=%�y��M��(B��
p�i#qKJ�6𾼆ȓ/���á�w$�Q��1����3��S�g��q2���%ȅȓZ2,e�6�T�$J4��,�PN�L��(F����d!4�G��=�����q�rLIՀҚ���7�T~���3 iH���q��N�~24I�ȓ9�F�p �
�@)�W�}�8��>�����Ѣ1�	7�O�H4����2�%�. � x���+F�P�L��鉓;Hjȣ�Ç+Q)֬`��.G �a2�ھm+$l��%B4!ۜB�	3��㱁�N�ެ���t�dB�$\�B�t%�&�TȒ�e��@˴C䉒Z$4�"��p�B���=f��C�I-N'�����D�f�3�n*Y��C�	�+���U~��ćB��B�I����a�̧[�"�׈ �^�B�	1�P\��f�&Ou&�`�+�*�fC�I3'� ���z�:䱠�"T��C�I�]W` �_,�=�VhU j3jC�	�2�8�sPc�g�y+�Я�~C�I	!O�|��ěR&zPS���T�B䉶-H��zDC�"SL5 cB�|�B�0K��U��N�*�@&L��l��B䉵d����tG�&C:8aKB�Π]~B�ɦq`��� L�5�y@��}�RB�)A�dx��)�)��IZ4���\��C�ɉ�,4�A�:o�x�J˙:!�C䉉>�ֵ�S��cڐyhI��C�Y!"%1ĪK`�@�F �dx�C�Ɍ�n(@&�Ϙ8�0) (�Of�B�	ST���Ӣ.X��*��%e�B�)� ،��;�ع`��kǊ��"O���Y�¼#�FLS�|��"O���c�=z�y��Z� $�4�u"ON([�M[{�XQbB�5�p�1"OP�R"<c�@`P�]�Vpju"O\��h���p�e�
H����`���yҥ$:� �g�E�KU����HE��yb�D/c D���ڮ�2'�Է�y�!!`�����:���8�K��y�E^5H�"qѵa�;�P�qj��ybn��#�����-+��-S#$3�B1*�
=��F��~"*F�?^��v�8����*L�y�]0c�iR$�Ж�ja`��S�^��Cf\�Daeq	���b�e˵9�\(�� �k���F2�]�,���j�`�i�k�~�p@����	o̱�fȍ�5=s�I��Pxh��?�����lR������LH��~BN�g��x�%�V�eE��9���\���JviG�';}	�%N�l�8T��� �a���ȓlp��%��C¦�x�+	��\����\�\�
t�ʋ6���K�y�djr1i�P�TQ#	��Q�rX���5������0�O©ҀDД6�n�q6l Uv�d�cE �L��Aq�&��e���	:Q��i�#lʰEҮA0��0	�gņv��	fAЂ�hO�K0��76DR�a1��-?N�qX4 _� 	������X� r ٲn���ɓ9�$��I�j�H}C7��6	hѱ�֥B^7��m�Hq����$2���h� 	�2��v��k*��#-K���|�F� � &8�jQ�˻3��I6"Oڐ`t�ɇj����� ]����%L�Az�T�1�W�=	�5(L#^Wܘpd��hd��� B�l��ռ�A+W��5�5̂��2L��WX�l��e*�8��@�<�DP��C9x|��H�$B�'��� j�"�.��g��qA2�YB �>�^,82�D�3j蛧l�;a�UmN�f��0;I>�u-��f��$s!�=~���S& �_���:&�L���� ����U��!�#�h�ڴNH����	$x���	�8L
7� �VY2� �>�@)�n�s��P���⥋^�<�;gj(8�J�l6M���4P"g�ϱ\��� �b��R�P�ѦjC,^�ax�F d�����7T剩{ᚘ#'�C�)d`� ӎA������H;t�&��R&�
�6� �Kث甄g+�*lr=��nRE����'n��� _k��s�/���PX0�O43_O��� ��	��V��q!�EGg��mDڜ��J����O�8#���d�1�:T��̌Ey�d��ٓoBԀ)�E�Q��C�ϊ6����2��!fL����%^�?&��̓/DD$2v�Y�����Έ2����2��"dJ������Z�6���3���dLYS��lB9�"�i�l �N�0���W1
kT��"�;,r8�ƅ��^>�[w&�-g䱳�ǁ�jY����cN1ue\���޺)}(�FE�.Y3�0;Wf�8(m��!a&�	G�z�s�MF�H}(!P��I�%m��)qfma�*V81�|���'R�'k�6�L)4t���W�aV�%p ��%����AcG (�v)vX��`���ɫ9v0�"�Vd\�@p �$ㄐ��G<%� ����E�# �hp�K��p�C�i��M�^L�Q��ͮܪ�·�&�
�ٴ��$&�8�
,�f�k�i�Ȍ��	V%I��i�&H5E@F���ba��b�tc�DE�̆	���V�M�qO2�!���Zn��0�*I�YÃ�v6v)�ՁE�$��dۦd;,�IGcW�|� ���,G�eb�c�v6N\���c1�0�'b_a@@x@e�"K5�1)����'M��0�_	~R�!u�a�6�@�L��$	c�	2n�԰����^l�d
J�1����.��	� U��FK��i��i���1!�-��@��9^�+R��LD�q������'�>Ix�k�9p ��
ܑCǲ}b��R����#�U�(P�Ǉ�b��`�7.��=�0��Cz|,�yֈ	~���X ��hE�B~t<�A�HI|���hPCJ�U�"H���5N��q�"��<k��:cb]�=��t��(�`��!7.ȕ�c�J7J��}�	ֽh��%b���|�S�	�:��a���=�]��	(?����c�ߵ9�.Q����$:�v���?��U��"�Qf:.��2̎, ҲMY��ݴA��9�c)*���R��[F	�yc�����i�5iY
8�m�)Gw�aR�ll<j8rw&�~B���&Tɢ����F#ve�#<y��?Z��iU��+I��I3��Zf��� ƫI�$�T͛!�L�z�Vg3+0��jb�	7R�t�R��<mu�!�RC��"�Lk%��3���&���kpA`2�F�Le�d����!�1O�h��ŗ�'�6-�օ$@l��4�^Rt�JB� h�p0�/�c>6�U��$g�H����+��:��4 5�ʠtY���p,�>V�h����P��j��I�M�3��A`�>�S��X�>)\43A��b��	�Aù'��Q���2Ih^wCx�n�|
�@�)��0"�A��Z��5�e��%'��R�ϡV*�u	�[��pa"�>/��Fx��)x�8-�p�
�  A @گu�����S���� �B���rǜ?���߆$H󅮙"R��03a$�"n�Eb�`�%A��m�Ao1N�5�fa]�w⟨���A�O�����`(��P��R�]�jl�4�]9z���!S>=���ƖN�Ʃ�W!#w�*�(b�S�\�tT��i��2���!S<]x�	<,X��ɇ���F�̵��/��#V�V:U��xO�u����<9�B5U!Uy(�ɇ$��_VL��L�,~��8��	'P
����)�h���[���x�1% �!Y�*�aK_:j6Z�r��ּӦ��Z�bH��+;"8�!UnM�n�Z��
��i���c�R�W�����T[��S'8�ġa2�+P2=	Q�<SV$�&a�7%0	�bœ���X��#m��)�ғ*](Y��I8T\4�=R��w:����ϧ8S�i���ϑ$��=g��J��X�C��J��$9*^ v6���j�8\�]�D�N%��	���ɲB��h9r�D X�V�JG�յ)%�KlM�&.^�UH5�ɓ* �z
�T��m��9� �B�MH���	��
 ]�؀�M��ז��'��4�o@��-���~ҥ��{ x`�v�QjA 9x ˍ�@L��"�$��F�Tj�y�D�E�@)椑����Zt�ۮ4FV�Pd)aʣ�R.�Hs	ƕ99V�9`���8�$�ʀ��3�hX���������`	G�?4H�YЁɪ<�.��1 ɣ!`��$�H��j���5A�c>f<bm@�x��ղ!/x>ͳ G%�D��_.��59�)��*�]{P�O�ˆ�B`GK��zɲ�дA�̠a�	�|�``	�)�QS �.�IPMh\���	q܆Y釀_;����<Bj�Hw����@�
�VBlT���	pҚQ�7 8	��Pe��>p0����K�x�\�A�["lv �C'���Ơ�ȗ/ ��'QB��g�K�E�s���
l\�y���lo$-�m���>�4&T0�,͠Vf�n��Lʷ.S�MaB�i��S�hg6ᆍN�x� )���3�d�DjO+�j[ ��E��8i�{� �#b`��|ߟS���� �o���Y��U�u�r��P��� $�5�KW�atȥ��BW�x�P�Z��p�V�\�|%j��X)����d�-Y���a箞�_�$�)�i])̦iC�oI�9��ͺ`�ډj���76��di�H1Ը��ݨȮ}{SO��8q3M��M�h�#��i�#9'Xe���l�Lu����W9h�3��Դ�`�����5%��Q���x�/n�{R��"\{��n
�b ӂ�_9"YD҅�8%��Sv 0*g�KB�E�Zv �S�.�>gt�b~!���7�(3��Ÿ
��	�㇕�x�N`Ca��0�V��p�9
������y�Nd�H��N@�g��94H���X���Y`��{�F��c�-��Pp(_��JL��V�f�0a�e'0��CD�l�ZG������+K:Q����C��CE��E�e��Y�cMT'1p * 	nɚqy�:^���]�D%@�6e˲�x���L�J��'ʷVVL;l��a&����E,D{�hC� E4V;ڔBŰf>@S�J�s�0�'�R9 $�C��$(��!5B� �J�Bw.hrꟁu�Bc!�2�>!�f�ݿ�e���+|檜a���0o(���0g��������3�(۶�\=r�Pi`��	��J�'�)Z�ޔ,p���d��l#2��!��m1�b�
��cƊη#�" � )r�ٗdY�F
,��rj��6����){E�UQ��B���O.���M�L���32��Jz`Y�)����u�Q�	�@��mQ$�u���1�O����T�^�Bnta���
�K'�Ƭ$(a�GœUaBU�#�5Pb���$a�"����?�t���̘���¬k��@;GI�MN⭃'*�)Hh�����Z��]�v��%��0)�@�,�EI$j^T"1�K�ff�� A�^��q�&%���� q&�'8�S��ȩt���sF%�$Ty����CйfӞ�
'(:eW�@b�G٩]2�6��v���K�E�Ws����c�9a6�`����1P�,�*�"�D������,�|9Su�S�7$�E�A�]?�H�R��]{��ত_8�4�b�%�,%�5͊jF���E�΁(4�x���^}Ό�DN^:�0��c �6�9j���pV�಄�Қ)���"�Z�"xG�ɥ5�� �c���7�ݙU1�l��L3ʶ�q�F�4�НiUÎ4YO�0@c�
fl�]�o��T1�X���4Ġ�Q���ؑq�㏜2��I��AM�)����(\*��'m�=2��9�xj�%�7���R&�!w�T̸S̮bp��達Y�h�����Y @���F��X�U��7��-���ct�ѩ��u���>h�h��UV����3>�����65�|�9 e�K����\.�yk��XL��T߲?���9��#��[B���$��h�I�G��;G���$�3MD �V(P$7��S�;�-]��H����l_ [�lY7]G�D�R�Z�cR�H٦�QǆU����ź���Y�4^�m!��U�g�p����n-tTydnY#F�!y3$�Y��u�F �G�ay����=���/��e`���3���R4�&(j�i	�%�s��Mz�έAlr`�B�\�&V``�.�%6������+o�a��� ��aB9%��,W��Ic���ղvז��3BA��iU`�r�H	+��X8</
��3&
���]���ʀ7�� ����8n���!+�Z�@SML�b�K~j-�3���_cڽ�c�T�^��ొ�u�X��E�ܹ>�ZͰ�O��(x'MT�Ziʗ�z��O�Z��EF6yk|����";�J ��)�>PL�gf�|�X�cnē[�~���A�t�'��B�Ú�Z��(A�j]nA���g��,b4������a��hN�����d:�ͳ�Je��N�bf��s+X�E�T���I�t�c2���ea�k�%�<��Z���H��9 ����81�o��=#6��Ac�8uV�kS� !n�H���"��<���'93	$���E���)S-sne�Gĉ?�ܰ;Q�ǝ�Q��选�,wvQ����:�̔k�,�
�"�W��&�r`�-D�;�^�a�� �k�B�!�-�r�VH�3�D����֨5�������'��)���VD�*�Q�GF2\���4$R�J#�>��� C :|9��Q�2�.��k�%�#L_�A��f,T��:^%�tр%�}��)sԨ;���RK֌Z�(�>��g��P5S�+Q�ߎ��Ћ�lxF�+�!T�t���AmY�
�H�̧\��ޘт0�U�irH���}[r�Rd�@�&yx��Ԁ�@]�e'<Oz�҄`��TuY�H�0l,�H��WC
���VQ�:�v�6�-��A��`�95��k:�(� ��uw�?q����t4-�̅�5�.��@�)ړ'_6�!\IC K��M4	i>�K򥓏"���@�Eu"����g�+�T(�i���R����	t��b��  �����D[��_+�nۋ-y1A� <��`�-�-2\�'�F	��H�ÞS���,{5�r���!R�I�4)6X6V�u�Y%�D+B%��M�V+��Zuk�KD�jF�(�$)���'�dq��
�Dֈ���͍<]��8P��f���Ct�,����L� #�`͓EՈ�-��_���@c�����;4 fhf��d���p��!2	��kS�� g��>I�����	��4rv�X������aO�.-5.X��[:?o��qU[,���R�7����s� #创�����2C�4�������Ng�XEA�`��Z��C�'FTx�E@&1k��BB��2C�
�'"\�|9C��9.�r�	r+�Pl�.Bn,H�'�W�(��.DL���2DF 0pH(��S,�R��s�urj�/|ޱ�r*�2+h�tBZ �P���ݚ,�.S�ǃL#��>�Hqc���4	�I�h��%�t�O9c�t�
¨Z�k*��-a��H����Q1l1	�m˷I�L{\w�(��L4�I?4����l�1� ��A9AFT�`�
�.X"�"��;$$ž<��� $0�47���s�����`+	tx0���dX��Q�K8�8�2@��w��X��>P��Gx�Cʖr1X! ��<��j�q���UB[�̞͉�N r�����-],�IR����8��	�A�}����B�'����SNa��"� H������dY�,Ǫ*��=r��	?Fkұz���4->�����ħ;ՠx�'��i���Z��(9>��S-
�}����٨�2�=ٴ<H�灻m�:�A��,?4��;(��Y��vi�%	�O�j��BAۙtN�	G�ݐt��h��Şq��x�v�.���s�̭p}��G�;ؘ��?k��rg@Q+Yxl����~�f�q u���GF�}D~�I/��)\b�����Lh������e�b���~%@����_
yNf�!�۴)Qp���4R���o�~�hڴ��'D⺸A5����	� L�N�U��
�P[�<��	17�O6�,�㥌�	=|���"Ɣ@EX��[�8� p�Fz td)pđ�$�2��:r�����Imr-�X�6��GØ}�d���VZ"�( �%�z�'��0i�� �p���A,!��O=2��qȊ50B� 
$0.X���3O�@�dɣwHl8[BD_5"��!�J43J�(R�D��&T���w�p}*��F�m�h:�ǅ�>�`$ �M�& 8x��V!̤7~V�����OxX��	 '�dYj��T�]d� �)Z�5(�i����{H��Ձ�p���H�"]6+�%	�GT�\�	�Hܓ#�N\��� +;�N�
��-f��]P�i�V��p�0�Go/>�����D,l��8�l+Q!��r���B3�+
��u��n^)?x@\;w�
�6Ɣ��0hw�'�活
ϟ��f��4'�����vV��� Àl���j#������IWE
~?�ů�~�#�]�)��9� �O��a/f
 �5��u��9�鉁��1d�1���}�D*R!B��Ɋ@f[��J�D�`}��0�P)�@h�&�U*�DM���dbʙ���:��
�O��@�D���?!��-�����)-}��$i�8vJ@!sL)$p0jQ��eBb��2�Đ��nR��9S�Jc��%��l��ѦOf%
`G
��~2��2����=��J������-zS�4�A��m\C�	$O��(Z��N9q0�x	EW�L~\B�	*���#�%Ⱦy@��p�k�* |B�	�e|�����De���Q�!��;�l��T�[M��,K�Y�!�d�֬T��]�U1��3t`Y.{�!��%)��g��G<f0a��#&$!���s����T6I+��Y ��=#!�D�$P�,�ˤ���"#|m�6�+Q�!�P2M�Xy;Xh���'��H`G"O8����SH�`�F�ά�&MRs"O��i���W����pf]�;�,q"O�L(�%�+=}N��`��H�,�"OF ��05.l��e�q@�%"O�4ڵ*
���x��J-r� i�"O,�����Pr���0d����"O,��B�j�b(ʤ�1&P���"O�a���K�w�����;O�S"O�)��%h���iןp,���"O6m����$�&y�C�\�o�P1�F"O�i��7I�R"�3
�X��"O �)"���r/(eK��X�NY�M"O��z�0@�5+�9\�P�A"Oh\Q��eRV���OGa�QI&"O����!_��}��]�LW0��u"OL���蟕C,�b'ۘ .`�Z�"O�9��(�3�|H�Ҧܼa�fh��"O�U�ԭ����� ��|���#"O���Ȯl�Nu�qm����] �"O� �I:j/B�Xa,��|0�#�"O؄H,?P  �5�ۋ`�xh�F"Op4�%n��/ \�(J\�u�f�X"OD��/�w�ȋ�d��Ωw"O�L�E獱\ T�J��P�C*<���"O�#� ��P�>�"��<���6"O�iˆhϺ+2d��S�C��2"O�mrSH��~��h��K�#^0��"OT5��ɐ*<S4�H�Eڵ<8p�:p"O�ZQ��@�z][`��U�<�P�"O�E-P�r�r��D�E��"O�<�ԏ��Knt@ ��sfy:�"O:m��)�Y2��bA�5�"Of͋e ��f�x���fX�eG`�f"Oڙ��(ܯ7΁q���&(>$�E"O e sL�V}.y��	�cr���"O� ܜ9����b@v��l ��"O�h2F�Л0��9�2��4��\P"O|Y�����!�l��Q�cAR�	B"OJ�)ÆJ!Z
D�ɥF�?Jn��2"O�����	X�m�7�� Azhrb"OƹH���%�:��­k DI��"O�xK��O���L*�n�a�sV"Ov�Q�[���j�������"O�q26�6�NŚ��3k��1�q"O@��t�@�E�@��$��hTh"OUv�����	�V���"O�J�ǆs>&=1�nŴH�$�R"Od���&#J��Z��+���`@"Oj����#l�%�Tk �:D�"O�<+Q�-[F�����O��PdcH��"��=����O��Rs�P0�(D�Ѝ_	e���$"O��@���~�@�m߈�␢r爹 V�=A!�e�a|-)fd���D64�J@�,
���O��	c Ϋ�� %�]�*o�L[g�Y�Cv���ίTvdD��.ǂ.Ef�+t
O���aK�i�sC��1Z�(��O�@�'h�QB䠱j��^�����͵x��������N�1j��C��<	@�8���y��O�P��ؙ�	��x�MЖB��K���J'��c��A�u̟@4���
���X�Q*É^��ȓ�:*�\���I:+�T�aPk@��h�{1kE �ֈ;�n�����oV?�BlI ���V��I1�����O@���ܔ,�DXy���/qh�U���ɇQ���c�%
4Q�QkE�ݘn��]`�o
?2�n���G_jz���� ��V��C����?�am[�v p!��͊�`,y`�K��i����/@sԙ	C� �H�փ۴;��:dG�;`�H��n>�شd�@Ļ�N���X���5v/^C�	}zz�� ��Fɨ�@"BnA�W�y�=:�,� />�`P��|xx��q���C
7�i�wް�������	Xc˚�{W����d��$�7�Z5Y|� ��R7a���*v�'cO�ȲGI�d�0Qc�
^�f_TQbV���/� `&��g����P��
��\a�7��,���'��G 	ؘ��φ^jX��@
�L�x� !�|ҹ�6�Xr�B�� p�¸ء�Fa؜p�D�	�Љ�w��#�r��cߎx��p��L9y��p �IV974��ا��"UظçkI�%�~�;�ߌ�M��$�r�d�����\�f��.��t��l���e�G�t�6�$�wy"�ݶg�a��h��׏�^i)'��,CT��փ�o~�ey�KԖrݐ�bąJ�j4xTؖG��Pט�f��	3Wk��U��[�]E�A(��3?i�K��-��X�Ѐ_���	��nU|�vA@�J��!cΖ�y��@�K	�d�ѯ	01�jE�'
ʗQ��FA��� [��W{��\)k�p�s�<��Ǌ>#T��O�N�VA��:y��ϓ(��Ű��E{� �3ǋ<'S���L�XI�K_+��gn
7����R��z�.���b��}�)���()v
��V
��-�3��,x�a'5v'bi�!A#8fB�1`I��sJACGb��9��ĝ�:h����q*xI�ޡ=lr�����YnV�ES�
'j%G�	2q&v����,Zd˝?.�^I��9:�
��Xj\���O0#N����ck3h@��%[��;�$�N6
5��C�7^ pt�N�2&G�����j7bT�u _>ж��d�.^ ��@�b��v���3��M4D�҅�^1!�ZG��=վ��tC�\'��c��*s��3ӡAeL�;�E�O#jݰ!��&u"=Z�FE=4_>���"K(uw`�C`��,�U�=�C⇇7/��� o?l�f�����;#lP 3"�
�Z��Fn�	k�����B�2,�	տi�|��*Z==.nP�0�ϩ_
�"6Hݹ"�0I E�ƭ���ߩf�ډ�.3���wከ�Ta�(�>Tҳ����(��"�ʮV�=�P�\m�D���C:)���uMP��!�6��6���K�5���"�:hɀC�&[3zq�� �2O��C�H�*A�(K�-˔$$�ڡKS=2�ur�Y0@Ѧ|Y"@,�&�������PKх�ӌX��Ӌnr-`1�	�Q�X��I-S(����� ��|A�Kۜx�-I$����Gi8�3��Wnv 0���޵*n�*4���p�t]�V��2,��}�ҡ��Cn2�#�K�m~�"��|�m^
u;`!v�VM��]��)W���� '��gxi��l�(�t�ҷM߈p6Ty�"�Q�\�`+pc��l�����X����m�73�e�`&�
k�e����g'�Ab�)�!Gzɩ�D=w<�"F� $:���P.�;K��A��> `F"<�7�	Bb(C��,<p�S�c��o�}ʣ��SV��v̍%F?�hP%>�ȕ�E�,l��`Þi�A�C�݊VS��v�M%D:����`�2�ӹ9e��
��+{Q0�<�h�*[��dA4y�6��cf�$�H�ҧ�@!.F`�%#� ��׬/Z�G_9-9� �,Wr��R%@#x��e�5�4�BE�+P ����Y2�f�O�B�Tb�=#� P��P����d���J-�+�I 4<����QK�H�D��6�����V�,@�Fk���ū�;A:q�E
�pK��P��	<^��|�cdS[���	5y(��A谔R�A�27�M��@S1P|��cnJ+fR�0S��u�T�Q�"�jF�4k�
T��@�l;�ݩ�eԏ 1T)Ae�H�N���ƃ�X\@� ��)Gr�"���h���	�AU4��ӽ��	�ɜ�b��h4��>�.�cA�����z���?��S��>��9�i�,c��h d�}.0Y9�($#f���#��'����a� g���C��J���R�[;�$�PL�}`"u�&��X� U#6I�$F~��F�Zc^���J�6e�I�W h,mȅf��Y�(M�.�!Jh%���� b��D���v�E(VO���ƹI�Α`��9�R6�IC�l�`��Ի���U�1����Q.R*Qd��+b� 4Xm����"��"5H<#�t��&�.+�Z�x�M�Wi��{©�[h���)�)��ь�c֎:�`rHɜ#��1"��Y�9|r�(���&���2��׀�g֎2�@��'��M�Er��a�e^)D�J�! ��$_f\�\cq�E���?SgqO��C��+6	:-Y0�
)�J�r(K�D)s��	q&����.V��8ѡ+U40�H�"��mhF�J���~�iŻ�US#j+@FȽ���Ѧ-lXs�� �V���yR��u��D�$�F�1����O���m�0R�~�JhL�i1�	H0Lݞ!s�k�+T�ʘ��Q�l��0��M��S�p��ȍ
e���1N�����<27v����?fN��H��7`��s�G9LB�ԯ��L��d4!�oA�Q�f ���͈�P�,�;��X��N�.8�X� ���͊���K'?��������@�1PL��8�qO̼��4Z���`�#A=�0IC�.�zd�͌36��cK6Ĩ��4Y���p3��|=�,	�aM)�b��)2�P���"D���ѡW�T�*��T�o.h�P�{R�Ŷ�f��U�
�@�����7p������~u�$��1-�a+p��j�>��7 �I�P�9�B�5z���f��zI��*��1/�uPK��"<{"��k�D�[T$���'��=�Ü^��hV�YӟX��# |"��n΋�*M��*�N��ak#��Bބ�
��_�����(�7S�5��̛�*u�e
�J��}+���EҐ�Q��&�Fi�GGR=g�\�*�OV o)V-⑪T�}s(�S&�E��Ѝ+G?V���%xɒ�����@�j�iݜ�!,ܯ@�ę��*@5o�`�	�(?���t)�8x�|��/����3Q윮C�ʅ��{r�٠�d�H�l�B:�=��҂#��: �W"��x0C*"<xҩ���f�X��D1��b�S &��):`�J
�D%׈	G��+gm�3޸ԙ�IU u�f�P��=ʓE��3W٢2ܺ6M��0�Ԍp���~h"���bn�qS��GB́��o⌐�QV5�ʸ`�������Jڻ$�|��%f�$"��τ_��\�͙���DyZ�X�H?�EJ�lǘ�@ԀB��4��/vzM ��l^�(�d@���R��фP[t��ƥA	$G
�h�j�pu}Pu%FoV�p"��D��ݠB�^[n��D�]*\��G�O"�������?ɕb/p����fêZ\`�QT)['p�"���	i4���f̸u���ђd6&�ș��Gdڬ�i�+B�U�)�*�l���p��#<��/da���S`��U
�*&��+�l�P�2�%a`���f
A��B���8+� �P ���]4D����ï'�$!s7(��9��mT�A(_���8���:C��.V����fV�.�T�)�+ʩT�>	�I-j~��Bo����Z��Q������v��[F��+�Bɪ���*"�:���7b"� ���Q�����"
��7�
�I�m�@(��(��SO�T��1�R�A )�"U��N��"�+��*����R�H}������-�ҋ��,�4i�� J��1B0k�O� &↔B5x�E�̈́W��ɀ1HK c%~hiԣ@&]��DhE(\��<P��G@1l�5��R����a��c*���fj����z%)�2(��l���q`a�.S��1q#"[�et����J>�}�h�sd�Y
)j�L:���K�r���G�@������
�F�ꑢ��W�~�d�Ktϙ�)h�D2t_�M�d���>]w�H'��Rw��o�td��'�wF
tE~��P�}�:���.;�|� �e� %i"V�4Lद�s�R��RF�*)c�NhB���(.a<A��3�N`���T�r�T��b�Uvh�".����XT��(D��O�SG
Х:eN���J9v��#P>q�
E��՜b�nuHU�C7*��rJݶ�� rf�ׅQ00h��@�/��msA�"c�l}Xu�÷+�NK�t�Z���' �x@�"ȭa�lAmƊX���zT"�!%��r�L��g�h���K�C-�L2"	,c��_�B���˺_!.a+�EM�h�tU:��5e�������WS�4�ȗ%B��T�q�x�'�p�C�J^`p�n�+P
D��rF� nX�ĥ�%E�@�B%@��u�o	�50u���;U�F!�k
���Dr�'�6TRE��F���c��$����R�&��=�GS�L1S�ڥ.�(��k[�`]d�Q�`j�}҂�S�:���	 �$�X��/�<颓kZ�dZt�AY?��UoB�-v�����(D�X�Г�;�I+ �8���ֿ ��AvJ�>?��:�"�j/v���eL&4����]�(z�Q!KOS�X*S�m[�1��@W�k�D�ĕ�����j��2��Sse[<G��\Rv�?U����=1_��#����cL��uk��4��k#�|ⓝ0g�A�(T�*1��0��z�0�yt�X��T���#[�vT^�7�ӛD���Y@�I�v��0U)��8£��h��sA���:92�,K�'7��1G�?��a�� Ŭ�Zw�dh��&N?{�!Ð5I��� *�j�z��W���6
Q��	�.�X��3��W(vL��ǟ!Q��R�(�#"2�cF�n"d�I����Q�f�Q��=c.�\�VB��!P��zu�!&4��O%�}[�U�h���y�l��T~Yk���5 �]�n�(n���1L*Q hq#Ѣ�6Yuz�'�?z���	Ga��a@�P�r|��G :T&����� X�O,��!Ԇ�_?�D�kQ�}3`�K%Gz��tS�7�(iV�Uk�
�Bp�-�N�5*@���F�_���'.Oꨚ�A�9}�Pe�� �@^���m�3m���7�2M�P4%ܭ}Ԇ!�v�+�.(�8�DH/lH&$��Ѭ�,E��∱XH��ڦ����a̓�|�U��hB.0��kP/�,q�R�0"~֩���#��Z4�<C�@�ABg\���<A�N�	�'݉��
J� ��H�
YO�^(!����
��H R`߈s��Y�t,�� 
 � jˇ&�@_w\���6����?v,�x�JɊZUl�=��*%E34]�Go��#Ԭz���Ljd�P�>�"� ��B�H��`�q�� a��R�v�:$�D�K���5@�W��ӕ.? M{00�P�� Ц,fݫ�	RW����'a�2F<�0� U���s�V� �@�f��aD�P��U��4P�N�91`�KĠ-8�����vj�+<-� )�eР_�K��O�iq�Ы��42��ٜ{�Z1v�\���rPMͣ��ّ8��n[�<����	G���+G�2^椡�7��u`JHJ�`Ǔ>G	��#�>K���pG�%6
|,�S�1�<<V嫄n�t��}9���R���!��E9���X��e��`)�kc=\�ɏT��]�.MV�Р	�#��:���x�Z�e?N��@
I.rǦe�e�ܛ;������,��TՄ׸fߪ��6NM]�$�¡3�� �K�?S��@#H���M3DF��fU���V�a�:3M�@a&5�a(�'}�|Q�p&���1ord�$b�iy�@�v��r���6��C'z����%o]ܠag�Hy�'+f�@\�:4�� �9f/�e�^Yp�*�)`���([�g�64f�U��e��FL#\��)v��S��i̓8=V�	��V2!lҰ��#ۭc�����#��P�j5#�&	O1���	ic��q'U�^ʄ�c�i�f{��M$�TÔo��;�0��*DJЀ�W6I�f,i���^�jt�4�V��
 !��i����Ǭ�����r�W�|�5J(��!舉$�8HM�)Q���P���@ҩ R�f�r�OK�[��.KK2��0qm��ba�ŉ��� !CTY��Tp�@�b�� �M|�"� �>	qO�'s�y�6Y�*��-c������8�>a�,XV��ɐ
0���z͜��p�:2�e�v���S�P�,�@��K#&U<d ��ʾF���)�S�D���b�Uv�.<��kfG��$�(o�)JN|���8ƤO֭���аu�����fF���$=扱HN)CLQ�Y�c��hע�	�1��;Q�ڲP�i�v���MBr��P<P�%o�MҨ7-�B%�M���xFvaI��@8p����Z%O�KT�&���'@O\�'����@�N �y�d�V /��C"�7g�����@�`u!RB�"?ZU#�쁋>]��i\��x�	�Rے1�N�@m��EȬ�l����G�=i��;_^�"<q�k��]�����'P��%rJ~�g����3��Φ*^j��u���yB΁�UU�T�e�8^)�1��n���s��,U~��bѼ��ߌkHK̗M^zy�#�|�@�b��4 "�U�t�V�]4���)��7^4�݉�M�/2�vT3��O�O�~��d#�h
�U83 ѵb��ɔnךH5Vu�����2 I֏�|�D��ӫ	д�ڗ.����K� }��.�~a��ǚ_$� ك	�lR`�ӂo��~bf��O�"H�f�]��	�^#O����ĩ�i��]�E�R��9��I,d�0e�p�$t 9�V�k�,18ԦX�J�v1��F��c�h���*҂@h��$�O�˯��9��4\�8��(B���)�t\	�gF=�4�Dz���#�z��D��;/q�d�CK(*of��R4[�@I�$T�Ti#�����J$*
% 0D��=Ų?)Q�[2LrP���%\�$�O�-�g�1��T:H�b>�10(܎$��yˢI[�M�����'�6ni�S�-�!���(��`���s�}��� =��b.���&/��T��ꋶ~�qO��ą?6ΒU1v)�1?r����n��yr��\��参�*^ى�=�y&J�66tU�҈ �:�A��ꆀ�y��J�5�vE� �+5��a⛲�y"K���MbpKZ/ �l`�FV��yb̂�M�0���(83�h�Ɠ��yb��>?����.:�jx��.�yrA�,�i�ьq�"�q���y��ɏ��8���S=Q�#���y���^�D��쉉zH�e�q��1�y��K$�dІ�X�}��A�$�y��F��4Y��"4zE0�� �y�7w�kg�^{�xٲ�I��yb��t"yrLG'M���P��y�j��*򺽘f�\�p�@a���y�%*x�Y��بsXX�� �
��y���1~2̸��;kX8�� �\=�ym�n����lO�w���8Gŗ6�y2�ε{�I0�	=4*�8[����y�aA�d2�˖
+�"֧T��y��N���c!J��!���z���y�D?��4;���*��F�W��y�1PQ��Y8x��s�	�yb#�bOx4�bHU?�`��噪�y���`\9�$ܫHfd�c�R��y"���m�dp��A!z4i�#���y����%�����f!�hQB�B5�0=�p-�0x�ٵA�I	������ #��+P�\pb�%D���
e�E�6]�E��i���0)��T�"� ͍�3'2%�/OPi��"T�7�̘�L��|bd0'Z^P(�fP&
�2=�SD��{��E"ia�`=OF�kt#=�矄�jZ��c�/U�np` R��;?�0O��H�{��ħƌ4���u�8�{"��6�x�'�v����S�S�O��q(ԋF���aj�(�D�ܴ�x5ˊ��iѐ<��<sѮ[�-��\����S�	�K���b��O*�?��O��
QJ\%�tD��bҰU1�drM��@��<�L<����=)Ȳ�GNN�9�0�$�Osy�'\y��(�Խ���J�Ľ�W�@�diR4�'��Gy��IJ�~\)�
�:`��-�0��[G� ���'F��'ڧYN���T�\�d/¸T\�e�%�$�8T]�a��{�~�c瓌"�X���KԿ#"�ۜq��O���{2ʟ���'Ul�,H���	V�@��4��Q�'�$\y# 9�)�g�? l��C��������&�����'��PP�xӼ�OQ?U�/�,Nw�Ap�Jΰ*�8�2�8J�!�ݴ���nZ'�(�������q�L���& &����቗V�fƞ�ݑ>����X�J`3�bў���h�gH���=&$}��ƏP�'���'i�K�.�D��0H��_p^��I����AТq��b��?����p�Ҥ��u�fy�������^&|c��}�a�֧16��A+�l1:x�v�� 'ny�@�:����D�q�n�<y�B댊d(�Iě�c��)�S����[�5C��1�凹��i��N�d0��O��	d1a�d@��k/��57��P҃(ٓ5� ��'o�$2'j�*q`�5k.�ɳ��$�xf5Zueڹ^w `��"C0!�$��f�Ԗ=&%��`ё� Q�'u�����1U��tQP�z�~X��'�����J��~�@�BE_<F�A��'Oh�{�/�Z.�h�%�Senx9�'����_�8T�t`R�߲K٬,@
�''�T�/	})r�
R�F�n�	�'�x�X#G�y�� n�('(�4`�'�ES��L:S��Xʐ/��%�=�'��qr�Ę�e\���l�d&\�'�$�zU�ݏ}�b�ׁ_<�4�'��yx�T= �8y`'�-�X��'��9��_�N��G-+.0��'�,����>�ؘK�B�L�0�Q�'蠂�a��l�����Ѽ=��'F�ea%M���z�͙er�I�ʓXm:��@#O�__�0*�HT�>su���ib�ȓ�x0b��7-�&M,\�ȓD���R���,��ȩ0�H�{�(���e~�ۆ
�����1�@ >��=��M�<�c �I(ne�=� `U�Q��i��YV���
b�&Ȁ@iV*v�����N��wF��M��ś0������Z�cЫ!�|��VJ7zaf؆�,�JQ�'8Sߎ!xTAZ#�戆�S��1;"��{~�P�Lri�M��{z���@��*)=j3LI�Z�I��q�P� ���L��7��P�t�ȓB7��%�ںx�<�����wrI�ȓI�f�b�G�?Jȑ����;^p�ȓj�����^!��ɠ���4M�2H��sc��Qg��H��h��o��Q��1��@���IN�
S��6N�Ąȓ;�j� ��E��}���Z2J�hm�ȓx� ��Eޮ.`B$`��S(��ȓ@.txzBă?�v��V�Q�Tq��ȓ\T�����*���
�"����5�ȓN$�#�"Y/ ��a�&��H���%Tr�CQD��5����@�"0�ȓp���в z=J f�]e���B�$��"�>�0�i����`��.�"� Q�O�Z��w�CV�ȓר8�D#�<4žx��F*2g摄�K?D1C�׋R�6�c��C�=�����L�t��b��AJ4��$ZC�ņȓ\ӂ�ud.P��@��$i�~u�ȓB��ʠ'�6�6P���9&���ȓ|ex��� �Z�0 IO�@,��KHh����Ǟ��pQ�>ǦQ�ȓH�(��菅~R� �g�� ⠹��y)��!�N�(U�(�q���@S@ąȓ��2�l�i:�9x��V'~��ȓn7(�9�mբr�U`E��n�.u��K�@������X�C�S-���S�? "d� c95O^��GK�i~X���"O0h���s��(���Z�#f�ʑ"OdЋu �7:�Z���b['zm:��s"O���LM�vfD1qȈ�4h&�{5"Ox��'CP�Kh�T�A��cQ�T�"O�U �I	Lq��@3Z�VE�q"OZ�E�	zhN��WA�?��Sb"OT��M)	4���`�f�D�R%"O�ᡓ�ܓ��!t�ǹ~ Y"�"O`J��L�):3gL�� ۦ"O�`Ӑ���
��}ZӅS#	��m�"O6tj�iƲB*8�a����8�E"O4��@�ֳ%9�aAE����,�E"O�Тũ/��zt��2Ro8�R�"O�S�N�V���dS�1"�"O����J¥(��K�|b�- "O�A�	�);^<*�[7D� �5"O�5�F6�b���[b2�l�"OqW
�bDyi�LY{�Hi�"Op8bFj�B�����+n� 0�"O�=Q�ωI�ف���3"�D���"O�9�Ꝃ � P0w�R6-x`�"O�IB$��	GF؁ ��Q���E"O�řg-�+mN�����E���sB"Op� �NO�H�䫌�|�"�i�"O"��r'_7>��ⷍFu��p�p"O�ݲ���6�>� V�s��3�"OZ9�dk.G��x�߾&@"5��"O�0���Q#�,�F�
M)�9�"O�9K�IǍ�	���Cu���"O8�x��C�N�b2�Ti�L��"O@�y���,H�$;2S"hgdy�1"OB�2@Q�$�������Jf���"O|�Q��uQ���bB�	B\�\��"O&Ep�T*Y��,�V�W5�,#$"O�P�b�^�B��X����fP�"O��ȥ�<u�q����6����y�i$r�RD�Q-FA�E:��E��y��S�6!ԥ.�F\Z�A�=���	�'�����΀$W�(`3�۝8m�	�'.��jf��&��e�q���(ô���'b�ʁ/]!V3�H���	u����'�tȲ�f�\���0/U$�,�(�'j!pF���!:0�h0ca�b���'���@#J6?����ٔE��A�'����w�B�Ą�S�ϻ9'�Q�
�'�� EĴ]z�Q�%ㅣ=�>��n���{��_�l�T�33��4|�ȓf�z�PD!ɍw��`{��\Mi�ل�o~��7��"��!"�}�Bu��T��D�	�'H�V8sc
�4��<�ȓ
 �����D�'� @)�̑(>H�9�ȓx���8S�B�v$$)	!�$��Ol)z�l��Y������(x����������3M��m�@� #E�|�ȓaG����er9q���"&��ȓz-`ي�!Ɠ�^���6tp�U�ȓ0�����ߞ7
�d�"-�'L������)0e%�p���+�ǀ�3[9�ȓ@�Ha0�Zn�#�^!3I<��ȓ�(�x�KJ0 ��0���}+,��rㆡ��[����)�t�ȓe�0 !1��T���W�9G�hT�ȓDHa�0D�:H��D�:�4ņ�S�? �H̯Y�\�Sn�ʹ{�"O�\��n��U�X�k ��K�����"O�P����5.�Z���.�U��(p%"O̩���7�Ę��K��"{f��@"O8�b���I������I�%V(��C"O����$V� �*A3�ÂD��� u"O����	�D�����[�h���"O��R��
az!��Ǌ���l�D"Obl����wՊ�8���C�`ܣp"O���i�E�v�Q�Y�<ц-��"O`�@!N7-�����
.��� "O��`��݇(�j͑�hC�#����"Ob��K*~U�RΜ��z�"O�9qԏ�My:!p�!U����"ON=K�I59���D��!^��"O�T���ِ&��p�j^
{��r"O�]���Į���3���0e΁�D"O�T��M�y��Q(ݍ
��8�"Oh�a%Y�%��Ǌ=�F��"O���pn�'}>�D�D&B$�v� �"O�=�$���za�!��"gw�ѱ"O�M�B���<h��q���&0D�0	��$S�:����׍=�4�9u�-D������%��v
W��"1;S�1D���C��zaPh��ԛ׬��0�5D� 1��`]lIC1e3 L轐��1D����di&"&�l����1D��!��;�P����U>s�h4�-D��Q*�(�#P��L��q��.0D������-'�"e�)J��i��+D���'�O�<T�qb'L=m���V�'D�X WǓ �xQQ��ƃ�f�8+#D�0	W��������c5���"D�xP��ea��j�ğ�}
]��,"D�0JaD
�|�Xwl�3E�*����:D��$�E�D��d{�E�4a18D��2�CC?�d�4�{d�8���5D��k� ��:�*�p�c�*r�Ԁ��&D�\���ıS�xQ�"��D�8D��Д�Y,�M����<��
q�:D���D,L9ED�< ^7�XЈs�#D�xp�&�Y�+�-����u��d D�XH�fJ4l�j���ڤĊ�yg�=D��2���?�H�
�H����AE/D���S�H� i�Ҡ�P�f�'�,D���J��P�0�taN [���`��+D�� P� P��,Y�K���� (D�Tr:Z�yT�W�!K�tsJ%D��7��S�B<P�.׳�V�� D�l�s�A�e��Ӵ�X#-!z�#D�9D��Sr˘�<0�e��aՍ5�F���*9D��3� ٬m�)RjR�j3.1Xa�;D�PJr�	&@K����F������Յ8D�ċA�yz`I�����R��Ӏ$D��*'�]4O�d,+�` �����&D�Hz`Yg�<؁�/f@f�A�$D��avMF�_��TPG��C4N�hq� D��3r⍑iJ�{���6�2!r�-3D�8�R�6*.P��&\�	 Yy�N>D�Pxgk�qnd�cN�Ju
j�>D�,�R��K�*ɪЬV. �����/D��q� '*nx`MDM�r�,D�Kp��$I%��Ҕ�8q'�Y���)D��Ҫԭ>\�AmT�"�p�ɀi)D�� ������:YKXy���ڃ+�)v"OH�ɢ&�Q,ttFf��d .�F"O� x0c��?����F�ٞl�Hb�"OL���
�[ nqٓLҏ	ސ�h�"O2��W�ОRȠ +���.A��u��"O���vi�M�f�{�߶9��!�"O�ŉ���-6����1AS	N$ّ�"On�qE��&���
�O #V��"O���ЅN�CX@)�/�1j���4"OX�(&P�8�0�9�ρUM2��"O4�����)$�����)QB�Q�"O�Ab��\��-�mZ*I۔�"Oޭ)pjT�i�Vupؓ
��� d"O�t���ǩ0�T�쎔r�09�"Olxdk�-^�Q��;?�8P��"O��{�   ��   �  �  3  �  �+  84  |?  �I  >P  �V  �\  c  Yi  �o  �u  $|  g�  ��  �  ,�  o�  ��  �  5�  ��  1�  ��  1�  ��  ��  <�  ��  ��  �  G�  � �  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@�>������l�'q���[��X"���y���t,de����wQ���d���y��G��pAa�w�*�p�(��y�$�U{�!�ä �jiv�X#ONVB�I�Y�D#�&ՙ"� uQo�)�.C�	�/J,�0cC"]�*e�0H)C�	�4��,�󈁓PV����ԆuBB䉦KT�xA�¡L�\)�DQ�%OB�ɼY�Z<��A��&m,y�̑@��EE{��9O�1ht���;�n\�q��vg,1��8�S�'O�������@�ry��DU>~�t܅ȓ���j�+��kW�h0�;[�nh�ȓt��C�C�|�zl𳨌a\���( Fh"�aJ2/��	�&�2fx�x��1��C��B=:]b���r��Їȓ �L[u�X2<�R
",�ȼ���s����Q�$ ���N=AZ
���.}��)�3� TX�B�C�X`9�N/ ��B"O.�@p��x�J�h�����]+���>���i>}s�GSF䀛�h� 
�b$d#��n�|���L/\-���k�.�L����'�?��$l
=n�^�˓��(R )T 4�Ө�l�A��;h�H�������}��>)�5�J=��N�t��a5����O"�����O�4a!IƷ-~�a�A�a\��R."�P����E�?i����	%g/�U��!���<a�1��Ir6
�`�䙠�.�7� a����UƉ,;6V0�
?�nP��i2}�'��8Â]1e.���)�&�DE��g��	�'�ҝa
��u`T1R�ԛP��B�ɥ8Q|����̓,
��H��^W��=���iR^�Ν��kʍ*r¹s�H5j�T��GO�u��m�4��1#��B��n���'���]~"��I
��4��(e�E�����y��Խ9�h�FN��XZ^<i�@B���'�X#=�|���ן-�����mܰ"t�܊�EFCx���'Һ�2�>)3��ίnnD�ЦJJ(EN4��(����f!��3QzY�Ď!_jʄ��`�'o�U�4nE}i;#�@�d���4!�D94/Rɂ%BD�f��	��2'�	X��^��~ê{��|p4�f/�i�s���y�Hݖ�N���hYV�%`���y��@�@�"X��%G`nD��s(��p?�O�l�6HؿF�L݀� V�H�t"O��k��\C�re"��)"��� "Oʀ�?A����Ҥ�=�5�W"O��1P��^Q�m;��-N����Od�=E��_�TqNE��������lO"�y�拜Qx�a��O-P�v�!�!�?1�O,�@��'ؕJ��Q�����ͽl�@���'7�����IgA�w�Y�ʔ�'�������H��܈�6M���'M{�I$j]옑�P=@�n���'`"XZ��ſo�����%�(hI���O��}�:;D�+�Ν�'ö��q�S�\�Նȓ�6�2C	U6!~�)�a\�6�>M��.aP��q-; B�0���~���3�+FNVgr���/��I/��ȓ*�RT��9��e�bڷUx��ȓ�8�x���+�B�!ȶ4�:��ȓ �b��Aҵ4cdD��ɳ�$a����+���g
>�3B0 ��Q��i�ŀg(�=a���zҥ¶��]�ȓw�j�K��8(l��e�5`�^h�ȓ�����(��t�T&̘qq$X���hO�>e1��41�<���KU�|ّb(��hO�N"J��%
*8Ip$�'u4"c���T�I�O�X�H���D�U/"C�	7:�j)�D�]�h�	�0���Z�>B䉏l�(�-�s�y��D��@H"<A���?0wEǁ=����\�E�l:%�#�O��EgaR3A��i�`����?Z�a�ȓk�m�7�Ƞ&:^��"c�>\�\��'#ў"}�d��A��`,�0R�0X����<��'�:� Q�B���!Ư5#Τl��'*����� ��;aba�tIWx�<��j��d��	;W��?�l85Cx�'�ўʧ�L�i4�X��D�v	S�xڂ��ȓ�x�����<?�P�Y��@�l��U�<)��A����q��N?j�`}��<�����,R^�!��ȹ1�q��S�? ���w`7.���D^!0o����"O"(��Rk��(��&�%T��"�"O}�F֕6]L-;���+{�.���"O�%��-@/e���A�vyr`"O^(0w�DY�Gń-z�Й�"O��k���ĥ3��ИP�|�G"O�q+g��1.����)\�gr�V"Or�#�;0�Z1��#}�H�A"O>P��σ�Zl܀��Y)3�:�@�'��	;
���1�=?����eL�y�jC��'h�Z��O�8��a�O�3%�C�I>vbNu����[�޽��ɶ��C䉃9�����)�,/r��S�	ʐ�/�S�O{�@���ţ6$��92�Ν!4v)a&"OR�A $�3���C6��>Kl�y��IC>���,~�@��a �V�RU�a�&D�,� �
nr�8��R�}�Ҥi�A$D���t��|z�)
�Q�4�y8�A!LO㟌i�!
� �(���p�&�=D�D��ґj����T��9z�#c;��Ɉ�:|��ʽj�dh'じ!>�ua�"O��y��tقt�D�6;np�7T�,�?i����>en⥢/I47-J�@!]�b!�ĝ�C��cŬ��6*�����R������r����;ʟ\��yr�32�#�5 �����#߯�yB��T�q��ȑ�Ĥ;��؉�y��'�0r�N�}
��J)��]�'�%��i޾Y�Iʹ+>Uy�'���
�42�	�g�6%;�@�	�'2�e���?Vt���ꁷ#���	�'h0����F"Xm.9[I��9*�'����&x[� 'j�qM��'��a�SO&�m� i�
���'�	gA�<yڀy�-�4N�!		�'P�!����:|2�Qʎ
���(�'c��f�+!o&�ʣ��R%��'P0@��0�H|��&�?`��'*�0�(��s6�A�eBY48a���'dd���)q��/�\,Kr��yG�)S�x�� K ?�0�i�R��y�B�0v���J2G�_�.����ѕ�yB�J!8��\��2T�ҁ)��A�yRK��vi"�8�=�b���y�욆N����^���Ed�
�y"$�lvx3J
'���M��y��-J�2M���dqR�4Ñ��y�D�'����$Z��<�T���y�Cs����)R	K�2��ň�y�KX�W�P|��bVNS8�ؓ�F��y��/<�J��d��6�4�*�M��yr���&}�-CS�%eC<������y"'F>k��@qg�d�F)w��2�y�Aةl�b(j'LEHΜ��X,�y��J��,hLҚ&i�����	�y2�$yȴH�a	3&s���D˂$�y�5����ψI "x�M���yB$ bWջ�/W.r��1�C�:�y���C0Ӆf :_�4���A
�y2�_7z���C<^\BI�R��<�yrAƦIP�}X��A�P'�x�,ԟ�yR�H>G�(5S�Kժz�*0�` 	�y2�
%d�$�#ϰw�Xp�׎�y���7e�P�%��m�6�K�EG�y���[�����폙9s�\��Gќ�y
� <�B0)	��L���2r}�T"O��B��E)oEQ�A� ���"O$H���
w@��΋���q�"O��"�|�|H:�K�5u��a�"O�lR�c��
�� � �Y��'>��'Wb�'���'��'V2�'/��@B*A���ǠѲ4�*H���'���' b�'�R�'6"�'���'���3L$�`��ϙeN���'��'5��'Q2�' ��'H2�'�z�	V��� qr���JIBf��e�'���'�b�'w��'Ob�'F�'������`\{�K�3<m,!�U�'���'�b�'rR�'��';��'�$tJ�JD�N��x�bN��EX��t�'���'�b�'���'�b�'I��'����B̃u~�R��XG����'2�'���'��'H��'��'�q�3Ǖf��Ck�Y�,���'l��'���'���'"�'�R�'bճ���[����M�*}z��p�'���'*��'�'Br�'p��'��M�T�ӡB����"�۾\޴�`a�'b�'��'���'�B�'���'��q��ԤX���xAa2X�%K��'eR�'/��'��'�"�'�2�'k��g\;_HN�Х���d���S��'bR�'��'�r�'^��'�2�'l�!D��
|������B�H����';2�'�b�'���' B�k�&���O�S�J�cg���o�-"88���@qy�'��)�3?�G�iJ ����(g����Z�,�������������?��<��iP�m��BX�5J�j�f��EN�L��7��O.M��������O$+@F��v����Û��XAm�
]CRHf�C�b
���1K0�	쟈�'+�>M#��>�dB��ߧZ*�\�d�M�MѧW���O�7=��(F&B:Y�(uP1m���L,���ȦECߴ�yBX�b>E�D�
e7�扛R�z���N-H*���/W�(%(�I5mO�1���"�r�E{�OoB�	�a�*a�� U�"<�B!���y"_�$�0��4�p��<�ڵSV��s��U�o����T����'�D�3W��HӔ�	h}�F�tĢ�#C5n!��)�n�d�:Z��1TK�;u�1�0�aԌ�]����ɖ^�$K�)��TeN��2��Cg����$�O?�ɔ\�p$��d�^����8)g�扽�M����S~������S�]T<!1 �c\L������ɣ�M��ibg_�ty��OXPh����U+��z������)�㣀T�24�D�%=�P����N�p2&H*Ir4��0!�dQH!��;W�Tr���*E󮎍c���!�"	TXE��	��T<!��xB�Q���	�i�̢�bΐ<,�����/8�����)@1�|)��8wb�ِ�`�#z`�l�U`˚(�8f�]�1b$T ��)t{������]"��`�L
�r-#�Fىt��Q���P�:�4����?XS�m�V��eRE:�B3Q��12�#QN����i&�����.!���t�)��6�'���'����3?Iw�-f�ME�	�|�*7EAƦ9�	���j���Oyʟ��I'}�O�07�bQz�#��6
L�a���M�w�ʯ웦�'��'��T�=�4��Y$c��\ia�u!�Õ�-�6<l�<b�6}�'���'��y�'R�+`�e�t����GB���La�P���O��Ď l�B$$���͟��I�E��q�b��)7������79�A�OL���O�X(P��O����O:m15��M�
	|�hp+=�7��O*�W�i>Q���ؖ'Q�z#b�+)���BT$h��p�y�F�$/�1O����O:�D�<�"��_�F��)�(>�P��&��0��x�'R�'��I��4�ɪ]L��:��SE1�H����?Y���U�<�	�p�	���'��1�iw>m�w�RNt��K���65J��t
�>���?������Ov���V���S��eHS���:ȁ8�)ӣ}"��?���?�+O@����y��n����*A*N�`��?M9���ܴ�?q���$�OP�$�z���"Ā��dB5����[�"0��i�2�'y�I�d�~`�J|������%�i���I�"p��*F��@nuy�'�R!�����il69[B�;�hP�t��6L\���۴��D�?ln�=����O���f~"� 0{t����!�<GƎԳn��M���?q��
��?��3��6g��	����6t"���Y�T��O�f�6M�Op��O���K@�i>�f
%#$<�ǯ�,�Z�U�S&�MKA�\~�Z�\&?����22�D9pŤ�PBف!Ҥ	w���M���?�[���Aa�x�O���'��E��P z�\�ib�ĵTⒼ��n�>)��?3�Wu��?���?��L)u�������pJ�c G���'�L��� �4�X���O�ʓup��$Q�	L�$�.J-Z�",���iV҇M���'m��'�R�'���,%6m��J<q�Ʃ��o�i��Q!�p�<���O����O��O��	�����l.1S~��j�.b�<ti#��>n�D�	xy�IR���'���'�N�1�{�r��s⇂Y���� �N��%�s���%�	ԟX�	��0��Myr�'�nl!�O3R3��bnV�������h�ct�b���OF���Oz��O�`[����Q��͟��u�È)٘��!'�j�ԭ*`���M���?����d�O�=��M�<9�'����#��/�&XHf�ȬL���2�4�?A���?���Bӌ�р�in��'��O��8��0{��	���4>\�`P�p�@�D�<���a�M�'�?A)O��  �U�K5�
�(G2Ty��J6�i���'G�|;�Go����O�d��i�O�Ը�] �`�HW,]:]��eIwaR\}�'A�����'��^��{���509�՘��N3AѤ`��e�%lT�ք���67�O<��Or�I矒��O��K2���!��S��6��t�ֽ�p8m.jJ�}�IǟЖ������'J��#� �q��9�C��JM��2�kgӊ���O��$�=)Ȇ�lџD�Iџ`��ԟ֝�?n����ʚ���!1��o?�7�O\�i��Q�S�D�'�B�'o�0�S�'2�8q�*!UU�!�rLvӜ���.T`��o՟��	џ��I������8�.�Й��N^�3�6١O�$�)���<�<��'�?����?���|4D�X��ܳg��|��̀�D��w��I>���'$�'�2ȧ~�.O���#~A.��kH�@s���GB����4O�ʓ�?���?��?1 k�t��f)��֒�x�DF�k�$R1�Z�s��7�O���O��$�O�˓�?1r��|Җ$S�C�P]:ĥ�&2��CG��� ����|��� ���LJ7���MK��?q���	9��`&�O�	�"3P�V*��6�'�"�'��ğ$Ad�~>�O�A��͏�B����왟lf=�ķi�"�'���'��	��{��D�O�����}K�E �`�A0Ԍ26	����ئ��Fy��'�>�0!�4����V$#o��*$�M�c�$��葈�M����?�"G�}�F�'�r�',�4�O5��H�.$�l�s�u 8:1�֧~[���?����?����4�$�O9Z�z�
.W+N)S�
b�0��ڴJ�ry�ӺiW�'��O��d�'���'��� ��̤���3��/&`�@W�v�$I�Od��<�'���?�p��!�t��)́Cd�Ԋf�(/9���'���'�j	reJgӶ���O���Ol���x�Y!��~5l�(v�0� �бi#��':I�4�T�yʟ��I�O�D��/v��g�0L��eI�bٹx�T@l�̟\���
�MS��?���?١U?���$c�p��Y1yn�Y�CF��J�o�q���R&k���	ɟH�П4��Ny2�
)\�j�5�!B�jP����^��	���6�$�O���)��O����$t�,[����X�`� ;��j�4O�ʓ�?9��?�+O��:W���|�S��5Lz"0$	�"�89j�_h}��'(|��')"�#B���ZD]�y
A+�iF�����Q���?���?1,O Ip���w��e[dT[�/o4�˶�Ӧ1�5�4�?�J>a���?IW�+�?�L�hx�(�?)&�ԩ�&�|�F�p�n���O8˓
͋��ħ�?��'M���g��D]�1��~C��xb�'���-@��|���Q冃t��Exe	D�0��BE�i��iAb�L��M#GW?����?���O��KGl9l�p���\2w#�m��i���'�����������%���˝By�!�@�I~ ���T�C�6�O&�D�O���^Z�I��<`���*�z1��^���v@�MsER��?M>E���'�X�䡍4S1Q�K�
��J��`Ӳ�D�Op���*0g�$���	şD��MW��fb�uOl�9��d6l�o�b�	�>v�pO|����?���F���:���.T:�`f��� �F�i�h����O��O��Ok�ܼ?�H�c�IԘ{�����ƞ�P��ɵ'4���Ty��'���'S�ɲeDЀ�4�������d���E
q'�&�ē�?1����?9��	�I�5�
�x^��r�ꘃ|/�I��߹�?�/O��$�O���<i7>��I�iqjU��ǔ* ��sGhM-��Iݟ����	ݟ��I�i�p�I�8�z�`hD�W �ͩ$ܔ4a�,P�O����O��D�<I�ظM��O#X$�мAH��j����K�`��v���+��O���Er�0��)��K+������L��c��MC��?y.O%��W������/K<Y�d�E�F @�A,1Ju�L<��?`���?qK>�O�����8`�4E!d��&{����4��D>81z�o�����Ol���}~��$z��9���G!g��HDm���M����?	��<�M>�~���ZXH0���҇~��m�f$��haň��M[��?������x��'Ѣ�����qc<40��"F�4�".v�&���L�OГO>���7R��}XRL�o`F�3�΁h����ߴ�?����?�Պ��'��'!"�'_�����	R�(�?��`��E��Q?���|͟�yʟ
��1"�`~B,�Sfp����8}�4�B i���y�8Py�J6��n}�ԁ�p=ɒ�,p�݂��ن0�\��mߢA�L������֍J/\�{��W�o�Xw��!.�h� �C��i�V����C��C��~G�	:e�E��tX�&�q�<�0�@H5k�4t��L�[Uʑ�I�%��� �6� ��Ap醽�E-Z���؃�T�W�xIڒ��^��a��:&b�'�����'��7���K���j��E����*��{u�:`RЁa��3B�4Q0�p<	SA��#���XP��!h���I!�NF�.�q�B�3 �^l� ���q!0�����c���'��-Ra�:^U�8Ia�4Kr�٨�'��'��O>��#�pz�k�i��J��z�)3�dS޴B֬h#�@" �.�&�A�'x�ɼ|�v ��4�?����)FB/�$��%A��
�T=8d�RQ�="��d�O`ي�GF0"�6H�&��(�moZ6M���|"��Y�NV����d�;o���A��y�ā�Oބ���E�WA��b1/f�6����_�Q^��+�h�<�۴g�H�z����\�0*���>��E��h�ID��y�3� @M2�/����� ϋ	|������Ob�󤊪N<�Ā�#RO� ��E��Ec֢=ͧ0@�����H�&ca�Z;N���Ä�Mk���?���	F�]yVE@��?����?�Ӽˑ��5&6p�7��U�x�*c�u�g�!�T"���mS�5x�lŅ�ēF�zQ�,�!p4UiQ�H/?��f�Z��b�s$FS&~T貀�
u��鹡[>IP��¡$��s�hĠC%lM������*�m���䟥U�����?���cv�1������C�$;��P�	�'tv��ԆH�0�vxa�h�0��,��'k��8��b���D>"�)�S爋O�$JS&�H����� �x����O"��O�-�;�?�����$#��V�R��0�C�Hg��A�Ə�K�1XV)�2>������G�P2���XU�
�
�!K�us������4����n\#7��D�QҖ����I8Fn\yr�G[�����ADn����O�dmZ���I��ӟ��	񟜖O~��ì�>�1��z�1R	�':���1e�딫s�IȈy�i�:��<��,Y���'#R�O�6NA�a�Ѕ
�FԮ�B�'zp�1a�'l":�ʉ����3���ƙ�-�kS�(d�p�h�:��F�ԯ�p<I�Y�ˢ��Peڶ��C�����x��o�>�:��#����yK�-�'�U�Pl&���a�	��Ms��i�2�n�p���?)K"AA3��2��	ğ��?E�4��.,�j�O�%C�<zq���O�=�'~����1:�X��i��k
��A[���|2����6v���.'HT�b	�&�HB�IZn�Pq� ��&aVH҅m|PB�	�hT�Ӧ�U�2�0Ġc�S{�$B�/��:�׀4$�M���6�<C�I�s\��f���؝8f�Z%Y��C�I�6v����L;X�|U���7��B��96���G�:7��A�D�	՞B��
v@q9u-��$وT�C�[��C䉇$��4�#��9C�hsP/Mh��C�I�9d�f`��;��2�NнۢC�Ic ��T)�&���Q�M4tC�	�#K4a��J`k6	H��Ck�C�;c�б��_"=3I�#��C�ɴ@V
 j�k�
��.<�VB�	�b,Լ8�Nѣ]qah�Q|||C�	�f���C��#]�)�JM%�C䉼_� }��F&d��@!��˪��B���p��SCF�#�����ȴ��B䉄J���#eR�f
>D	C�	�r�HB�	����p��0`�ʀA�F�P�fB�ɤr�yi�O�i!�ܰ�)E�;�C�I jI���Շ_"x��L��D��DC��/<�E�e�F%�f�I�AÙ��C䉽d�~i!��#{͆ȩ��4:��B�	�4���:"�/D
jB�I:�<!H�"��T��54�:B�8R*� 1T�r�L��7��B�K����Ҍ:w��b0�ȍ"�B䉚��r&�S�@�`$@F7A��C䉢�<	���R��nq�f�>'��C�	�lQ��H (X#K��-��ϼ6O�C�	sh�Qy�Ș��u��+L�n�=���iw�=I`D=��3�0yy7�](� ��b J�+H6B�	�@U��Q�]���x �M�`�:7��*�!��c�U��@G��Mk 7|y�av���GQL���_�<)��t8��e��<��ݲc��2�.�n�6b;�񀔟|��?7-��`�R�wp��3�qT`��F�1 ބ$
�#��K2^�1��<4#��C��"�E߻������ �A`��7�qQ1o��g f%�q�&�'��̳u#��>Z<HCA�5|{d��D����ظ��S?m������
^��Z�)V��	�A�X ����Ęf��PI���zpN�IÓB΢��Dn��X��e�5,ڹ|���I�dh���J�C�����]^��|R�I�\4��Cg$̨�@��8�TK�MCI(<a�F*AjT@��ʘ �
�cq��&锠�	�Y+��M�(C!@��|nڜjX]��;�l	��0G���/	61T�X���'���D	S�m�r� ʨ�$�*y�00�+��!O�P;����cd�GoÞ5�r
A9TG-?�'2�8�T)ۿ�|H
4��m�F�A��D"Y�h���O&�$���V��AKP\&��k�6��!��.AҴ��mR�/06IcwZ?��� �'žp*�CJ&������)����"���c� \?m��0��I������7E�\�`J��,�AaG�v7�Lr��ڵI&�b�[�
Q"� aK�JˇJнOƸe�-.@����4�$r��S���<(��`���X���"��)(�'˫[{�<��'�ZlQT&_����E/	�rp�5펻S̀=��K�^��hV�� ���jR,S�9��8`�U�{~��Ǵ2+�}�5H�%|��hJDø��d� -���!Q0�~RnU���116�2_Dd˳��cޔ��F���*�MT�|���8�EY1`��Ph��M�H�f��A"H!�	fJ��h�h��y"��ј'���3}Ұ�5�&�aw*YaΝ+=�h�qi�?j�X
�q� ��G%����3�0:��U��4\�Q7�>Y����ؠ8�'�P���y��0��1�4D���
>�9�j]����Fxrh����Y2E?B�}�wZ?���-D�@�"�
і�R�-�<8>@�'�U����y�	�V�b�j���Y��E�U	�S5� 8kWa�)��@$�:QK�c1v�4�qO�	�\w��YUJ�=z&,b��2uY\=��`߽%�ݡ�i���>��E�7�y���;C�4*��:�2E�G�e_0M�|B�<�P��)M8�A�`�"cQ6x	��'�D��-@m��h �gr�1K�&H u�tD���D}I�t���c�$m��!�+
�6�$�q0
�'�^a ����3��!h�"=�dų/�`�"9a���y���*�dlrp�C*<V��������O��w�ūC����蜧��sQ���Jf�Q�t`=���Zڒ��ϋ�$��IEƣ��̢�%Y�q~��l�c�'�eE'\"O0���_Q��`�K���$�	�k.�-M�LVax�=@��hP5+	cn^$h��C�j�.��'3�k�)�'�ڭ�u˟rČ�[�c��Z�< G�-lOzMpPCsaD�������W&ݖ)ȃ	U�m��@�J�S��OPT��IQ���LF��L;Ǯ7t.fm�a��0�R����M9æ
4�fl�i��p!R��96_��A�T�}�������
K ���}¢�2Hn>|C3(����X�F��ē=(1���W�FM��C-*��nF�r�b��)?t�A�S��z���O6�RĞ�k̩�w*���s�f�*%���;�Ό�<'�d�P[X�x �fR�j��
R�*� j���' �&����i�*G{��T#"�Fm�4�ԩ_�Ɋ���Y�Ї����K�
�.f���IĆ��Q���c
`����A� ��H��aX�j�6[?-x��Rz1�Ň�ɪ۶���`�+�щ'��G	0�B2��' ܬX0$�!V�����#.��Txś�l;�@�[�hX�,�'B4��#�.����̒!Ѱ�Q.O�!�c?sˆE��NɡPMz��4�I�S(�q��8V�B�jt�Ì,�p%:5�9'J��a	�{OpACn�K��}�W(�%�b|���0td����'�>��+B�z�"5���c�
�f�ض�<���ȖCn<� �נ#��[q	�D(���Ѣ��86"?)q�Ȫ;Ȉ%@%%ܮVM��µi��U�-T�o��� *
;9N�	V1ғZ*Ƀ"˧w��E��\���'� �*��;�0����H���`�'�(��iߐ�xDH.� �jʍ��>�4< Fȕ�)��A��$2�fk��G@��3�4u�@��@� 6�(O�	�U䘼���*�D��攡wL�ZA��~����d͔4�X�\���ƠЪ	{�MK��z}��i>X1i�)) !@/z��/�M��頩)�O6H�R���f�
I
��ˆ�������y���q%�A��(O7헷M�X ��ɟ�srİ��B����dԊ8�N��e��!��hǢ�4�T᱋ֈU���P1��Ֆ>��a�3~�f��PB�%>5��I�<�#gK��HR��@ �����i&�?^����_��yV���I����ʑy����HP�'�����:��y���  21p(N"{@�x2�AP���(�O�%���.4-�8[SД+��|�� �N�@�J8}�x�>�s8O󎝻kb��u֍Zu.b�Xa}"�L1,�q۴o��)�ǤQ��ʌ����!�����T�)7��Y�R���cO��}®��]cb�ՈD��<%~4+�B;k�A:7�5ړ�" &�O^�bgog�>O`)yQ� /
޸k��y`�tƓx�*�ϟ�� �e�j�A��;�?�$<?�.��,%����[b\T{gIk�WUޘA��Vئe+%%U P���O����������j��0hNLHY��O̺�x�D��&>��̔�5p����	(��0җ-�&i�Jh�	W�n��F!�?�r��p���O�$�H�p��=�9�#&E�01ĜZ"�B�,��1�7F�C<�� y,�N� �(�YpE�8aO
�'�2&���XAaܢkj��nP?J�ԥ�#J��c=��.)~�����g�ؤ ��i}(P� �4��E�+����e�����8?�a��>Lo�Hץ\������n�� P���
�
4��mZBL�2g;���s�D��]Tf黅��4U�T��f�2"�'*�����meu�v�3�Nm��B^�*>>a�R.@�*��8�$��6�p<IVG�/�"}���hA�!HB�$�p��F"�_(h �Ԇd���'��x b�$���)�$�� P�I厨�p=I�iy�%���K���$!>o��\quCќ'͆��<q����-�5��B�$�*$	3H��Ht���P�F��r��(?ۮUJn� �M��/��i�']z��FD������+!gL�ȍ��	R9��h煘*}���7���I>��{�G�Q�,]�a�\oB�t�јw |e�ɵ\�f���.4}2B�E��w��q��*�4���A�0�#�e7����C�H�Ecu�0<Q�j<+���v�,9x
Ԏ�1U.�͓�?���G� mh�'U���;>H0���h�}���K*�P����I-* �贈F�d �zB��" �:,��'K� H�,O�~(^��g�C#|0�b���`E���ꕿ&�4�5�O�.Y��~��ܧx&a��bY1D��e���L;j(�eˠ2J �X��	�%��d ����R ڶ��'��<H�씲J��h�K�O���y��Ӧ��I٦]��J��D��(ٓ�:"<�6.&=��T� |>m�4
^������� ��Ӈ-F��e,?޴J�pX'Z�uI��@@�`;�q���{<:����B�oĴH��;���$Ȟ)Ҟ4���7|�)q��6q���&5O��h�%�ߴc�p���	7*�w�<}��H�$�P�R(�pF�
�!���4��53>��qψmtZ y�I-D���E,\2�ଘƷi ����">��IB��Q[�B� �*���Ojxأ啗Lఱ�"���_ND���	�8jyا텷`���&����D�i��Tl�ǲ7Gгb���J��>�(��s�'�I��t �/�0<�*�,� Q��j��ޔ`������f ^-v)��])6�j,�"y����D����I0Õ�G}d����&&�(K��P�D�\Xy��'��T����U���b*�#�y�CT;8���n&��x}b�	���9���Y���e�l�{�N �U-��۵�'PV��gǢ>�EGK�o���X�(ȗ7��@XSm�H̓wN|W�>��eƳWk��OU��O[)������P+U�@y�Ex ߀r�L�q�H��,�R�<�M�Oi��" ��k�\
��M�'(�[,O<�sw!��w����bI�68A�v��+z����j� p]��{�Y]v���ç�z(v���$�a�i�����,���+��C�౉�͘�+�d�;r�;<Ry9{X�(�FI�=	���Hu�L|xg��TT7�M:���%LʢPP��dc�i�mQ� jh�F�W�3�*鲗�!�O
��PA��l4��\_��� C�,Ӕ@b���I��U'�@�'��i�#�r٦(���А��4P����Bh�F��	���#`Ey"�6^���F`�2�	�����+X���K��y,���`�\c��ɘdZ��!u�M�c\L,`���$E�]�h�* �[5Q�vxi��	�;���
���p�"c�4�̽�"?)�GQqV\q���إ_t�|�����B�dc�'U����O�E�A��	�6(jm�WȪA�����v�jl��w��M:��Ņg<��b�˦q3T8��cf�r�o�	<s��Jq�
߽ekX���4OH�OX�����7�H�S$�T0.��Y���P3�x���� ��`���8ړ"��M���zi<8�De� XrDd�B�椙wk ��MzQl�����" l^�97A&τWE���C*O������+J*Ҹb���R�\��:O꼠�*�VoM#���j.����>O��D������ ��2�s��םB�"���S�J�J�	ˢ�0ĠL�y�u3����!)���m�'Qn`T.ܜ���~�t5	�ό�A0\)Ѵ�����d�/t�X,��玎!"�C�ܒ5�شZe�pv'��k��x���0d�(~и�l][��O�s�%����a�j�>i�#퉈~B�x�fh��6֭O��BnD����H�d�R</�m!�nQ�o�����	X�P ą�	Z�m�� �eBM�i�Q�<��K��a3�)�SO�h�qbBֱ/�.0�s	%Vo~�ũ�'�yRhч^մ�kQˎ������ ��=-��OzT�&�I�y�Th�An8��\jv�Ԧt��ȓ8P\=�T$B��0�PL|��T�Jm�Ԧ�$$ �q80/�& ��ȓ��E���F�I�u@�N�<�"l��by��8�[�
�	���@ B�=�ȓT��Q��N_�#�R�#r��F(^����lMؖ&��W(�`g�F��t��,	"I���LE��x+S$7����\��i��9vd('oW�S*��ȓ-���'R?���a�&lry�� %R�	`�*� �A��B
(؆ȓT��c���8�ʼ�K�&���S�? #�@O�/��\�Unפ>��QU"O���t(�,(� ��#-�O���@"O*�xe���}� �j�A�Ҥ�h`"O|=�c�*V�XR�M
�Y��,Z�"O¹Q�CX+�6��q�ŎU��8�"O��sAN�hC�1	㥇�"M�٠"O�`���6`j��e��0�<��C"O�sf���]ѷ��z~��"O�P -Ǎ�n���Ȋinv4��"O��&Z�zܬ�3�#ώ#��@+4"O�\��ݿV_�Qbt��
�"O�m0�Խ
�t��͵'3p���"O�$�A�J����%��5�u"O.9Yr�"�\9S�i̱V�H�Y�"O�ͨ�='�:�i֘ &<���"O ��@!�?Y�D�0�H&����"ODD��aظ/�49��(�w
�a�$"OjQcRd�Z92R*U._�\0�"OHa�gۉ�B���n�9�nT��"O$���A�)��Ǫ�	���Q"O�����+դ�۶�W�K԰�R�"O��b��>[�.,(�e\�z�����"O�E�� �N��E:ÆD_�`0�"O8��5]kL��k����H�"O��q�4uHN�rW�B	#&M�"O�4˳m�'GƔ��2�?�X,p "O�|���%(��	�A�/ir�"O:�ɥ���\4C���-a�Zb"O��@�. � 1B�����0B>�	p"OLĊЌ_�_�H3gT�b3�k"O�!��̛�QRLa���\ ��C"Op��o�!�at��q�"O�1�a
�U�p�م���c�"O
	��[?�*Dti�R�f%�"O�X� �X*;��3�)T&r�dŻa"Oh"���9H��X��X+!��(P�"O�Q
TE��n��H�6�! �"OȈIrJ�k�NQB�WJ
�"O晲��v��pa�U�~�X��"O>�鷉��b��ɺ�E��ll�R�"O����P�>��i�#�ѷP�u11"O�)Rl��3&�4#DP3���"O=�Ռ ��hBD�� $ �0�C"OV,��g�%=�
�z��Pf���f"O�H�eD�t
��ؤ�ZM $D�u"O���CV_�j�OS)'�J�@"O�y9�Κ9L�ƥ���X��{�"OzM{pl���ш��W'Oެ�A�"O�,p�� ���8���8��<�f"O��`�įM*�����h�Dxx�"O0�kAd��Y�q�pbI
7u&��B"O��+��D�5���b$�6njɶ"O�4Q`@	�,�	�V��4Mlh��"O~Us�'߄[���֢{G��S�"O�����%?�X�R%��]c���"Oؤ��I�)[�ع���xk@Tb"O���`��:�XeC��ז+�ԍb1"O:A�F*5f���*�0��"ON\(,SRU!҅
٫q�<|��"O\d���ȋIܩ�`��]�҉��"O�%���#�q��DN�p�tBV"O:�hv	�.i��R��7�<��"O�{0�X�-C�Dbѭ�0��騧"O0�PO�,�$��#c������y
�  UX�"T�\' $�U�}�8�p"O~����O}�f!��a���C&"Oh0�4ۇi��8��)
��"�"O��n�g��Zb�CY�j�n$D�y�G5xA5Cߔ��[0�=D�����-4\��� H��=D��Q�.R6w��8bp'�$/��dE?D�HB�������-�J�%#D������%>�x��.tFĉ"u�"D���T�݈$qVZ6��+s�H1*d.5D�0��C�)�j<�Vm'J���gD4D���$eԡF��Mq��]�t�1D���*�`Ĳ�p�$��O��@C�!D�<ȣ�Ÿ�D9ӡG|�܀Y�F?D��x�G�(H�\�qG�/_)¤�7�=D�Ȼ�D؉9f�y�p�-���1G�<D� (��ǋ#n��',�y`���;D� J�ȏb�&��UB��&�:1��$D��bc�L|��1QaWeKR���m$D�X
Rɉ2���蔔m�z�� �5D�H�Ђ�A�v��Acѡ9�L�5D�@���O�_궡� ��1n�npA�H D�����?��|8@�Ƣ�H<�"$D��9ЎH�w�<��
:'�>L�g D��v� ~�\��T ��@Y̍�r)?D�d�ӀD)VF�
U��4V ����*8D����	:�.���� %�5 ��#D�ȡ2B-�dP���+	n��Zv%6D�|����\V0�I�;:�`�,6�񨟰����O�\p9�F�"�@"Of�e :Sll�"AAM�p1�"O8�9�R�pk��Z�8J$Ia�"Oִ���5&Y����`(B粰�4"O$�I�D��쒐���E�f��P"O�Y�"l�|ZB���)� J�@ô"O��B��8�J]c���,5��|�"OԌ��'� �����L���0�"O�B���Iz,J�'P��Z��/�yb��>���3W$��"��I��N��y�$X8+Y���D�%��̣�J��y2�%��0���U�칰+�yB�"nb����L�C��ܛ�h��y���l<�ӓkO����V4�y�\�,6�����rS���3���y2�"u�����p�ʲE_8�y��_V8D�ר��&�X=3�\��yr΃ldh��I�"-�}�����y�	�4�8(]����+��yR �CȪq��aY7$ �IJ��:�yr�@&�`a�$J�+v6p����y�N�(~z���Ħ'���׉J�y"
N�S�0� Q�2N0���cۣ�ē�p>tnG�v��� @��:�H���}���'���d��;�=S�._qTJ
�'̐DY"�خ�ö��C9�hY	�'���@E��	]3v�r���g��=�	�'�6�!Ʃ��t�@�{p�'-�:�	�'	����/�4u��a�m�<1�T��'!��Xw�R+���C�d	:#����'ݤ�gDJ1B7Bt��"l�ġ��'�V8���^�	W�*d��B�s�'�t�ʠ	[�ң#�5)6�H�'��<����>�(�+À.	�|��'��zQ.��(�D,�RI�F��"O� �m�7�ה
Y�(�+ϑU�~e��"O�(Z��l��d�ĸ) t��"O��@ ѷ)P�Վ��~n�!v"O.�� �){$�������;��4D�( "̋,��A���Y�� .3D��:p�X�+T���t�V?o.��"l0D��['oG_|��/��Hb��!4"�x������,h�d��I�נ	���A#�!�5"�d�[�k�>Q�X��C,�����l��!x�Yf�ƒ\S> �C(��b*B��!F�H;��]"��ѩ���B�	.IꅻCL��� �% N�O��C�I<O��`�Cj�3�(���&ϳp[C䉽m�̴[�����t)�/��B�ɬu���єj�3Y��d���шkm�C�I3�
�K���O�Y@
ӫ��C�I�8ǐ10�ԙT0�%T���I��C�I1`N�q�D� 3�q{3ΔߤB�Ɏ	��C�n+jɦEk⁑�?�fB�I� ���H��#0Z���($�dB�: �Xj�Ͼ7�Z�J ��6�C�I�h�^����>x,t�u.T�C�	�P ���G�.9�fE:'�ͪo�FB䉫6)s ��"�E�%"�8O(B�	46ƅ����\�\�g"&��C�	='�8�1���.Or� "Dj��B�	�+s��b��P4O��u{�D�CW�B�	���P�d�� �1X�L��&s�B�	5L�[XV�̤&Zt�{%$H��C䉚m�6��EOP�T��l��iJ�z�DC䉅&��%�ԧ���l�(D�̟
4C�I�J0��ÉZ�/��4$]�_��B�H�B��Q�۟8���{"L�!�B䉇r�p���lS�o���*B�^�P^JB�	.-�`ܙ�K	�^��X��`�|B�	�uz�YSӅF�qu��(�+�R`>C�	v�М��-��U,�Iw�! �|C�I�Q����v��5r� �╆E=B[�C�	=�6� '=a�eIB�F�6��C�9~�Qsc�_)>�R�kF6c�pC�ɓ|
6�J��h�h͒DSLB�� W���It��4�:�"u����C�I��!a��E�jy�ehɜe��C�I�U�t��A��bZN�s Ff��B�	V��=�FZ�O��gD��1C�	$+�@�#'�^���DѱCW2C䉷qS���3���0��:	6B�	�<lh�C��d��h���C䉩z<n؈c���~��ly���.w��C��*~�å��@���*G��8y�C�I2o�Ȅ"\:}h�ԁC&��1 C��fS(IQ���.9�|8�#��ƾB�ɷ[�
g	M�J�n��G� R�vC�	($[�$Q!-��oȬ`��KO�m�C�I8���%ޒT\��C%�ѥ�C�I�{�vasц��
�<�ÅS�1 �C��!
��@n�wgj �+��W)tC�I��q���,z0�1�*�7S�B�	�C*�����.hjE��ɍ�_�6B�ɈO�t\�V��!�R-�BKH'*N�B�I�/q0�@� '(�lR��<��B�	�sV��Y�b��pK��u�~B�	��Z��6a�:FZ�X��Y*m�hB�I%`����K��n�0Q�� 5��B�)� �Q`�־1g�5+g@��sB$�1"O�|���XI8�
�[AWV��G"O��(X��4 �)1I�Y+&"O����O̮7���EG�H��1"Ol�Cc��)2|nT���hN��"O@��r�ؙ�EP5"x���"O����kU�U��E"g '��A��"O��R7$@�:q����;D���f"O����J=�,�1�"[$*Ԕ�E*Ov�8��^�8D�X��D96'�y�'�&|���J'z�t0K�MUy%��	�'l�3�!7��k�B�w{\d)�'���V�9c�����I#�z��'�HTS'�D�0�/GȲ���'������3d�h��� FId���'��s���[C,���'�3�����'6
� SY�h�ȜhA�VC>q��'���o�6[7��oV�\,��{�' �Ua$�P5`>�S��� z���' m�d��2ZXB-�V�Di�n\c
�'�XXD-F;&F���²ZV��	�'���Ӆk3Ǟ�	��1a���	�'����ej29�i["GϪ][VA��'�DY� �T����Q�D=�LC�'�Z`c#�L$6J��GԱq�<a�'��A�cԪ]0D�&�ץep�M��'���!�B'���ZW�$R��B�'<�#[�(�t�A'� Qx�E@�'�J�R�	nͪ����B�T�2�'#p� 6S�\�:�7��|K�'9�\	���sP�)���Q�)�ĭ��'�x��CJ�-��M�DL� �x�!�'��q�� A�,�c��0a�'�t��_z���{�$�|�����'��!�cAO��85��Ar����'��d��@Q \ܣ� ��lJ�} �'L�M�ӂV�=��U�0�����' x+��-�:iC1�Ʒ��y	�'��5���ђ%g@����/K��"	�'H.0��e�-]��0`�$s#��K	�'OD
�c�(&�x����r����'|����ɷ
��T�����lz�1�'lx+��y1����R�i�<�X�'��AƄ��(�^th�.S�ve�'�dЈ7k��b8�&'SNj�J	�'�!����RͨU'�%L�=
�')���A5r>	�cĂF�8�X
�'m�P��L	"}z�:@@��?D��+�'��]`q��3����`�%JzHQ�'�<�Ȕ&A%���:��^�QH�Y�'�bp��]/�����GQ�W`�\�	�'��!1�גbXH���� 	%�>E��'��%�wO��@+R����Ś�R0z�'j��˰��ro��)4@!x:�d*�' 	ID Ϧ#�Dл��^�����'��%�f�E>f�H���ُYv"hi�'A,a+���)+��RFm׽J��,�'�h���ԛ0����ʼCǈ��'�fdpbc
y�2�bi�>H�a�']6�cTc�n��9	�:Ax�	�'Rv�C�e�C���k�=����'��`�/�A�@�,i���)�'.��c/=���r��U�b���'�r����K�W�Z�DO�R����� ���Q�>�iQꚣBp��1A"O���af=A��0*@��(�����"O�з+�u�0���ў}P�@�"O�Xq3�����9p��:*c�`"O$�	`��zh��[�lџ%b
��W"O�a��#� -�a���O&bY��"O!"g��<��ġV�ęY>Pm�"O���gJ�};�Y��\,����"OLř�;,���ֆY�O,�!�"OB,Z׃�1���إ�2��M@�"O����N' j�;u�54���I"OZ�7�U��^�r6c�P�� "OL��UK�[480qV��=lF�88"O��[s�@B+�-\vFR(�1"O~I��>'_t��eQ�ED�2R"O4<`�DN�?<(�Ĥ��	"M��"O�x�*�{Z�x@�QaA�"Of\���Yݞm�Q�C�qPF`("O�Uɇ�9��|��"������G"Oh<��#��E�f�x�!l:�Ȑ"O&P
��؅F(t-���۩LujX��"O.���'%�9H6�ȁEF �3"O����Q���L�LTyr�"O��r��U�œ %��+�"OrXK��V�> ��� *y��z"O���R-7;�)V#M�O_�D��"O~�R�5�t���A�+BD�=I�"O��Ѳ�șWBv��G��k b�@�"O���U��~����S�~F8p"O�MH㮋�"�4�u���B�����"O]b0*��'X�EgH	4�%��"O��)ƏA�j"J���GQ�8��b"On	��ޣ����,����"Ot�S�U�0����!��\~���"O�@{���%\?�!�@>P�*E"O*�Ԏ@�I�ty��ϟ?JR���"O���@BT%H@4ls��P$FLB�a"O���D�/��q�%C�D�=��"Or|P�H�s5�(�eg��i�|��"O��	Q��<"x�q�h�>�i�"O����h�F��h}��Ip�"O�=�+�W�Z� 7M"V�r��"O�L�O%j�PL�l^\��@�"O'HIz=2[(L�J��Ʒ"U!�d�z�(�b'�Z
	y,a!��3�!�dûf���ʇ��&<[���HI�C�!�G�,����5F�G���Ap�N�p�!��� hP��1�-�; �!F,]�!򄎵1��cv)�n���J��W�`�!�$�(n��8�	G �|�clɁ+!򄋑B�P���F�w� hc_�M/!�[1Y4���'?��Zw�{�!�,�@��rï&����S�M�Qx!�P	|��� �[�8��f��$g!�ĉ0bp!�&�/6T�X��%�v�!�F+�v���#�s7�P��
�j�!�ٜZ8� �T���4k��M:x�!��7;J���oӱA�v,0���4!�!�$F`qh�"�%Q�s��٢a�
�!!���N �i�3�R�W�	a� �( r!򄚹33��
3��E$>�R��C^!���<1GZU���w`�+����
Y!�W;oX���U�*�*��f�!�d
+ni��#�&	|-���-�!�� d!���$WI���S�Fl�c"O�5��y�0�J0D �O�d��C"Oм�&i�X(����B�Qi�"O^���%����� �9@8��[t"O��3���/M�4��bb�;e04y��"O�`a�2踤 v+H̘Q+�"O�œ����m������%|�D��"O(X�@�E2A$l��Z�^�:�rP"O<�fC�/�.iq󄇭=����"Oj�Jdc���^��$H�Z�U��"O hx�Q�)jJR�CC�c��(�T"O��B�J�U���cޤ/��ě�"O�x@��J�|�&	Є�b���"OJT��.�V*ͱ���9�m��"O�`��F�\L0��B�X�S%�dZ�"ODD�Vo�\e��8�ӎ-6���Q"O�1�%LJ�o����%6�x��p"O��Y�)�:��h�% �:�x�AG"OZ]�e�B�TKV���CY�g��m��"O�l��U�6��FC�F4�"O<eP�Y7�r@$BE4	��	�"O6`�GT/Y:��0ြ��Q1�"O0��kc괈i۾g�@�؃"O��2矼xP~MsF-��F`x"O� 0gX�UDdI�톑+��db�"OJ�˔�F��SF�� �pk`"O��p�	P��c�� >.����"O�H�rU�H�j�ӕ
���ک	B"Oؠ��KU.E&Z F�ݓO'�p�"O�dX"��M��ٳתZ<'jz�"OlyjԪT�}	tI#��0xT���$"OZ,ha��\�J�F�9Vn��Q�"O�P��̉���'%V"P��Z$"O* Å_Zs��Co��]TX9� "OR��� O9�B�[H��"�"O�����д*49Pu-8,�	�p"O@T�j� �<)����=�M�"O��3�Q/f��<�AL�3��t"O������F��%�2,�D�t��"O�Ѱ�\-��H�-�"|��"O���!2�i�C���N�"Of�+p �s�,���k�
+��{"O���׺<���7�ӳ}����Q"O���ac8�е/L�p���"O~4ĉ^�L�c���wx���"O�1h1�9�rI� VX4Iq"O )�P�����rF��5&8�B"OLd#$MH���DF�}�:�"OLT��߷U�Y�@Ŏlf�0Ç"O��ڗ��n,`��w�� �� ��"Od�!5C FZD�7I	�M�D*#"OB�@4��,e�6��֍��G�AZ"OB���Z�H� P3��L+^�ۥ"O���%	V/gz	y ��G��+�"O�S�AV�2t�ɇ�� ��}X"O�T����'r��R�*s�|Ős"O)a���`�"�z�D�
sn���"O0��P��al��V�ҌSf9k4"O��˓+Ȫ+����*L�9�"OĐ���2TrF�{҂[�C��M��"O\���̧bZa3D�-y�S"OX �Ee�1f�kt ��n�1F"O^�ҧE�B�D�96���"u�"O�9Ƣ��tI>��$�{���s�"O� ny��#��R¢���*� p� e"O��	&d�	"X�'��$K H6"O҈��EB�l��|��$ƗW���"O�dRÑ&�qxcR9"����"O*�mבE! � �hX>c�	u"O.\C�"�:Z ���&Z�~|�m�c"O�A�q
��,6(�Ǡp���"O�	0W�U6v�b�Y�_�҄�Z"O�̢K��	l����G�.�*ɑ`"Op�³$%�����/
�9!�J��yb��$MUx����/��J���yR��`{"<�Չ�%�t�q"iR
�y���eV�T9���%�����m�=�y�m��%��5�`�3:x�X䃖-�y2gӝxa�YS�/��l��s#ET��y���)��G�����SSI0�yRh��U�V$��	�:�	FjY?�y���Z�aPaH�P�������y�+���%��M�D�ԣς�yRG�7O6���ݻP�Ƞ��热�y���K�C��A�w���Z��΅�y2�@��2� �#՗tK������y�g�=��eۀ����D���d)�y�ɋY8D���9L���[�y��Í,@��w�&�@�zEL\=�y��:*�ԠU����MH��&�y�� �;�x�V���}ȴ��֬�y2߿G�:4�c��~Z�h˶"ܥ�yrA̞p�����ʌK��+�˪�y��˃y��Q��=n����ɘ8�y2��<&T�Ѻ���i�Z1���D�yBB_�j�j�Rp	�b���P�,��y2�0�V�ҩ^^C�]C�킎�y��"fI�#�f҆J�Ѣ�����y��+0j�|��J�0�Q�%g��ym�3O �]i�'Tx�����E��y2iL'���`Ĝ Rq����y��� NAND�`&�*8�Q���-�y��R%I0�h����. D1�H��y�F�Z���{��W�},Is�]�y©�*��ŊE�A,|��uP����y��%Xp�+�!�	p�+q9���ȓdy�qX�I���Ds�Dżw�(%�ȓ.���`��1y��1s���7)����{t��#S:����E�2-���ȓ"D�����O�H)Ղ�/n�����R��JU�� �i
�:�Ԅ�
$48��`��O �,*AaB�1ݮt��qP@L0�-�? ��uȓ��|�i�ȓMrh�0�T�,)@ap򩚾����ȓjd�u��ћ4Մh:��97�:T�ȓ��}ڲ�F+LPle�a���zm��PǢU��m[,5�<���	98H�ȓYM
��c,C�B��B��S	n����I������,l��l�L�&̄ȓ��Q�E	J�n�����*UOd݄ȓ*�R-*��TGx%�����R5�ȓLT`0$�.�����yAș��OD�(F$W)���zj��dTPх�O�P�0��gp�QO��c�L��K�V�j���s/n5:W��y�I�ȓx�b�Z�n����7�Vƶ �ȓRx���@�+j����Q��5)n(���3��b�M�%{��`��
Ok�M��S�? lt:uP"
�
��A-m��e"O��렆�Q�n+7E!t{R�A�"O��!,ƶ/����
@Փ�"O��5��$5vl�b�ݶ%��X	�"O��ܖWИ�cUj��Ex��ZQ"O�T��<o�\��D�o]0*�"O���u��	2.��e[SN�=+�"O�ɊG`�ys>%���rϐ�y�"O>�0FΞg���S�X</����"O�*l�	{?fD��ΰ:��	��"O�a+���`2py�	�$V�0�"O�e�`�ɇ|���&G�6*��2�"O�W&L��9j��N�l�ش�$N�i�<�s(G�!擄z`�sq@HBkYb�<᧬��7���`�LTh��@��Og�<��#�.{ΆHc��S��V(���`�<����5��ua�T����"\u�<��S��v��  ����EJ�<�3O�^�� ѣ�4N��h#k�<Ѵď�q~Ą����+-?JP� �Q�<��.Mg�,b���rJNm8s�YO�<�-�f�X�R�m�@��)�"D�v�<q��	�3�ΉRچ�Ƀ,�n�<�QF��*�&�)�h��"���G�T�<�	N�)�=�Ө�Y0����u�<Y�l��F���2�k�X)wǈ}�<�+ڑ:,&�a�`C
Ub��F�Ne�<�׎�g�<d���M*o,4�q��]�<�'f��xQ$���&�"R�V���Z�<�5��4����)N���	��Y�<1�.�L����حwZhE��B�<�
Z�J���IXʺ<9��Xw�<��CT�h�ReP�kT�U0aa�p�<i���;|�!	�-������@l�<�ud�hD��#^'}R��4kGf�<!�^+Y����IT�n&��s@b�<a��� �H�`�.�$@xx�!�B�<�i z(��H��X�����<��'����0h<A�H3&{�<і�<@�$�A���:��ū	}�<�# ߔl�Z���Cg;t y㩜v�<!�ς7Sj5#��.,H(�@���m�<�U��H��a+�	Y�T�z�g��n�<i6KV0'��`F��:-�!�QV�<�0Ȃ��:�AQFv��9� �]i�<�`��;0n�e�1��G�d 2/^�<I�%��iq�X�2��e��/�Y�<��i3�l����1�b_W�<!� ߦ}>6���'�1�5x�
]V�<!��K��XX��������f�U�<��/��F����#�[��R"�V�<�rāY���9c%�z@�I���_Q�<���O"���AQ@�4�HAK�)�r�<��A��A��d��m�pJ��Rt&�z�<a�i�=�>��^�>14("`�{�<���c<� *��+}��f�y�<���!wH��dQ�@ 'g�{�<�b�/Y���YpoŜ|��8���{�<��aL:T�Ji��hMl^\M�k��<��Eȯ
�ḷB�;����IB�<���2Q�:��Y�QH8��S�<�1�^�:�΍���2��%@t`HV�<�wA�4fv1���S�0~Ȥ����P�<Q��@3���N[��aGw�<� �=�cH/�LG�V�t(��Y�"O\h9 ���9Ō���	�xB�H3"Ouq�f�� ��ؖ�5/�3b"O�%Q�k�q2� �#	Fe�e"O������59�����2���"Od\��&�C�1 �ȚI�ܵ3"O��y�ъ���H�Gf� (�$"O��`l� �l��2\"s8�!��"Op����C1\a`9��ė+��H�"O�Y�s�g�eګz����"OT�A��
?;<����E�%bg$1&"O�djC�Ј+x�4n�� L��"O�B��o���c#�bRF�HW"O�U�v�_G>�#�US�NH�C"O�qsħS�aK\��苸�ұK%"OT�Ӆd5�*�	��۵9ш09d"O^@�V*
�M�\Y�%ŧhˀ��"O�H`�A�R4i�!�#����y2�0Y�8((i
�N'"��#R�yr��4��5�a�Y�І�SU$G'�y�ꟓV�hc����� D���y�)rZ�ܓ�B�KYJ<˶�y�lXCA���	>�:�p#,��yb�>!.iy� W�:��|@�f��y�I��rS�{��=6��h�4J� �y�d[�=?f���M�,�d��)�yr�6Wh=�(�(�&���O�y�.���� )��((2�3�]=�yB��u�B(r6a�3tn�I�sӀ�y¤�.s?��wB��q�ؘHsɛ��y�E�)̨����+5;�$��ܷ�y�#["pM��a�I�8/�2@�,�y�(�4_	��1g(��1�X� @��y��G�k~N���s�Ăg����yrVWfT��cBӶz�d����6�yl�A�z�(_ x����؈�y2NظC��tB��	F$|H�wA��yR��*$�����b 	1����Y��yr��<NB��*��џ X��&�P��yB��w����KB�/8`�5"J��y2�3XLԲ1bu-�;dn��y��T�<3<���EY�k[0��TN&�yb�ms����Cf7�	sĎJ��y��x��-CȎd��a�ǚ��y��_)�`�%T�F�a�d.�yr`�"?��-�!)թ:�����y�E3HWJ)!�A�:U���g$-�y҆N7���3$�(<�����y��gK�L��
=�$q�FL�;�y���z�|��`�ȥw�M�&)��ybjB�'Ҵ��.ߐ32<�����yVG�D��9�� ���y���p���0�'I,јsEɲ�y"� $�"}K�"CI���;����yB�\�?����'�	LD�h�n�1�yB��X���Yӊ�*ێ؃ nN?�y�>H��R�Ԩ,��<r�+���y��N?i�ԁ����*_h5�ϐ��y"�BU�j�pr�L���Њ�yB��H2l*G.$X�ر����y�(�`�M�%�V�OZ��MМ�y��޽xd�lx"�[�;����F��y�L&t��a6���/�
D���y�� ���'g��p9b�Hǘ�y
� "hE�	�vL*�싉��"O�u[)��}wRa ��L��q%"O�����Y�L��ɋ�� $�u"O^��V>>�]���s�!f"O�0����MɂJ6)V��B+D��z4�I3B�P=��%,h�j̐�+D��B��U�k�VIk����b�"�*O:���xԾ�%MA'T���"O(a����5�V�
0LI=\,j� �'lḀ��LM���) �V%FD@�'�Z��@	>u�%f����'�\����Z-�jP q
�-�25��'?$�9`蛸8����`���\�(��'7TlL9�]3.�?e� ��'�,,�lJ+�
� ׈�T�vY�'�ܩpWo��N�n��#�b�8h��'���Bo��(��%\����'����N�3��<�(�M���(�'�.�G���t:�4�0J�=u�-��'i�����W�dy�.���%��'�a�%D�O_���G˖x��|	�': E����C����6NQ�y�~D��'�ҹ�2D�G��4�u�_0j]�!��'����Gd�dH��ɷe���k�'�@q�@��Br$9�Eh��Z��p�'0�5��01�(��"+O����'�X����ܧCD�̂�፶@�~=�'���&Ё��e�G̙�4�Q��'4��6���"fl�F�L�<�:���'+��3��s�h��7�L+[D`R�'Q�	[���:�``�����'�����١8��!��h���r@�
�'�X=�TIХbP�����(�*�8�'zj����xJ����K�<�{�'J�)X��)6��L&P��ɠ�'@����Xɾ���$�{�Px�'�Z�7���1�i�4��kX����'�൲�Ȗ���Qs�ƆZ�µ��'-��S".�O�:e�B���U��X�',��*�2Z�2%˖�R�Nx��'�#�ě=��ɇ�J�z�&��
�'�ȉg�� >�(�ŋ�^� �
�'t����FW�0z�ώ�Zd�(�	�'����%�¢5��Ek�hϫ[j�5�	�'F����@֯H�P��)K�)�����'݈�h�&�|` �wE�
L���':p#���(�*H�7"�;4�ָ�
�'�0�A䃙@���@�
�<B�H4a
�''"��Vr0΅��ډ4Dt�"
�'�lA¤�_���E&�<>꬀	�'e(5D Q>��9T�F<>��\�'�D K�CY�Sh�<$��>C�y��'�r�yW��@�ѐ�-D�>�9�'��	g�V&p� �g��;�H��'2tx�	��LE�g�Q:5~N1�	�'�"`a��S��Ha�M�`���	�'��v�+��%�f�Z$�
�'������(�	ыF�~��HQ	�'��|����	�h�`��O*�\Yq�'Dp԰��5t��e�B)�{*�k�'�����%J��T-ɡ�c����'f��ڔ̕P�J�!qD��a��A�'<�IB bEF<�0U�05��Y�'��XUO�i�uPW*
������ ���G
�Y�<��BÚ�D�9�"O��!V%U�3N�L��`A��I�"O,y���+2 x� �cF1\$���"O�a0"V}-h�K�"YX�ɣ"O�<�3�4�zreC�5-nP���K;�y���*�a����2�����y"�Ж-�`�ȩ2�@9:7+ҟ�yr�X(Xv�p�LF,2;�����	��y�@�,3�T@�E
#������Q �y"A�r�9�0�X�j$�1+4'�yB��Cрi�T��M��1�8�yR��Q���Z$�GO[ta1�°�y�'��1���zp�D�P��A��y2�ہO���F�<���8M��y2�ޙ:nX��������
�y�dU�U�v��P"Z�U�IP6
M�yR�7�69)��	�RX6��σ(�y���<��C�'�>Hl���Go��y��ޠ���z6:Gu^y��h��yR�H-Fg�%͕0��D	����y��,8\�VC ��eX�,V �y��S-=��=�vc��k��]D�� �yb��N��b�Z�9��A�'+�y�aU�UNX��Ra��Hq@�z˚�y�ɂ߼����N�k+�3�L1�y�aա{�B�,�;���)e���yBlB,�nP��J�!���!��yBO�8�$�x%.�8�����|��'������0Y����N�m��#	�'�����F@�
^d��&EM�Z�����'��us���Hw���s���#E6���'o�Y�
�
~�8\�b����8	�'�|a���%L�)�gT��^��
�'��(���[_J(-ے'֞=���'0n���H�
oީ ��s�*-;�'�`���柮jҀ�Z�\/\���'�� 	8/��a
���Q�Y�	�'*�,�U;9Ɖ#���<I����'��e���$�i�ȍ�02Ɣ�
�'�ƌ��#[.H���D�$�&��	�' ����P<\�j=l��)0�'2rl)���QV`�R��%rYd�"�'Q�\�T˅�ucL0@5̇�lQ��P�'Dn=���ȴ,r�x�̈́V���#�'���/0T޼HEǐ�@m|[	�'�.�Ja���ؘ�a@=)~@��'_8��Ն��O�:0c���n�%�ʓB�0*�o];��A�(�/  ,P�ȓwl��V琂l��lˇ���|���ȓ��iB�&O6@l�x��Ş�I��t��t�
�R�:p���8��!^?H؇ȓ5�h0ˁ�7P�ըC�H�PE��;0NkF(W�yP�@�呧y�\��ȓa�217K�%s�r��R��vDH���"I
x� �1U�&	9A#H�~�,���C����ث$c:�x1FT
t���A��-I�
�O�JH�$�P	����'}�ك%�@%R=4���E3?np�ȓ+���!�_�'������Q��ȓ-(�]�G��MR��Pg!�)e�&�&���ᑭJ��� EA%%X i��tʦ|aB�� ���0ǄK�:,�ȓ*��%��cO<X��,hW&�P�^ ��hM�(AңL/o�`�c!��K�bم�S�? ���sJ�,,��o(8]Ҩj"Oڑ+V-�eY�YBn�/x���"O��y���<R= @�v�k�zY��"O����<P��`� �W1y	�"O�� �����A(b�2��8B�"OR�:����\:����C:Kw ���"O�ݻ��M:8�-ʤ�!X�5"O!9�l�12~upB	۲P�5�G"O��
G#׮A��(�6H
?8J��"O؄��j�p��)�@-�1
Ab�"O
�q�L�5	�h�*W�&Ԍ��e"OR���lhd!��@�$UJ�"Or�Į�>�z��_�>��'�Vyc O�o�6u���F�n�[	�'b�!C���/O�j� &3%�K	�'����H����Qr%��4<��p�	�'�1��e�,[-PL�fË?a��x	�'PX�p@�2������	%@8��'��ԡsf�]TDh�c�;�6���'�����	Q�0~�t(t˛�x�����'���
Ş]p�P��YT�q��'�!0a����"i�d��Xq:���'��������!�]H��؋?�����'Ĳ�؇��2:&��m:f�#
�'�
)�gٻ�`��)[�Gϒ,i�'J=����}���X�if����'�(�b��v���xǨͨw:��'����8�D�8G+ɀq$�my�'9��pv@*=�ȡ���f��]�'�4�EìtJ�B�WD�0��'����w�<����V�ǆ[Y�\��'trH�c�<��P6� �B�y"�'�v��Dc�'8JSƕ�o�>u�'���� iR�
��]R!O	�_��+�'��9�@�0i��!��NL�E�����'[x�"�c[r+�_#|�*]Õ�7D���ȤFy��0��\$��;D����,I=F^�M;%�+ka�\�ǧ9D�t�C2����O[�^1�X��#D�d��]�>u�|�ė�g�ސrЈ=D���'�?3�i�$LB+%�5��N/D�0�rL��Nݘ|*�E�^0�}�"&-D���rɏ�\�,�E��,���ڃg*D�D���=o(�,R ����|�c�5D�4�Q�_J�
��O���r�&D�̰a��8�8����^�{ fL;�f8D�D����5]Z�9E�;zQH�1'�9D�hPwd�%X�J�+�@�N6D��r0��,@f��]	� ԁ�+7D��`!c�#w�$�����i�Н㶉3D�X��ЬH���%��_<��Q`�0D���	� m*�����)�<�A��.D�|�c�'?~�(���H���P@l2D���D � 7M�y��ʚ7%Z)�!$1D���FkӕV.��!싦9ߐ�H-D�A�=D�J���2�Z�J�6D�4c�l� '����6gP@!0D���`��C�v�X6��e|�q�`�8D������_��|�Æ�:��F�$D���2QǬp���09�g�c�ZB��671L�9f���5N $A�X?|B���v�p�e��D�,�Qѭ֒`�zB�I#~sV���f��1`�dk�oZ%E�C䉮f&���GLY2H��ġ4�!g��B�)� ƽ�'��3�8�$���@�0�g"OV�)�̄Y�aׅ��$�x�c"O<��"A6�d����׮��2"O�q	XMCF��b@�B�h� P"OR��+�tE�02�G6O��X�w"OT���(_t*�2�ꂆT�,1�"OtU��Fo����v�D6|����"O�$[6�WϪ�E�\�n�\)Q��y�<ITZ�
��0�&v|d����a�<P��1i�&��M*v�0�y��^^�<�g�Oˊ�K��ѧQ�M�eZT�<�$y0u�g��&�Ll� 
P�<��BC�j^��is� 9}ٔU
���J�<q�θR�����͸%��:�F�@�<9�� �1�HE�W)^@�<����.Jo�9� @O�Rؐ#T/A�<i �/�F�P���C��t1�l\}�<�@�;s���A#/#E����!�|�<ه�_a�2�J��7.\I1"�y�<��&^�m��x�W �0Zɰ�`@��]�<aSƁ1@h�a[���S�����a�<٦�E&r$�0���*A��K��`�<�7t�T1��g=.�mK���Y�<�#�  Z�
 ���3-oz3��m�<Q0ޗMTfH��i-e��r1�j�<�'b�"����)JZ�=b�@O�<a%.޺HhI
�αGS|�e�q�<�7�A�3:1���I�$�Xl(��q�<�BQ&+4�CF�,_IX��&�Gm�<aUɞX�v`zū�(V�\A��g�<��$Cj�d���M�{a��Q��`�<Ap�7<T݈"
�H�ޭ7�`�<�tmr�Na��ȈJJTI!�C�<��8����$�ȆhL�M�G��w�<a
S3k$�����?H:2�+q�<і*�uP��E�
�8F��a��n�<�ΐEZ$9���1�2��B��g�<yaۦeV�	���`�\�[3Ώj�<�0I1\���'�e�b��&A@�<�  ��R0(�JR��a���x�<���A�,zĄ�	!�,#��^w�<����vP���%ΉA��/Zq�<y��	�RI���"O��zċb�YT�<I���=K�=pbC�q���C$iZG�<�-�oj ��+�,�0-�ʊH�<#O��D�s���<Hik�IH�<ir癳$=셢��<>RV����B�<��$ @�^��;a;�H��G�R�<ismV�!RN��V�L�8~�4"�of�<� 'B�h��͠�iE(��Q"�	d�<��O�i�<��g��o�<�-!��B䉰���ȡ���Ŕ�P���%f�B䉑,X)��ς6S�r"�H$W��B�8v[��b���*%�bH	r�9+��B��bR1+$�V�T��S1 	�7?�B�	;y�h{��!gL`Qf�I�1�PC�	��`����	="ؑT���
ЈC�I��;6������ǁʹB��,�!�+�&�x;��=69�B��d� !7� �����rB�%h��B�( (�÷�4�P�����I�.C�	,��4��(^�S^�11�!ٌ[�B�	�
G��:�J_�e����%i�;!�B�ɜYQ�=�R-�7 
zE
r�S�e^�B�)� 840�������A }j�Jv"O���m�L�f���*� /j$("O���&��u~��Ӌ��2�X�"O`=���^p��CJ	�`� "Ob|r��"ZL�q�I����w"Oe�%)��$E@eP��ϳ,
N(�%"O��*�%F$�Is�?5�tcS"O�����P �~���f�	e����"O�Qq� ��7V��S�ՆdK�A�"O�Yk ��D�`b̀+05v�S�"O�8x`�ܹ˶�i��.%�u��"O��R� *\���SD.�A�c"O:�k�����Z'+@�3.�l(V"O��i��V���ZD�#&��"O�EQ�*	� ��J`�V��2"ODt[C��(W�T��,%$�zPz�"O����ǇqT��΀*y�\��"O��ʧ.�2,�u�E8���Ya"O�8���`4��RR3 Fu�"OF����<f�ƱӁ%K-�"t"O]�B�{��� W�O�	�6"O���ID�B��^��Q�,T�Pz!�ށQv�;�*H d��%酊C�$o!�
�^�R!�sǝw�2!I$�6o!�Y�
��<!���nv����@�!g!�d7�0�SE�ݓkj���1e�V�!�D��iY���F��)p���$ f�!�d�^y֐Ѓ��n&<)p���R�!��K�t��4D;ujV)j���.*^!�$6���%��!��H�0�Å`�!���T�t�a�r�ܡ��阋o!��Eq�����R<l�$�G	O	,�!�DH
��E3�i�\���] a�!�� ���$/�=���!E%�j�!�$_�}0 	J�J 9B!�f�HR�!�HB�~x�O�.jA� (��q�!�[1'Z�{%�E9?�2T�⨖"b!�dO�5f�e1`*Ď	���Ș�X!��
�D�x�#h�.�{d���!�dK�{��y�@��d�L�(�!�%� ɔ*�	��iJC"��a�!����  �/b $�	s�����N��c(
/ B�%�S���+D���sK8L�L(��ӡt��MҪ2D�Df/�6k�� ���$= �0�0D�d!ck���l�s�Д=x���.D�8��΢/�4EIE.T1M���&�8D����ʱ!U$��p�Ѯ?���* �#D� ˷n϶o��`B�a�t��2�<D����ʎ?1C�+�#ݐVw��f9D�l ����"���覠��z���0)6D����S%�X�Yt��o�tA{��5D�ĸ�AC�u����+ׁ"���"3D�ȃ�aĻoɤ�*�F�1DJ�I��/D�`�ЯZ��R��4��bu"��2D�X�uX��B�E�6X�:œ#O/D�����!�P����E�{-,D�ԁ��\��,ʓ�T�,+�4��+D� 0��S��P�t�R�u�� 9�f&D��)��X	���z�m�`d�Sր"D�^��M�o��V3 9�2'D*IOBC䉋RǄ ا ��$�
Ѡ���QgC�>hO&*�Ѯd ��fK߷�PB�I�G^jQ#�n	�C�2i��n �7`C�)� �P��+�x���YX4܊R"Or`�4�B�5Q��"ÆZ�7R��R�"O�	��/�&lUTe�c,��jWv0��"Oht�A@K�l��6�	!nQ�p�%"O�b��85��D �$7JPZ�"O"(b��H�8�(��ƣD�T#Bz"Oz 
�`D�	$���!��N `8iu"O  ��֭lGV҅
*`��R�"O��%� !c��i�)�5��"O�x"�U�.a���;b�ސ[�"Opݨ �y�٫�HGF���"OT�;f�Y�<	��Ƈ"t����"O$���+T�1ִa1��[�$���"O�hz�L�"�9[���j�6͹�"O�4��Ⅲj��x�0R�Uך�	'"Oas�\�=��,��L�"b�,�%"O��%�_*W^d�q ��hP�T"O��!7��k�葱�ޮ*	`�)�"O|�(�@ �	�8�U�2J���S"O�����-R�<��'�?	�|��R"O�p���Y�"�1�@L ����y�F������%G�m>�ٳ�b�.�yB�5ZD�Cf�ōu���5L���y��C��8K�kXj��4�Wj���y2 \a�T8+%�@!b��87���y�+?IH��R��TܬĹ5��yrM��fg�����Lpv���A�3�yB�C�NEΕ�A/ʐY��A�Mͬ�y"�\�%�,���E�~��H I�y��E�0���Yt��)��!�:�yҬ�>G�"G��gj�QgcE#�y�i�6����ŁX`�飖�&�y�i6/����ֈ� J�<���x���	Is��?sɸV�<$��A�&"Ot� aN\�WX���4	�?��|�A"O�2W���� xء�ھt��컔"O0��- ���)4Ъ��R"O�8#Q#F/D�����	���!T"O
xg!��G�<�D�FL�G"O�����_�| �B�)^c��-��"O���\7sE���i����a"OFL���ޤ�hd��G�2��h"O���c"rIC'��X���"O,ya�mH7V��@�Z�V�W"OT�(�Q�#�Dh���\�;��=c"O>I����%N�t�ʁ$S3A����p"O2�i�.���"F߸b�d�u"O�����+�dI��w{ʡ@3"O$�ׇ�_�pC��3er�I�"O���R��\���cDpD}k"OV�`cj�!v.�,��m�
Qp\�"O�8�V@Y�WAN=z��.GB�)3c"O�u*�+�	]�ҽ���<d#j{r"O�����{rk��13pLB�"O~$�6���@碵�`
�L��"O ��[��Y��]�\�0�u�4�!��8[>�Rv%�h�޴���'�!�D�1����6׵�Jw�V�o�!�O�]�N���^yM+�F��@O!�D&(hKQ�O.{2ֽ��؀SJ!�ĉ���KJG�vٰ���97!�5��!��M�/��	b�Ѿ^!�W��e��[�z.��-Z�!�$�ih4B�F�3e��B�ŦJ�!�� ���jB�.~u�0f3I%��Z�"O �ٳˇ;ܸTS�G�?V���"O��)3�^��p�ХbD�� ��"OB�3�̉�&���ے���6�Y	�"O��I�XP��`B�G�&y�ej�"O���E�=!�T̚&�ɶb[<��"Op� ���skl5�W�� %Gd4(�"O:�y���
p�(u��+(	��A"O�4�!��4g����0ə!����r"O��3� efp3R�����0a"O.0�e|�k�l�
^�@XW"OLT#�	�Ncz5�Y�*��Fc�yb�֗-���� �	�q���E-'�y�"�����`�S�Q�L��EG�y�$΄xD�[�J�R8p���σ��y�W�C{0��e
�x��C2G��y2���
�X@�$JU� .n�0_��y�lYr�}SfN}&:��A���yJ��.N���5K+y�DL�Ʉ�y���<�6̙c�T	[)%B/�yV\*IAP�˕<:���?�yr)ި�$(��'H�xPp�ig�Z��yR�U�N($H�w��pBg%V��y��
&6��r��p""��v���yR�׈$C�,a@ȋ�� �X���yҦ�f�����gg����l�V�<!�/�e�0� U��JL�q�r�K�<��Վ0ZEA4��[�",ؖ(J�<QďB:8^��� )�ٜ����_�<�f�/c
�u��I^1!ĉ�!��A�<��L6<��܃�,K*t��@`�L�<��@�� �v|�֪$BE���R"�D�<!g U�"�b�㵬Ŋ)�=iw/�B�<�F����6�#��	xY����G�<�d@�BQ����,PºZ��Y�<	h*LCX�����*R���q�fZR�<�c� ��`U�&,�D�4�Oh�<-UZ.x�A�;H�4�دL��B�Is-�݋BnF0}��l9,�5��B��;�p�FdW�/��h�- 6U�B䉍h��yk`J� t�a1��t�^B�	5FgZ�`7A�(H�Dß7U�B��I��5	׉m��Ks���AVB�!~���9v\+K������1v>HB�	�M��M�CY�6�*u���>@�B�	�n��c�@��� c%K9 v�B䉔>@5���D1�#� M��B��8)N���U��d�jr@��6	�B�ɊdZ��V��Yt�=IՍϖtC�	����7�4����R�M0�FC䉌|��d�`�v��A�a���O��B�ɕNtx	�ϙn�r�Ԁ�K�B�I'5X�A�-[ kόx��Y/_�C䉱��"����x��`E��5*�C�I�Wg������w,��Kq';iҴB�	�&J�uHł<��Aqj�~�:B�Ip�:d�T'�C����	�Ey�B��"F$ r +��T�@�I6��kzB�	�B�^������r�%��c=lB�5 lȐ;Q'ʇgQTq�a�4B;hB�I+}�U�d�D[�D�ƀ29�C�	��J=���9<����-8_"C�I�u�N�cG"��A%�̊�C�B䉢�����͊I���iR�ߢ{L�C�)� H�)E)�pl�����)K���T"O�K�M�Tʨ=ʃ��!!�jT��"O�yS �'#�$�y4��w�i�B"O��Y��>�$ ���&LZ�T`A"Oh����_�W���0��0~���
�"OVX���K�J"|����?0��M�a"O��3W��~0���E��:( "OF�!0HA� �$E�$%�6'�bu8�"O<���僀N�!�d�c,�x0�"O���dL
W�v!J�h�:" ,���"Ov@��s�LY'���r��ې"O`��F�ɺZ�����j�I����"O�m��Iޟ]J��!��6.�x�IR"O�CR��Y���Wǲ��"O�D�!�B7O�I1���G�9ç"OLKB��IS�=`@���\��|��"O�p�7!��|�,!�� 	a��8*T"O*��֦Y�7N���`��]�ʐk�"O��z�C�.M� ;��^��h@"O�e@��m_숀#Bڍ#��"O�IP�.�d��R���4]-�y��|���m���'� P�Q����b(6 �,�"Od��.=N�b5Y�ȇ���IEx�,�fn�; 5X�e�6b����/D�8R�a�u��MZ��̻O�أ��9D�d��h�`�%�R�I�<x�yp9D��곬�>�9yՊ�9ysBLRl9�	o�����JƤc����&Ĵ�6<1�7D��3�J�[���ET!"���
!o5D���u��#��m7*S�ae�h�1D�t���GoLy��յmg�њs�.D�d���>T&��$*���]�gm.D�,2d*K�h�,��
��I*OV�Д��IJ����V0� �"O�M`��ږg�©HK��?��lsv"Ol]��n�6c�t���
]9(�<�"O���F���h��8))6"O@i��P�(��A��Bi�v�+"O���F�a�(q��9�� �8�S��y�R?@K�5Ӆ΄�$`�H�C���=Q�y2�@�%�P1�t$�j �Bw℘�y���*c�z%���([2�#6׷�y�K�~�������"�z)q�d7�y�%U�<Ŝ%� �͂1��R5!���'�ў��.1z��י!~�ԙ℅�$�� :U"O,43���88/��{S+%�`A"Ỏr�H�>r=R�U�'y�dqu"O�� fkV�(o8��c���p�(V�'�!�䉘vLP,��7.P�*��3a{��Y��/;�`��i߿P�Z�[5��9g�C��6y���-�}�680dB6Y��'���O���'��~J�#TJV-q��V�(z�����E�<�m��I���dD�<�Ls��J�<�R��X�>PE�������UI�<���|!GJ	3����RĈm�<I#�,K��QS��_�2�r�`Jl�<9��	:O�MiK��Vg�l�#�Ig�<�d�V����K�.����%IW�K[!�Ď�4��)AM��a��AE�
�z!�$�'oܘ퀔�ǍcKa�u�> n�E��"�g^O�]���?Ku�T�6�.D�8��-Եdk��صl\�B��hGd"D���)��kbVh
�/����@��?D�@� +L�]I�p)�,ڨQ��4�N?D�� ���6�Şc�0�Q��2"E�9�&"ObQ�����@e^�a�I�}'&UZ�"O��`g�	3np!�	��.$dM"OD�qj��L[�HH�N=�7��Q�O���B耡w�l��$�~u(��'��XR�S��V���
9xW�i{��&�S�t�ûl��3�jίiS�Qy��أ�y�b�(E �YA#F�9K���VG?�y"kE�f$� ��8���y5	M��y�Pp���P6���2sZ����C��yr� �:y��JV�,�����Ǉ�y�^���X���*ph��3�yb��d�$�xC��5q��x���%�yRm��J/T��'߰!�ܠ���!�y����X�����~��j���yb
T����r�Ǖ"t�8�#����y2��9�@i1
W6v��,r�н�y��-d����*�h�B�����y���>f	�PEA�5ن��O[��yb�Y-~���+�' T$mr�����'ўb>Ea�Q�
���a&���l"T���)D�|��*�
�m'�@�D �m4D�����~F%�P'H41Xr�R�.D��Av�U�En���B�4+�``��C������
��a��@.D<�2pΟ
u١�d`��M�D�ϛCk(��`@,u�<��"OP�C�D��D�#���j�<�R��D0�S⓪*9�E�En��V\irC�g��B�
��A��=lH-��g��B��(,��5�q��=_������J������<Q�M�'s�:��d�йl����\m�<����Q��k�-K�-[���1�Gj�<�i���`=��A[� �y�*�f�<����	,�޹At��5I�QA��N�@$����T�q�X��X`����&D��aQ+łc��TnV�b@�R��&D��p���4{v��w@@Q��2�Or�')R1�@	85�9ҭٝn��B�'#,�ʀ%}���KaO+;=�,��'.�Ģ�$m�I2�o� {@\�'x��O8���e�ЦNaJaS�'*�S��?���ߞLt4bՃƪ��p���<q��t���;qC�)MO�PVn�p�<�ǋU�|Dva���%:���]q����>Yq��dQ��+�-�$��<�
��UtTe�~�=ٗ�
�G�=���~?�d�X$<��9��K�Ѱ��Le�<�A�ßM��x1�	QSt�0���e�']�#�s�N0uv�"o�W�&%h#�I]�<� �] $QK�`Q?xXN��&s?qJ<�O�>Ie.Ҩ!K��2�[=~$�M�D�2D�`�e�܊@u.�`�J�&t���8��0D��Ⲇ�5Z�*��*��+T0��l�N0ܫc*M]�x���݀�C�	�n�^� �R$EXA2�ڤ����&��ߢO��lS�&ЁT��,!O; �!�$����!g��w6�$E�3n{!�ċ�y� � �9>=���U(Gj!���%���)��̰x
�BA��!�$F#��@gZ�Jژhsa�2\�!�Z0'�%q����D�c Ӵ}f!�ē�n��[�"� (�V��N�zO!��S�u峠��6#�J�X!@C�RD!��V��)#T8`8&�"���'�'Na|
� 4��" *�n�r4#�M�pic"O�̚���N�6�+�B�J���x�9O����܀_a�9贏ބ�E�ꙍY��b=O��;Fi+�0�3ra�)a�R	y�"OPa�AJ�=y�c�@�L�����	B;B#}��f��� �Țw���bv�<�v��3F?��ۣa�]�>�م�|�<k���<)����2�̠z�kL}�<�A��'G��[E�D�%oH	(�fw�<�ҥY�#�fJ%���l�@��Qv�<��ۑ8,z���m�.�����|�<!`�*#�T��EڍKQ�lʁ&�A�<�Q�ׯE"����%*�>�mR�<i���u��Xï��e�0�����M�<�ς?D��U�s*X�7�t���hI�<���CY*1(S�L!'�, ۂ��B�<�o,8��1��Y��@k1(�e�<����4k�d�R �F|A��Jd�<�PY%@����eH�^)3!��]�<�D�5\�r�Ŋ�,/�1��T�<���Q/&���P��45�!���Q�<�r��v:��a�aO�aĨ�B�Er�<)p���n
��х�*J1�w�k�<)G�St(��	]>����Dd�<�WJ�!T�ѺAFD�h���X�\E�<9�k��Lv����X3.m���r�|�<I���<o�}f(3H��ffy�<A�l.Rp���p ����l���}�<	FFǑ�j�2�M�4,�]��R�<��Oȟ/�V�fˎ	@8@&�Uu�<�F�A;[��+��՘H*���kCr�<���q?.	�ʅ28$�[�NXf�<��b�l��E�7AX(��3E�d�<)p�1*>A���ljL[�h�a�<�-�X���4~'.PsC [�<� Ů9�jAS��H����J��Z�<�'�/ ����W`�u�ƀ�6"�R�<�V �:r9[� ��;\Y2�D�v�<q�f��dl�@p�W��4��f�Tz�<94�>s
.X+Da�G"T02HGs�<١.O��$KG��jCV�s`m�<�!!K�5S ���hH�kD`1K�ll�<�P J�=����W.�7-L�5�ǫ�l�<y$ꈏU��!�n�2WwVy���e�<)E Q?Fy�H�1s���� f�^�<Q��O�K1��^��['�a�<YT \�dx���ƐdrB��Bd�W�<)tb�@�� U�"r����
L�%}��hS
�E(������8Ni�<��A�0!)�&(F8+��s�B�q�<���A�k��8����0��c�K	l�<�o��i���R�1��L�`�<��,�-MH�ے��2p�B��g�<�G�:C�Uՠ�/
��W-�\�<��aVO��H�*�8'�a���\�<!2�ȟMk��mƍB)@���)X�<����]��Ր�-_s����1�L�<ADFQ?60��i���B3�FQ�<i����w0�-s�d��7��AbanT�<a��-��5:���3e���c��U�<��o�|Y�P��d�tE���H�<	@!��W("�9b-Ԧ�ݙ� �R�<@ʓ�K<�BD�D�Ig��L�<qW�� |8TP�%ϔh���bG�e�<�V-�7������6����'ca�<� ��F�O3.R�I���FԚ""O2XnSs �+�nԕuͺ�[�"OX�&�TT�T��N>��Q�""OP�8��CSY�\[7f�06�BQz�"OΈ��H�i^��1K��JFHQ�"O�����a<�P�D��Ъ�!�M�:ހ\HÎ�0D9�X��`�s��~"�ܣ7S�ps��Lsr��^�K�x��E�J21��C�	2m6�j�(X�f h�ȵ�ݬDc�">Q���RIk�l�M̧q'6(#����L˲�i6�n��ȓ[�.�D�����a�I�~N��ɹ@�Zp{P+�U�\���O?����/8�YS�b�[��)�1��G�<!p� Q�r5)��Gj�s�־�$P,U�|dAD@��4`���HO$<PR��6˸|ZÅ�ġ��'JF$ ��V����PNpR��@��\^��K����y!E+�Ò��I��E����S#��t�J���.Z �)_@����#����z2�ԢG��#'�ńQ�"OV�/������Q�{�M	BjU���`	��)c Y��ؕ!�Q?�$��8Q8��:'V�,�P��7t�!�7@����s�"Ql怙��Fo�4aܴt|��
�*�7�h�pr�?�=Y���	%$P� �8�:�f�p8���d�^$��H����?�1���8V�2ك��\��L�S���p?	�펬 ����`J�7�L]�)�_�'���1e��/'�����-��4�H�O��<��!�$��� t���F��p��'�`�H&��y%�ِ3C>�޸��H��g��}�b^�>^&���k+訟r�S�b���&�7z�8�U�ӥ�y2�,aPԝ�#������ �x�n�1Fv�±#]��@��qԟў`��	̡;�
\� �J�t21(#�O8٣�"
.Dz��ýQk.(B���		�D{�]y�*�#�fb���!BC�$|q������n�T<ڳ�>ʓ<���i�Ì�z|��%cl��'^�d)��M#�y���Ayc|@��`���PD�1̪�㑠�.�6a�I0�T�As���ȂKv��?��k@);���#�J��t���{-�l�<�dJ"xzT�b�RL�����N�F7M��h�L,ê���L����hO������&(Ӓ	�"�P3hp����'��z�E������T�NzV���d%<t1�uB�@T�L3�H��h�X�;� /�l����<l]�iF{�i��T��]�g��9� ���	Z��#i�@q�fЎ
�r���"O�		&�F.?H�Se��-f(D
 :Ojx���;W�rԚ@��"~�B����#ݔk�Ddq�OKC�<!�	�ny��@�KM%�D�$(�z��ך-H���%hz8�P�Qe��B�����ȵ.?��U�;D�`"u$U�B�n����< �<D�<��Ό�"E<��f�O azT�a!@7D���-I�er�BE�7�B2��8�Sܧb�܄�#J�}L���A;@x��Z��jiڶ6���
�	�"^4��?i�E>x��%�$7��H���D)K���Ɠ3��6����� ���ۀTDZ�	�'7ʸ�U�����t��Le�U�I�|cG��1��x��On"<y��׉0��"  T�xD��D������"�F��*��dI�eAgFK�k�T�"�A�`�&ʓ�hOq��,�ۛD��|����fx�� 3�̝Җ�84�(i{O~da��/���kF�7DMJh�C��Z�<Yw��Bjjycu���|2v��%�צ	����l��ɋ�F� ��)�禝zЃ��[I�<{���$W��Ub%D�h۳�̱_\�4J/�sk�	´�7<�����E��A��N̵E��9�g�'l$�k��'a���$L�>��L:�`!��(�'�3������H�=dD�>25C�Ϫ[Ś8�&�Q���!�	�4��ٛ7nO�og�1i�b!�I�'�V0�Ӹ���N>us�d3��|����3;�`��P��6ڲ�1G��~�<�U�ӻ�j�B���Iq(�I�?_`4� ̇�c�����Ùp�������9���zx|!�Ѕ�L���2�9D����T(K�lQ����z,9����@��d��(4�c0A�U���Ti��� �)����=QN踁��V�N��m���'rx�:��X=="\+��=���XU&ӌk�%I�i2
�!K�Vc:����nE2Vk��<���!ͥBB��=٠fҠ"�	��S2]t���ֲn"
�П$� �i)����ks~h��"OΩ	c�ڇ7�H�K�o�Ho�`����5�I Sk�?s�<�D�H�*/ĥ���dC�yW'��1����0�2k�����

���x"�R�/��\8Sa�6��@��5+A4ق
�7L�YA�B8��a���R�,��x`��D�t|>�Ê�v��i2i���y�ꘑu��1� ��J}17gW3���(B�ʮ+�f��􆔭jh�I�
&���
�:z0*g�����E:�-�U%�LqT�(�a�Sg� u��BQN�'�\��N�?5�⦛KE�,0����9���Gj?D�����#Q��QT��	ҺT:���� �ॉ�B�2}��
'%��7��K� ���]^?�����8R+������.T�C�	1sv� �LУFF��ɥk����zw������[�����jJ.qx�xq�1ʓ;�|-�rk�"�@�AGDG L�牬 �N���͇H>p�3+�N�PŬ�]�0�A��_M&���M�SǨ��I3�O����eΣ6�4͈F^d/Vq1��|"�ޅg&@EIr�پ+Q� �Nk�m ��՗����F>j�.�\G�0��킎��B�ɃxX��ؖ�ɴ@�L4�6����W��k��psD*�k�,�p�*�yY1�:�0��n�Y(����&X����@
��X\$��@�j��H��$ʟ7f�z�jL?BX�6
�6A���f�* ��p�Ca�h��`��$_e�䠘k�d3��D�8�y���l�@{2�E
>�a8��� �U��J/.[4�3#�0RQ��IP۔K����dçU�С;FF@�Q��hA�e��^�1O�da��S]�"P�j�8fo[em��U\�S�oլ��	Q�����z>�U��"O�,S�	 b, �fn�@��X*��!�����$�(� �
6(�E��¸�h�e�h%�0��*޽
	 ����'D��Ҕe�y������2��q�D�)L[�Ű���M��1�1��6BOL�=��}hF.�/xs�8ѐ�H�_�HŅ�ɓ��d�eI��e�S�������
XY��S�#49�	�[���q�`ɯI1Jٰ�KבgV�Ez�
N-Uf��K�d�%�hb>�#�H�2���G�A�p*p��+D���0BR�-<>���A�8��3��O&1��C�a�h�����0�ƥ�kV3c�:Pz�*�~Mfц�Ez�f�G	=>��I'��vb�:(O�� C��5m�ȑQ�?#<���a���6A	�W�����Qx��	!E�Bg��@çιb�v�0Dd�s�.�A&�L7y�;��'��0�v)�-
|t����2)WdiɈ�dC50
�}J��^=<1H|��'ϰ) �E{��H�7>��Ї�~�<2�O � �� �� �(�����A ޥw���3��c�����iPt�34i:So�Z��y��}�<wƓ�%[�N��:e@[@��?sd>��2'�D��� �8���HO8��!���O�٣�C_���	�'�����b�%q6~�
��ؖ����D�Qp�	H��ګE��y�P�'7R�hbE���qc���[�FM���$�5�~�r �s����:����SjYH�mH�\���bŔ�y�j����nI9[�ܘ2�+�M�q�?1��A�KW!h�c��sӞ1�tkŤjs�hR�P/N�&	{�"On�Ս�	.�����TT�d ��M� �?�B�>�X)!�G�>��3�8�~5���!��a��IV>|�V���ɬ}�&�2��S�#s�D!�o��'Ch|��̣N��*�'��P��]����V��XA�ǅ2f�J�C�ߍ��=�.�;7^ �1!lY����L	��G�	d j�B˥m5���"O��b'48-<�d7��� �'wfL��S�C�\aF�z?E�dGӃ,��
e!%jENM�b�Z#G�!�D�1] �j�@?y8����0:�&ʓ ���8��/����O(��F�H�~��i�Ga�3,�,��' H���ۉy�$��!f��	uB�s�؂��`<���t֡%�$P8�ڷ�Md�'�t�I�&�T�c�H���� ^6��q�/��耆ȓY �;6O\.(�x��0V&�5�ȓ_�H�(�fO�LN��DƶAjȆ�.��U���� ��hIgĉ4��0��U7�Pi�OO�I[�]0F	���z���S�? V�C�G]�;4�����;��eq�"O���� <qtt!3�=	:y�S"O�5���J��A H�U�a�"O��R��'m�.e��Eh�A"�"O����5IM�Q���C>}H(�@�"OȢCo�d�F�ۃ!N=H@DY�"O�lA"��fDn0`c�S�R9�p��"O�u�T�#���j``�,9|@�7�d.\O�mâ�Q�0���5o�;K�,z�O��3V�8�l��	�1�T�+ǭv�<Ad7s��1Z/�0J����1�mX��GybB_�q<��6��^x���&���y"��3Gdt�p#B.���s&�.�yҤ�8�����͔�\�(�-_"�y���c��䈒�Ҭ��"���;�y�I�&�.`�	S�1cڱ�H��y��]���0똹.ZD��FE� �y���\��|��)L�#��\����y���0'<р��v����V9�Py�dJ��=��E�4r��C���O�<�qA�:Ğ50�jW(iǘI����J�<QE� �:Ea�O�%9��-����K�<�K�4;z����S�o���΍C�<a�mʭdozѫb䑀wp@��W~�<�@�>�b����[�e[fu��y�<Au���a9����T�%�mhw�n�<�DJ,K�(h�@	*"��R
�g�<���(g�8�����@�ʈ\�<yPG�"3h�P���'�I�`�_�<��Kܝz�&�X7(��HR����Z�<Y6�[�?<��3�"����b�<���3yXp {�$ơY���!bD
F�<I�FҤ*��p���Yr�ybk�|�<I��3c��9��#��4�D�c#Rt�<��f��K�hrSZ[6���⠍r�<�0Ƌ�_��� �ؚ��=1w
Th�<� �S$\���!`�M�*QTči�<�e�=w{(J���3,�����L�<Aw���-R$�e�w��m2��W�<���LxD���S
�\�����E�<Q h�Lf�T�q.�.,x�H�L�F�<��ń*���k`�G%)Z*Z���|�<�����x�J��� �T���cu�<��KړG[�,�U�X�q��\�%J^o�<Q��B|�s�.�N�HT��i�<���6F��U�`��-&��]H���\�<��T�"b�K`N�/>"=�kOW�<�`� A�b0�%)GJR��w��O�<��H��g�h�b A�{dj�K�<���W�}1\MY`��	D��3cRF�<�r�ڕ*:n �s�
���Z��YG�<�G�U(`���˘o����E)w�<�A���_��h�dS�3c�A��j�l�<AU�_\��"�G�8Lό����o�<ᤨ��6���!��M�=����b�<����?��������|���F�<I�$�-\��I⣬���%�'d�<CEy��a�0KT���Y�c�<���ϔ{T��4@��M,,T���s`F1cf����F�~?�!�F�%D����9�������7�P�/#D�Ds���1;`8;qH��<h,��pI>D�� "�s!��G.=�ܙ;D�8PpKB	px,�g�ܯd�V��C8D�� �(;2kX�,��"�O6p���"O��`�����qO]2L�G"O��b�qJ��Yn��d�|��U"Oj}8���(���Z�.V �yR�S�D6�:��M�c�`�p��W��yR��E�4) ���X�����aۘ�y���JP��9D�G-P��B�I�6�y��
G5��a��V0BΘ(��l���y"E��5<@������F�e� /���y�
ޥ��� N�5��Y�%W��y�+�#dy"t���t����N��p?Y���5��y����W!$4I6��JY|�!c�(Z���'=!�
".��ںܸ�R�	������D�XE�5�� ;�$Y����0�S�H���r��Ͽ�mC�6s��=rQ��4�����և����#��Ts *
�,�juԧ���5xw8:��/]:8f|eH	%D�4�@
�km�lk��,Xl<;�A�3�y�fηU|�պ�&0 ��g�'	$9U�
?6�`I8�l���Wp��C��MGTAذO�4�q���׀'H�r�F^�	��P��'U��X(V�L6�a���;��`����R�� �H�:I"�Y���D�����x��Y�2%���C$I��!��8n��SG�(� ĨV�@9ur��æ��;y޹����n2�C'��OTJ��O�������-< �tP�"Oj(��-V)]?�­̝>*��f���M;�+�gH���#��:���3ړ\@��n�q��(L��Ņ�ɢbR>As�ޔW����U`JTh�s�ƣ���r���|yR5�cK艓�&��`8�����@��~9Eyrj�`B���4�Pf3����� ���1���*�)HTB�hB�F.�yR��V�zHZ5dI+SVbd[�^�"��`Xu�F&SL��J�E4��-)���'�t�!eg9b�1"}"�9S	�'[�m���l�h��1�C���Х^Ʀ��_�058aڑ[�&�퉔"�U�3	= �}ⱃ�9����=�(��C�}��� �Q�@�(����" �@%Z7*������6N�T�*FO�n�= ����D�Ƣ<Y��J�L�B��8k�% ��~jA�\:6����c	�UJ��p���<�Đ�9��Ж	ߺ�T�L� O@
-���[�h��Cʁsʖ	F��!��!��N5�����ԅ�.�T�bc/&�@�3$�������i�d<ҵ�Q�u� 3ÒSF{�R*��em؏.P�)lF4B+a}rL؍k�X���eJv��0� �<%���y�%�.��Y�@���?!'NH�/,u���
�yu�}h�Md�'�Ι;r'KH��r,>���5~�0�"E�L3�� ����G�!�D�`�$�0�d� <��r� S�B���Kΐ*��_�&�)�',��x%̌ |?�t�ei<=R(܆�/�L���b��e�,��hߤf�V�O�tI�Q�H�h���ɶ<� %W@�7b�q�EחZk6C�	;R#��F�&?�v�r��li�B��0v�&Dh��T"�fܩG��B�I( ���q��>�"��t��$i�B�;�<�1A�R�c�jQ�B�	�6+� �NbBٱ��Ђ!��B�ɴx�8�A�o;j2�/�<U�nB�	�{�zy�D$@�:�� 
��pB�	Lؐ��rC�"��@�vʹ*�,�'/<�D���rT�����f�b�7�:iY�d	2��9ya~B�\�
��%�ǟ�;�u٥�4"(a!"f	�~����'�� �(o>>�B�_<w�H����t��g
M�V�'?�C�X�X�Zp��煔m��]�A�*D���i݉5�*��@b�!^ܨ�#Oh�2��&�}F����{��s�������R���7Tj�qY�"O:5�g)��y� � cͅ�K L�[�!���M���!h���)ūwl8�3�r��\���+*��6
�T܇�	6P�0�` ��;A@8m���Q6��0֬\2;@�%c�}Ӈ
,�Oj��$�I$L��V)�D!"����*B��z���$ �x����Vĕπ �C�
���TW��r���"O�IY��ˉڠ`�q����l��`*�f"��@q�˅���b���:��#}:�w<��Fg)&@�+5��s�R-Y�'B<Ȼ�'��Dl��
U�@gѠ�´$�xy~U t&J-V
�	ƭ˫����ɯW.HeBA���"�q�'�a���d�!L��$C�S"X�B��7�/ ��IZW�i�R�R��\F�J �%ta}�㘘^�nakH�i�����'�2�1�HI�����_L`TH6�C���� [��3ׅJ�K鸤�w&��N$B�I�j�^�&���s逴��/��H������fm�d@g�(	�\�4�*k�q��H�?�h����8I�Dic�c��w��a*�O�S�%Xh�I�K��z��,;5��"�eZ�r�J�Ї�1Tҡs�mѧSQ�813'*w+��0bE7'��0&7<O�ĵ"
��a��V�4|<4r��[%0�ƱceٳD���Z� ��`��aZ󍜺2T�|§�hBHLKS�M�kr.�*`��0��jv"�b�A��|st���d73�Ę���S,T�'@B�,y��Nj<�IQ�D�U�(�ȓC{&`Sb���5��I�˄��^A`d�c��aS2��u��+��By�'"���Pe̻��ӥ���i#(M�
VpH�Ɠs���ŇĠO����h�&;Q��Z(�VqZ8��Y�?��T���+���Xu'c�'���c�16]|���Δ7-\�h��7Yp��WnU�*S�T�(A*>�~���LD3$R�iR�I#4��t+9�R{B�f8��P� a+���sa 
$�L3$�D'�^$[��E�r<�4�����,ı`�	�1y>@�Y0eO#j�`��@��?�!�ə^���&ϔ�*�*��g V�u����H�h�R�Ѣ�yx�[(	ޘOj�cw8���Ř!K5j�Sҏ�G���O����̽%�% ���8W��p�MZ�M���B���6唰Ո@�Ұ���M?�HO�4�3@��l��!fE�4nmȠ�R�'��Eȶjdސ��� =�`X�I�R]�IX�8|Gb�:�Q��	�>�O�){S���c�̐�`+׾rߞ�8B�d�pِ� ��^02�N�bV���~�3ם?�/�
d�7�TZ��҅Ԣ C!�qB��S悊3^�C7ʌa�i  E�:l<�p����w�� Q�S�~�g��7��ԫ#OR�z����fmC�yr�0�w�A�/���#�OS�c�,�C���x����	�q�:��(���u��䗋8l�#/G<Z|� s�I
U�{҇��V�>�`5!�>r-���f��QHu&�8j���C��L����� �L� EZ���^�<Q"���^T<jp��k���|1��y���b�Քh�$�;�d�<����0b
�7�hz�;��ޟ��xѺ��=�)�' ��x"�)*T�i��f V�*�'LA�fhT%v�4�p.LUGڥ��'(���C	NU;�I�	ڒ4��'oe+�a���t ��
'��x	�'кŉÏ=i;�Y�v���8�	�'�ș�B��[����a'�'�@0	�'m2ٱUL�zdn���OΧx��X��')��hS�R�\o�9��R�]l�#�':"�A�@�]��D��Mũ֊��'G�$!�#�zM�B$V��t�c�'�&$3�Fͨ@! ��ca�4Z�b�'��Sm%�Va�Bd�JJf���'�8��K>m�z�Ą�%FB�
�'���[�cC4"�܉��NS5=+��'f��Y���=Z��VJ�f���1�'�4})4�ڔ[wl<H�L� a=L�X�'Q�"�̺t�h8��@��k�8���'�&�P��շ�FtSE��{��	��'�����-�d����!��7"Ob9hA`�Jf�����9t̢���"O@�˱$R�x0��	�(U�Ȅ��"O�IP�]�?� (�E�Ve�΅K&"OƑ�!��.�N��!/A[����e"O�T�4@ʕF��q�����	�w"O| c����|k�����ˆ�HtH�"O*!
�G2OH:�BG�Än�As "O0x�5H���AӒH�=�"O� ���@�H9�F�z��S�IV���"O��	�n�&݊`��U%}玈aQ"O�ѩA`ˏ)wZ���
�"ڵ��"O��b�F�UC�D�W��>|8*u"O���uN�)a��3� ���pҠ"O$0�"��@6" �eH�^�\E#v"O�q`�� �MR�-�="�4�B"O�!�u�pd�5���uIĐ�"OR�[��1X�dY����2TaW"O`�:�E�:���P4KķK�Q��"O��w��BM�%3`�
�a_���2"Od�pƋ�� �J��&��"OJE s��fY���
�
R�|�z4"O��{�!��@�0	�+ӗ7�&e�c"O.�cR��n���:��ؐz�� �B"O��r�M8-n� ��I�-Z��`�"Op{ƅ�(e���T��b|@=�v"O�3#g\�pج�Ӂ��f����"O8@�œ�l��Q
qG> �#"O��62A.-�2�O�c=ƽ�B"O�SkYn�0�+S�60"(�@"Ox`+��QB��y�èٹQ#R��"O8�����ç��,H�"Ol��@'=N��2�HY�DŶ��e"O`xJ�0����þf]̵ۣ"O@)94L���V�1�M%|F<�;v"O�����T�S�J��Lx4T���"O��h��%-��%���*QH�"O(u�R���,��@)/@;P���"O��+�,T�����Bm��V�C"O�h�T
ȎB:� ��+}v���"O��5���Q��蓋۵Jƌ12"O`� b�_w;�0q���~��c"O���Â�X�irԪ��fX�ˣ"Ox�26C�'v�H�� ��I4�Ca"O�t�T ]L����8X��!��"O،�0�AA�Ԥ�"Κ�U�&���"O� ��A��k͔�Z㌅�{txU�3"O m Q�t�dZ��B�1i�P�D"O�{g��]��ː!���,+�"OJyVfZN!X��*o�$�(`"O��mP��[�&Z����p�"OR頥��;O>zq���L<��3�"O����P�xa�!��F���A&"OLYWoէ7�n�2���1[���"ON�fn >n�Ҥ���}6<��"O��uj4��P7x/>�h�"O2Q#G(	�w�$�퉩-Z�ہ*O�<�D��9t�v	��M���a�'f�i��Rs_D��EJ�KyA	�'�x	Y�m^�k���%$	R`��'2xh��늂y�x諱��B8� �'T���lh`��!GQ(U]N}Y�'bzC'W�pD�]h�O�05�y�ʓ?��X��A�`:�䓷�S0��х�L���`e!O!Jb�d΁
���<ɔ.@���8��o	Q�iR�}≒�-r�P7^X���F���� h��'�u[��ki�a!��O�?�95��M�#���x�N�p� SҺ��A�b/���'���iA�_���y*�VY�0AeF�g��
���͓Tb�qV_?�Ik�I޺�#j��}oR�Rd��*Ђ�Ee�Ay��i��Q�V�*Z�|�'�z�Q�ϭ~���2N`��j���M�A��=4�6��<Q���)l�� �*��b���q�'fM���P�
>m!&�Z��t�'*P�@̟�i�7�O�Ȅ���Ԁ>;�U�"!Z�c%޹�t��I*qO^m��� �I�Ӕ��4:aC�7RDՃH>1qcַSF��A�π ^�z��ȕN��r��]2TH8�Z��x�"�;d��t�J?�g}���7�tP�!��4CP�P�Β�~��lriG�h�I#$�<E�dϔ�H؆Y�q��#`��Q��O�<d�N}��M؅v�I�}���iM[��!�B��-� :jG4��й��Qy�\(�h�}
t����H�?��ź��'r
AòȒ M.� �'1�IE�lz��U�`�D��o6r��Wd��6* }X2dL?��d�'_ج��A�1�B�|�Ӻ��J�U�@Aӱd\peG}*�%����'a��ӬD����6��YKX��B��2�M������<E��哑ޔ��aFM>[y�=[��'<_<��m)?q�$	�Ny��>%>I 7�S�m��TfLAd�΄�����,����0CJ�t$�G��D�	U@sď]>u��ai�8��$ڣ~��k'� ���)�'wI�A��g\&��`#�,��6�q��\�M�$ߞl���|�#�S��!���)iyN���A��F8�9n�bX���'\1�A�O������*>���7IE�yC����mA�<|���*�V��'$)���]�'FK��w��=l�RT��l6\8TEi��l�,ѹ��
*t�+�*���g��?��g�0?���kv�2��$�B�ɼh &}�C
A�`=��Kd�M�W�VB�ɰL���igJ	��LhaO�k�0B�I�zҶe�ť	攴�"��Cz$B�	�E�p�0����7�2� |�C�ɳs'>� �a%}�Xb��՝'K�C�#�]Bu"��?)")�tK�<�B�	�p���{�*�/e��J�A�6o��B�Iqw�x���TM4����7�C��=����e&�T ��BA�C�I1Dx��8�dDlc��ޒV��B��a*�A�·�4���NVA�B�4F������/g���;A��!T�xB�	� $L�!������)JsLB��0����$�pHZ�Rwd2f�XC��f;�	C��D&>�P]B�ڇt�B�I2&�(@r 
:2�i�ΐV:�C䉘��h��گHԜXj �	�lC�ɲ ԭ0k A䚈Q�#��3��C�I�A���@#*�7H��Y��B��B�I l��E���k��#�͞:��C��%=��\��.ڭV����%,ٗ�C�	. |�e�&��c�P0P�Z�o��B�	5NH��àB�(`���ydC�0F^�i���<My:�ôDW)�BC��o�,7K�+q� �X�? �B�I�;�,�P��\�'u��	�-�,8�B�	4e�xPt�	�:V�0�֎�rw�C��.c��A�fb�8��, �S�/�C䉀Vx)#�khu��ɱ�LX<C�	lhz��i�(4H�Z�̮�XC�%�Y�E�4=Z��#7 ��
�xB�	q͒4��n׷4]���,K�sabB�ɑcf�����j�B�c��I#��C�8�� ��*[f3�������uXC�Ɏzt�HЅ��9}ҍ�C�:��C䉥�n��&)l���ÕHY�/)�C䉕V2 ��,@�(ƪm�ԅ�!o|C�S�޸�f?c�l�契�Y�bC�ɶ<fH�pb���)G��&�G�hC�	(7g���JW$,=(��,�E�zC��	{U���§�����D��tC�I!t��%b���K�M�%(�jC�I�\i�Q�ȜD��z6��!;fC�I�:t�S5%�,o���#��R&Y�C�	�ϴd4͒�~���A��/'�C�$i�J�����Q��`����w�C�	/M��b4g
q�ɦ�O�|��C��:Y���`�)�{�a��H�K�B�)� ��xw
ҺJ��E��2�ĕ��"Ov4K��P�P@2G˗�k��p��"Oxm�B���(��	뜭m)�0I "O%��j��D��ЫT��rpL�1"O��y���(*��$�FJ�9s�ꨱ�"O�xR�ؾZ���K�"o�TibA"O�]Q­�� ��X�� v��Jb"O`<;E�@�&��%m�����"O�����E�L=�N%2���
�"O����i�+`��91�@�B�($`d"O���o�$�S�OSڴ�q�"O��	�I�
` 4�9E�:m��, �"Opܠ֯ӑi�n�$*�F���"O��0�h&.��\���*E�r�"O|0B�Ϙ~L�b=10��c�"Ob��c��!KI �G��Fn<	G"O�Q�)ߩ�2yr�	 V,[�"O�Ja�X׎ ;$KE�U�q��"Oxcg�$2�t���E�7�|\��"O��b��
�k�6ș��� [�v��"Ov�y��iHq�VLP�8��"O�I�D!�:*�9Q+'\��,[#"O�Л�@��[�*��*�!?�|��"O����N�/6�P��Cc��;l;�"OVb���.=�=r��_n�t�g"OȐ�wHG� �Ѐ�`��*�����"O��8�e�@�� .Ղ-�F�Xw"O�qb�����\�(��?�����"Ot�KCN�	|���`S�_B�т"O���0���)p2L����	6n-��"O<HW*.f9��N�'*��
d"O��(��+͊-�񭝳��I s"O0��q�R�b�F��B�bF��g"O>=D�~�N��� �U?�)B�"O�5� H�O=�dc�.R�:����"O��9׀�#j�[K��ָW)�5��"O�|XE�Z���
�� %KGDth�"O�2���F�Ȩ�ĭءY;���4"OH�a�t<>��eF�$t',M8e"O~!Ǝ�	
ʴ �A �%	�!�"O�᫂@Ӆ�p�o\�ic��Z�"O�m�@Ȋ98��	�%.��1B���"Ot��wo9�
��`�\,�PjF"O~��7�M(M�����·��a��"O�c��Τ|��mŚ.��X��"O����I�6��5!�\�g"O���A�)a؁���ϸ��"OV	�U"�=� H�͊?Ek0�*�"Op�൤��x��E,|�\��y���!V�HP��0k0� B��y�}�����$��yxBH�a���y������Go��3��[��y�!��H��KL?_���u#��y���a4	����,��"u�K6�y� �m���`V�%l6��Tf"�y"�P�_����`��V�	���5�y�kp�H�#�ʀ���a�mڽ�yRh(^��I1��E� ��ce-!�yrG�<��Y��M�r����8�y���&�,а��C�و�B��	�y�^�7[�ĲEg��>�"��`䙂�y��o�Ȕ��ė�4�a����y�bʮ&����;)���qg
�0�yR�E�E�P]�N�; �6h��y
� �슔��7j�H �e���I^���"OB�(G���e�#㘧?��@@"O��V!���R�#�������"O6�2���y>�����jn�}��"Oҵiq�E+L�\Z��Ie�qc3"O6��G
9(��C� �1yfջ%"O� �A���?�8��ů�>�
�X�"O�$��"���3�^"x���"O
a�ƃ 3F���)I�e�ly+f"O�lr�Q�0���g����\x�"O�X!�둻M�e�$��	�8u�3"O	�`���e
fd3��7/��9�"O��2ь�]�J ��k�d�r"O�ەGó3��E�"N)|#fH��"O��ء��r���-�8n�t���"O���I��}��1�+ֵ\��ň�"O��8�-K+/'��c���5(p���'"Ojy%mI�r�ҵ��&]03��UBG"O���5��F�Թ�a$�'x���)�"OB9��^�l4\Q !�$:�4q�"O��x$�T�T����J1��YR"O>]�W��!��:���e�Z�F"O ����"<r�E9FJۀ=��eA�"O���h��t�E'�3^B�+$"O� �g_�-�Yx���4D@�Y2�"O4�VNԆ���R%�W�Li�"O�a"�`�hѸUc��!� 1q"O�P��.�9gtbE�BG�
=�q"Op=�1dѹqR041V��/Fq�H"OBXJWD"V<@���R�̡��"O�!�CҸr��P���	��u��"O4�%�R� ������3���v"O�q�bO��_$��У
/�B��"O�h��
*vʮA�@DK�x�ԉ`"O@��G*`�GU
1|͊r"O6ٻ��3&�Hآ'�]nk�"OVI�Dc;q�b}�����4)�Q�v"O�����5Y�����^�<���"OR���ǉ$'Rmy����S<L!�"OH�s�l'���bKޱ�!"Oh� �!�<*�� Ɗۺc���`"O�e�ƞ$e���K)�B��"O�E����9 tEI�gH6q���"O�X��i�*����'��V$^L�Q*O(ڀ�-�x̛r��N�1��'D6(YC��2H����}
R ��'i�@��mR�Jn~��tg�����'��Ly�!�3��x)$%�G��8�'l��uDǝr��)���*EN�-��'�P<��آ-��Ɂm��;�E��'���ȷ���~Y��j�I� $=r(X�'�2��ŀ6 �NO�nK>L0	�'��q#,�:=+MZ��ٲV����'�M���]&b���N�w��	�'j0�W�eZ�Y��hL{���Q�'���W�:�D��L%��4�'���@��\�z&�h�H�`hd �'T�*U��HD@��\�r	�'v�4h���6����H��a7�`@�'葪���#\�D��C���X����'��a�3�C"6]8@n��y..��
�'�D��%	�*�D��&�z��H2
�'d�90C��	P�x�Hց)�6��'��h�AD;L�<��)W�&d�i@��� �"�m�_wyA��b!x�"O�h�Z%Z�s5�H�%߶q�"O��ƅŸI�����=� ���"O�AG%�Y�BijÍu� ���"O�� �_�pB��A�̿q��� �"O����P�}�p����=!��ȋ#"O�����jvP�ƀ\Z�Y�*O�i�NC�G}�}���D�(���';���d\�J�B�𓣜�G�x͢�'h���:iduړ�9Q|\j
�']��ҡ�F���C� �|�I
�'Ȇ4yc �@��!@��L�1��+
�'��xe�Z�M��� #g��*|���'�%"7�E;l�b�k�Z�Y����'��R%W�M��������=H�'��{�耗`#�S�g<��Z�'}.-!�!7�8�w��..8&�H�' bA(��ٵVB��Ǝ����X�'�|�㴀��7Ĥ�T�$[z�A��\}�]x���I�FR����8@��K_1�H�k��+�:�C��p   ��   $    �  �   z,  67  �B  ~K  gW  �`  g  mm  �s  �y  8�  |�  ��  �  D�  ��  ɥ  �  N�  ��  Ѿ  �  ��  ��  �  ^�  m�  ��  �  Y�  � �  N �  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b��=Q�����] ��k�O	d}�E��y@�ZY��qE�#�N�@%G��yR��5 ��ɢ�NkĮ��<�p?y�O��ҡ�X���Š,&f~�JG"O�q�.� rL��סέElb�;���x�O��ӅV>u��`�0gx�	�'A��Б���<�J�¡$�� s�D��'_(���)�'�PU��l�EtfP��I�`�Z���4T����.�^�	���;��'>a~m\+A�
�Œ_G��a�� �p>�K� ��-H/�l�Gc��(����D�v�<i)^�M��H��(�&Kq���B,�N��'�x�V)�2%��@�+���-�G�$D�4xP- {��8S��#��|ɷ���c�|ק���+��: h+�:HZrE(IN�B�	6#0���ᢕs>����U"�JC�I>{�t�z �Z�M�<��"c�B�2iG{��a	ٟ��I1@���w;/YL�r�ƻW8�C䉿)a����)T/ HT�{1���H��$=���E��s����ÌGp0��%8D�<�ǀ��ܑp�i΋��A�ht�(D{��i?]��y��ä6_�Z�L؞�!�$݁�l��qB��.�!PW"�+s���>!�H�a?*|(�bC�W�5H�g�<�E��64�p(�+6���+QBIY�<I�G^��D�4��m�7a��<q���'��?Vh&~h��a�'qN1c�$�O~�Op�J�F��S �� 2�ȕq�"O6�:g$M�@*8wCB<&��e�v"O� �-PuǓ:B��TBIvҕ�Q"O�8�F�: vz����^-1�"O�k�ͅ� cFM���"O���b�ƞD�q�Wf��$���p�	E�O�d}qdUI��Ӓ�R-DE�
�'�`x+�O�+�va���N���'�T1bH>	���O��1ѹ3���a��1f�t�j���D�O?�l��X:Enu���ŲG�\aP���~B�[�P#$I�E�pL���O�-���S�����db�82搗0����!-�;2pP�"O��4��s��˕��G
�E
�	y�O���clG����᛼�����'	�!�ď�KNq0# G�	y�,��'���#�
+XQ�2�
�xۈ��'�'E�FA��EGΤ�z�ȁ�Q�'����	�o��|t�@!8�`�@G�)VvB�	���YGNΟ,1.5�5n=,$R�g D�h���H�p�Qd(��U$D��k*<O
"<���9B�=�F��Y6~��F��l��&�0; �+�@,���B	=�������<�'J�%�"~��E�ikd��E�?M�T�� KC�'�?� b��r_V�s���0=���T�"�v�n��dϹy�%9���B�QdnR<P�!�$�	m�Ne(Rg��{a~�z#�J!�!򄉏W]� H��5l4ع���<��|xr��p"�U��N:L<S��C�C�I�md\#2�ώ+i��A�T3iO&"<q�)"��ʧ(L�}v�ϑ#ĐqR��AU�<�0�^&bQ"�Q�%�1�����A�ў"~�I�j�( Ze.�V�����E�d�B�I�;3Rg�F�`<Cp��7Z�*��p?Aq��,#��J�!Wq��ak�)S^�<�&*V8tx�e[ ���m����]�<�g�S=b�
��, ��ܸ��D�'�ў�T�r�x���o�|�ʵ ��w�ɇȓK4��ӤX'\m��{$� <]����z���.b"Qj�#ҏ	Zvԗ'8a~���"��Q�NR
C���Q�y���C;�`��eG>\׼�a)�"�yk�0e�nd�0�Z�N%P$GL?�y�GT�#Ȭ��`�d��HT��ON�Fzʟ��*D&Н��4J���kVы�"O�� r" T(�[ׄ� (&"O8�8�oG�7Tbp$ކ&JD���'%��>Ʌ�>)�bh��B�����c�Ux���'���)�(~�4TYo�&ֱ��OB�3�'�ɧH����VC�G/PUAbv�9���	�k��?�ɥ�;'���@��c~(��mx�	8X�$]ɦc>c�,�cI�c�
� ��R�c�"�O�MDz��I�p!b�+��U�J��N�	$2�e� `�>�	�>8���Ĉ*:�Y3�	5��l��	U̓_U�f�ÖH`�	�QDŻv5fX���Sy��:XtE�r��_�X|1�%���y"+ĘuK���@;g�T��bJ��ybC�Xٌ�qM�^����E��y��>n[̹`��ϋN�k@/�!�y�I����-
���9J�b�[ nO5��D$�O8��/�q�ޤIą�C ��B���y�����c8gԭjvnG�-�`	J2�A�y2ǏGJ�"�+ę�dI�A���y�,"[��ʶ#6J��]?��=aF�g�D��dm�cB�؛U0��×�^n��)�6�p0v$K)�ma��^���M;�'�x$���I�\*1�f$���"AS-O4��� ����%��U�|�X©� �X �'��dŭ)	�H���V����!h-�!��ߙ??Ρ���R��h��f�-o�ў�ᓑ�0|(&�Z�В��Ƨ˩>|C�I9+��\tNC+k�P������:B��8L/n���+�qdb���I!N�BC�	�qO�L)�L�7:B�8R	����8�����IDЋ��T7WZ�����viB��U��I�"ҝ������rИB�I���8c#ؗY�X ��iH�">ь��	�p2p�@��F�Ѹ��""-�}⟟ ��l�/Y�����V����}�ܢ=E��47�ZM13&�������3P��ȓ�2i��с%�(��$,�4v"Z��'�B�'+(qe��(Zv|��kY�/{l�j	�'z���$aԳ=�v!)���@e��'�L��T�ۅ<��[�fS�r�:�H�'p�,���T�=I �����pn|��ߓ�'Ntx)���Z��H0�"c�� �'�H��W��Z�'�@�Y�H�'����dB�2e^R���*֢!R����'�f]����o �ݪ� ǝ�H�N<����?��@�Em̐P��$Y�/* �ȓa����1́�\N�pJ �V�u^D�Fz�O��}b3S�D��Q�BC�(t�� ��.^^h<�M�w>�ܰ%@ K�L �&���O����	�l��X�K��d"N�1%��B�B�ɢb`�6�;G��]���v�P��YJ�Ti֊Z�[����k�le��J�@xg�Y4]�@�QKտ,�ͅ�d��Ł�$�*	��!ED�����j��V<MzT��Mud!F^�5�!�<���"!F�-W�}j�-t�!�$�~VPYt�\�Qr�JճB�!�䓔vzN-ڴ��kE��r`hG�I�!�I-��p�dɑn�M��	C�p!���c��0�m�P!܄(u��,a!��
��ҹ��n�]k6x���N;^=!�d�c��a9悃�vXz����ɤN!�$ߡ~�b���ӇH#����d�3�!�Y6B\�|�f��k���gY5u!�_������8 ����v�X�"[!��ڵ;AZ�����k���	!�")/!� �g��e��PW1Eȗ`��8 !��mZx\)��
)N$�}��L�in!�DT�ĤI�S��"�Ed�Ƚ\!�ĞO!��K�(�b�y���+JW!��)V�j���~>A�'j�:-E!������v��C��p��IǦ6(!�DF�6���%��d��q�R◩z!�[�F"8�;Q��E�*%S��P;!��"�������%�X����k���ą<x%�cB�B������y�&3E�,(b�W3ЦY�揇�yZw��PK�='~vѴF	��yBJY��h�!�#E���B*�y��!g>�M�3#��x�YW.W��y�N`��(r�KܢE�&�[3�yknt�U+eZU�U&���y/
�͂ؠr}f�jE�M��y��T�=�~�j�F�h�6���.���y�oA�Z]��Acb۸n�rD��J�8�yb(ה�*@h��מe�D�R 䅲�y�dܘY����Ċ�T�֡'�֞�y
� �x�ȋ�A^���(ݽF �PK�"O�Qk2̛g�x�9�H�����S�"Ob��`�,e�Td @�ƅ8�,u�"O��{��	.��e�K�(�	"O��1((HX����Γb������'�2�'4"�'�R�'��'�2�'Ю���H�>~��-�!��}p��'���'���'s"�'2��'�b�'�v9�ĕ���ݪG,X5M�^��'F��'���'�"�'���'��'cXH����NK��`C�"7�(�k��'�R�'��'���'.��'���'��-���q��w��=|�IV�'Zr�'��'�"�'br�'�2�'Q��"�K>X{F�1�L�j�$���'�"�'��'��'N��'�r�'�K�i]jPz�&
�=��f��?)��?i��?I��?���?����?�׋���1	s��7Ŕ�Q���
�?Y���?!��?a��?q���?����?�2�#;u�8J�M��eHP�i�&ۄ�?I��?���?���?����?9���?9t��i����[�9����?���?����?���?����?���?�q烫
��%P����\d�c)D=�?Q���?����?����?����?1��?!��Sc�
�s ȶ'�$�����?����?���?a��?����?����?�vI��ٶ�+��<JҨHV���?���?��?���?���cK���'E"��Xe2��=2�q�Β'A���?Q(O1��	2�M�VCP=!c������ i\7p5F��'{�7-"�i>�	�Ms�g� p����İFn���D��@{���'�4�ɧ퍔�y��'��s��]��P�O�2%��[���xAR�FQ��R�$�O���h���Z��
f�(�3ŉ�%f�Ib���@Ѧ7�}��L&��w�`�UOA�[,�$��jЋt���$v�j,lZ�<	�O1��L��0c0�S�i����H4 �rr�]���] �zlS0��/q�=ͧ�?Q��X���;����J�A	t.��<A(O(�Op�oڽ'dc�(��	����r�N�@��`7%�B�8�����M��ih�D�>�G��o��I7m�$����L�H~2l�&N�(D�!�آؘO�<lRB.��X��@D�	�l �цCy�RJ'O��|yB�����*a�rQ���:i�8���-Ξm��Qզ�R7'4?��i��O��  m�Y�3k[;0���s�s��$��m`�4�?IE�@�.�5�'P��� ;\,���B� �\�Ƈ\�*<H(��\b���3Ň�P��q�7{��U�։�3$(kt��k�S&�Yv���[��J�a!.y;��T�w�[� 5SuV��Ue��9�E`R�_L2 ���Ef�m���W*ra���G;OB"<p�v5
���7[��Q+�	�E(��cW���X�4D	��-����;`�2�*�L>^���k0�Y����\I�vxR5) i�^H���2E1��:c�Z�3fo�!'` 	��Qe����,6}���C��	�B��F�|ؠR�Zrw�:�m�+�`)p���T����@�M���?!������?��dCx�d(��A���w����U���I�阼���ȗ����'m�ٺ+��xPզI���%!Қ&Dj7��	J�49mZ�h�	ӟ����?��	���	&(�
U*aȇ=R�#2��??f�e��4t�N�������|�H~��E% !Zd�رN�:��Thڦ<���C��?���?)�i=h&���'c��'���u7��.�X<���p�>D�kS���ı<��(Jm~�OVb�'b��?�UӀ�}�8��Z6��OB@1C/�q}�Q� ��~y��5� ��b����F)�2��QH���8�MK�� 1$�̓�������$�O8�d�O�̪�nµ_�8жmF5]�,z�݈o��QoZ՟��ן<��>��I�<q��A������Ͳ
�t����h{j���`��<���?A���?	���?	��&~����it^�ܻl.01�	�~��8kT�j����O����O��D�<��������!�h�#92B9A�<uu��e�d��d�O��$�O��WW��×T?=���em�T;2*/eo���!�:�P��4�?y-O����Oj�D��Y:�d�|R��W.m���+#�	d���AƆ-Z����?I��?�pgY��F�'�B�'���l�E�hܙ"��F威�Ȳ+W7M�OZ˓�?YT�?������Eu>7LfeJ���w��x��)G�h|���'B��ܲH�27��O��D�On�	ꟈ�dF�9;<A��ƓO��U���B�mN��'��C(iR�|�O�1E���2��=b�9�S��#<*1m��K��x�ߴ�?����?��'����?���;�1�т*rU '�>s�1
ҴiRW�'���'�d���O5�O{�����[��U��7S\�j4���+�z6��O����O��C�ŎϦ����t��ß��iݙa g�1_�HS�� q��`�Ee���ī<1c��<�O�r�'Ng�,����&��"C�\�8J6��O"0�$����U�I�|�	ܟ���d�I�M��1g%�)�1Q)@�3�86mJ�Y(�#�2O8��2��?���?�#Y�p�<���@#������ �Hʐ�icR�'r��'	��'��D�O(��EҮN֌A�됞'@`K2"�)^��O
�$�O����O����Ox��"A�Mڅ������GB>,ܝ"�l���M����?����?�����$�O�M��7�|0��]h��C4��"׾SR�Z馵�	Ο@�	ݟT+��:	���Ӧy�I������_�HYSC��4���ò,1�M{��?������O~�c�3��ĸ��I$L��an��0-F!<�H1��m����O����OxdpgHEЦ1������	�?Ir G�X����"�[b�������Mc���$�Ox- �1�(�Ġ<��� Z�R1�P2Va2Ae�t9Đ�G�i+��'P0�3CgӠ��OD���)�O�M�b͂{n��iDq�Ќ���w}��'�����'/rQ��SZ��O!	�B<atͺIrU��g=Xޛv+�* A�6-�O���O��)�����Ob�D�%kAd2�5��d���L �eo�D���IП������$�'"21���U�D�
ͫG�U�0�@wz��$�O����_��Mo����I��������>1� p�� C��
�a�t7�O�ʓ2�ĸ�S�t�'B"؟1�%$-{�M8$A���YqP�i�B�A߄6M�O��D�O
��P�t�O,� E�(e�|EJ�1}dK�X��
nw���	��I���IK�4�DY@� �ǅ�M���*�=��l�Ka���d�OL���OP)�OD���KSe�f���S� �RA0&hM2[�	ӟ����}(��	�4��ٟ�yroS��Mk�L˰Q�d�p���+4���V��X��6�'b�'��'<��͟HX��z>����Wn�𜹃�%�(Y���K�M���?���?���?�@?!�v�'xb�[�+ �<y��l�b���	(-�87-�O���O<��?a����|���?��+��2(��J&��F�ȴ!4#���t����?a���?9����F+���'���'[�T��o�����(w�ځr�ł���7-�Ol��?q�lN�|���?)�.�|nZFR�d��(�$%����ny�b7m�O��)f@lZ�l����0���?1�I�96�,[e���VR2d�dk)oo�D@�O�$��S�J��O���|*M?�YW�S�z�"�8D4�xh��n�&Hٗ���!��ϟ����?��S(����x�/:: �D�m�1.�*ոe�D0�M����?!����4�������Iπ�jG��:7�-�Bj���]oZ���������RPo��P������	ş֝5��6bX�k�|p[ ��Q�n7m�ODʓojF��S�t�'���'�<��#/U{b�r�lJ�0IHj�l��б��m�ҟ���ϟ��	���	����ე9�\�%K�����o�>���<i���?!���?����I5}�(�����(MP6拑7$��''W¦��I؟T��ܟ�J��<��?qDBG�@��@�ƞ�v�xt��
7�q��?y�%X �I��?	��?�AI�~4���H̠�t�A���C�J�7-�O��D�OP�D�O�˓�?qs��|n"3ɰ�
�f�	���b�e	�듨?����?	��?�W�R0ě��'��IN�8��Ő*T񡲥���6��O"�$�OH��?!���Ľ��8�i�rt��e�$��!�m����O����O�yP�
��I֟����?!Z��N�.T#B�$^�V���%�Mk����Ox@�C7�D�$�O�y�&8���ޟ7;FdB�R7,���@"d/�M���?YE	�dK�V�'u2�'���O��?�*aӐ�3r����6 F�B~���?y6OA(�?�����4��O3d$AAW16\�(����q�4v^��b�i���'q�O����'\��'qP`S��#o`M3��^�~�T�e#dӒl���O�$�<�'�䧇?�u˶&8Y��
k�Tl���8:���'i��'��ia�.gӞ���O��d�O����So�UKvJ�k��U�V�ix剝"D�]x��g������?�S/� K>0���n�r�F(ݚJǛv�'吵�C4�Iٟ�$���]�Z�("�.knzh����,�R��<I��?q����3_��H�((N���@M]��llbq�Qd�I����Ik�	zyb G�d��䮊S�d�`CO����y��'XR�'��	�\���O,*ԑ��T6b����j��J�O��d�O��O��o�@A�'�ܼ��ݯP�
�7FJ�[�Nq�O4���O6���<�&,����O� ����_o�L`g+[+v�:�{2�jӸ��)�D�<��e]x�s2�����U48�=�C�%$*m�ܟ,��~yRD�����$������=d/6dp$��J9a��nM�	OyR!K'�O��6q������B�D�%���߯�^6m�<YBj[F���~b���"⟟���J�m�����`��bI�`��cӴ�dGx��4,� XQVyCJ6hQ��	��
�M6m)J`��'r��'$��e,�D�OH�b")Ś/��J�mٺ]�̅�q�����;�4�S�O��`MdF�dhZ�$����gމ~$6��O`���O�L�%�A�	��	s?ɥ [�x����u��*�HM�I���<���?���l��Qۧ)O�.%4��s�+[��C�i���}�(O��$�O"�Ok̃*,L�����
��Qے-F:`����3a
b����ן(��Vy㉊KP��#��8$�Ԛ��6;h��R0h5��O��d4�$�<��&O�A1��Wx�d�Qh�3�v]�<����?����䊹T	ϧ+�����×�T���D-Z�ZrB)&�X�I|��oy�
 �����di�UO��_��%���ZeZ��埬��ܟ,�'�,Iwe9񩙁Fk �V%\>|�>4�� �1�&�o��'�H�',d]�}r��R떄�`-F4RE�L����M{���?�.O�`�uǁi������RT�:D��>=v�5lƵX9<uPH<y+OL�u�~m��^Op���O�䠺�Ȧ��'3����mu�΀�O�r�OP�G�y����
��D�Vi��:�p1ltyR�;�O��R ��!>���Ǔg�6�'�iMlI`�Ed�L���O��$�$��>I�Ɛ'��5bg	�gf^3�/b�������O���O~���O���B|�? @����
�-�dq��%w�樉Ӹi���'��n[�2�c���If?�Seb�jl��Ē�0��5��P_�e���<A���?��iD���6)�_�l �Dǁ�1V�����i����cP�O��d�O��D�<��9�.EzG�K�!3��q�/��l�'S���y��'R�'��kR��t���M�'nݨ��ٛ������?����?�)OB�2"�P��%6ZP�Ź7�ןV��"���t̓�?����?�-ORAf�A�|�6	E�8@t@Z����<���"�N}��'���'X�	Ny�����	؞��I3��A�K�HD�ҧ77�	֟��柸�'�>t��6�i�8V ���Z����JX(p��l����I~y"_� 1N?�'�ҜH�Üe����EQ�v�����4�?����DN�f��%>����?H��N�T����e�3~�ij7O,�M#.Oʓt��A���4����7!b��@�O/o�����1�M�.OL��w���㯟��D䟀\�'�*�p�޳u����w���Z��ߴ��$�z��b?5�Ə�1bN
�a5� �d�9� r��l����������(���?5)H<A��q�򄐲���@��<���6+�����ig8�����S���"��4
��9�L�>Q@��`��M���?I�p}$19��x��'`r�O�<��
U��VJ!�6R�A�#��K��1O���O����+V��@��a�!%4�K�ON3INxn�ٟfI���ē�?9�����`�؞D3�HV�� d�2ga}b-A/��'���'�P�����P�%Ih�huc����ar� ʄ�xb�'C��|rX���P+�6D�r���@�l}hy�q��A4Db����˟4�Iky�N���ӱ@�*��B��X9�`�!!w����?��������ڴ��	�VT��H���u�|����&����?����?)-O>LTnBo�p�z$@�@^(�hk�N�p�d��ٴ�?	L>)O���d��;��4Q�(W����bJU�nC��'_RS��!��ާ��'�?���+�Xp B��+��)q�A@u`d��xBR���Dk/�S��lݘu� ���ٔ[��d��Ĉ�M+OlA0&�ߦ������D�|�'�~�
�"�#[�H����e��$+ܴ��1l��b?��cjش����UC�P�c��nӆ��U�C֦]�	�|���?Qӊ}rh�0#���a@>gNN�Fā4A6��#}�"|�\OJPq%��.oQ\2�ě>��y&�i���'B���0O��$�ON���|�Xs*m|���5�	�1�c���&�,�ן���ǟ�IՃc� ��d�*W7X��o=�Mk�b�Ӛx��'D"�|Zc�d,��%/&ڃ�b�a�Of���$�OL��O"ʓ'j��0���DJ���_�0�Ν����9j��'b2�'��'c�ɐ;�B� �Τ-�I���X�S�q���-��П��IڟH�'��	GKj>A��	�䘤�?�1 ��>���?�H>�-O���@P����Fؒ1)6� �&R$v~�z��>Y��?)�����Q+ I&>����	P�8���);(� S��*�M;�����$�03��O����,6���H��(��i��'��l���`N|2������e46\���8hpj�+�i#'��'��|"�_
����-�=�^���-3�M�,O"�;ʞܦ����j���|�'�t������*���2��;��s�4�Px�/�Qxl1�o��������M�%].o!���'e2�'��dA$�$�O��B�@'W9�!8�*ٱJ����-�u؟��I�N���X�i�,8懟�qBD���4�?a���?� aZQ^�'���'��$�e��U��8MJh�jb��+Fa{��'��'$ʌ���G�XC�E�Q�+B�Uh#b�^��  2%����៴$��Xi��P'��I�`P�$F�aT"?i���?�����D�'��c�⁩cAx�`ңM�V�9 ��~��ڟ$���8�'j��'E���%��V��G(#����N@�ژ'���'�2P���$׀��ԆP���B����D���������O6�d�O�˓�?��NJ��O�,�w�>_�-�sJ�3R':P��O���O ���<��Z�qy�O����$)ΦV���&�?W�v��A,v�����O�˓�?��>Đ�����SnA�� �*s՛뙘G��V�'>rS�lxb∓��'�?��'[����$sr����u�*颣�x�_��)���� �HЩr���Yb*�'��MK+O�՛�c�᦭j�������f�'�}QWk��X`�xijT`�8�4�?���_T4������S�';���b8w� �aϨCk�n��Nع�4�?����?��'G4�'��m't�Ib/����q�N��j&�6m�<�d0���ȟp �L�Jh| ��F�r���@%���Mk��?1� n�̀��xB�'a�O���`�ԤM�ŀs�Ơ)����v�i�'�������O����O6Xӕ�ܽ>$hy���+c���0�a릍�	 l�@|yM<!���?yJ>�1C�����s��/�ʀp��h}��LMbV�t����`��Yy�@/� @,X"g�G���+�'%��K�I�Yq�'<��'��'=��'^}��E�<'��᠍V�M�0Pqd�8K\RR��I���	Iy2͛�@.(��)��!@���Y�h��.�*���?A��䓕?I��M�(��Y��K�<׺ݡĩ�]a���DW�������gyBD\<|>���*���+x|��x�b&!j�	�d�æ���v�ğ���0���r��H	T���$�Ӫ+�p��g��&�F�'�bU����L��ħ�?��'\�niʰbيI�X5�Eə��J]��x��'�5g"�|��H c5��T��uK��U-%B��#ӱi��ɔ_#t}
ڴ'���<�����S�*ӂ���0;��P#��T��F�'"�(���|���(�� ;�!YB�ֆ��@���:�M�A�ִ]H�V�' ��'d�4d)�d�O
6��3-��i�6�B-�h�PGƅ�M+�#�?�M>E��'ִx��c��;�Zb��>lرf(x�&���O��D� }��'���������I0�5$)$N�&���h
�nZf�I�b��M|���?��OײY���s3>M��e�$&}:ukݴ�?����ܱOj�D'���d��A�+_6�����3t���Z�T���p�p�'��'��Q����ڥU��{���Y	�%� �G#촽A�}��'~�'���'V2F�A���b%hS 1������10 1O�pbU�H.S�(���I	6���;��~~,	`�/�[)!�d
�X����N)	���LkqOb�CdCL�6TP����Zq`<�@�=N"����#jQ�2�� Ҷ &g�:���bd� g�h���	'kf�����32��걁��F�ӥ`��(HC�b���E31��Ee�E9 G��8�n5XBl]�èy��_�	�l�����8�"rjT�v�h��Υ��\��'VUY���X����O��r4��'�߱S&���K+5i��V�j��3�O�哆P��ɠ1g�
r��Xr(&G,�'�����]�{P�x�,�+.S��;&�������<}��!�)0�P����������ɯ=��D�OT�}��tw"��Ď׽4�b�����/2"2��EZzx����#D>�Ё
�+�=���4�F�FzReǮTU1�L$dP2傸FOt6-�O&���O��9�-P�e&��O����O�n���}qゎ�v(�r��5q��9�r�'}8�A�^8-��6J1�3�d�n\*1Єo�m���k���I�1��c_]��X��.��y�t�&�Q1^2���O��(�"g�伋��.aP`a��X&6���C�W�,�6�'�&�:}��O���'d��'���r�܉b�BA�h�5�G���\�y�X����&�����Ť'w�D�O0}Fz2'o���D�<b��!t�9���>f꼊�B�t�� A���?����?��&��n�OX��}>D���p�����5�F��f�^�Z��xDI��_X��²��7o�2�DR��n���&��K�fH	ģ�2Nڔ0�l-}��Ŏw[���G%`�eЫA>[�*}%�$��@=aY�e鉘%8d	�ey�a�'���I_�U��UA�>*�u��LM;a�����	m�ɟ3�jmk�Aue(ܹC�ڮK� b� B�4�?9+O�1z3�R���	ӟ�[PN�. x�c��qd�����@�|�	�����	��DϧR����H��Cdl��|��T�@��'CD/F�N=��S�eZ1����q� ��mɒ��1"�!t��ib�І*��$�u��:,D�G{r/���?	"�i� 7-�O��X��R�pΨ�%��5t�y�rϹ<������|�	��aQ��LSZn��zO�-n5��mRc
���%c\fБ:4��O2�Ng��	U���4�'��5���ɢuZ@ �gZ6+K^�J7�K=�
m�	ܟ$3@b[7C���P��?E�x�S��V>�v�Z��Z&@ҿS��ڠ�3}���9KTzر�G����P�1�ӔoA<ْ����-���X�NV�," �'\������?	��	�O�8�2iI*|'��+ �J�(����@"O���Ad@2hP0cǔ8i�eh��'��#=�Ч�)�pIf%� ���b��|�F�'���'M.Y��c��(��' ���y���&��R&��2�,�v�@+[j�*N�N0�n� 2�`���%%�3�t�"5�`�%g�+ � D�0Q��\
 H�s��Ӿܘ��G�D����O������ݼ���
Z���i]	g�H�!�I0DǛV�kӂ��C�*����Y�0�ɋeQ��;Q
�3e�N��L�Ɠ@E@�p �u�Z躲���ڼx��?��鉱B}tY��[y�L�=^�:d���A�P=~l���$-�v�hJ�����'K��'�8������|��dؖR�)�1�۷/� 8�%�^�~��(l\��$��1�'�\5��#άv�R��ꜾR_*��P��fp�D.AJ���D�n�Zik��4G�HG�R���1���'���'��Z�D��g��|�:��w���8�4�0�X̄��d�i��S�D^�h���ql6��<)B/݋�?!,O���H��#���?�����+�2� �'X�?B,-9ץ؜�?9�l�b����?��O��(Y���$lX4��^$�HtC�p�� �@gO! ]p0C�k�p�"?it�:J�ف!P2iz�4:C��Bബx�căXaQ��p}vh('I˂/R���c�O�.P����ΟĔ�� @���(K;{~ ,RTl�r�fTq�2O����O:�"|�գ��G�dd���,*pɁ��RJ�'Nў�S�M#��	
 HesFԶ`rT�sP�[��?���9Ov�
�Oæ ��E� �T,>|��7"Ofax W�])l �T�˵f����"O�4y�H�6��4�Ū�;0���"OnDU�E���,�b�_��Z)"O&���.U�68�"F�Zx���!�"OX�z&�6T�$��%�a~�`��"O$1��Y\�@�k4D<_8�"O��i�v]�8:�ة��-�b"O�e˦͓u9��q��	�I$�(&"O2� A��<Fb�y�� V����1"OJ��%#E7dk���Q�F-%��b3"O���_f�Xp��̘�z�T�"O�)s� W5K������{~Dՠt"Ox�B"�G�q>P%𧄈�lhd�j�"O� Aڞ��FI�"��R\0X�"O����߸,�l��a��]3�*�"O�H�6m�%uVH��I::���s�"O4�8`
��QcN��r��M����"O�˂m�N�õ@N�b�b�I�"O�q�H�8<#v��C�9M9��:�"OL� ge:^~��BL���X�j�"O\�y��3~#���e�P�V��"Of3��V pn"�H�+
�yd�@��"Oȡ��կ[+|h����QTt"�"O�Y	�B�8d���DZ	so��"O�cB&��RXX���%~c�M��"O�1��,�XJd�٨�0�ra"O|y�Ve6�,�#H�$MR9�!"O<-7FT�k2�IM)M54�ˠ"O:�Ӕ]�f`�q� %�X>�]��"O���+Ωh#X(��ةm>H�#"O�Qi��Ɩtj�`���^�bi(��TA	�6�lmK�n+��*��B��?i��ʿ�6OC�a���P�[T�(��I�yr�')�A��.��5_>�`���D�?�aȳ,���m�vV�C.�Q%�l�rF����ӯ#��>1�Q�
'C� 3�IO�^�x�Ao\U�q�5�c�%Ey��px�Egq�Y#���5��8&.���P���T����R��(���O/>�3�,�b�"L���-{�|y��}rÎ�n����H�ֈ �4i
���uz,J �G�R�Ѷ�zu�@PQ�ׂD�|U�5(U8-+ɧ��+Et걃��wZ$�钪w��j��%<�����U2z.�x�%�6�Y��!,�)"�a�O挠��R>C�R��Ì��|���>��93�\�&i��Qt6T�c�@j��q"�K����Ƶ�G�M�*�#�0�	?P*���X�Ow���I"�����)}E���w�J!q�8��,B�Hў0�dBO�c.���>
��`4�>Z�HY)����m�����O/Ӫ�OȢ}"�O�Q
B��K��X����t`��$�
���`p�?�x<�֋`]��MU�
e·�>d��U�7m�"��f|�(�[�xq�H%�$��bw�h���Qk���'{��� M�-<�Xm͓\��s��X*NP������6Hu�P���s�|H5��h=�UqPԖ*p�SQ��O
���I5G�@l��UU�|J1��a<͂���gH~���گFSj9���l\˓+?L����S��A�W�\��OK�>xa"ざ?2�5y�ƕ��=�C�i�1�o��*b��;wɓ�P�l��� }vI�&��Z�$�M� �ވ�O�"�	1A�rds�ؿU��m���P �ؒ+��{G���SeӀ8��E��ZɣD-��(��<� ��~X��䢅
T�H�A�O09�������z�5�5ev.tb��^�~�4=��1�(�w��]u��٠�	��5e3Oq��F�#�q����&~����mߪ�M#s̑�8ؠ��9Z��Y�j�'�4��!N�O �!�_�p؊�bQ�^��h�'}�|���FD�,O�O��.�G|�q1�X�@���e 8``2ن�I�~b@�p�S��ň-���Y�_5�TУ	�u�X��.O��QM|b�'~����9y��H����WiL!,j*">!��Fgo�X�N?Tw*�+(�����]�����F�!\΅#��i�r��#��T����0�ۙ0��#nZ�2��@[�!z��GJ�&[���	�1,p�/]1$Tl���I�2�7�SE��s��/^��X��OCLY�Un��=n�9����1K��h��!ۖ
���>� �)k]&:*q�I�f�-RGM��b0�d���'���h"��5Ta�D�����i	�AE�|�����Χo��H�5#�v������k��	�JեPQؙ�ےq��� S�۽p,T\�� ����+rU���)�:�z��HщTpA��#II����ECp(8��hr%�%�O0C�@�=N�R�2@ʯ<(�W�� A��=)H$�G>T}2������LJ%�$/;Fd� �O�1��D"r��dLV.Rz��� ����8��"�˜5!� 0$�L2�@�ORS��I3B�A6����8���	;p~��&߷O��u��JE�ر�ڞq����䒏WPf��ʓHpA)��˛(1.�zm ڰ=y-v����
3+���j�cN�����#1�O�l�SO@�xX{!C��I���#b�]5-0�T�d�X��3Ǧ�6Xê�I6A�+Y����4%_�W\��`$I�#Zj<�9�D�>c�j=�ɯ��x�mK(qOv9�m
�h)���G�K��|��d�NX����
�?$�X��G�v�?Y�ޤb�16/� vK��sB̆r}��ѐ9��Y&��3"��,CgB��HO2��'�^�_�,I���)?�R�Xf+��?�!��˒h�*��#n�5e�(��a�-+#�-���+zb�\��䞂{�&ذ6:�� ��	e�H$��
�T)y1��M����>��(�%pnhЈPF[�4�&z�)бV/�q����N�Ѣ����tL:��C�#-���Lt*u��'A�2�J�Q�	�6�Aç���?��/<Aj2�H� A�I.6�CǯC'o7<�Y��[&�@82Sd�B�֔�w�C�Uȼ�c��s�6Q*�e]��~b�� ���0?)��Y`�!�F8R���cUj�Xy2�LXaHX���E�Q�
�Ãl8�(O�����/�^p�2��w�q�P%�;i�����=wn�Iu���C�0��	��ŉg�0E���8�7���X�z��$@�Aӄh��3�~��U��b��82���)���c�'U�W,����g}b�Uj�*.!�����T�'T�0���>F���(�D�t���։2Ϩ�nR-��	N%M�h�b�'��̗'�O��� ���4B0������p�&`ٿ:-$�b&�%Z j��$�|���J�&���R����J:��OJ�-�cV$�m�(���[Cm�'�8�3��.�S�e&Fk����d_�+��h(�\@m"d��G�Q���6���~���T��B����i��u��l��o�teP�*�/<xf�F}��ky�aH�w�hxq,I�t��-C��܃Y)h��4M��$Gx��iH�u�d^�d@W�]-G:���gԿ�O���s*ٜ�~R�M7m�:���S�I3TDR�?�v�Ӫ.��z�%	�&(����b?i�o�˟�|�;j�R�B�
_<����q�K�B��� �D+�������eӑ>睄������^m�!.�
�pIZ�������'ȋM���?ڌ���DpxQj�3�ɚ�F�	x���7u!6l2�HR�
v焮3�6x`# R���`��{�t�K��	;Aʅ���OB|	�#^�'��A3㜘L\A
�*ķP��4	uJ{y!�����OΈ��-a��i���D�b֚��TYx,� ��Ւg��dƺT���P������E��[�I���m �c^����Z��͑5�`�\s���)���E��8�΅b�>T">���	]����'�L`�v�A!꓍L���1'B �og��,O��P���2=��J�+��?-���T_��R�"�8������C�7t �`�<ʓp�H�2��A�eS4�_�T��3���H�v1��I�s~�S�O�� �#�'����ܭ>�Xt0x�r�s��P�'1��������y7�+Ce&�h��/��եЏU#��3�OTx�������'>�'k�=ra ۿ,/��3!�r�$qA1g�� `�L��?�^�cJ�)ld$H��j~����#�;G{�`�)\S$^�+�*�6S��p�#�V�Be�?�ǂK�,&H��SE�-&(�dW�yf��KdM���y	T

�nMd�ʙT��5��&�� %��C���$�,�HhU��5�)HH�P���j��>��4q1�Q"�*��^���������d�G*Zd���0ʓDϢ$��*�x�3��K)@ ��J�$Z[�<��X(7E.����)�'k� �*��c�^ѳ1�=�)�����,|3B�%�[3 �a���ۣ޼T��uV�]�2p��ʇZ`��pg���W+
�OX8|���o�4���Ƣ������o�D�������Ox��6���y�'�+k_8����O�I� ��|ZtJޜR���$��E� ac�����'��<��脜y%T�9�A��Y��E��8h
�e���N"ؐ�T�Ûc� ����K�K���� �9%<�;��8d����*�X����TG�;Y!�x ��P�JѲmR �I9��P��*DɲA�ge��FF(x�Q�|� ��d����O1����W�÷���K�KQ
�`4R�׿YE��i�Oa�͘�g��e(�P�ɒ�D	��ˬ9��[���`�'�4�!�vށ��W+`��(��$���r��3�8h-��	�a��9���1��g�d���hc��z9L��f]�R��\cӯ�r��tC��E	ர�SIA�x�l&jX�M�p��Ѓ��;ݰpkv,��@�5��?O()���&G�	 f@�-|p����d��rtT
���_#j�۱��% ���B�T`t�Ucή-,. �1K^	d��JBߟquf�'e�)��)��Ҡ��<q�d3ae� ��0Mв�T���/���&�����S{.�[q��w܄0�&�\��8��B�U��r�E#)"�O�D�� v��F!�O�"x��k�%T��d�)�"9�ד|e�4�;m����!V<5��PF�H�+ʾ �=�T �E��ĺ��V����5h��D�s/N�p.���K�I�'1�#�	�H��ī�	ޥy�t0�2��9��X�=Jid���e9�5��Č/��kԫı�X�[����r�i�'5�x�NTC�NP9��\�K+�i`�'iD�2�����$����&��y��S�O\P`���'�����C� ��q�Vq(	y� O>N�<U�H�?�QF}�f;D�Q:��Ȝ
�.���⁣J�&�A���?��?N�9�çg�=��˽� �$��~,x���
o����S�_��<9�J�V�<ȎMRp;�p�є�ы`Dʇ��$E�а!d�I1�d�IsB��:� �4'�j8��W4O�<�gF��'����H-'�b�'��yQe(əVި8R�����m�o*$;ׂ�;U��Y�Eʂ��ȟ�V�Ѣxh��S4L֕�����DS��y�N�Cd\����<�4d�T����y��''�p4��fјV�T��v��u{�G��k�A��.G�qZ�/!�O�)�K� S>tZ��Y"PL����h0�	6�O�f*���Y���9���r+ <) !� <���2bD�)PnL"ۓƌ�fFj_u�\��hڔ� ���Y��R#��<-
�����(���h1��)Gbȝ96W�/����I�1DL8G�ܑy8�}1�@4SX7#YX��h%�LӴ	��nC#
@1���I�.i�0E���4��	$�Ӎ6��	��x�kF떄.AB)��֤qeX�I7$uB�6&�)ǂ^*���)��'骉x��L�-m(3!�$
Ḁ��4QOR�밫��M�&��@)��T7�TE~�������$�0?2�bpR*3��ɡ���)L�H�3��~�!� �l��x�)�3G�������]�
1ʒ<\O>q�C9�R�X֋B)L9yӤ6��r�*�%=��#��|���K���	ݿ
Vm(�#Vs�$��U��o����sKъM�rňf&�$u6���b�p h��\"��JכBH�Qf��Oƨ��-(Q/t�C�����Fj��~R��XOBH˦/R�RE�	�a��zE�q��,��,z"�+Q̋0 ���<�Ou�$�RPy�DدR�9)����_����%qVhA?r$��J
/��#< m�Ht� 4z����!O�ARqO����/c��퓆]Ѽ8[�-�o��EQ�i �t��h�ś�%Xr���Lt��R�a�44��]&�V@Q-I>}�����)s��d��c$QU����ORPG���?iBP��dX@m�81M�Й��&�I3j�&a��) U:!�1h�)b�Ov�3ç�;"�la��KF7[��wi�s�:�!&�~<du%��O6�<�����a�4��_Mx�JeE�Q�\̚w�J��ь��9�Ռ��S���o�W
��
'�"J"�R2B�Z8�'ĔEZ�l��u4p@�B�A�E��b	�1��Is[6pW�1�!-GP�O�0�%�u'LU��H����4`�Ȫ5+&-�t��P�̉�����J�"RB"=�;*i0(���m��b�C�0����m��-�L���/��')I���F7?�I���ԟ�%%�0��Z�T�X@p��
}��C��)�B�8q�]�B�dp��(M��C�	�'���)W�d��%�nVZB䉭]���� Z��-C0L�;.FB�I�!:���(�����/��C�	�.b���B>c�����<�C�<�z D���`ҒYH��D��h%6�!���`�q�e�1F�!�Œۦ��G�L�<��}bU'�h\!�_���;��	�3�dx��/Ax_!�Ĉ,�(�h Ҽ��Ax ��Y�!�A$j˪�:D��E� T��i��g1!����"�SÈh���)c}�0"O��i�gL;�>�!��X�\��1�f"O ��L��0}�D����#tD�"Otq�1%��<��mAw�]0M�p�"O�i	P�K�*�Q�����$�"T�a"O��	�sNX2���<^�l+�"O�q���U.f��z� *$*A �"OH��q ���i-_*/k$A�"O8p�Ӈ�-��iy��o�|ڢ"O<0�m�2��1�VLɋA��S"O�$��P����`TU�HD"OL9BE/Mrzt�;'"�!� tH�"O�0�
Rd$ՠA@ޑX3�r'"O<�2D�B�fa�S��'{)����"Ovуu���i=�D�R��nk
D�0"O� ����Qu��]�#�~@H�"Od����4C��)�1LN�w�^ K�"O��0$I�:Q�z��Qk^3Lb@���"O�E��"�>�顠���rJ��ұ"O�����,@|����y.�T0�"O���#KC��0���p+\��"O�AH���/׊��o
�z8�Y"O���B쟠B�d��ċ�g6@�v"O���Q�07B���%b�-���;�"O(�J�S�>�X�C���(}�Ss"O��1`��F~~�i�U"s��d�"O�����O<�I)Gɗ!$�@�1�"O��aY+~E*�0(�m��IX�"O�$B<d�ˀ��\L�#��J�<)�B�N���a����+�e�q�<q��ɂ�HȠQ��08��a�B�k�<)a��J�
h�c(�'9 ��sd�<���S�l�5f
��Pa[�<�e�@�1X��q@�6D�`p�OZU�<a���/������Ŧ4D4,��o[�<i؏3Q��J��<�`��I�V�<QGc]�ư8�B�ݝwj9c�S�<­�/lM�w�h`Th�0�y�<i�B�5P�Ȱ����Z�L�z�<��MW�#ud��V�N-)�y�RM�<�G" �&7�MaQ�<�ء�_x�<qwg�R���IBj@Oj�q6-�M�<є��-c�(@�֓^Z����b�<�SF��J$y�.Ƨv1����v�<���� �������Qi`�
KDs�<�w�/��} �L:�Y��Br�<7$�)�0Pb!l�A%���T�Sc�<Ab��/W8B��G60L��1��[�<�T�Ik��-cnC�OkN!C���K�<GhXj
-r���I@��TCWI�<��3M��$����
(@�9 b_H�<y�BB0c��`� �'+����I�<)��G��`)�K@�L��tR5ǉm�<A��K���ڕg�Q��S
�l�<���H��XTA$c�0Ң}���Ut�<����UY�Й5+XwĘQ�\r�<9K�-,� ��&D� &ԣ�eH�<araG�h�QX�bˠmg�`�CD�j�<�4"\�n�B�b4�
�c�0��Ee�'�a������D(G��$��5,��y���0��q0�`�K}0��¶�y2�Y5�N]��KH81v�q�4�y�kžW@���Ȗ�1p^�iv���yҀ^0?�����!������"#���y��Y-HU�T�%�&F�&��g��y�.Y)ި��a��>��i1�,T*�y�	Y���:��TLP���0�y�O��]e����#ܗ�r�ʦ�ڈ�y�-�	[��5�	��R��B*�y�˞O�L�$�~�.h��B���y�N�4�c B�w�ps���y�Kʨ 0@"��Y#�hK�̓/�p=��}�A�9;;d��#Ú(��\�` �y���`�N�s��ȭ�.�q��A �y"#�����	a@B�� K���y2�ܓE�8t�g��	p�) �۩�y2d��h 	D����E����y"�؉c�v-S��JH\���Ç�y�εs��ucC�,8��D�v��y
� �!�"r���Ƞ�֊nМ<�"OҴy���0W������*�0�"O" #�b����~�|�)�)D���I�Mް��jM|[x��A)(D�tˣ��<{8���.��a%r]pH&D�Њ�T�{l��s��ɺ'�� *D����"eK��(7��]||8�)D��ڲ���>��� ��D�jrX)q�!D�  ��SP���DYBq��%D�ĳ��ٚ%�����nBW��`Ն"D�1�R���5�Êp�Ҥ	s�?D�4("D�;c��j64���"7/;D��L
5* Y+G �\��x+gM:D�| r���F�&�;&�#1�� �1�%D�$:'�߳H���R�� i���H7�O�˓k�r4YF@M,C�PDX���.��DG{b�'���	����ْ��Q�b7he��'�2 s"ːa�x�$ F9/�xx	�'!D�eo�:t��� ��,��A	�'�\DYe	���R�)6Oɘt�:�'BZ3�mҎ4�m�%썷f�v����$5Ot�`�a������`!"O^AcpǄ\cXQ� ��/G�H��"ObA�3�An�L�g�&m�̰p"O�(�t��D�.��&ˌ8[���6"O~��iŰi���6z�Pj�"O�ECaKF+��$�A���2~��zR"O>��㌈�4w�u�S���_�Y�w"O��Ck�%6R�����]S$�B"O�D qA�>>6��gžkބ)�"Oᚅ/�!Sd嚄K"�F`;r"O��`�(�5h�h@�e��(S��0V"O>�;���:���ir��cREqp"Ol}X�FP"�6K�FŊ>��8zV"O���T��m��k'Z2Y��p�"Ox���ī��ή*j��U"O��PU���M>����e�>Z�R"O��I��0yo��6D�J@���"OhP"�`ڈ&�*���ŉ%!�6��"O���j�)o����&f@br��A`"OF�@�mٓ	�HM��&��=�n!��=I�ڵLI�Y�\Q�e�D^؅ȓV��5q�4~tz()ѠN�6�x���G.�=��b�#4��x�'��OA����?� A��W�w�a�E�J6ZA0���4�n4P��N�)�, A-[	©�ȓ�찢jҚnsbHSUIQ�?rV��ȓL�����b	�2�ɴ�0<�����F��豄݈^+�@�A�"�)�ȓV
��9q�W�o�h�q��_r8��ȓx�	��A×Ŝ� g�~s�p���?�c��/�)��H��p�+�*U�<�c#A�B���� ,䠫"*�O�<� �(���Bf
\�Z��_O�<	-�_vbp�G(R,b��֋�A�<�d#19k�\�ʟ���Y��,WB�'�ў�'6��X��9nf ��I��" D�<��#�'T:��{�d��Aah١e�(D���%�@�h�1���K|�}���;D�®D�A�h�SV��A�}��O%D��ţ�	m5��e&�r�P���6D�x�B��?jJ�#�*�atXyO4D��k��j�[3ē�tzj�"�k>D�0`1d�?.�v� �-q�(�xע=D�� z�s���#�qP)M�n�����"O5��B�4R���VM'"���"O:S��	5<��xKg�̸.d  b"Or(+䍜*H�`Ȼ�K��7�~ܹ4"Or�B��Hi"I@ !��$��r�"OD�
�dI	�x��p @�9Y�x�g"O�X�ă�9<nBDش�?JT��"O����-Ұ��P���?v5��"O69:�LòL F��AnY�X"�TaE"Oڈ��À�z!���g����q������	�bʪ�5�L=`�$���DB䉯#���θJ���/*PB�	)Y�h�EJ��q*�Mb#�U�5:FB�	�Ȧ��Q�H�&��1cR�]�wwB�I +<9�E�V*��=H��Y94�C�	� Pf)��sp�9���V;l�&B�I*5E\@�Fg��*�ԅ0fe�RC䉈?v�@Idk_�o������B�1X�"����!�?a�B�	7w�`�
�� ��#�
� ��B�ɨw�|���جa@�0��%u}�C�I�(o�r�LI�z3�����JW2B��&P�X�Ɩ5K����w�׸��C��.�9���H%�L�"nU"PB��1;�V���Ʉp�4M�§�I��C䉻o�(�"���KN�y�����C�IoRrZ���5ʐZ�K.v�^C�I�b�u0"��)�lu��	=_NtC�I�fi<�`v'B!�@M�0�ȕQ�\C�	�v��j��/ =.������JC�I:*��sۥ?��T�J��J$C�@��%��֚p?�qb��qg�B�I�t�8ͩ0�*v&�]CC	�n�,B�IhФ,�r�Zt��]:	+#ZC�	E�5��
V�f`�5J�O�.:�TC䉱c��i�*K�1�EH�B�!D�d��w�B/d��7턘g�
B�ɷ�*��iM.)�J�iE�4YJ�C�Iu	*իe/R��0�*��۹[|C�I�0r�r�B�C.�tD�:H<C��#m��Mq�e �c��$��?�FB�I�X�D����W	4ִ"r�¹ �@B�ɳz�ɠ�V�*ѢZ���.9(B�ɺ7��d��-�L�L``�T*��C��&"8�@�L7Xr�\��œ�3�2B�ə���+�6_>���C�	1x����7 �)o��U�t,ՓbuZB�I�)���t��Wb����G�'�^C�	(I�� `�Z(
~�mA�3�`C�In,~<C���h�i*��9�"C��-_����U�4'zi"a]%fjC�I5Q�� �'�F1U���@*()��B䉛+mJP#b�(x�ԡ�D�;+��B��=R� �	`�Ae�VEH C�	�3
�dm�8� ���׬I��B�ɮ[Ӥ��v
�;vB���jH~��B�Ɍu8H {ᄤ\ф��l�K��B�	�U��pC���z����;�C�	"L�	��Q(DF@ps��W+l*�C�	�|H� E�ŋC�0t���Ȯ9/�B�	&h�D<����`4A�wR�B��J�%gW�e+��ZF�ݬ5ԪB�	�"�! �8	���3q����B�	�ys��!쁕7Q�})�O�Y��C�)� ��@��;�2jT-W��R<��"O䡹cу*4����+�0 a"O�����ʚ
h~�8�-G������"O0d��V�`3�)�g,^�kw���f"O�ɺ��5mu�p�%�	1gQD|[�"O|tA��8X֝�F�@�5S"���"O��{�R���̀��A�o��cW"O�xӇɒR�僒
PZ����"OA��Z�t�P�@�L�pZ(�JS"OJ��%)IR;��v�P:n05�U"O���bK�<b����dBD�p�:�9�"Od��"��'�B(S�
�T`Ҥ"O���b�pP�8�����R"O��"�k̔=D�\�A� ��"OfܢWÊ8{`�a�C�$Z�"O ��Ξ:?[̨`����0�@Y�"O�u�Ʀ���0��o5`Q�s"OJ�C�A�%	�Q�ˑ�w"�Yu"O�M;���0y)��E�B�S"O�,RՀ	�c�x� ���B��Xc"O(y���W��9���W4B�Ġ��"O�M��DQ��	ыS6a�B!#*O�5���As,�8E���F�J��'N�-���2U 4ƃ <�P�i	�'z�ْ�<�4�*��F�ax�Y��'���`釲5��Uc�ǇgBڍ{�'�����B�z�~��I7k��Y�'8^���|�bR1� �`���'����w��v4��P�B{�}��' �T�1fO�U4ꩫc��+o;d)!�'��ݳ@�?X����G��kY�t �'�(������d����B
�i7�$��'E�y���z0���6h�4���'p�\w�X�Clz���Õ7�����'�@#�Z$C�Xp�H�1�,�
�'��C�),��xB�� �H��'��T����$	�L���96NŻ�'�0���(��y���	%�<\{�'�LdP4')w��hh�7�8�'5�\;��[*h���`��I��'�ư`�mǣ����E��/�x���'+\ݙ�"��i�e�J"�0�'��QCp
D�z�bnY�P��M;�'�"���0�YG�s�����'J����U�I��%��]�r���j�'8���#x�$�����lbx�X�'A���`KE/RQX��U��պ�'���B^�F��+nBK���'��t�w�� ��}�1�J��8��'ќ(	"X%+�`��A�.dxhc�'�0�h� ʋ'���;�$98��	�'B��x��P�4h�MQ,g0��'ż@���#�.`0F@�$5��0	�'��
�A����8'�U*I�(�'^���; ��L��&��<��I��'E�PAC�Ǽ�j����:�l�p�'h��e�ŕp�``9��9Gor%�
�'�e	�/�7!�T���$X88.J1a
�'�
t�%�LD�i�ր_�`���	�'�H���J8�\�"Ɗ�2_�\�	�'���UM[�L��f+V�.}C	�'�J��c�5@��y����L��	�'�F@HT�N���F@�-Gx���'�J���!���������N�"��� �<�/�co��*�E��:B"O��d���9�q�I�p�PxP�"OltB����ꄋ�IR�*�T[�"O9���:U�
}���K���'"O��;�KT.D�� 1%���
���"Oz���ņ'�f��J��F��+S"O�� ���J��@��;V� ]i�"Ob�0���-m160@�f�4�4�Ѐ"O���f�<�T�0��V��u"O���E@'L�H�7 �t��sv"O��B����[#���Unۡ_��A�%"O�q3AZ�+g���9l�b""O����(Y�hn�(�l�M�rusd"OdI�D M4'e�E��#�V� �"O��9�JP_���cL�>�:�@"OvE��OL(��%��]:,�� p"O���b�E��w��%,�Sp"O���B��R��Qф(��`�-y�'x E8Å�!�@p��D0䜅*�'��Ս�u�q($B� ~�P�`�'f�]��\�[����F�{ ��	�'%p1�!�ֺIܾ}��߈x�����'eX,�0s>)�Sg�"�~�C�'�~L����	=��"� �L����'�ܸơ�:� �XR��9�6�+	�'s�A'gI�_FzC2��	�'��,�E�6\����řyi���'#D��)�����)��z*����'�F���Kƃ5�-��*ю eZ�J�'��h	peUu"`���ٜth�a��'�z�Վ�I���6f��䑡�'ۖ��&�hyl�J�"ކ4����'�0����ۅ$E�ยX<ӄ(Y�'��P�LK6�θ�%��;�X�'�X�1�E�/ =��H5�p�0	�'��`��>,����I���#VB�<����y��xa ��NN�Phv��v�<ᗅ��w?��˥��<gF%f! i�<��)�i�4L�Q�R3=��!8��n�<y'��J�(��W.W^9[���k�<2�D�)_@�� ��<�8����f�<�`m�P����B		gU�ȈG�Zn�<i Z7-�0l0���:/�8�A#�S�<)I`�!��U��$SceL8�ȓC��1�2����v��>v����Y���0n	k��� �!�\��ȓ	� 
��ŘY�ܵ��HQ��i)N��%+_� �H��I�j!�ȓu�rx�b��M&!�X�l�Y�	"D�zG�W�,���%R�+@L�7?D�\4Ń�h�:�F��`���S=D�T��,P��0�� "~/�d{�G9D�H� !��_.�u���2{V`@&7D�0�T��@>�"(Z7*�Bӧ�5D�t��M�
{0Qᣭٚ] �p�2D�xӀhR�0谪��V�,Uƀ�T�%D�h��82��l����d�Δ��%D�|�cJ��nct�8 �G?�L��!D�xJG�M>b<��v)ƤG/.d0� >D�dsf�N$w��`1π�#*(�Bh=D��r���O�4���^D8�H�$>D����D�e@�����Ł���v�)D�#��,4ܚ���"]�� #5E4D���G��$@�Ѐ��0u�rTY��3D�� B0ӱ�ӣLu�`3�%ަa��exp"O��Xw��)�B�#Ȥ����"O��Z�(ڒ$ȴ��&��n+ �"O\}��b�;h(�b�D�� �"O�i� �b*���!�0�ڱb�"O>�����1�>}1�Ƙ!"��h�"O��gbP0-,J�"$��k�`�0"O��;�A��q� ��7�� �dͳ�"O��cEH�D�䅡5�J�k�J��"O��RJ�>V�R�č�>��%��"O�k��K�_�V	�2Q��pC�"Ov�[�3oU �3�!	X��I�d"O�4�B^�S�N�ZW'D�C�nTB"O�`��ցV�"Sä �8��1aq"OZ�"��?DĲ��UD�^��2�"O���!�I3���cᓨQ�)AU"O:L��ꉶa6��/T8-r̒a"O�eɐ ��!�?䢨B�"OX�{T�A�p��i@-w8��"O0��$K�er�\2$�4S�d=6"OHH��H�"]�$��ʆ(7�T�"OV��LR�]��@�;�Pee"O���4G�4>N}��b#9�࠘�"O8�ڃ��n`�t�T��$�"O���IY�dܶ[�@\����)�"O(0����
"�q�'eړ1����"O�xy�4o$��cR1-�9��"O�	� �8FBZ-;���/�$`�7"O(]�bL=t¹s�DW/w�0q�`"Ol4&!��N�aJ���<�6U�v"OV@��� %p4�����^�6Y�t"O^x�6"ݓg�`�e�=^���'"O̹�DBE^z��E����4"O�QJ	�^�\8�$�(
�b�SF"O���6���dvb���
��<֚�kE"O,�X$���s1������"O�d����:+��Y�T�L&���Cw"O�}U��F�@�d�G:D��1"Oh����J�W1D��
�b>��B "Ov���!��U8�{�(A*V,�)�"O�)Z�n�&	�^]���=��u�d"O��9e,MD	�ZV� h��"O�pr�⒧&�&�e@6��"Oy�Cdƹq�"�l��i�F�z"Oԭ�'
F\H��s��	U�<� �"Oڡx��P��q�f,�3Њ=�c"O8�MږHR���!�u�$=��"O$"lѬ
$P�P���{�:4I4"O��!
	wj�<P-�j1�"O����K��m"l�1s�N��� "Op������� w�p "O���bj�HXԕC��([�7"O������*~�N��VF�P�@��"O�|c���:��iB����G��9��"O:DK���I�r9j6ƌ�cuX�"O~�Pp�zS�d�腀WҠq3"O��b%��v�ػ�HL/<H��2!"O�x3 ��
l�J�� 5=/80��"O�M�'͟H]a閬ԭ �*"O����M,m��� K��6�.=I3"O���C�\<&O��c��4��\��"O��ծX�6��"N�0�̝CQ"Of<��/�5աá� `�*���"O����C��7��-y�nÂ,Z��Y�"O� h���烻2$���-�4SpK"OR�j��	�F�K�A��m@Z1�A"O��k؅'s�i��A�:�]bu"O��D��,]/p ��a�0tJ�;5"O�`ᯖ*�@;���	IA��F"O���Y�0w�U�R*�,u���"O�σa�:a�0J�|��t� "O��s��eh��aa?&�F�!���&�*����E���T@�zY!�d]4��Ѣ!ɘ<WP�[0��8G!�$^�C�Y��dG�(Ғ�Y$!�D�9bҜ�s�֊8��c��_�!��V�J�0�ᐏ�P�t�P7���
�!�$G<|���ӳ�Z�2�t$K�>%F!�D�mɐD���#pfy�Ae��t�!�]>2�\�b�Bg�Q�%U�Ns!�ď�"����(O�e�
�+��6�!��
$�4��r��b_J���@�!Y�!�d�K�ޙ�� ��C������	�!�SI���"�%ҡ|N��� �&@�!�	�o[���ƂS_VPZ!�՗n!�$�*2Ih�IKi�B�"0�RTj!��o�n��"Ǐ�҉�V��t]!�dL�P��#�e��I�.�!�D��浀�� g�~����ϱx�!�$0k�(�c-Тj����l�!��D4,���)M�	�&�p㧟�zl!�D�?Wg�!�t��9�ލ��>`!��6�8F,� {z�lyT q!�$Cx�&�P��H��
Y��s�!��c"b,�u�I )�b@
Q%�!�dW�/�X�wlO�92|"W"�4�!�Ą�<�^�����-�*e��ٔ_�!�$�>/x$�`Fʎ<�B�r�GK�!򄚓\��Ű�lM7���DF�I\!�Dϵ3ȌP�������ʍ�!��vzM��%��>����B�?�!�$�9TS����g��l�/�M�!�Ւ.������+b��������!��T�@�lX��Ok5�y"
�u%!�$N���!qG̑}�m�⊑�A!�Ė?���� q�0���˄)7!�$��JD)��\g��%ÔɁ"LM!�N�V=�H�㕘Ӵ��d�!���H�0��CL�G̐����S�	!�ʀX�g� '��1�C�,M�!�D�M�dA�"������.�,:�!�dF�(��욦F�$6ڦ�*�.��!�D�OCP���Qh�tf�(y�!�d�0(h��=P6��Gn�49{!�D/z�$�rb�0s�D}(C��mv!�$�+.�z`+'㇦6�d���(_!�M7�q����]a���>m�!��!�갑��DQ���kK�!��J�kM�샆��n�)��'M �!��>L<p�">�TI��A.�!��Ʉ.�2Xh�$	Z�B}�� ��!�dE#*��qA� .�HԀd�أv�!�$^?��q���̩b�*�3 ��x�!��8S��Yi E�� �i:���4D���6IP
Hb��Z�M�:TtH+1&D����� &H�ǁ9az�pb�&D���M��q���E��.
tz��.D�P@�o�p���1���G�.X�)'D�� ,-H�^8.|��@�$��А"O��Q(F�l\���ڌiEet"O��l�[(�����'B���"O���g�ϴ%Y�id똂?�>P�V"O"yb���!v-��f�4��h�"O�X���*@�д��a��&����G"O����Ĉ�����pt�ͨ�"O*���\v�,�
l����"O��x!��'C�!LHwޘ�'"O*x ���[j�\8B��rh�r�"O�M։��6N��� �O�]�a"OL��r�� ',䀶W5X�8�#"O�m�۬cN���WN��]L&m2G"O������xS�, h�,l�"O`��'fA�t�z�ᒁ�j��`"O4�ZF
��l �
H�(�ʐ"O�� ������ [-^.���"O��h��@ E8-�0%ژ G��P"Ol}s�āF�4�`E�tDYh�"O�pk��J!gen$���V+71���d"OPuBR*�a�0 �*.IN�HY�"OV��7HN;�Z��F�_Hr�"On���V�(:���ȓ�.�a�"O�-S�ȁ�v�JE�F�(a�8hW"O� �h���(d�-IJ�T��"On�k�䞜@@m9e-pI0�S�"O,�����&"�e#X�hD̬%"Oڄ��%~�(��a�*St�#�"O�i�G�A�E�0٪&�[�m�=�d"OZ!I��\�#!F�0��;�ެ+B"O�m(6eYͨU�A��TujP"O�A[4�_��0�!�+�椳�"O��"С÷L�x�ݜw�4,��"Odm@�Z�ip��:��G)^�pa�"O�Q� �R"D*�ro��ږh�"O� Ä�֦E���k	�[���y�"Oy���;! :�Z�GX�A��"OJE	�F4K��{���@�^=@�"O����N�h�6��p��h岰35"O����ۿB�j���Yi�P�"O���fG��<��@D�!\g�ȋv"O̥ڵK<i�����D\t� BV"OUz��K�#j���C��Z?Z0j	�'�Ĕc�,� ���?�f���'yN��e"a�"%y5l�7u�E��'�i�F��?S� ���HG�*�*�H�'����"K�`YLh�,��(��<�'R�A �J e���O� `�`��' ���2��;3P����R��xX;�'Y����̖'��l�Ǌƨ#��9�'74	��P�X4�Pq���0�J�B�'��٠$�;^i�)~�8���'�
]`�͗/N^FH�0�D*|�)�'o^����T��j|Qu�_��eR
�'��|)B�ï<k�`��G�Y�*�Y
�'�l���fS/!궹��ƃ"<�F؉	�'�t�Ѧ $����f�4.�pP	�'�jx5mR27͋�7ϖ$K	�'G�@��Ã�|$�yɦ�>�@-��'N���e�8ow��q�BѱJ90���'3Ιp䐟4WVԲ�m�	N��z�'=��J�N�'vـ����A�Pɉ�'� $��J��%�.��T�T�	c����'�3��_�yTb��À���� �͂�"��x�BI�wE��"I�xy�"OX�2�M@x6]Q��ԂEP�4c�"O
���ԫf:���Ĉ�927��"O�E���V�2�<q�PF�THA!"O ���+GNx:b�W<>М�6"O�١3mH�	zl��`Ă�0�@"Ohͩ�'�D�@��f`��6����"O&T�wk_�[�l1�ѮD��`���"O���ƻn��8��ĮH�T�"O�����$:o��C��	4�&t� "O%`��0n9�UєN <z�E*�"O�w��-�j��͒ue�1J"ON�����c'�F�(��z�"O�5J�Q�AҠ���[�LA�"O&=J�FG
{ `�a0T�j�1"O�8"%gׄq�J\�'ᖚD�1"Op�����A�v�(ƀ�($N�"OfL��Ο�;3 ���"#*��"OL�)��ԛ[�L�hAŋ�}2�"O�=jᭋ>/#XL#�o��ۂ"O9�W��](�l`�I�9��ȳ"On@�T�P0dk�
r阘x��"Oȵ��AU�A, �n_�#�D��!"O`ڥ�߮^����Lܵf���B"O�yP�bՁ~u���&8|��'	��!�,�dI��S�l��iS�'pr�YR�A�$dB ���˵��� �'�Ni�ȚsMZı�d��X���y	�'�d(��%�1q��]Y�d�#�b���'��D�,�9w��u�`Q��D8h�'���I �ҎQ���S���p�'�|@;�`�~NXq@��[���H;�'���Q�I�W�}��[:vW�	��'�lma���Y�\�{egƷsv���'��X�S���eir�ӤL�,]�X!k�'�2�R�I�=-#J�`����'��hb� �8H�0�2��!
��`a�'u���D͔5&
�7̝�y�pp�'�HY�֮	)�����.j`��	�'��[ �ܠ"it��_�����'��XyC�z�:G�*"���	�'����v���K��2��� ���b�'�,y�I#`~���(�2!	�'᠐b�c�i�"��V�(�@�'0�URSO,�@
;�� ��'}�@�������ʀ���u��'����!י*�^�Ұ�Ȟ0�����'�ڠ�Є� @���b��V��y�'�B]0�jB�8+ a��-��*S�'�Ν�G'.U�=Z� ��j�)��'!
Rb���g��R���~0����'�F��¢N�lw��Ё�a���'��h��-��"A�i2��		�'+�!m#|	TH�(�);� �qG"O4�
A�@�/vl��0&H�  F`�g"O��6�^�A��� ��3����"O\��&'S�e�`��t|��"O�i�cȬ�AQ��8/�(x�"O9j DF,}Kl�Cre;MK�P�"O�
%N y�O�?fM��"O䕉ulN�� ��BQ<0J@���"O��q�w��@�����x�hD"O
�мG5#����(��"Ovɔ��9�\E���݇Br�"O� ,�[����Ō�30k�A"O��k��Y��x�
�kɢ>��5��"O~Ѡ�G(E�NY�V*�q� �B"OP����$�X<��n������S"O-��	�v���M�0)�D�"O�!'��� {������E�0��g"O�l��,E//�RIzC4�D!"O>���,Y���E�ؐc�{"O��� ��S��h�O�h }�W"O@XXE�R:Ժ�i{��""O杓�A^!W�AA�E�$�C7"OrЂ��<�*�F'TO��#w"O"���$��2:�٫WӪ�䊵"Od�%"���0�A�	� "O�e@Z�M��8��O�<,�A"O���U� KN���&�"��"Od "cB���̳�F! z�`W"O�u+��
4y��%N�za�pZ�"OB\���D's��ʄe�gpˁ"O�+�&.
֊�
��7nY(�8�"O�	*�@�� {:Y豌
X�~�*�"Oe[�A�1OP��'�
6���!�"Ov 9A�3|��	��҉~:��"O`hq��5� �LˇBnX�"O<�!�]��W��Eڔ��"O�R�nE�Z��h�F)Q8K��q�f"Ot���.h|9�Ǎ%X�����"O� ��T!dX�H��
�t,A�"O�Z$jՂY��0Pd��� ��"O��b�;y�Q�%��=����"O���w��/8�2ܰ�.b���R"O0�I� ��jV��e�ݧ@t��Q"O Ai4���cW`��}�8�3%"Or��!.�/�����Y�Q �RU"O�H����
��*e���1_*���"OR5!���%QI@M���?x?���e"O (q�E�;B�`FJ��7���q�"O��I�nӐy^���	�.�$b�"O�i�pAQ�V��Us��#��e��"O��ɥ�Y�4@�� ����x�"Oh�C�ζB�&��M�q>��f"OJىvf��?a�U�Ɠ�o�����"O��Zu�M�a���x��G�.���bt"O.a�l� ^�<D;��z�n�(�"O�ɫ�&�.?.���F	7+��1"O�St�`!Хy��ҦP!�Q�@�r��L�f�H���`ѣe[!�dY_�䅑&L'G�^@ʧAJ�4[!�by�i#mZ9>����抈�"T!�d��X?�5�����T��T��!�G3~�4-u��A� � d�$y��'#�q(↟�3S\0y1LB<$�.��'�.��ąoFD� ��"+ ��'��ǀNh]P�s��A�L
�'��y�#6fNNjc�� �]��'&D)c,X�/���&BN��'.��J��X�bT��X�KP� ��A�'� ��l�]�m�s�&��'��3n�>u���Em�c�����'Z$�����}*���t��H�1k�'Yf���Aݴa%ҁC��N)9Dv��'r��Q,N ��$ 䣕8�0��'؂A��!��IȠ[�F�J�'�^Y#��ف=%>�:�W������ $�*ƮE�)�,�h�( +�Jp��"Oh2�ǟ�
�~�`FG���y��"OD����U
y1v�*��w���"O>�B �	�"9��gϻx��s"O�Pb���)�����9w�$ͺ3"O�Y�t��tz,�!KV�`�b�u"O"8��B6�(�0��� ro�\ه"O�U��/t�l���bڦ#Rm� "O~	x@�ј>�6�H�!�%�ڼ�d"O���!����J'��A�P���"O�yG+Xf̼���E
n@�g"Ob��҄�#D�Τ��S�J�S@"O�P��C�X7����ō��EA7"O�%艤x�+Fc 9/˪�)#"O ���C#��d�ł���4DK�"O��h�A��Cj���� ������6"O����Q�1��Ա $f��Ը"O� 1��O�2�Ƹ+�Ő=�9��"O���d�N33�*Axw��|2<c"O�5AE#M�(���-VYi:E
�"O�1����
L����UL0( "O�8y��׆3;b��+ۀ
,�5�e"ON��%�/��K��F�Q"O���A>[��C�`�`	��"OL��H\*_a�{"CW8M�N���"O�q#�L�p��t���.���"O�����5H��3��
Z��%`u"O�41�:eR\�C��.���"O� Y����=x��CBT�\�
�Q"ON|��n����2���J�P�a�"O`�����$G�/c0|��"O��Q'�C�(�b���#�^���Y!"O8���i�2d�HyW��3�
i�"OL�!';Y��%c1a'\��%�V"O(lz�%upвF��
N,�""O��YɃ4{V��,�0{�a��"O �ӂ�5}X)q��U�t~4�B"Oƕb%�P���2�B� _m�Y9"O�-b��۳/'�Dz�c�h˱"Ofd
p���8�#�
%9=���"O�}i�M�^�Zȸ(K#82�`��"O��1��Z'FpCF�F�U�P"O�P��M�<Ly����6�j�"O�HR`���? <	s6�=���X�"O�<` �T1�
lY���$K�F=�p"OB��� �-�����S(�� "O��*��4y ��� �pqfL@�"O:�H�A�X	&�QcO]
}��"O�e��$Q-c����Q߯@Z|�	�'����@(^�₦X����	�'ؔIT#Z!Q���E�/���'����d�͢�͌\Na�
�'B98ԥ'uj�Mʄ�V e̐��	�'3t<�S,:�
h��^Xl�	�'D�]P≅��Ќy�cM�[�8
�'��<Q�o6!tr�Acj@�*^��	�'{�q��ɫK��H��h @Z�s	�'����s�S'c��C���H&���'X
 5�)d��:B�WJ؁��'��ղ���\2r�M?F;�,J�'�xPɥ���
��,�Ѣ�%E�L���'�!����I T�j�FB�5��'RH���ͤUT�qЯ��{6��J�'�عH���+h�5���Ff6����� l:��yj|=�'���h�"OD��BI,(�N�[�1V�&"O��+cfU�:�2�r'�1鬨�r"Otl�f�@[X�5A	��u?�y "O\,[�F�0v�QI���'j(H�1"O�AQ)��,`H�C�E�2n���"O�̈`�ٸ^b�ŏ�[4��C"O���Y�������.+d� @"Oz��AKH�7��0a���
y�Ar$"O����&�"h:@!���2`~�3a"O��a��  !H�
�!�4�4"O0�	��e���#�+x�F�(b"O�1�d�O�3�@T ���Z�:�"O���GM)��l�db�y>��zU"O�]kGDB�;�~I�㞣EQ�]��"O\0����>)�Y�¢S+5.pIc"O�X�$�yd�����3����"O�HGi�5F�ڭ���䓕"O ���M�7��0��c� -�� �"O�T��ǆ	j�uB�L��&�6a{�"O�ٸ��jYZ׎�2�8Y�w)D�<)W���:�-�w�D��*e���~�<��"�a��lPLք�6uaf-	x�<�b�T��j$�!׃j���ǎr�<閦�y8�"� qK��'I�q�<��ȖZ�]a`�<���ȕ�y�<�Ũ3ha$Ÿ6F3s�����]�<qG�#Y28.��V�@�t�<Ɇ(�/h �#�{�bA��%@[�<�A� �,����4����M�S�<Q��E�
�"�i#�Ç[.��#��O�<i��z��y�gwfx���CO�<���_t� ����b��<HqEJ�<��@O5[rL�2A�a��MpfI�<��d
�,��c�J�6�i+pJQ�<	3"�=o�I����;9����dnH�<�"�:-��Crm�8J� ��ȌE�<�'QWy�`A,��d� A*�Jz�<Aw�׀"bTUH��T�* �1dw�<�C �91N��#N�hȼ�Ǧ�|�<�P!L� �,i�↎'���jb$_|�<	���"�^P�1�
o��MB�]q�<�0�U�8� (�R��>k~Q+r$�q�<�w��6i0���,:M�ڵہf�U�<��N���pE���\Y��D�S�<Q��k��[�D߇��%�2%�P�<i3T($R�c�țy�5aQ��I�<9tǙ pB�BQiR1@\np�D�E�<.Æ����U��+#�D$��<Y�-Am���+F��A�J}�<q��.�Πs҈�<y���m�<���:9$��X�(
^f��84�o�<���0�#E�w�����l�<���CG��!�Ģ�;]{�`��b�<IfB��FG��ƀ�1f� ��"�^F�<YƦ��s���7I�,;r���#FA�<R 3T_<AQ�M ~@tsT��A�<	ĭ�7^����P)�+,le�Nz�<Y�E��]K\��Eg�ui�ĉr_N�<�š�:qu�UeKS�C��i`�_N�<ɦ��{^�		׭��P�(�H�<��&�X-�56�I)9C��Q�_H�<iC��:��BH$+0ؠ/WI�<�ƨ�R��wpP�飬ڴU
B�)� \yKS�B$X��<1�! :�t �b"OH�2�N�m�x|z#�E�u���F"O�C�!=�(�u���GD�p�"O`t�� ؇��d($�DKC"O��,ͨ~^-r�i�?{r,z "O���VGxI�%��� bh�l�"Op�v�B�޹;r��UD�9�"Ox��W�ۭBjzU'G��bc"O���BAO)7J2mYg�#�p4�"O܉ҬݮG�N��W(����"O�p��d-5��1��&[����"OhLk!�\��Aa�-my$�5"O�d�����4X�3��#/�,@YT"O�!����o�4;v)�w���"O��[2d�?^�<h�U#ʙ1Z �[�"O\y��� 5����!
(Sl��"�"O��vܘ^҆Yat��;H,q�"O����W `p�0�Ε�ON�s�"Oj�X1dQ4~�l�4��"G���"OP���D�r�TX���º^/VɰE"O���&8�B��&�R�E�"Oʘzqh�;^\���d��|#6"Odّ�N\�lA�ɹ�B(%���j"O8XQ�ׂ(Ҝ
t�Ӿ!�� P�"OrT�f�X�NZ���_$-��"Ot��䍂%�s��A"O�2�"O�2u�O42��*N�&�l��"O�@�B�*�pA6J���p�9�"OpP��S�=K�pu�3~��`%"O�U`Ut�򑀓蒏e����q"OV�FL4^p5'�`F i�"O2Hap�ϑ;�\�85��w�`�2�"O:X{���[X��0&\�
���"O�<�1�N��]*F�G�����"O�o��:�F� R�ڱ
��}'"Oh���FC5�ʬZgI-���yb�V�S֤��Ɗ�r
����bŢ�y�	�r~ॢ@C��c��Q0���y�Ɣ{F�⒄І_�N�����y��M�]�6*H�N@�1���y�k�R�t��a�2T���³�yҠR8ct82H$(L+&ʞ��yJÖ��T3q)\��;0l���yR
�S��u���M|T�Z�F��y�ON�IPv�ߊNھEa�*��y"!�q&�!3%�C%��B�3�yc ���(�Ġ?q�F�X��y�IA	<�J��o�����]��y���(.�� H7�
�p,�څI�9�y��7kXX�2�(]�ap��'�yR��2%��8�e�ǤQmRyp�G���yRC �ܩ�7�� O�f�A�۾�y� kN2�2�Ȃ�M̴`�0���y���^�>��ҡBs� �ՠ/�y��[�y�
�cG���76n�It�ד�y�G-�$d��˲2�ha
��2�y�U�@^n�S�i[�Y�^�a�\ �y��Ҷ#"�I��}	jU��'���z`iܓ5G��r��M(�0�"�'���Q�@Ѣ>� Ez�Χ6t���'�n���P�4F�h���,'[�)��' ,b�l�.\����'�9�^LB�'V�j&*Ȧ���H1��4&��+�'��!��эBp���&�:�I��S�? �Ġ��39ΔQ�K5p�ð"ON�T��.ׂ((T�9M�Y�"O���iԕ4V � 3��J&"Opq 0e��"����ϻ#+�9H�"O*�x�	�:d	y��(��2�"O.T(�'�3|��a�G�0�`�"O�����?
uPWGN�*~��"ON�R�N�u�`����	���"O�[7b�=:��`<@��� "O��#���cM��Xgʗ=־�z�"Op��Ȇd��r&O�h�L��"O������dܘb��h�$�Y�"O��#�+�+G����d�%g�$�
�"O��P��jO�qB����'��E��"O<L��n�\���Ga�[G"O�b���/y�^A��J��!��"O~�q�3k���RW��o��ai�"O
�8�c��"*,)WH�66���*�"O ����-	z̻��(3�V��0"O<���ٛ�Z�����7��	 "O�y�e�H ?+.%�Uʞ�(~�hc"Op�CDZ�m�0�T�ɘ
FI��"O,�ଡ଼�>�����w����y¯��6���@�$k�=3���y�OSR\p���	�7{�B��&@=�y"'�,��Y�&�t�F=�Wh���y�X*#�`T�"D���b���4�y���-Ʀ��W�О��\�fQ��y��V�.l���o�с1fَ�y��\�v�f��  ��O�0��g�L�yb�E�OH)��`��K����6�y�/�<{q�y�$�A�t(�듛�y�K�='��(�N�5������yBG�VT���	�-v  �8���&�y�"��!A6�L�lM�<c�˛�yrN�$+�Ĉ���O���� J��yb
W�6e�LZԘx�S*�7�y� Ǥe_z}�sQ�p����y��7t��1#��
�) ����뉅�yR��
p�ّS	�/OR����#�y�C�6_�6h�Ջ����I�����y!YvC �ɑ��>e����ؽ�yE�5��|��I�	�0�taJ3�yb��&Nݰ,��m�&�Ri�&���y2oU�84i� �Ӹ1D-"g��7�y�h��?�L|�o�%~�ك3���y�h��5 q��	O�iá�6�y�45يP����6RB�u�%I]��y�o܊6�䡋�o�E������ٔ�y"`F(��� �>��)�IV��y�n	�Rc�Y��ȑ;E�Kv�I��y"�I�pO@��e��'8G� Cvn�)�yrG �lR��[W�ϳ%f*�YB���y$F�?�DTR�h�v�uن�Ǟ�yR"�R$�P1R��=X�Z�t�<��b#���M�'Z�����-1�I�ȓ����|�"�j�@Ș^[�=��A]�<�Ai��b�P
 #Y	B�	�^�z-���
�OϘ4b���=?��C�I+&H�����:]�D� �'f��C�I9�zi
ġ�~6I�*��.�C�	��2�� ��ZHΥ b.��C��	u��,�wnN�m�������.B䉩
i�<��G�iN-�V$	Sj B�)� ��p'۠�:8��IK)�t���"ON�saa[%��8�h����"O��Dـ:�B��'��#��!!s"O>HAr&E�%���[FE�Z��*T"Od�@�N�$E�^�y�C��^�zl�g"OZ1�d�(a�>ѨPCA5��C�"OXX�pkG<$�B�cPE	�:��c"O�)�얮|7xL�&+�=�����"O^$���?��!Ǐ1��)�"O|��El	5>��9s �M���%"O(����51�`��T���;�"OP�w.O���(��̛[hp�*�"OR�{��M�1���7n�Ph�l�"Op�`/N[0�ql٪YX���"Oj��ۛ=����p�dX�3"O�u�1�tќ�X�զN��ixd"On��ƇO�Fox�%Ed���"O�M[Gi�Y+,��.��~ƙv"O(9 1/N8x]h��͉	2c�"O�tn�/XN>�Ð.�@��M3b"O���E�ׄ\�=Z欐�J �[$"Ox�u��*x͎E�	*a��*"OL�˜�}�(��%��G�
��"OJ�8��_�렘0�M��~�J�b�"O6<�sK̀" ��L�;�Tԃ"O�ݳ�fXO�ݱE�#�0�C"O��CN�5 P��!���6+qr�ȓ¼1�ӪW�u~Yt�3ke:i�ȓ+�p��h�=Є鰄�R�ń�pڍ�ч��~K��c�oF�b�>��E���dحS�BT�6�U5��5�ȓ*z�f�.6��;W3�X��y-�xB���:��D�$�2m}�܅ȓK���r��
Cb�t`�/���z��ȓX1��Х͌�Fui��"9C�	��K�Ʃbh�5�d��-G�h�6�ȓbe�a�f�-D
h��@.i�����(B@qBf0s��,O�Et��ȓc�nб� �eC"}����At�d�ȓ,�X��@ vzRMJ��F�R�8��6G�����^���Y��QT; B��=\1�պg�����R��%mMT��7ѾK�ԭSl*%Z�,E7Q2���/�����\�%Al�)�"���ń�i���4�?������C)�4��ȓ��1�Ai!C`�� �T�H�q��?����B����]i��VIX��p�-95�Ǭ-,P!��; N��ȓ,�da���[6��!�K�.U"��ȓq�����P�4�H�� �4�PՄ���4b���[z\��F%O5��8���Z��\T�]JaAN#ZE���[�@@���2UK�PRiB"FQ氆ȓ��|�5�+ 4M��z	���� 9U+t"��:y���F5/���ȓ=����¬�ƌ��I�2��P��.rFE�ܜz����,+ְu��uD���禍��ly�$�&ꌱ��	N�e7�ܤ'u�@+�80��ȓjv.}򄅰��8����;}�	��[v���/��^����g��ȓ/e�9����R�B�H��� c+�ȓ3%��ڧb��Hp�� ��>Q����>K���r��=#�@����~���S�? j �D��V�~���HY�6=�a��"O\���L%X�x����$��9�"O�Ļ���}�q����4���S"O����[wp �3��=�v$3�"O�a!���6�0���̺҅i"O��PK�\��԰'	<-ّ"O�!���|�4��֡�?�=�"O��S��I'$�[�f��5�B"O����Щ�N����5m-p�А"O�ٛT(.m�kpd��#�TÐ"O)���x�4\����r��a�"Ola�3 �Q��
��^�c"O�4Q$��s�t B�o�j����E"O~�rl9/�1±�C�(�����"OvA0��ң|d����Ə`�T�E"O�,.���l��;8�V)��"O�Ay�K�����7흴
�<�;�"OD(p5��4�
t����.�
�A�"O��� ��Q�Ҵp!_�o�\t��"O4�`C�8s��g��C6�Cd"O��1%���.΂�� ��+0V���"O��`d@�<9#�h�I�F�T�"O$�r4�	|[��+���?V�H�d"O:mȕF�m�|9$�8�Ni�f"O� "����!�2��&2~�£"O���V�ȫe)\���y#����"O<t�r�еh������[�`~ ��"OĘ���Kg� 5�`!����"O���u"O*
�\���%��|�b"O�����"f�$��sn� |ԙ�"Oʸ�f�����y��u���C"OT���'^�R��B
���#R"O�	�׭H�\�V]�$	�)��j�"O��������(���+2�q:�"Or��C�S\�ux� �G�=`a"O�+��X+"�.6D��+�,,#@�(D�,�Y�&b���1a܀1��@)$4D�������X&� �6��&i2D��b�
�U�b,(�/X�K�z�ꦏ"D�ȓ� K+~��eJ"�X�M�|pf�4D�0�S��"�虫�	$	0�(I��>D�D�"K'@��Mjĩ� 먩{��>D��I��#��PY�ھ:�`�jf�=D�$�'�B/�]k"�ұ&x=itb:D��d�N@T��ЖG1& ��7D���$҇!�ic��!q`�3��6D��`#"Ѥ��xP	H�z<nI1�n3D�̊©����Zg g �QS�1D����0D:޼��d�D�� �-D���3�*U1��0ըը�\JR�/D�ظ�A"dN�2�R�w�윚�,D�8ۢ�D�J���iC�Du�@�u)D�P�P�T�f@��	�'F!��\�W):D���GoD;ޒ����3'� 9���;D���goҁf�N�����v�4��A9D�t�
���	X6�CLԤ|�[�y��"?'r%��8�t��	+�yB�u���q��?.-Ԉ(An��y�d��?�\hԈX�ӀM���(�y��{���0���Y��� �F��yrJ^�ol^�2�ń�J�P)	pI!��xbjɥZ�8�V��1eމ�`Q#{!���=$X1�f��X�M+3)��H1O�c�lhC�8�I��Y8c,WD��f�U�d�C�)� dlU�Vv���j��Աsm���i�'� �S��M��/YXÚ��%a�/xn<g�f�'�ў�"jN�W�ʑn��h>숇�D?ĩ9ì%f� n��9&���$|d�Sc��H���d�͖��ȓ��Y2�˗sA�C�('E�b)�<�	ߓ�&��j��j�Z� ��9AJ�ȓ
�P��K7v|�Z��Qp����)�(��F��	7傝z�+ӽB��ą�igL���lC8j����G�LnLExR�'!�a�a�� �J]!t��.N|�)��)��<yU'��r��/�Y���[�	d�<qGD9u�lC�+���L�"��D�<1�隃 5�M�tC������A[C�<�1��U�Ҥ)b�[�6�8 ��|�<��)<�h`vDK4�( �I�x�<���C�`�v��c	��P�#���\�<YšXs΁
1�V�.�<�����n�<i���q�Ef���`�f��~(<q�4r^�`�u�'x�QW�E�δ��	a�'��� 8��J%1;:��ѧd�,�Y�a*D�D��2�Д�� G:r��-D��:S��G7���UEI�L"v�P �7D�@1s�#��8i��þ7�ZT ��7D����N�s��qG���Om�u�0�6�Op�.���P��kL~�dB�Y.L��6�L3��Q� D���.ɪX���G|�F*�tsb���h�qf���kZ*+ె����O���c@�!�rt/�M��y@u�Oԣ=E��`�c9�t"ŋ�{b���d���~�0O�O�"�u)۬ %�b�D�EK�)Rg�d�<�#O� �,��q���t����a��p=ǡ���~��s�S*>�8!`�N�A�<Y��X�"�#L fe ���b�<�ˀ�p$P��g�փbb�9+�v�<�%��Vh�̑� _�h�#� �G�<a��	?� '�\�YTx��"��Fܓ��O)`��	��Pd`v��.����'�ў"~����%�D�4Ǔ/ْXpU�PG�f��H�0��LF>(�v���R�K�Zdڷ�'��	�X�D�%L=Y�d���f+� ��䓹h����b�b��"�s�r�D#G�azr�O|�'������B�����]��M��4a_�=E���VV�b�
#T�W�F�+_+��ļ>	�y��4�'���bE�6��͹%ˆ�Ryl8���d&OΘ��bή\�f��$+�ig>���"O����z�P�((H�F^�aSO���Eݲ5��Y���+��MY����hO?��*#f�R@$�+n�R�!���L�B�ɶcn��CIӤI>4�2/�8"�p��P���i
�O��@ /�@�P�	��!�$s�fE�&A�5 ��3�+Łg��ľ<�I>�Ϙ'�@��!E:e�x�Ǣ�[{rr�'��\B�Iѱ%�6�KƧ�?� ���'�V�#E�D2C��\k5�H�1�R�3	�'Ib��'�/�D���\�/-���'>V�`Q��vEL�F3|��e��'d��i"�ђ�L`�v C��Ne��'�>tSwF�30y���M�*�[�'��s��Wδȹ�)N?z(�
�'^ �`FW��3��C8"���	�'(�K ǃ`z�X!�*�**u`�;ܴ�?�J>��T?�+��I�A��:%D���:)��*�O䘦O`��p�Ɨ�"����
3z�3�"O� X���J���:P)#�-A1̤1��	
�0|�C�#�F�.J���E斺��x"`"PF!!��Yl���I���y2d��u�@u)Mc�ļ�O��yR�K ��9��nZ�sb�J"��䓘hOq��1fވM
�qt��/G�5�"OBX��SH��\:�F�*v<���'��PD{�O4!�7n-t��	�ԯ3P�\0��ēT��\��N�09�����5����7��Pt%�{Ъ�"P	����Gx��)�tIY Do����NТ6����alu�<1�ƶK�q����.e�h�0D�=SIB��3�g?ɖ�Ϩ�����	��my6��n�<��	�3
t��F�55�t��Nq�<yw��-O6�䇵BY��Q4`Y�<�3�@�%'�`Y��1G�=s�b�˦-�_Đ��%U1x,�z�熸 :��'�ў�|�!��QsY�so��a��hK��E�<y��R96|´$T9�V�҄*�<����4S�:SgC�m������M��C䉺9�<ъG*�2-�dI)�J�=@��c�H��	�o���q��Z��9y��ƃq�v��d0�IK��3�X���qh�k�: �R�D{��9O���c(K6en�%��C(��0"ON�Te��NP�U�#��S � �"O�Y�mI1ł4���d��p��B34��9#m�3��p䁂7���)&D��$ �
5��#��&�Ҝ-�"<	ٴ�h��D�=�t�ɅBH�v�Zd�%�-M2Q��F���þD��2%��i�L��B�֥�y���%X����B�ΰh�LK�b���y�@��U#4��6M_�Jt�=�6��y򮈁4�~l��-�ul��a�,Q��y	�z�*���g�Z ��@��yR&�j��p���	*`tde0�k���yr��8�*�.#G;���c�!�yb�i��ؖA��F�`��#�rў"~Γ0���4�V�%��xi��\��n�v������Ձ`M*�s��s� |{�m���y��
�QD���a�39������y"�Jm	�威�R?��pA朱�y�Ð5򸛣�%	Y�b6DY��y2�Q���aY-$qI���y��ÙHh�!2�	��~�Z��T��y"��"Di~	�cE���.�i�4�x��'�Y�eKi	�D���B�(����	�'T�(G��]����D^�	�'�"��E�Y%$�#��+���'y�����@<8�,P6c��RQXQ�'ў"~j��Ӿ9�]��h�M�l��H�E��hO�'�TC��{����&Z�H2z ���Z�9���3�����S�2Q��T�� �"Ֆ���cјv�9����}0V�\��LhW�A�ȴ7k5$����J6�xP��4~�B1CB�8���D���D1���S $\H���7:��y�IF�'��?�F*��8�цD�K�*�Ѥ�"}b�O���?%�%�Kx�*�5�P{�J������x�\[#f��Y��⫁ X~C�IZ�r�bC�x	�X�lT&]�2B�I�6��I������WlR� �B�ɻ&��w�ӷxt�X�4��"B��Uږb�\v�,�Dw�C䉆(�]�v ��m��l�G�>1��C�)� ���4��d�H���b@�/���"O@�
�ލ�pL0��-d����"O��X�I��/kz
���8�[`"O�͑FL�*^��'!��I�n��"Oj�����4�č�m�2�&Yxu"O��c.U�K|���,����,8 "ON��u.�G4:���� X��"O��B ^zD$r��_���P"O��;5cš�N��%��?/�lmQ�"O�܉�BN�?��aYd�����]!�"O��*���'�������N�a�"OjMkw�\�d����g�'j�ri�A"Ox裶��S.���5%��y�PR�"Od͚C��K�6�d��P|���"O���4��+�\]!PMM�w ���0"O�͒�%�.&�y���,��%��"O�\�F.:Ϧ�z �֤m���2&"O"y@�ŉ%�8�@ȑ+w�,
�"O�؋5M���#Aٌmp��e"O0�h4![�<�D!AL�Y�-�s"O� c6�>I�� 5 ݱ+L�c�"O�DaD��?j����X
SL��G"O:X�ѽE�ά�d���O+�e�B"O��z� I�>�lx�4�+��C"O~p��ŋ YJm12�X��-Ct"O�}�GE�%�4aC����%�!"O� �#A�C�=�Q�ʛ*���p�"O�|�SCQ�M���"j�QàH�3"OI�E搑~0��F��&9��}��"OrAZ��*g�4��LI�r���t"O��v�҈}��������cVI�U�DJlHu��e��f�2����h�1O@!*F�\�z\JAs��Q�t��Q�"OB�Q'�K�:H	X��m)�t�'�y���HG�R�o	�l�b9Kj�y���cAZP��I˗eM�]J׆���yRI� Cz48s�o��n\بH����y2!".��+�"L�f����a��y¤%5�<I[w̮T:�c� ̳�y��ۻU��)3� ϴUNv��.ɉ�y� W'$��p90O\26�Aڐ*I1�y�Ja��F�����r�߼�y�)ӶI������2a؁���y����H�����*�|������y��*cE��b�F#��^6�yr��;�T1[P.
�x�Ȑ�ܜ�y��(l��x4��x�$�r�ȟ��y�0�jQ� �r�dˢ�(�y@85SFz᪂�h֮���E��y�ȁ-}��B��m�}�t�K��y�]<z�ɫ���ZD���dJI�ȓ+$Y0!��@�ڕ��2���ȓxf�����wB�3�_ lѪ��ȓHZ��-[��J���N|���_�R$��6-�r:��6���!��U�ĮRBh`0�M}�h$��ZK�����	�r��ghĽt������rS-45�\C�Y�]T��SȘ���$�< �#�83|��d�M��O	O:���@;`�ny��a�L��$�'H��uN���Ƶ��=E���%	�P7�H����) ���;���QA�{ ��QC�H,</����\���g^�d)�F�V���ȓ�� $ �x��D́x�����S�? ؍hk�7G��)�C�G)j\���"O6!���&����c3Tx{"O�dH�NV�4��D&�J�b��=y3"OuS����vꀫ%���HW"ON�rc��E��p��@�?��!1�"O�A�@���'�ZU��@�/Q�%k�"O`mم_�?��qb�,G����"Ob�+7k�� ���kV�xQ"O�8cD9tx0Ż�� �E�6"Oj�RS*R.�8��s��*=�ɒ�"O��4�I;"��i;��B�[�|�ZF"O�H��ɛ;����BTB	���6"O���kW
��<+C��.
Ș�b"O�m���yF� QS؉�(E��"Op����?y�z�YU�ѳ`FB��6"O�����&~����� ��,�#"O��τB�hm�S�I�A����"O��qL��BH:dm[�_)!A"O����U�0����A�=�h`�$"O�ۖ/R<{�H�1 �+rw��pP"O����
T�*<t�%ݎt$���"O�e��Ş6I�VE��.��ڝ��"O�P1�τ2O|̪�N ��`��"Ot�[�捤�L�v�]�B� ��"O��G���m`ÀC,|��p"OƉ�� �!��$Q�Ζ<MR��E"O�k`,.:���ŗxM���3"O-�6a۽^%�}l��RFi
�"O��D��/t�j����Ӳ`�����"O �1�B�<oj��R�ܷ�dኖ"O�hy�Ģ.�L�8r��L���"O����i
�K��3���1�ԹE"O�
f�#zyDN��	�R�;d"O T �D�9�`D9t�V9(�ʈZ&"O�}§�"936�S���;DD�R�"O��lű0�5yv��=4��!�"O|�S�gI@}m�7��5h5���"Ot�j��J2i��v�S�49�0�"OM�uLZ �hL�F!W�I�*1��TH<����S��y�T-��x�	��"}��P�>	��V�ڰ�(�(6<��\�bʙ@�<م(1Ql2X�cf+#�^˷�Cܓ�hO�O����#��;��d��N�e8`8I�'�����6W*|�f&j�
����0,O(����y�P�T�{�B���"O�8+dH�E.�6j"�HP�
�sH<���#I,$�Z`�ʥ} �}
%��\��\�>qc@H (+����ze�$�aO�B�<qd��U��a�����R�(��N�d��hO�O���:3��!��q��V9�	0�'L�5�T�߱a�v���F[
^i�X�'J��'&Z�G�`xh�]���8�'�=K�d�.7��\�2#EVoȸ��'���P�&��$�� %�D��	�'��S��ܿJ6TlkA�ɴ}� �	�'�$�*�iF&@����NY~x��' lp2-R�����F�Q�
��'ph�$�6��DxҀ��H���'�h�y��ە)^���b������'�0��S"ĩ�R��p�
-b}(�'V�%{u!)�U��A�&z�}��'����x�H���,<�~T��'$|(�w�R !��EZDl�4ś�'(bP̑�7�f�"��!r� ��� �pSU���v�l��vǋ&����!"OĠd`_�kVt͑�̐5,q2��"O�T����V�ڤɈo�"�
O(D Ȳ��x4 ǘG�������$�(S	�'�,�b�$.�^�0���&���D
�v���c傘���'A󢴀ѯ��(#� �I�P �ȓvf�����M8< ���6���'��`2�A�{9�1�'�ڼr�˗�c"�͉�ɑ�@-F����'��r!R�H�f��J��@7ȟKh*$ �A�%h4h�I�@�z\j��(�����1ɍD~���b��hӨ�k��py,���'�����a��Q�]$�ٜ#%��!����!bu�R@�2��y��[������l/�uR~�KǎLV��X� �ܥ%�rb���=w��b�ZeW>w���1�L��u�UR���OY�5���6"Jv���iv٧x��	S�/�O�]�`.�l�V�`�N�6W&(�A�'�n��/Տ�E��e3W���F�i�T� ��:�IK�#4�P�b��ͪ��%�A�{�L
�7P$ta�'cj���k�	q�M�5�򝐱FV:*�fW�6������iGRY�t�Lzy��ʮ� ٩���L��h,��H���	l
�H�����5r�ܢ`D��-���ڤ�,DX t����oK��B��,L���6L+�lK����F(Դ���;w�6Ea@LA�eʊ$R��*��'��s�G�\��-�d%�1�?��
7UV	x1�x�JPc\�;�8���@W�(� B����4�9fB�^������h"@�	c @Ÿ�Iڨx���vb��|*V�T��O�@�!w�YkOܵ�f"O�u���	�'� �B59 *H	�pP��Z��������:-L�M��Ot�����?���� J�85T��b�'�����k�8�6}����"Z�Y���A�-[���Cm�o��ą�Ɇn���@Mt\��+LtB��>���;� e9��Ǆ+���'S8��Hҭ�8�t���ÝAD�ȓn���X�HN(�h�#�T>��';�|b�H20���i=����ƈ�,W�Fd��V�MQ�"On`�%��Zb�����28n��r�FF�$ʵds���S�<��U~�j�	�+^1Nlq8q"�
>��K?w/��R��K��%"�љ1��y�b�!�xr@�'H��(��r�q3��ި�y��G�gT������i�l$��fI��y�[3jɑ��@3Y������y��ad��0,X'P:e���\2�yb�@���T�q>;\��� N���y�h�@H����AmG@�� �%�y��<Zz��ƪʻ?�z=�a��y�ԱJ#�!�k����3&D�
�yb/�E�@��l0O'�TSU��y�[m`��eQfE�E���y���fL HY�Dą^�2�����&�y�G�5N��"�`�^}r9���ۥ�y���ʮ5�@�R�V�F<K�䐱�y��X`J�k����ܘ03j��y���	��Ai"MX)d~	�BNU��y���,�����	*_���2���y��M=[�53����g��$+"�y�d[�z� <1C�cC����EO��yr�ނ{��4��H_#�r�χ1�y�
l�ܕY2H˗]���Έ$�y�雤V�r��㛥Q�LAxDk��yB�!"c��yW�@&>f|�x�j@��y߱iЌ���ӑ}�l�st��y2�?J*�=Pb"У'��Y�Hۢ��x���4RNi��-@N�1�dX�"�V]{ 
O�X��d�0_��r�=j��|9�'�v�s7hIG���)�V�&"ֵ�cţvM�ȓ�6%��S�@V�U:&*��O�J���*����O:��:��L����c��7�ؙ��'>�� �yްQ���J01�{��
�"����Ij̾�K��_DԊ��T'����C�ɵe�rECFL����R_��t"�Nֶg�!�� X�Rb�'*J�b�<���'�v�A��H̓$�LaK�M�1W��86�\�X�dt����r��E.y�)X�C��_��&�xK��Z�S�'<v���F'p�䁓u̐��ȓ!0JqS�Y�P��y�7L�i�<���t7|)�aJ$� �#�$D�^>�`�ȓ8�ƽ���9ڸUq��;��y��E�wil䬍a�-�0n���)J��R��N{͜<P�Ȋ|�݅ȓ{EV9�3�H�>p����UcЂ�ȓf�Zd�&:�`@�S@�@��$N(*��^�ļ`7��
��I�"�S��yB�A�h��`��6Sv�����ۭ�y"��-r����w�Q�Iݰ�� 
N�y2Ξ�`J��!��LO9D]�( �y�)['k(�y@w�T�`.Mj�h�&�y2jΐ��:B�P-yƁ�B�E�}��a����O�\�v�ڊ<S�	G�ȱTS�|�'"O�����>��1`e��PC���P"O���R�� �r'lR�KQ��B"O�	ʴ��^]ʀ��+ԛfMr��"Ot�J����o���A��=m�D"O�9hl��"6>`3�
�}�(K�"O0m��O�)�t|��W�YB�"O �����gi��c���;`��	5"O�e���6���k���6A����"O
�s"�M3NMu��Mp5N���"O��!�`�O��S6��>(賆"O�-@����l��
�?(�e��"O�EZ�J;e"rLyb%�OV�:"O��٠$@-��"%\��b"O
Q0�,�v�sC@+P"��u"OХЅg�YbN����-e���y�"O�D�ČV94B��6��;Fz�1�"O���sJץiHJ��ƍG9{�t]c�"O�P$�M3^��Q��з�y��"O��3e����T�@HÑ$�Ų"OH5YpD�%e`����R^�H+w"O��ѢZ�Upnm����:TVY2d"O�<2�bѼir
1)Xe��� qDj�<f��-F��n��>���^�<�a���W��e(��?��x���U�<�boQ�*���w+�=}�%�F��~�<��)��
��2r@\9Q��xǞ@�<�ת�'Xڨ!�Aѵ]�R���[x�<Y��R�!�V�Z�Z,`[���H|�<�E�ǮR��PQa#V�f��ܲv�V�<iB���}\��cݘ�e,�M�<��E[�ڱ�	nŪ����E�<�P"V���!���D,'����MD�<q�Ѿ9�CJү��}Z�k�A�<���H�֢�(U녫�p��p�P}�<��.�
.A$�BnK�A��e��t�<���+�(�2���1f'��1q+�t�<��4*�tI� ��䙹�Jr�<�����θ�gꜭy�t���	�k�<��ꍯI��hXD
_$5��<g��b�<��N'JD�!w����)�7\�<aį�ľ�� GJbʬ)�kT�<IGHC�)���K��b��MA5�UR�<���es����n�RwN����I�<�6�V`���ȗ�\ܘ��Ĥ�s�<��
�0:����o��D����#�B�<+�W�,H2P��uR������<� JeZ��X�srl@/Ŭxz1�"O��'N&Hm�\24N��$^�p�"O���s�;4�¼[ㄆ*c�����"O򉀷��,�>�ť˱�t(�R"OD3J^.��b�*D�"]8"O�@�A �x�TĄ�ڈ��"Ob�B`"W�uI|]�� ��2�6�ɶ"O���!V���%��鏢�p䓰"OFcG�B$.�
Œ�W�joިs�"O��CVȎ	@D>���3{����"O�� ���5K/���g� �[�"O�����*R �i 2`$mh��"O�G�Jg����5Z~У�"O�q�͟�z�$5j��*U�<��"O��p�J2:߂]�҈�;`IL�v"O��1�kɵ?+4��gՕP���"O�A2�oʕE� �"�٪^�A�"O��fnW7� �3m��󆽚D"OڑX��.p�m�Js��i��"O*l����x�R`FDL4� "O�t��.��-?�x`�$D�+3|���"Ox�Z��	\�1{䀆4A8|�"O0('�q�r�"_�K�˫�y҃ �p�rP���B�	���y%�"~,�r"% ��*��L5�y¢:v���6��0W,��y�'�TMX	�mˉ{_�%��1�y�I3@ꟶ��T:��D��y�i��
9I �׸e���Bk�2�y��E73��(k���:�<����+�y�	
��04Ӌ��
UR�1
R��yB�t��u��憷
�b� 5�_;�y�$��S�I���>xA�A*C��y2�P�qj�#�eڂM��^��yB����%z�bZ�G6l@�aK*�y�NT�?$����m�a�ئeB>�y򍙱T$H=��	��5*`&M��yR�_�e�>�HBj�4,�c%Ō��y�T$=�%�pm��N-@!��)�y��)<	���G6zJ�j0�9�y
ÊD�08C
ށ[4�T���$�yr!BW�x�J#�D�U}����^��y��K�+R�	����.=]�̫A(ӛ�yr��
�4yk���'�f� 2�S��y���,�������r�̅��yb�����ą�E�0�[S��y2��oְ��s��0!@ҫ�7�y�I�>����+c�|��E�y�_!�a���+�f���V��y�T�A�&%���@h`ȿ�yR������h�/�r�`NG�y��Ǝk�P@9�l@}G�i1���yR�6S+ ��WO3qV0�s��y��Ѝ[�xe���Ϛ0�besc����y2���+��薨�(k"%���	�y�a��F� ��ᨄ�&���!�4�yb��CX�D����5>���$l��y��ݴb�.]��Ө
�&�`wh��yrݎR'F�ѫ�&]��E��y�!ۨ$ �%x���x�8�!(�?�yBh&BZ�=��c�tz�A�yr�Z"���w(��R���:�$���y� �T=b�CT��U1��Q��Ժ�yrfM�<h��Dq̕��#ց�y
� ���N�[�di�@��)A�`��"O���ܢuŲ�3��ڶs܂ؠE"O�I��iZ�%F�����=� *�"O�|R㈉1���p%�خw��Ih�"O�aE��!;
��&"�(~Ӣ-��"Ot�*�N@�b4��fB�.��E"ODzA��$�0� ֥#��,s"OJ�˦��M����������s�!�1q��9&.ݽN��U�&C�?6�!��-7��=�s�'V�q���c3!��C]Բ���a�1�ت�ȻTH!��ڭ[�� ��H�e=0XudJ�I?!�d��o�ȹŎ��XHvؙ�DI�}/!��'9�J	��K�4�l(s���,!�DD�f
�����ψ8����ƍ. !�$6iX�0I�S�9g�J�#��}.!���� ����CTi��W��!�$ӗJ��8C!�/\�N�P%����!�\6g�ι�[?.5ԭ�� N.lx!�䐢`�h`�$-H�p������/�!򤋌 ��A��(�l�.ԎL!�d2u>�P�d�&  �mL�R�!�ֱT6,�L?w+x��Ċ�h!��)�
�Rr�<��"��G�n�!��`�rرd�,T�l�S'�h�!��,V��-�eݭ) ��鐽�!�d̡M��!J��B��@k�O3~!��ʃF7����kL�B�0@*�gA4Lj!���L�>����${���@�P!��ף>�R�
% ̨|�����HN�-G!�d��r�|H�
^H�a3����k!��	)N\�-`4 �c��L�V�ثi�!�C5"�E���s�\q��n�U�!�D�T^D�����<-���a�
Hd!�ğ�%�t)5��Q˶�dd� re!�dض'R<l׉�k�ְF���
!�G;�n��c�[8�8�d��)!�"�>� v䂥H�ĸ�Q�!��Z��`���Y�t��y��ƅA�!�d(yʅ9��߅c�0ꂭ�>�!�D=
YJ�@V,L�M��b�C�c�!�D�|������4/t��%�t!�d�6\w���& U�I�%"P�NS!�D��be���Q�Ĺ_wN�P/J0!�����`)5��e�'�B�e!�n��)�!E*�#�)�W
!�@�p��F�~�"c�\<"�!�d�n�Y��낖gŌ�:���z�!�N6T�@�g"�� ��<�ք�/8�!�$Z Fl�㴡�-����e�A�!�DF<rY̐�����x1Za��7�!��n��h{�͈L��d ŕma!�d��	�-i2Ǘz��x2�	>U!���4���&�2QZY�'O��!��E�v0Ƙ�a#	bXl�G�^�e�!�dƜ?�Hl)3�,�v���ӳ4%!��\{��AGki���O+�l:�"O0�U��0 �|�&՚?n�2�"O�HiA����fy���a�x)�"O�
� �U���X�
	3�X �"O0Tb�?��|����;a�6  "OZ��+J�'���VL~��d�"O�Ku��py$H�ЌH86�8E0�"O�Qt͙�L�4ɘ����Mp
��w"O� �A���������q�yc"O�E2`d	�y����Xrve�f"Or�+�:~�����g�2p���"O4�H���T&RԸ�%�>fȈ "On:D�����j�N�Z �"OHU)�쌕 �^�R�P0D�h�D"O���7.�-j��[��3 �z�!�"O��H�e�:\���V#Y
Z�v<�#"O�a��d�X���:�����"O<8ƂԼ6�(Īq�M�:�Ip0"O:%TI7�j��c�{�j��"OX����J'`%�g��*�r2�"O� ����g���p6OܨSc���a"O��p��9*��F�1E	�҆"O�y��X�YՈ�˃��5�eҶ"O4ux�Ȃ%�2TjT!؞1% 	"O��:�*+��A#. f���"O^	"T�<[��7`+	* �h�"Oj��ՐV5����)[ �C"O��ifƻ?�\�P�	�.pQ"O�P�3�My�����䘒p����!"O�s�>M��VI+R�脪!"O��C�-ڭ�z\�DBˏ}5���"O�k���12��`�ުpO�]�"OB��A�P2�:퀑��"�dXA"O,����U�-��rB�L�y�(�bA"O�L�F �&6�-��1���"OH8WB+�\��b�HV�x�)s"O������#`�� FKX�$L&�I�"Oĸ
�.ֿ=��k���K�f,A"Of}ha��h$�`�1�ٷf����"O��z�,Vp���� �#��=�a"Ol�	��O(_��C% =��,ȱ"O��x�M=(�2fc��=�P�"O���V�ښl6�(b� .#��H��"O�re�^�5��tad
U[u"O2 �3.��(}8��-冩A�"Oީ��[-A���1�q:ٳ�"OX8A$kD�+�M�v��Cy.��DNDw2)kUCC�Z܋Q��o�@$�@y�,�Q��-1�51V(t������n����'���|:Q��v?&� gߢ|<�t��c����mDȽ�%�R�!��PB�͙7p�$�Ў�uӶE������,<�W	�.���B����'���i�Ş�^a��!�[�`Y���D�Rh�'���6��m�;�=ٔ��-��p�'�(1�E��j�	�"�'
Zr�R�L�L���<!0���i^)l����1�vd��q"$^�#<�T�+�Z�!h�'P�����м1&@ĠR�Dl��<%>���!��k�4�SDM��-��}ob�I�;Q�b?aYiY��D1���Z2��P��>Q4�1�S�O���!V
,�]#�$b1�D#۴=���uy�̨�?���CK�S>%��@�>+X	��� �`�Er�'YV��醖I��q0�׼ �T�+u.۬"5�OH�Î���nN�P�������R�b!��T���L�<�~�u�L'A�t̉�(�,Z�]c�Hc}�Cd��b��A����� �%,��P�Z���۴���Ҍ��ݺc��1R�D�&)�*�V��2M�51gJ�`���:�g~�%�1O4ڶ�S�b��y��'^��HO �=�O�B���u��P2�m�0D��]j�O��p�S�O|�g�J�<��Fm�2$BQF�<�4�'�4��v��xG`�#L��?d`�`eCB�MKR���hO�>=���^�xwB�'-�B"�dx�K(_
�#<	���D�$�ٕt��aU��=f$,�,�'2�7�l��|nڶYͬ��� 4v �@�/N�蕩Lo�<� ���n�&��KE	,R��"Oqd�X��:Eڰ�\?z��"OZA�d���2�p	$HZ�yfI�!"O��u�_<$W~���Q=1;W"O��
�ɝ��j�����<a "O|x�p�ه6���D�i.�(�"OJe�6��e����E���Kο�y�G]%h f@�"�>�`������ybNE. ��S�E���@1�ACW��yҎ��MI����%}��8�R�Ӣ�y�NE��d�A�x�`=��,ޙ�y�/��&������n�>8ᄤŕ�yRBX�<G�@c6^�mg�i�U#ѽ�y"�48ÜT�+m������'�y"��=LT\�)Q
]�h���.@0�y���9]��BM����1�~0(�'����4�ǔ.|�0`�J\�`
�'Y��gW	p��9���R�Ř��	�'�@M����r��ݑqG�M�	�'oLI�����=
�ɞj���p�'L�!\�@�J�b�P'+�2���'���u푡��-�B�%��Ua
�'��5��J�~����C�%d,X�	�'�^Ű�n��g�Ɯ��fS�))$$��'��TB�痕vTXaA��&8*�'?�Q)�B�	��H����6���'���M}2�ek�KJ�@ϰ���'b�Iʳ*�(SHأ �5�����'�l�aFyl����8{�@b�'Q��&�r~�h���*nB�
�'�J�kB�	�!Ŗ�: ?�hm3	�'Tl��Õ�bV1j`E�
�	�'>����z(F�8��y"ґ�':�|I�G[�2 �j��]��'�� ��"3*ԂD��7P��!�'�HA��֘"N�(K��Y뺀P
�'m�E�q�6����%ů:c��	�'Kjh��e�o>pщ_�>�)	�'Xh����~�D����+����'xb��s.JA\��$��|�����'�Ьҗ$���U�/@�ro�h�
�'Z��V��&�vLqT��A�z�;�'�~H��,�6��%36����'��T���3 ���e�݁��M��'�t�JT�"g��� ���y�ف�'�2��y������iF�}��'B������I!�躧�
a�ޥ��'|1�䉢�^ +�c�8%:��C�'��0Љެg�zQ��*�$�0���'@5���ژ͖��	fD��
�'��Tx�?nHH1,�&'!�)�'�Uq �s��|9�B2!� b�'7�dZ�Fɫi'��IdG�G�P�'\�Y�@Ƈ���C���&!XH��'��l �d]%��0X
�5��0	�',
5Vf�H㬨��ݶ]&=*
�'�6t۷��j����N��с	�'b����ן_D��P��u��!�l�<��In�*y�Ɵ�4�4(É_l�<�RdӯB�P��H6lQ,}ؐ�L�<�C`ج�$�E��@Jn��� �J�<)���
��eK��d	��Ԡ�o�<A(�Sd�ћ��,��!3'E�i�<qթ�t���j	6Bc�ðml!�� D��`(�t9T�P>
�X�5"O�]��џ��=z�ϕ����s"O8���@�M�6���.2:���"OB �F�Lg=S�J��O��1S"O��TY�V��3��6n��E �"OH0��!��w���P�����:\"5"O��z�
\�#�
pB��4޶� �"O^h3�!ԾI&�[1�R�ho��8e"O^�٦	�^Ĕ0sނV�9�F"O�5K��Hxؘ9x$�Y�P��8p"O*���"��%�	���+A�0 Ѵ"Op�B4j[2t2���-�!�ĩ�"O��s���3k�l�""�_4*�"��"O�����:
�P�d�)# f)�5"O�ِP�M7)�T��B�H�$�hT"O�cѯCn ��ҋƒQ�@\s�"O����/dg� �a��V��2�"O�؈�l*ҬI����P\��6"O i�3���9[^e`��?9�d�#"O� r�N�5ss�Q�J�=-FJ�"OJ}����A�eH ��!\��"O$��g
��ETJ)Q��	�& A�$"O2��F�H<#�
Pi�!�*-��"O0���N�x�$Ke���b��PQu"OR )1eI�84v!����v�ڼ��"O��	�;̜D��-�q�D� �"Oxu�n�p�p�F�$p!"O�Ѹ����y�`D���F�8��"O2` 4���O���:�1�0J�"O$�f�ʇz˴9���ꨡ:&"O6���F'-�`�YԬȰ��H4"O�dK�B9(f-Y`+�)�ι "O�yz���`��%R)�RCR q��B�I�/�ա�%L�"UyPϑ0G��B�=N��2��H���|0�~b�B�	@���S�j�,}
ČC1��E�B�	�9f�@�'�� 7^�#��Q�>�B�I Qh��x��!<�x0�D�A��C�	�#P9��P��:�1����}1�C�	�r�2���O�*�TMJg�^�l��C�I�9L��2
�3�McG
b�TB�	�<��a��W�\�)a�"�:�.B�ɜT�@��f��b���&���B�ɅZ����3t���DE�.�B�I:�4�PA��H�$�Xk٧@XB�I6Jx	��!ƾ
*b5��nK�kW�B��+k�ݳD��*S�i���ƀ-�B�I�l��7���VpR��7ǎB��CU���\=Ja<��gj� K�TB䉨U�v�8����
V��1prC�	"n�8*��sA�T�q�ƢjjC�ɾR*��S��GJ���PB�. B��$M�u�ǃU<4`�ɵ�A0�C�ɱ#�9���ðy�+��C䉺a�
��u샅2�+uh$��C�I�0� %�W�b�OQ�@�zC�I<�J=H�*�(+K�P�QN :��C�	�a!&yyuP�_�Zx��#��%	`C�	�+��%RD��;(��웢�Z�<�B��By��q-S'{� 2F'�Bj1D���عpU��1�_2��dA#D�`{�LS�D� ��W-��D�ч!D��rb�΃pr,�oۉWݒ�r�?D��昞L7R !����!�&9���<D�� z�huC�.h�l���D�_���c�"O��+��A�Q~�8P�X�/� �yp"O(ъ��U�q�n]�"K�$p�s"O��S$��+0�Q2P�ˎ,È&"O�=�B�U- ��X��	�~����5"O����.\��,1��ш\-Αv"O�Y�c�1G�\"Va�0�$�R�"O��C��'-*4�A��Z�%te`�"O�	c雏`��仃�	)oZr ��"O��V-[�-F����E�+Z�-"O�y���U���:�iΚ%o\��R"O&�!o�u�p���h��8��"O��#���t��Bf����Q�"O��$Ght��H�"]�"E��"On��P%!X�*�	��b�b4bf"O���*Z
�b�ևL�|� �!"O�U�E�W�9��5ԦW+x�$u�"Od���ۛj%��a�S06~x���"OX}bF��0��Y1Bѕ/��!I�"O�,�Q�b*�I�l���8y�2��V�<aU#��qHn�Q�@� �"�[�Qy�<�Κ�O��=h�j��y��@�dt�<AF��S7,�)�Q�L)�X�Yw�<���G'b���N&o6���^�<�𤈚�D붌K�^�a $/�d�<���C�(^����ߙq�1��WJ�<��M�;G�¥sP���.2�Б�ȓ;��@[���28RD�3�j@�a6Ą�7�Px�e"\�˂��-Xo���ȓ|H!��9Pʠcb��-�Xy��Z�4QK'�M�U�4�	��ݪv�,���G@f H��
Y�Z�!�ʚ6��4������+�O60� @ґ7 �P�ȓ;�l�I�dT�J�T	he�҉*��L���V3e&�%
~,����L�$Vh��.-<�Zs잃c�L��'�YA�ȓ(��.�=	\���t�ӷ�؇�f|�B�e_�1b,|	��S;Gv	��nr��ʣFӳ;e4Q!�(G	x.���0���: Ƃ�tuZq �o�9��(�ȓ$�p �W@V�T˕�'���ȓ Y&p�pM�/M��4��čS���4��E ��C�s����@F�0�F��N*eH�P&W�n� t-	�B�4�ȓG�ę� CK�G�P�KB�T��L�ȓ���i��B��4 ��al����"m��+0+թas����#�"�e��}���Z�zQkb�b�\�ȓ[�1��9:8�ۄfQ�
�ԩ��HZh� "�y8�,��]7�Մȓ}|,�9���/Bՠ ��f��{1�%�ȓ<�j�2-j�ƀ���@��ȓ=�މ�6Ǝ� ��L�j�t���ȓ ��@��Q
�l�q�*X;f�4��_�TU� ���e�]	��5����|�<l֦��CuB\�Kg�4#��AT�<�v����p�o��8�rMáGR�<QW�ڶg%����7�R��*IQ�<iU�M�#�t�7Β��j�"6 \b�<�e�T:�3�#0Q��i�i�W�<a'�O6����dC� *y�Â*T�\qD�D��s`��z�r��!D�h�d��-��HK��G>�X|�$�=D��Zt�GK��j	#Q����9D�� ph5	�%�qz�#����E[�"OL�T�>�����"̃}0�d"OR��C�8g�ڭ؅�Y�����"O��{��أ#��XqJW�кP"Oa��   ��,!r"O�9b�6%� ��b�Ӵ�\��a"Oްh1���F^D2�k�t_<��@"O� ��t�G$Z���S7@�wn���"O"�h$�Sz�R���M� ����"O�P��i�=v��"��*K�� &"O\��KI2���v
'�pѩ`"O��R���;'2��_�-�䌓"O��cPe1�F,��\�N��)C"Of!0�.-�A���.F�>��e"O
�"��^�����!�j-�5"O�� �c�O��� �эU5%��"OΡ�V���<�JL�~@��Q"OpP���ŴN������O?]�"O�ydc�D����@T�5"`h�W"O��)���
�� F� 8&Y�"OX �.C�~<��Xc����p�U"O��$H
�T��)��B��t�2x� "O$���$dk,U����U��b� D�̘G�\["�!���.?i�/*D���F�H.a5M�gJ�����=D����)F�o%r� �c�0������<D�p+��=Wƨm`�덄yx(h�l'D��!�#e(�	���3z � vb+D��j2ퟃ%̚H@�J�\�L�A>D���HѺ���r�	�U����$>D��H���QѦ	�#\D���!�<D�L����06��)��d�L��%:D��s�I��jz��	�͙�i��z�'*D��cg�A�%��8h��Se4D�T�f`& >�7e�t�^ �7�0D���S�VK�tQ$��#j`|�2�2D�$!" �[UBM!��'&�H�"�g0D������&~�,�����'+Qd0�H/D�����N3L�D���_7�j��U�+D��"AF%p����F
�^�}@�K7D��S�#=�n��IHV���C6D�41d�ޅ$�Vmf�j� 1�rN4T�T���ٞ���«բ>��ՊB"O��c�Ij44��*KB���t"O���/I�g�^�0�/��u�4���"O� ̉-Y���E���i��"O�ӷk�8�&8BVfR8 �z<�"O��qc�)愤XD�Ν.�H1+�"O�K�Ƙ;?B�pऌi��I$"O�A����)�غ��C7tD��W"O��A���Q2������>��q"O��)��+AuH�3R��L� �;�"O��2��ȩ!��0���$����"O4��
W���z���T�l�bU"Oh��ME:?�©�V�7�P�@"O�P�^+V�6��ԁ،ZN�2'"O�i9��8������JN �"OP=�ԏ
�H������	WGR!�&"O�qJ��ѱV���Z���6fN@k�'�>���O��!�ĸ.y7F��A�<9�j�i��Tb��
j�@(�&��z�<�R���:���a?,�h;��RB�<��O�UBN�H�C�u�p��J�i�<9�o�FE<u���EWV@����~�<i�̛�Fax9���ͼl
Q(���O�<��O�c[����W51pٻ��u�<ia
\����".��V��}3u��\�<�ć�/��@s//R�DC��Y�<	�;�V)��֡(�A����`�<yf��2*��Ћ��2p���y$�F�< ݝJ��̋�
�`������L�<� ����	�2mlH`�M�$��CD"OR#�o����І�;�E�'"O�pQ�9.V��+G�~Df�{�"O>Hꑤ��dj�`"��D@���"Oĉ��$�;NaK&�5Ĕ=k�"O����d�md�l����#����E"O����鞳!�l����>!�n��2"O|
��%`��6��Yk�"ON`{ċڄ�M#��T'(f,u"O��&�͗$��Eb �. ,	rB"O�<�f�U�%^��@	�)(� �"O�	R�LϠ0�;V
W�l ���"O�᠆fN�L7�E�E�9��@���'��O�M�@�� �Pq��	G)r�$�Z�|�	~�S�OB�]�@�`U�����+N^4��'�
`(a��%�Ly�E@�@��';���f��@��yt��#Gp����<<O�遨��~s�Ġue�!0;2�R"Ot-ScO��v	���Vd��H2@!Ԙ��D��>yc���y-��0" �`���`��Etz���$t��Oൈ���1w�,�@"��=��1@"a8�H2��D��{W0I�A�J)h��U'*o�''0"=�~",
<@�|�V�ͦ?ްX�kLA�=���b>A��
��P��Ҫ.���=�T�IN�X�P�!��\ D�N2Xu�c�D�
ӓ|V�[�͚�p��I�֕��ʌy�Jz�O��>�2���cL�P� �Ĭl�-k��@�>AqK�W��塴�̪J�䁋1`�&��M��O?��@4RqP�EN��:��7^�y"�)���M�2ݓ�b�*o�&�1g�.��B�I�{��!� �A�P��E��B듔hO�i5�ɐ���`�P:pj�d�6-n��9��R�^��Œ��\>�$L��N4D����d՘|y��[�ڪ ��T�0<O�#<�p��?^��t�Y�P��K+Z��Z8�Di�L�i�Z<aע�p���z�/��1�S�'L��aE,2_�j���8'�E{����F-gN�)�i�7���gm��O���
�U/D�2c#������]�<q�!XPB�(Ȳ�W�g�L�j�/�Z?9M��A�O�>��s��$>h�i�f�"�8�	,D��J1%IO�zP�ǆ 켁0Gk*D���Wo�& �.q)t�ĳT�H�j)D��S��O�Љ�D�Y8�1�D?�S�c�p8��^�<H�J!!��a�ȓPMJ!��J÷6d���D��f2�<�ߓ�<yQ�jS�\=
�Mʬ?d��	C�^�	���͹C��HRq���XO6]ʥ�6)8�IE�@�U����?�D�O������g�N��e˗�t��In����?Yv��8}�����2'��� �ɟ����<!�~�zX��B8s�ĈD�P"H�!��IP�'1�x�݂KO�qb���&e^���'
�e�H"Q=��R&T�X���{R���D{ZwZ(����)4�ш��D2��	��HO����
ˋ1�D�)�R�A�'AQ����A�?j��pGf�5Q�L��j0�n�'2�O:�!'�]�n���dƝ
�@�'�.�;e�F<��j�	��*O>�����|�$�>�c�!s�R X$��*afRI`0��o�<WDI8m��]x6%�%C_^�#�Ii�Ħ<���T>)s3芔i����e�9;c�t��$.�OL���'F�BU��/L�zl�&"O�yZ��8e���"!��%��Y�"O� N��!�M��Lt�Cę�D�$�*A"O�H3��<3�\��$��C"O�	����{�0xv��-~Ly�p"Of�Ң"�N<lZ�o�#gF��"Op�)� 4E�\�"b��0.�����'#�����F0�k��{q�,@��F�!�dAU�@�
 _Yc��aQ�Q��'�ў�>})॓�>Ox����,n�0L��2?ib�E��hO1�yq֨Q-7��u"��������'���G��8�-۱A�`�y5'��#�B�	���9 &�
GQ��� �R��ru��&D���ףL<�`�� ,LP}!d.D��{p���|����ID?@]�tU�*�$?�S�o%��Z�H7#�&]X&���9���ȓ}]��i�o������ ��$� �I�'���=!��TF���AI� T��@�_rܓA�<�����2��ѩsJ0�[W�[����I����Ұ�
A��Qh��жQ��$C��(�O��=�'T3�( $
�����JĶx b
��y�/Z�m{���<n���C�F����0>��,Ӹf��k���%-�<�K#/�e����j#�������%�5q�}22p�1b<�S��y�M��,Hd.Z!)1�hö�����<-�O��S���=7��t�M/oL�'"O�@�e
�'m7��镈0q_�kdo�L�Ix~��	J,SI,�0J�
�-X3)��/�$��'�`Ia��ZG� "C(?q����$JT8��Y��w󮍓��T�8=Ƙ��	�m�<��G�X_��ɇ�E�o�2l�ĨJ�m��:��aJsZ�Fs!�$-]�%��E��Ur ����Ae�p��Ճ �l���p?1�D�v�h�WcՊB�p��\
��	W�LF�t�� |��sTBS
#b: Goݬ�0=1�^$W��H6�ۊ2�D��CI��O0�=�OخqcaE=:�<���g�|�r�y��)�8������`��,Ƀ&�$ut�C�I�d�@��Z^�\z�� ��C�I�o�4���V�yN�Ӑ���dڮB�	5;O�}Z������F?-�P��wvT���`�|h%kјB��q	�'��$����])�K��4��a�{�lU��O�O���gF]Y<�	[e�ӭ-��	s�'E��pW�?�D��4��6{�Xxp�'�a�۸^| ,��g<ob �'�<���үR������Jv�r���'TP+NVbi��j��p�<	H�'c�0�`��7��aql�D��'�hda�V�4򸈀'MM&��]��'t�2GH�E!|ɧL;eX���'c �Y`�/t<h7�� �d��K�|E{��D�D�b@X�@�'fi����,�=�y�`�	f����u�U�\<�8���y��6�J��gV�*�4�Y��xB��)UJղ%+K�B���[�Y��dC�	� �f�y�[d:tܐ ×>�B䉮F4�Z�$ǟld!���V;1?B��  �j����=&$Y�dO� �C�	�|r29���t�D�bkGR�C�I�O|p0c�OLn4Y�-ė_��C�Ɉ&�
�m��/ς�(�K�71.C�	9X A�F�Q=Xh�i��E��C�I�s��� ���\@1UI�0Y%C䉓(���I��oq��ʷ��L6C䉴 -�aQ�A	+!���S0`ͧ5�B�)� E	�(��6�(��J�u�Ԩ�"O4E 6���t�����[��Bg"O��;d�:x�6�'qA�<�c"OF�PBo�1~�1І�T���M#�"O(��2&�<Q�ػ�m��I�<�0�"O�m)tŔ�'c���5��c�^�1�"O���V�X
N��cS,u�`9�"O.r&�P|�B�d���>�b�"O��4	��EvX��a� �Q��"O
��5�Ú'-J��׍Y!��9��"O<�i�jɸ���I�+V)x�Ii�"O|�Q�GP!v�|����I���9�C8D�@[#-:�J��V��̕2��+D����Ǒ:o�-qs��=.ڼ�Zנ)D��FN^���p
D�NȢ���!D��r�̴B�T�pjm��� =D�<Ze��-#�H�s֊Qf|�y��:D��xG�HhP*����.J+§%D�d�Y�V�Eqe���[Z����8D����2;(~� ��Р�o�!�(�����O� F�*�3QH��!���Uj�`��+�Jܔ�*Dw�!�S�J�����57�މ���a�!�d�$#���	wb�[���qBE��~�!��'VvJ\�r"�&��ˁ!l.!�䖐!�������P���C.B�YC!�݃~�δzӇ��
���[捁`b!�W�ru��`((3�8�1,ҹ"�!�Q�����{f"�0���/m�!�D�9W$m�@��,�� #/�}�!�U��X*3��#O�4�rmH#�!��(3���#�3x��Qq�+Ǫ9�!��0� pfW�gV����D�!Z�!�D���)�ID i=H���	�-i�!�$��.u.�I�cZ�6@�����;�!����x%BrKLk4
�ED;!!�Dbz�0*� =4~9��#B5`�!���|�xQ4.�V'�e��A�!�
>Ĕ%.�"l�f���b�r}!��$%Y ���͆�vy�)0�Pm!�֖&LȽ� ��Wr
��� ��>�!�d(&����:�́�T�L�A�!�dȞ3n8���l�8H�h�eT�/�!�䛃 H��Wa�:p�T�%��P�!��;7AP�G�<�$iв��SG!�D\>��6kG�!q@82��e:!���75t�Q�	:"\\a��!!�$	�
�`h����Z��mh��	�C!򄋼2�B| "�S/MllypEW�_!�Č.	ʷ,�FR\��W�zP!�$%p64�cԃs��U��D\(!��E�O��m�q,�r.��H.�!��E�x�v��ŭQ97aΜ�e`�+\!�dþ_�:`_pA��A��C�!򤐱�(��A�t\i7���!��|�d��a#H�8�Ĭ���,�!�%%��Q%%���A���!�D��A� au�MyHB Z��D)!�d�\'�<[��4]��0�6�84!�Ǯ�.t!��+CN�����/a�!�D܂*����3��MXVY�'	T ?�!�d�h�	���J�Tx`�T�Py�!�dJ<vz��2mG�P(�`�E4a�!�$܁v"ػGn���3� ߖ4�!�� t��a4A�̉��K��K"O�I��n�X�\Y	NK /�6�#"O~�:��" 3��HG�/��P��"O�a�艾?kRh�.8�bt+f"OXt�����a�R�s"Ф_���!"OVq� K����3f��n�f�`�"OB�Ba� ��y�$�y���("Od�2EG�jh��z�@�	�<�c"O�Q�GŐ@ 8 Pׅ֡ qx�$"O��)t��(��ms$A
�WШ�2�"O�(�$�˛�Xu!4F��l��\�*OjH��ʞ:�X�!"�U� l�	�'��K� �/�n�� �7I
1
�'�a0�B���d|��HF�X�
�'<��PB�_��8"�$Z�N�6u�
�'��̓rO�N:�����E�ī	�'�$�!�*��xc���v.
8tx*	�'�ab�ƾ\�d��c�'5��	�'2	r ��\$h饀]% <D�ϓ�O��R�ŝvlLATl"(O�I�w�|bj�u؞��$��� �Ⱐ�j�+J�fh��C#D�X"���1�ʴS��U
4�T|;2�!D�����5��-���R�Wo�cv ?,O��<9�Ӷ`�B����T<[��x�v	w�<)��ڮg�Xh�7D��7ry���t�<��'�l�$ः!�����t�<��h��`H��F��/"J鐑�r�<$h�,M���⣛ �>x�Ć�m�'�?aX�/�i���;g��G]f��`#3D��I��UB:=��b��f�H��0D�����_�S�&q��%Z�"R��p�F2D��
�gڄC>40�X�5T艀��o�`%�(秈�@ �bT�b38��aK�?P8�"O�-��wǂ"z�ur�oM��l�e�����&�^q�n�6J�:D�)��y��)�Z,��;�# � �u��s�\��Oh��%�N>���hǇA-Q��H��"O`��ǁ'N�\P�"�L�R"O�P�Q9��1��N�5ߺ�@�d�>B��?a��Ѡ	Z�K�x�hB�Lp�X���,�.�Z��C:U\���9��������w%�2�^-ISl�3�
��������#�,���B�":\p`v��Z��O2��0Fʜ|��8@�B�$
ĀZ3�I����4
W�$b�l��AS��Y(�"O�hp��ڼ{]�i��C+k�~i)f�|�)�S�Xo^<�#��@g@8��q�ZB�	�`�C	����h��� �vC�ɴ[2�qK�$��x�KZ�V#=Y�'�ўq�J��v7
��	Hn���f�4D��@�%l
"0K熼I�<���!2��{؞��٠S��w@Y�,Pl�y�O:�O&�^���̳M�2h����Rg�5;޴�x�M�bH2� �W�,1���䓄hO�O=���*K��Ђ�D(g�&�O��y�-�:����j��k�xze@��yHܪ6����!�-]D�j��K��7�O�#��H6��uzr��v�8��7"OaZjӃ�6�q��֣����"O��ӓh�F/p�	A�L���|��"O@v!��yG.��%�5Z���j�"O`�jI>���A���"-����1�	YX�0(��M�$�Xy�7�@(B��Y���1��`�'��	�f�dURk��V��������vؚB�)� ڵ���ށ,*���lT& <�Ɣ|�x��i�b�O,�H��"�W�*�k�J4D����R#�@I�͓# ����O0�IF؞|�c��XM�h�G�PH�.-D��q������@�2��_��=*+8D���DˈG�
���A�#d�U�u�!D��*���.Pj)�M�=6z0 �%�3D�4�a�4N B)�΁�o��=�u@2D��@%�Z[� �+�H��>�TZuG<�O��v�2�B`��	�I"��ʣ_p`��) �u�듞pV� fh�ad�ԇ�Z��Ur�R]e؃��V�k�\��=��^Z�!W�S�?�����i=`D}"��9�TU1���
d�ĉ'��	s؟�L�-2^|1��ۛn,h ��-D�8�H��TizD @e�=M�2�0aK*D��+s���֥����%�L�\���6�0?��R�z�،�&��k�^y�<��Oʒ9�X����_:^���@^~�<Qp�K#6�dH�A�$?�!R��d�'�ax�N���] F̊^�nlr(���y(F6�RŀRGI�P&�rѭŪ�~�M(�S�O3:��'mH!Kz�I�.������'���J���*z����CݙZ~^��H<�v�'�PA�6Ś�ل�I�L�^d�	�-���Z�z��Y��L@�6ՠ�( �hOh��$F~L��O�*EL��(/!�$�%B0��KO�p|��̷q!�d͊z��5۳ƽN�p�Я�t�Hm�l����Bc�7����V�؋z\����T��y�b*{����O�����vnH���dJ���>���˕S`t\`� ��a����4�Ixx��'?�� ���LDhB$��l�:���'G\	���_jm@2$]s���'�x���k�f�$���B��\y�y�
�'b���&Z�M�pb֚X��'L�'K�)��������v�T\0'K� G؄��nUA�<���4I�dY� C5q�
�1n�X�<9SnRE� ���9DAv-gF�Q�<Q�gB?U~uhp'��V�]r���g�<�bȈ�*��ZQ��-z�B�DF�e�'{�;O��>��.վGu{�(&C1�;T(0��<9���?/��3r�C�9����Z_�'/a���U%���	���"W��S���y"��+x/|�!FHmyt���$�>!�'���W�'��(	�Njk�����.:�e�
�'#�Ժ��R��Ny
�i�4 �dl�*O�����Av4�&�^�nz�9a1���T!�߫}F(� ��U ?��%���R!�䌠G�Ψ�"�D�ʌ{�Z�oK!��G=EY&}�!�	?_�6L2��[%�B�I*�Y7H3)`98f�_�D�(�?��I�9t��P{t�F�h !aŎ)!�D��z;�I��.\�}�vP��@�8?�!�ą�0�����ᝩ��t�(@-�!�F0%9m��L4'wJw!FK���;�OIi�n]3L�� ��fJ-��պ�"O��Uf�=D����+L����'<�N�"{X���;L��Xau!O$uU��D{ʟ"E����?E�p���_�(U)��'�0و.����GܤK�"���mV�<i���tD4hp�FGX ݹ��Q�<9���$x�����/���E�C䉐9���J�+L�ZQ�U+�
j����S�? H@�WMż:��jAj��\�q"O�틆�YZ�'�B�v3v��"O�QA�J�>3��)�O��/:���"O�訂K�7�>�I&�s{^�"OtM�S"�6j�l�����:��	�"Otl�K�
���ā�{q�d"O�!�2�ۓ~^��A��ү#eЌk�"O���7�@8I!(���O+rT��G"O޵٣h A
�%�%�\�d�T@"r"OZa��֥&��91b��/�<��"O��K�d�m��與�T77�<�`"Op�:�a��#�~	�'%�)ʜ)�"O�![�\�%w�Z�J�[.�s�"OF��eI0�0�B �4�3�"O�litD�4H�5����w>kV"O�	P�J��@�� lU����"O��FaH�{3D<+�#��K<x���"O����|flH�p�@��814"O��@��'p�@a"�R�(�TD�r"OĵJq.�PH"1ʷ�P�2UN��"O�r6�3>#x�br�J/7�|ӂ"O 1��˾`�<)�#�R3�r"OL�	,ѽN��BQ�W$*��u"O�`�����DJ�jW�΢]�X�"O(Q�Doןc(�H/Մ !�)f"O����
E��p�ՎN./����"O��i!���0�n<[��F ���8d"Oj%�C�H�#�!YH��N��iڶ"ORT
Rd��}P�$ǠL')
v"O�L�w䇚I�����`2��"O�0J�C�n62@R��g�s"O��R�h��q�1� 'φp�px�"O���Ȫ
RA�%�'^�\�c"O,�	F�B!`=j�1%�N.p2�Hx�"O*�#�j-���YPe\>|��K�'4x��"�a����E��N<x�'\jx�P��.%��A�!v�n	��'At����֓�*��a^��'���ǌrb@Q��f!\YRl��'�>i��h��7���鷆	�'�`��'� $�ƥ:ug� ڤhзujV���'V-8'd�yY���3:�8�C�'����6nޮ(����-m@-P�'��M����
��Q�@�F�Ep���$�&���f Rr���;!�
QA�4�p͂-$TXb�Œs�!�D�Z����AQh��Yb��!�[� �`X:5�͞Hr��KRh�M�!���AP����il���R&�!�:�`4k@��x7�����9r!�B�uT؜Q׋$.�Ec��g!�$G4G*r��4��E�Z0�!�M�o`�	�e�7Y�Qȁnr!�DK-E�LȂ�Kâ>��l��M7t!�IkAT�I��#O�>̚��_�]N!򤄨o��E���>��U JŬN2!��c3R��(O�B	{��J97L!��"�<4RH�]�N��[5!�ҏz�^(�VCO�?s����'�(�!�D�-��}BD�1�z�@P�<�!�X�H��y�]��>�� �X�,a!��ޱ^��X���*q�$I�� �R�!�DT�ld��s��'8`��Nz!��:���IPM�6;ph�� (�s\!��B���J��5c�!13�&S2!�� ,D*T(c�ٰ7�S�n[����"O(����� ç��V�4��"O ua�bq������1d����w"O
�b��H�3�|P��M�U��т�"O���x+bɒ�K2^�9�d"O��XBY�\Q ���;Ch�$"O,���tԵ2�]�T9���u"O`�	�H!ֱ��݉r
H	�'"O�4iأS�X���F_H�7"ONa8���tH��{Ҏ�^����"Ov�8��x.(]B��"%�y��"O�	���
/�Eӂ��'�+�"O&�ASC;Wqvl�'�@,��B"O�@a" E��`�xR@j"O����),�,�@P��!"O�ɻ��0vԉ�d�
�=�V�C�"O:��䓃A��0tW������"Op}�eO�8q
d��-շn�X� "O�]aࢋ�'<���Z���m�"O ��c�9�|��A����*�"O<0ՍA-n2�#N�B�$�@�"O�h���0hgu[�3|��*�"O����͙|r
�XB�W����"O���+]�Z����,NX^h`۵"O��",r�H��!� �Ms"O��)ߌ ��$��x�9�"Ot���$��)#��7�4"ON������0V�Ņ6K~bA"O�iQ�oC�U8��_3>�6�S"O�x�!ᄞT5��?���y�"O ��eHbb@���5U�ؘH�"O���dƃ�=K	� Ė)����e"O֥�a-�}��h��
.��8��"O��b�^vD�=ˇ��1M�~�[�"O�iPrI�:��px�K�{�-��"O$��#ƫXW��x�NH= nZQӡ�iRx�h5��?��'SQ���pL��]V`@�̌dL����'lO������A�Z��o��e1%G+f#�Q1���ԧ��'$�i�So�4:�&]���M�awN��y����csD�b[&9�����s�<�5���r�B�	�̓@&�C�I�QPty��ڃ{5RD�I@8)��(��Ŗ��5��O&�y!�'�s�Z�ͻΠ�1O�{���:݀MΘ��a,(�6��� �>٣%B�c�	��k5HYJ��X!�̕'O��D{b(T�
�xX� iӟP�P�b�9��<�@�S�T�D4���Z8}�DQ�P��zP�y�b�]T�M+�e����L���>�CQ�*L���c	Ǯ�֘ Pk�r�I�\=D�y���`�hZ �IW����@�$`F�����]Ӯ�:���	qvL]c�'�i�4��7N���rK�-m`��r��߅K�~\۴	����vf�(q������o�>a`� �ꏭ��:�a�FH<���� ��98�55�^M	KI n�q�h� 4xCJՕ��D	��hO��S'�)A��s�'V7�
���'��u���6�T"��P1�N�n-� ���x--M����T��b!�',�����6}�;0탦,�t-�N< HP��:m�'~y�H+�<i�/�Z4iR4F�L�𗏅�x_^E�V"OΜ���-K���ܦ0��у��M;8��l���?�Mݼy���>�ɽ�y�)޽�NP`����{�NS���x҂�2S�8(q��Պ
b�QS�[d.9;�)�#"N��PA����d��hO�u��G;q$���ł}��;��'�Tlz��K��	��s�&1A nUr^����̉y0��X����'�Ȕ�&�Q�q)P��cM ,]r�;�y�#� .Yx�$��oS�'AZ�ʧqj�A`�c�0\$�Gˍ����ȓ�* �ӊ�#JU��aB2��H�P�?���$�,���S�y��Y,�$��lM4$^�p�IR��y�G=,���)���f�X(�M���Y:?�B\�<���)� v�p���3Z��-�C�݊Qذd5"OB�
�현}�Q���1��ѱ�_���V2Jd��A�d��s��<,�E����<��]I�D.�8�;�?y�C䉒?�j�2�.+����d�Wl�<���T>]Q�л]���q��M�v�R�8gL8D�Ȑ��I%e�zC�H�9�|1�6D�A��.� Y�W��L��7D�d���Ь[�(�j���|F3D�t�D̙?g����
]G�����$D�Ⱥf���`��p8�iQ5\Q��jբ"D�P�'���3����΋F����6D�|ڵ�ʪX��-�Cg҇0-�Y�Č;D���B`��Dx����пf�@���;D�̰�L�
ey0����� g:D�x@��ђ9W�U�O�+[�(AV�9D����MX�1���@��vGx�o;D�8�T�ƌ|rn�@���(1�I��8D�X�GL br 4�S�J	�ᙂ� D�t{��)l�(����g!�t�Q(?D�x1&�"HU����T|�&��F3D��#��6kw�
��i[�	Q@B�	\�л'�+�xe)��:~�(B�)��Mt/^�\�������irpB�	�e&�����0F�r��!��C�ɴ��q�dۊ8�&�����xC�I&��ܙ���V��z#GOQ~C䉠l�pQ �L�	̽K$n�	yHBC�	!2��(Y2�N �����`�i��C�ɴ0�(Y��Ǎ39cL�x���j�|C��gp6�fb�O Pa�Cl�W%*C��+-����%�F�Yh�+K�~�C䉋!c\���нT�^TX�ӫ��C�IL&�x�ML� ��i�2OO#ϾC�	1���� ��&��+K�C��8|b� ��a��#Pq�3��nC�I���	�-%�81x4J�b�B�I1=p�(!擯R���ӔG~��C�I�t�x��fX��S�=<&�C䉱N��XgK�� 
0mP�-}�C�I�;�������+r� ���8�rB�ɚrI�Dڕ�
&�FE���O�U�NB�	�A�
���A�X���+7B�	�ى'�ŕ}&ȉ��A4!�B�I�L�f� ō�;Tyf,��K�R��C�I1_�&��ޙ]�\ȪÂ�k��B�I�Q����N<R',6f�*_�B�Pwl�
6*ʰZ�0C�YILhC�ɻi��ف���
	�5S�x�8C�I8;Zh��aNC)~;�t釃Q .C�I.R�:�!d��u��h�DN:*��B�	�2�`fD�zA�����͉<��B䉲.8H���%<||���ρ��B�I�s�x�k��4�8B�/Q4�6C��
4�̍��
ϣ=�h����)~C�I�Se��%�PDjWcG�>C�I�l�1cߣT�*����G�B��2�¥��b�0 p��[��CY\�C��<.|�2@���W]ƵZCi�6U�nC䉃2���`�{��5��N� bC䉧!XazQNB=Zs�ѐN�n�"C䉲_6D����"7���6 ̂=D,C�	�MG|�!F���k��H`�!AC��ؒ���$J7a+�4�ToI3y��B�)� �4���2�����ȣN��a�"OH����ƋRg ` S��L���{3"ON��b�k{ΒիFCH�T@("Oj���N=>8Fm�فM����"O�����L���v%ʎ?t�쀳"O�u+2��7.4Ы`C�.|�PJ�"Ob�)��ˆ1}ƈYФ�-f0�Z "OV���@�x���G��i�dX�"Op��DAӎs����"�
G
��p"O� ��.FG�t�07+�u?�h1�"Op�#�.�5>@M22J�f�8�xt*O�M�Ō̅9lx٨s.P�v����'�>m���F�h�~�z�b�y��Y
	�'Ml4C ���ry�x��u<���'�&Q��P�/���3�Nߐk���X�'!H�xW���/P��q�d��]��'P�����Y͸���HN�r���j�'�>e@aJ��b�Rq%N�"{-du�'y�٣`@�W1L��`��d>$�'�T�	�	���	h1�R�Bh�'�$1����XD����$~�`s�'����h�)� ��8^ѐ��'�l(s��Ѹ@��2�F�XJ�]r�'|�q�+`>,�x�-RR��4;�'Edy��D*-0L�S�C6'��s�'���݌cI���'K����j
�'	R}C2��-��S��� &z�pJ�'h��V�_: (�N���yb#�`.���Ai�Q��U��T�yb�׷]��	Sc����D9�����y�.�#C-�ԁuߦ[�͓w	��yr�Vw�hh;�.��l"(���<�yR �3ʨ�a�l��mP2Hr�����yb�V)^
�Xs����@V�D,>�B�I�{��8�ę�<x��Q�@���C�ɼGqڡQ��8VX�g�0��C䉘Z�.Si�']� eU,�+BC�I�Sں)�/i#*�zj�B��B��#l��q�'��1��lPG�#�nB��)aXP���1�v�7�� _�RB�ɑ@�n���h��H	��8׫��foB��i7h��g��k�Z�h�/ܥh6�B�I�&YP����+�l �Z�
'fB䉥`�`Ԋd�Q*.KD�K4LV@bB�#=��$��	 HnU��� a"B䉒��9�e�.u�@u�ql a |B�IJ;�����zjVuRՊA�:B�	�F�ݒ�S�q�M�1�Hv�B�	�tN �#�J��E��ˇ!{ C�I!v���p����H J�C�XKC�I�&EKr�;o{����/�C��$TT�
���N$����Q A��B�ɮ0D����� sJA���ss�B�	G����j�m�T�
��T:d�C�I�sG���L΁!��BŦլ��C�	=�LْD!97T9��MN�`w`C�	� ����]�
���7m1�B�I.vF��9`�N Ժ���㚵S��B�I���<*@�Y�H5�ta�ݟt8*B�ɑ�dq(�F@vz�s M��,TB�	�_,�	��A��IwL\;�ɗ lB�C�I��q��+�
U4�<��.si�C�({�ʈ�tf�,��H�SB�(�B�	3UezdE Rhl�{��@�B�)� *�*��F�8��i�1��R�4`"OZ�P��1Aƴ��iƇ^����"O\ �K> ��ӗb�І�j!"O1�#�P���i��ɨm;�e#�"O����J��J١g&[<5����"O0����%z~�� �D4-F��A"Od��$�J&�֭1���#l,ƅ��"O��j�_�U�����O�8hd"OV�{2�� N-"Ԩ,%��}��"O:,��'M��A�F��~�q�!"O��@�,��nݢ`��ǘ
^�#"O�Ī�Ƭx����U1[�&�A�"O
M�A� h�5c���~���Р"O`��U�ې4�TQ��ֲzG)h�"O�4���\�J��%�H6\3�"O��x�,W}'�M	��p8�a�"O���jA�.H�d��) ��p"O�(ç靍<jX{C+��c|!1#"On��� ��p+[6ꄜ+$"OD1S�����qh� .��ؙ*OP@�֪�<:n|�"��=(��'ަ���N�f���c _(�N���'��=2uE�d~�DgA�/%��@�'a�D�9Y��\C!�BO~��'X|�r��$�
 ؀#��EheB�'@L�HЋH||6�j�
�k�`��	�'�4�ɱoU�/��௛Z�Jd{	�'�Bi���Ԁ~)�\�pK�V� �j�'/��j��-ז���E�Jfū�'/L��  2`���j/8?�y@�'�eB�˞*/�=�E(i(Ě�'�:��#@V�^��EB���!��lq
�'�<� �#p?��3��Pސc�'k� X!�P�9�����I9��0��'�"�!$&M�O����C�I*�Y 
�'4�4�d*� AE����݌s*���	�'�Ա��U���(1B �;o�nxQ	�'�T�`��,u���a΄^��J�'[���[@�M�aL ��,��'�T���L�:y~���;��B	�'R���c/L����f�:�'G
HXbhW�����9�ԥk oZ.�y��(ՠ��F��uX ᘂ�y2ōe�d�S�A�9<�P�+�y�(>
N�"���<Sh�@�c��y"c�S�S��<W�t�iB��y�fB+w�����4!�8��G�yR��3C��\�s�ߞ�2�̿�y�n�2S�E�7�N9Yy��i�yr(��?�Ψ��%\��Yb�O;�y��98|,�K߀X���j����y"�9b��H̘�V�Lh։���y��"s��䋵�L&Cx��#���y"��@�����R=��-����y� R�TO�Qa+ݿ,D����R6�y�� ,���JP6���ҏ֔�y��ۻ~x�豯�%T�(��	 �y�aԚti�������E|�<Q�,��k�xaؾC^���f̛~�<y�h�J�����K�1�e�{�<!�D�"�0SR)���L�u��q�<Y�#s�����g��J�1X�fi�<�6oN�v^Z�i��Ah��C��m�<y�^*u�������P�$(ժ�S�<� �Т�d��>.ތ�Fɍ�v�N�Ad"O ���S�z	8�;5��x�(�Zg"O,h��m_����-Z�rb�h�"O�uS�"�Tu ��5��� ^H���"O�-��h
����)�2vF�1D"O�,B�'�1��%ѓ	K/I>̔(w"O���ǑYZ�cB؄DÄ"O�MYU�<	xH���cWR��"O*���-y� � f�ϠR6<PZ@"O���d�n�h!�X$H��E�"O�]��4ޡa�W$��522"OD; �р�ΘK2��4�3e)�y��E1ta���4jbC�	�%�(
!�Q�V#�]r�fR�X��8�SҲz�!�DY�j��$Z��Ɗ�u����L�!���e�pCY� � �!	ׇ/!�$�%ZŊ(�mBнR�)�"6!��Ȳ"�v�"��])+��$�3h��!�D�gܭ�Q��vc�����C�R�!��+Y2�����qc`o�=�!�dU�y�|Q+@oX�bu��sΆ��!���R��& ��V��0`.d���'6����фe���kv�J+��b�'$R���E4��1ZeI�� ���	�'�49��>W����.�� f�H�'�Q"�#��9K�mb��C�f�S�'��-��M����R�=h����'7�p·e��FȄ=Ӣo:p�.H3�'��ؠbZ"o���h7J�!W¡��'�<�&�=��HJW߫Kߎ���''�(k��\��p�sf�>jx �'�������)���Rn3�Ys�'%X��B�3J���VI��_x���'��1(��зi��d�E#)W
=�'�4��TH�I32��s��43����
�'�@�`�V�E�����0u�]9	�'�Qp�(I:g<X)�@/*��\�'��ؕFE/	vM�g �?d��'~�Q�J�B��U��I3�'���rV���A���# ���"O�\i�eg��}1�Z��@�"O�X�]䢀jGF���\�"O�\js ��j=�H2���a��9"O�8 ��%-
��@����9��"Oα����p�>����8��I�"O\X��`W�l���z�Eט*^���"O<��aƲY�ҐZVJH�:���"OF=*B͖%2�,�����/�0 ��"O�S� �'pT���l��o�Z���"O~�,�.�LϝR�h���W�?!��(y�@鈈�P�����+%!�d��a����Eo�B�@� �_>!�DD�e�ER���YgH)�r�͇L�!�D�;%ޘ��ኁ8'��pX!K�4�!��ѿ�ްx�iF� �+�k4�!�Q' ��@`Lα)l�8�V
]#�!�$��f:JPr��'xjȣ4F��!��n��M)��fc��R!d��m��X� �*ͣ6ʚ�|��$1��^�y�Hϩ�����ebb���\$�yb��9�A�VP�X�d�#���ybž�`��/څ_cT�c0� ��y�C[(P�&��f��0J��7�y.��#|@{�L�T���(V �y
� �A{���Ʈu�0f��egR��"OF�"�±7%~5I0��0EVH��"OJ-{ ���� C	�=�����"Oz�"W�]�uU�,HBb�<[���"O�Ya͋�I�Yh�� ?pX���g"O+��4 h���#�Xqg&�v�<ѕC�(s*Py�v�ޤ`�����d�<)�ǖ�"�͒�.�&P7��ɧ��M�<��)F�X�~��ML"BZ�|�eH�<���8w�]E�����R�nTJ�<�7"�ii��q��ٵ	��9bΜA�<�Ae9����S���i�NB�<�3H��2��2�m*�|c��x�<�lY Sm���T��5$�M�
�y�<���ԽzcX�1d�8a
��d�m�<"gCr�*p2�"����cXn�<iҦޣd1�Y�UCƈbDX�']o�<)�j���|�a����(���^�<9��LT���c�K�kh�3��s�<a��ģi��\
��țu[F��e�D�<�KP����"p�^�d�
����n�<Q��_9����Y�C�D}y3�Q�<A!�E�>�.�kf#�R�� �M�<Q#���m����D۫z3L}[�Q�<I�Knw������{�����@SL�<�%2T���W�(�B�H�<�r�N�1�y#0���D�c�EK�<	$K 9Y��iD�B�:3��Kl�<�2�ʲA&@�����A��X��j�<�J
6j͒��э	�,��@Tm�<1`�+[ϦmrD�V�&��q���q�<��J�:%�ܡ��F���e� �n�<�QC�2$<���<ał���]o�<Y1�Ӕ>�ɂ��
�hlH��!�[^�<�P#�?R���Q#K<$�� 03c�F�<AgGU�4�6�چᄺ=&(haM�G�<���י=��tc�Ab�8��FX@�<��B�=�*}��e"G�nեB�<yԍ�<wTs�M�O�~��O	}�<Y#�&8��I��M�x�2ԡ��p�<� �کF:$��V'!N�A�c�G�<�Q��2<�`��Gk��I�!�k�<)�Y8�� �b�.���'�y�<�Ǐ�>E�*Bh��vYԪTN�<�MF�/z��'n��(|�P�C�Fw�<ه�_���y� O2W{
��W��U�<1��-�B��NA,�XÂ9T�P�C�ƟQ�F�a�T�,���N&D��8�����$�h�6����%D�D;Չش=��ӅQ+�n�*��&D�h�a)�
jk�C2'΀ ���e���l#�O�>~88Ԡ_�,����$ړ]*�B\�VZ<�ۓȝ�)�Z]l Yj�wW����|
���� n:�v�)R�R� ]�#�~AyT�YA}��ר�?���'�➒�Rq�S�>ZT@��M�-k�b��>�`�'[���?Z7"�@>�xc`�˝~�¼(D��<��!�S�Oڌh�R&�Y�ĩ��a�4q�Bq�-d@�<E����
P�4���k��&+>i��<�çb�Ҡ��"	P��z��	�N&�d�?I��)��.��=�n�X��D$�F�����9ژ'�ўb>mz���8������JPx@zs�4?	���ӈU�f��EM�*�� ���ŕ-��o����J�#Z�1��'�#4*��ː�$�IZ?�OQ>q"p�E+� ��i�0@&r�hi����~R�O�?��+R���<)��}���3e��>�'rqO�>� ��+�Y%u�"劤�T�"�� ��@F{��ɍ�7�|���^;�"�q�HY�~���7�S�O�<U�S�US�*��C=��#t�)�`��`�ŵ������"KqV!��ቪ�HO�3w��@Ö:݊�r���~���O��z���I۫r�
Q��)ߏ"&�UA�r��'|>Q��|�T�@�.@� ���12/������)�'O 2%Elϖm���A���G�� o&ĸ'�� ���,}�2E�F��s�*���1�Z��z��?a��\>Q��P9�.�1;�DyG��n����'� �	�MK����b�?��';Bݑ�N��j "�Rӏ�0$������I�6����7m<E�T�	���т��ę7��C�I	R�hafc ����3��'IbB�	�~"�q�G���:��֪�DB�I2l�A�#��`Ծ���/�bB�ɍ?�~p���̯f �!�sGޝX�6B�	I7�$:V(�3�$B�j��z�B��)h�XC�cG�Q��P"F�Z2r�B�I#O^�h,ւt�� �-�.��C�	�r�x�w�
p.r����$F��C��r���T&��V�"h	g:R�C䉉l�z ���W� ,QDeL�.�C䉀P
rq�f� ���0∆Ѕ$D�\[�ó|Uk��� 'l|���1D�Љv&DGW��"BmP��tE0D�4�6`�'Y2h!:�D[xZAE1D�����A2f>uY6��21R`�.4D�[d��s�|�"�jH1M�����2D����e��X�@����W�"D�x��F33�E�%�Þ�l #�';D��@".gbu��@�$�
9
'5D��ѣ�mF�ي$l�)h�܈��n-D��vf�8:F8�p�	�rʰz�.D��� (�G�&��H՜Q ��9B�)D�Ty�H��Y���QE� ԰��G�+D�X��e��Y��_�<ظ<�K6D���ϵt� � ^�[^R�kb�2D��@Ģa쎥��N��<rpbg�1D��@���(GH�+P���M/D��� ,T�Utb��G�*N�X�I-D�`��!X+���b�֓X0����)D�$�$��R	,Ma'��/(�a�G�-D�x[dܝu�X<�SC��i���hA�?D�pA#Ð�W�ȉA�(N=d`R(�0G:D� )�G#;�X�ժˏ�`��.$D��&���a2��C�JϽ\3$��т!D�P!E�WK��C��t�Ҥ���#D��;�ɔ<P %)� L�f���'D�`F��v��y@"� ;�� �m;D�|st�YX�Nu��(�T�x��B6D��:�1/&�Q��u�L�� (D��k�cψP�̀j���|V���C�#D���-��y��e;P%EM+�UF�"D���d�]#oFXh�#*'� %�%D�l�!������a\��r-8'*&D��B���#�\tk�Jݼn'BAA$D��ӫڟm7���I��s�1�ш"D��S%<|� �x�`�X�2���"D���r)�)%��%:�G�B�yjЉ>D�d�c"*����w�|��AI��=D���g�./}�93�#X/L�|ᩔ�<D� f.��-ob�8R��MxY��-D�h�7a��A�����H�Z�rd�-D�xxT-�d����cMV5�*D�� �Hk��Ȳ1.����P/��T�0"O���@ =wЁ:��>�B�q"O
,;aEűrZm�0f��s=�� "OI��4��Fd�$(9�YS"O�px��\�'��X[#�S�#:�Z"O��eR�C-4���2��b`"O* H���:y}بWǌ�N�^q�1"O���
��" �Q���X�~�G"O�����X�0�W;]��=�D"OZ<	���f-�E��!Yd��˒"O�(�$�11���i�/�g�&y��"OT�膣G�4��D
�M'M��t
S"O��� 䃿2�A�+X{d�0p�"Oؼ��H� �8p�j%H� s"O��K�"@Pp +U�Dԥ!d"Oz@�'gT>���уP��x0K�"O�*wi	�4#�t�vE�/=�e`�"ON�:rgA�c,��C4�=#34��"O�p{��P֮�#�m
T1�Xbp"OH%�1�؞*���.J�Xqg"O~h�߂<]dI�Q�c�H�!"ODʠ�Y�7q&�G$Sd��9�"O� 9vpV�(�`�9��3"O��
2(]�6�2�Td-DE��"OP�3VC�9D��,��Y�T-��� "OX9�o�>���g�L�z J �1"O&U�bL^�2�\) u�D	`��Q�F"O��I��
"4Q'�_�6�@���"O�Uc��^~R�)�Ȟ�<�p��"O�E�5�P�%Q"i�IӔ<ܽТ"O���e�^�>�J P�؍U�(�"OMa��Ӈ(�F5���\ 0x�"O��@�'Qx@A!�D�<@p[�"ONukU�C)S
reyt���G0�]˂"O�P�Uj��!<�b��%���#�"O>�A`�ĞSzXX�l�o�|�"O�1`qCD�������~j�YB�"OЕ
$�lQ�����h��+�"O^��	�,~���O�ur6p�f"O<����k�4T�ԍ�����@�"O1X��8@�1�*�n�c"O��(��?�����b�$$�"O�P�u)M�	A��¡��l���"O^�JR���oܺ���rBa1�"O�@���P�Ipь�\�tC�"Ot\�D݂��!�q�Ax� �	�"O��r�P	k[��)��#��y�"O���ح:�n�GG��8��*O4�c#��>�<���H����'ʑ�#(A�`-R\x�M��\�
�'�P@#1@�-|T�P2vL׫5
�đ	�'/ ��0���j��;�O�,'f�P��'�*�/4�y@ ,�J	C����y��> [;Ng>�!�ЗE+�x�'WxL�1V��<��L��P���'j�����T�8"$Q#׈�#D�<���'T����S�A�h�B�J�9d)��{�'�vKǍՕ<��5
Y6Y�нK�'�f\`0޵��c��W�P�	��'�,��Q	Cu��!)P��Ne=x�'���
� {-�8�d֞2�L��'���E$Ɉ	��eكb��� Ѫ�'�x`Qɖ"X�yY�MNx@@��'�D��u+�$OP�mj2C�o�t���� �3�i *9�\���%��q��"O�ɻD�ڟy�>��`Cݖ,w��H�"Ol�6�˔\�^���GH�0ul�`�"OBpk�*��+r���	O7n P�"O]�7%۟���BDǇ�*e�i
7"O@����%D%�A�HN<eg�4�v"O  ��X���h�ϗyV�s"Ov�:�LR���P�j�ؤx4"Ofa���ѡ~�6�3_3:�H�d"O��R�����*�JҚ��a��"O%��e�]�u�@*�3�Ɯ3"O��A�*Ӄ"���O_�L{�T×"O.��E��UG��r�OÎ}{Dd"O��;�e��r�Y���X�w"$[4"OP��NC"D\���'Z� �$"O:=C`��Uu�� C5:�B�b�"O6j�,D9B��x# ���ݠ"O� i��ASJ]�.Ԉ[���;7"ONt�cBǴ/�(k�ʱ}��<#Q"O�}
Wč(0H	��&�V���"O�t�ܘu���r�]�|ih�g;D�J�¸��E�LO�욑�=D�pZ��2	# K�
��Z܉K�
=D�d�v�]+Zϸ��4	u������ D��aW��-i�}yNĝ>���#�� D��A��̅Ph�|�T� ����h5+=D�\�q���i�p@��Ɲ��Z(	w;D������U�Zt�5�'A]N�sf�9D����G_�n�,k�+�[!F�`��*D�x{EkC�X���aC�N8���rP�&D�Tp&�G�,զ0�怌�'����S/*D�C0��-D<��9w-˗;4f�"e�<D��0u	�?D=(��d(M�]�{��%D��J��H�-2ޑ�b� 
�.(0�#D�<p1�
�@}6Հ�,�ڽ���,D�LjPI�`�2�d��)�e*"�,D�x�7���=
X��Q�&��3С8D��Ye�T)�n���eN�)��R��6D���A<i εh �V=H���1 D����U�:@k&g	 &N�XZcL<D����6R��Y�
$� ��A9D���"Ɲ��h�F��^5���� -D�2�)[�%Ǯ}�7��݈� �'D�Ђ,�b̹�e+B7G��M�&D�8�W�dj:@oM2m��py�i"D�H��#Ӥ���v��(Lj��V� D�Ìɲ �6�)u�3`bՐ�:D�PS�	_�_��M��d�^]�9D������&��x@��Pr,u�U�7D�P@ �B(76�ԙa�K��3�6D��jF�;;e��z6�Zs2�1i��"D���")L�n����LY�(���bq�?D��He�D�z��=v`Ý!e>;�A>D��#�D
]�\q�k��9";D��#1�ʳBW8e+�o�c�0,���=D�(a�ς�kO�BL�$^hkt�<D��J�R$$ր���(x��U�G�5D��k��b���0�cI+�M"ƭ2D�8�*ַ#dq�q�&"k`M)aN1D��AT�H2�|5ph��m�T�4D����&W���e
1 O|�k��>D�P�q�[���s��.'�J$j��'D��Xb@�-�D�&��:B�0RA%D�X�V�znTY �%G�f�%×n!D�� ������a��M�6������3�"O��Ս23退@�HA��=�!"OPB2&apb�����%�pD2"OFh�ԩZ*Rоi�`Ǐ]�����"O�X[�*�� ٪,��A��XxY�"OVqf/��`�Ft��� ���I�"O��5��l�� ��8�4�e"O0��cj�V�%�։��~>�Qb"O��H�g�j8 ��/Xp��	�"O�I���xrpE��7s`40"O�P��ǜ%�>Y���-E@�Є"O^�Q�T�zi���#�5*��E"OZ�!�#�(4�q�֧}+(�ɀ"O䔃CK-$�H�Q���-'�H�t"O����"Q�@��)q�޸8�a��"Oʀb�#�E��R�����\5�D��$���-�(,�D�i��?a��"ش�Si�|Ȥ�2vൟ�ɚl2ZpB�Aة9�z���LH�[������P=�˧ke
x�D�����zp�($�(%�tP�� �4���K�/���p�d̟s}4 ReI��\؜<�ࠂI(�fHR�O ,���'f67M�s�r��7/\���cY=:�.ɑ�AL��'��'�'t�OȐ�F���<���ߪ$Z̫�'�7MJצ�&�h�֤�\��E�q���g�|��P8dE��':B�'D��$ķ�2�'�B���3 ��D�C�U'%�6��'m�+�YHCd�+!���Q	׊{�| A3X>�ӸnE,�����OpQ����2:�	֍W.HC�3W��,(��� b&��Y�x)��č�AJ�Q�0)	K���X�J�*<x�Br���w�Xd0��ֱ5;\��ְi���'l+�S��0�	ʦ�c�:64P��Ïc�t��e��?)����Ob�?�.�$�l�^!]6i(�A�<��?��i��7�)�$韢���>iԆߝ6��� ML(qprʟ�Ftf��1�F
��'�B�'��]�������C�4.d��I�B$��Q!��(恤t�!���^9s�b�D�¢<�F��+�ݸW�ޑ2dDCR��6ςq�r�Z�{�	���J����R�*ܪkde�f����i&m� rI��ʇ�7V
���i�ӟh��"���?����':4�2<En aw�( ׌m����O
��M+�S�''��H2���� h=�<+�� �j����d�'�7M�O8al��M�+�X<�4HĦ��I٦��0q�Q-W��PlңV夸`��?!sO��?����?A0 �n|H�Ȟ�d�npa�Ŀr����1IB�x$�d��<}_�IR�iHT�x��d]!�q0��B�K�f̊�/��LJ�����Ġk@$�;-���W��0z�����A#70  �I��q�e�O	l�1�~҅�x� s�'�2P����~��'�R���1k��8��(�(DE�	k� H��DΣ:���]y��i�N�r��p"AJ�*j�V=�&�C�i�'F ���`�>���O~ʧA��شE7Z���p� ���-B��X��'�B�w��]���N�dR��� �Vp�j���b_�\�c║u>����������0���_�6J�U�@�[� K��iT `�ٳV�F�(>�ؗc�8q��'S~��盖(���$(�S��TĐX� *� B+Z�d�H��`y��	:m5�t*1/��
�Õ�A	�y���'��7�Q��e$�@����q�L}�e�;`�Bd`� Q�W��1"��?i�Z�@ꖠ"�?	��?!��X��-��N�2E&�����%"��0�э��Z���RFړ
Q:]b�����N��.�����>��C��'Ѡ�"®V?��x��K+�tHP���&��1��B�~Ib� ����#�|	#"H:"B�R0*�n:z&TB2/��^Px��Q�Q�ƹ�۴be�	#�.�������'DkL�����r�L1~�8���R�sy�h�ē6��i٤��`!(�.�"�����?���i�,7m?�4����>1j^9I@,bc:P�.8 �l?���c��`  @�?�   H  `  �  )   o+  �6  �A  )J  �V  �`  9g  �m  �s  7z  y�  ��  ��  >�  |�  ��   �  D�  ��  ʸ  �  P�  ��  ��  ��  ��  ��  -�  p�  ��  _   E � %  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P�����hO?�ٳ�.J�j����XG@�ʂ�����5�O�k�`ܱ$ڀ�S6K���~���"ObL`�NӘx@�"iU�)��|ʒ�'
��+/�HM��휡*D�H1�Ͼ]x|C�	$To^�C2O
"����+8����� �tbX�Aԯ�'(Ԭ�� m��'����'\�_ͺ��I�$�Ry0BGP�m��K& �Ƹi��'��s�\i�sm�/,1�A���h�d$��o�o�������i�գ'�'v�4�yT&�'���U�����#��������c�f�<aP�'4�ΐ�A4@x�$�)(�Z��R�	�����l�@��2c���`���F�=	�y�gl��ʧ)��ջ7aҏ4�@�����)�&h�	$�HO?�S0/$o�񺖏�P��l�i�<����럜����fw �:VGNAtvl󤍿>��4��>�2M��-8����C^3����J��������s��l#&ǚ�tg����>�`��*O⤣�I\�,���u+��e����fmj�(�?Q��Ʌ�f���C�i#a���P�	�)�!��F9`��ʆl��h��0�7+Ԥ�!�۔l�<򢅄�j�&	ZQ�� q[���|Z�}
� H�+����M��8��l!c"O�5����2��ۆl+Fv�`�A]���Iy�80h��}��m����1Q(v��K؟�K�#�0euh0����$4��=�� (�IF�����ʌ6J؅���'D�w#�0pͼ�ɓ�Y)A��`�H���Z�<۷�R���0q	
�p�L!�!"D��2o�6u���hgO�9%QT��T�>D�lI�I?�$����/7lX��<D��j�&m{�@貍ŽP)T�䉥�����>�ɦ��(N�]p7LH�MR���D%�	����q�S7�$H��h�!B�C��?�
e���)�X8�"�@�	,�7-3�	�<E�ܴz��5�S 
(��'hE": lGzR�|r�'��P6�X�J�F��鹲�	*��ȓM>乻'�H�W�I��n\&.��I�	S�񟤤OX�	R�W��9A��(t.���A���C䉘%�2�@&`ɂN����'C�M�
�A����Ob�#���e��4�8Zs�d�a�'
�'=�����>�z������-�jh���:,O0Q�Îگh P�a��c;�SU�'�S��y*��~�2��(e��� �F�D�6�=E����p9ԩ�Kpv�㖜Fр��'����S�L����:6���A����0�7D�r!�ea�"+Q�z���A'��d"��1�)§a���b�n�@ŉ��P;$���In��w��|JP�L^F���b� ��<�J<����5}d��I8�}(�'ܨX�C�	�T�15�@�=&�i�gW�AS`C�I���
��4�j���`I0D&C�I� >x�6�Q#R�b\p�H�)_�C�IQdLr�"��-=����$S�Y)�C�	H�����U<�<h�Iˀ,&�C�ɰQ9�,��R�'G�4:���<t��C�H�W��_�A)���x�����'��>�	�Ru*!i��V�4`��L;<RB�ɒ/J4���L�H����e��-�R���O࣏}roZqw�y���F�<��q�
���;�O P�@��&p�bI��#�p�u��2�S�'U�h�b���b�8"���	�NA�?���~j�C�9:�p��6T$8KPԊ7J�}�<ٴ�S�7�@0��MU5'����ǯRp�<��Ίs\؉�7a��4�Ř"��o?�	��qC�L�8��{4&�-�����O���d@ӑ�N,�1;��*DE����<!�b<}[�f�I@�aܮV4&�)�)� èO��q��i�4v�\H�S�jy6�C�pQ�HG{*�]��FH�j����ޮ`��h�|��'5|"=�����u��ud�+d?�|b�%�=a�{2E\�8r�e��Z��2ꌟ�y2�6eH�a-H�\�`)������'oў���q��F��a����t�#j0�����&�y�$ ���1C�hQ�Q�
��=�P�)��8�6DW-q���i�q2�,���ɷ^�b���j}E0ŉЧφsD���	y���I^��[�/;�� �%̣t a~BL�>!� Y�pA�y����-0o�|�4�EF�<�LR�H[�諣&J3t����{�'m�?�*cL�"Bʡ1s����pEB��;D��Ri�y{�	0���̔�� L:O�=�!i�6�LsB�ּ<eD0�5��n�'�2����3D�0I2EM3�`�� �����nX��O�>�v@b��]����Y��#�(Vޟ G{��i�z�>� j�\�ꅻ�\=G��O���� �FA�w;�-	�^�A��|��V�d��ɇ:ܑaUb)^jv�U,�8ӨB�-9�н�R�]�d��Z���I'rB�"8Ӗ)")К��xơ�'̨B�I�>T�H�$:c���Ą�BG�#=!��T?Q"�K[�2����ȥ$M����>D�����,Q����%Ⱦ$�N��cJ ?q��i�����H��s��0�ZH�b�>D���Ѓ0iY0�A���6�(hJf�.D���2�ޝgWB�2%�u����M-D�pk+�$|v��`l�Q���2��+D�� d��0F�����A-AX́ے�6D�x6�E�0�F����87
���%�?D�0�:,rz�	���5���!D�p3��ؐG8jQrI	�X �Up  D��r�LA�'?��`�]Ɛ`q��c�@��I�|�!`C�T_�4�f��*"~�C�ɗF�\1rCZDإ"���()�C�I� �`r�얍�8��hՃ"MУ<1��T>x�#E��1�dO݇U�JH��:D��qu͘Wŀ�b���% �M��,D��1�Ao���M&}��x6�*D�t����NL�{!��
�q"2�&D����!�{�r����)d��9c�%D��J3��?�2l��mQ8J�\H� #D�$b���7tP��w��h6>D���o��{���2�np��=D���b [�QZ���~��[��%D����%�O���p�@��fՐ��(D��2�d\$z�XP�w�X+L��l �L'D�� �N4RF�r�Wbr��� &D�Њ��%(��*@JSG�\��a.D� �#� (���G� c\p���*D�Q��^2I������Q-�92ր;D����Vl��aO�&Ŋ@�SJ$D�<���Q�b+�� ϗ�6���"�.D�����Q�t1/X l�����-D�ۄ����H��	�q��M��(!D��0�@��"��0���	c�����?D��dC!mb�<8��@�"�tM�f�*D����I�n�H�7eݶ~Xl��T�)D�8�R���.pl��ׅGdQ��2D�|ж��b4M�0�����A#D��2���8:��Ȩ֪%/_ 	��)#D�̉"o�/���3��8r��k�6D�<D�:��(+�+	i������5D����e�
~$�18�OYB��PGG6D�h8�$p���H��h�$3D�hIb��?H���ʖf5l��m1Uc3D���v I�(;�<����3��yh�H.D���쎥 4@:!@�;�.8i�!)D�A!�p�Y�ТٵҲ� "-!�d�_�����MfM�|0�PW!�Dͮ
�<)��m�6��s�c�>�!�D�Q5�V�l�^4������!�����i� lE6�
����!�䖀pt-�4�R5')����ʀN!�d\��4ɚ'y� ���OL!��]�N���Z�DёE�8��E�`!򄊔M���XK�u��p@��E!��o:��3'� � ���i��ڣ3>!��ʚ0t��5�װq��%��Eک?!򤌡6ZЄ��i� >(8x5%U�g�!���XiV��S� ��ۧwq!�� �a Q��,�%���N�+��@�"OX�Ic�]�q,�M�@N9x�$`Hq"O@��$�6W��1����T�x}9v"O4�@�f� j1��B�@���97"ODe
��]�M
��R0(�4i��t�'cb�'���' b�'��'x��'nr��p�X2@�@m����/
B���'���'�"�'�r�'�R�'}��'�>e��մw$r��G�+|�p�٢�'(R�'P��'1B�'(��'�B�'SX�S�B�!�6�ڻ�lRF�'�R�'���'���'��'�R�'Ɋ�['k��=	H5#W�M�G<8T8S�'D��'�b�'m2�'d��'��'�B�P��˚!���h%��bP9z��'���'�b�'��'��'B�'����`E�^��+R�WWd�S��'�b�'�b�'w�'���'\B�'�:�E%�4AR�q��EB=zX:#�'y��'���'��'��'��'`UC���00 f�F�h!
��G�'���'�B�'p��'b�'���'=<	���)K�D	�� �wĄ�'u��'�'��'���'���'{:3bg@;UG�)�mX
y�꼒��'I��'���'���'q��'�r�'GJ���k��AȜt@�Ye�]{t�'�R�'��'0b�'�b�'o��'����b떈�<7��@��(%�'���'��'U��'m��d�P�d�O$�	S�?��A��ڊYJ̊��By�'*�)�3?	��iC��e�-o�>�:F�#{Є�2GZ���ę�I�?��<�5�i��m��Ώ;K�0�F��l߲��d{Ӫ�d�E��7�`�d�I4?N2�C�}��C��IĥL�GI(8��
]���<����1�'AU��R��SkiB6��!�<�Qŷik*DI�y2�	Yަ�ݠdtZ}	E)ۓ���2�ެr��A޴O���5O��S�'�=Z�4�y���FNp)G����8���ǵ�y��?u�́x�M�4�ў���+���U�T��5R+����Bc�D�'`�'�7�H�6�1O�80ҞB�`i�	�G9S�@/������ަ��ܴ�y�P���$Z;F��Qh`��g� Y*?���ܠ �t����ç�`)�_w���$�(�~��VI��5w�����*pʓ����O?�I��ӕ͘�R��	J�
J�J�ɻ�M3R��~~2�����2Kz��x��6Ocԅʓ8�.��>�M��itB��r�V��x �<��8��BϪ|�u+�iP�	���9��F{�O���p�O8v�k��ƽ!��$�2�A�`���oj���J���'��� H��SAJ4��2�@��r�
P}R�y��mZ�<J|B�'�?y�ק+ǘ�cg.��[�ty�#�6]y�0P�SN}���9�	�s����ў>9w���z!%Gq�Y��C\h��@���'��j���M�@A��<�$a�
{��7AĈ[2E����<���i��O�9O�imZ,�M{�jZ��5��6�(PwJE<
�!�����M��'��%���v����D៨�1-h��+UC�.S���˝%B���?9-Ob�S�O%��� X�p�
(S`G^�
���y�'b�n>?�B�i~�'���5 W<G�")g�ߪW>�L�@1Ot�����o�>��C� 6Mg����
fY`%�b�
q�je��b 3 P��_�-܎� W�F���X���I��x�{�����ˀg����W��
�Mk�B�X����F��� �	P&u:�a���N������V̦}��4�y���\�M��&l?��ñc�!�Vq@�	V3>]X$@=`�'$���ЭJ��� ��74{��Jz�J���Y��M����(�-��*àJX1�ڏ���+"��W�\Za�
u�@-�bLE�UfIQ�5  ��U���Zϒ`���?2�h������S9b){��&��H�1�M�P�1�ߏ'[�X9wb�;0��l�BV.��-����v裣��_4L����ԙF8��g�!��QDY0>�fy��9����ƴ0�� �=�>�-W<�Iw%?0_��@��U�к��H'`8"�"�6<:u�vg��mZ�Y@���Q��XRB��f3�p���̒y�'���'��'���'�"3��mt�5�a�9�E�?��'�2�'6��'|r�'��k��q�t�h��V��e�q�P�6Ҥ�'��[}��'���|�]���	�>qqnQ*��,b��)Rje����Q}�'��'g�?`ab1!M|J���7ux���O,�<����!E���'��'C�>{��c����Ν��v=���d(�]�@�dӐ���O6ʓc� О���'�����&B7ޭç-����|r�"f��H<-O��9R�~��F&h��<I£Ls�~����Ք'�T�6�h����Of��O���T��h����1�Y�P�i�
�nWyb@�O��.@���HZH�Q�%�!7H�dcv�i{����gcӌ���O�����a$�4�ɳGoT�"�M��0�nӉ8����4 ��Ex����O(������D����d�0���E�ܦM��ȟ��	�t��(�K<y��?��'�H1ED�?� 4zW�%�B,�}r��#��'���'�B��{� Rt�D��#G��"e4�6m�O�T�&�W������ȟ�
��z�IK堨��U�f��Ŭ��_�*�|�>X��?i��?���?y��?��$�<|Q�G	(��(�v^)?!�,�i�b�'���'�ꧬ���Ox � $���=Kɜ�*%�.U�������<���?����?����ɔ`�&�n�du<ة�ݫj��➒C�Rݴ�?)���?����?�+O����2w�iHtm�ŋA&O=P��V
it���OF��O��$�O4���-j�Υmʟ��I�[�:����� Q[ŧF�hw&�	�4�?Q���?)O���x����O��I	��\�Q��([rAb�Wq��6��OL�D�O^�$P�O&,m��H���T��:$O��S�_�PhQ��F5]b۴�?q,O��DH63��I�O���|nZ�c`��*� ٸW�R��>�$SQ�ia��'�h�ka���$�O �D����O>M����	j��{�eî{�����G}��'�8hKU�'�ɧ�T�~�q��2�(��sm����]� �w{��d�7��ʦ�������	�?��� �	�4 �)EgƮ��]j�D����G=�M˥�U,�?����4��������3�ċ7	rp�9۳K�8wj�mZڟ �����G�L=�MC��?y���?)�Ӻ�b�P &ndl�#��)Q�0�;׃CҦ&�|��)m��'�?q��?)�C.h�T)�)3����U�q+���')\��
f�"���O���Ot��O��'P��}nP�SN��0R���uxp�,����?���?Q��?9*�X����'X��	X0�A7	�ʼ���av`qnZ�����۟X�	(����<���N�@��d���g�F�A3'X;N���a��<Y.O���O��D�O��D��!�Vml�'#�ʌX�k��B�h��J���uA۴�?1��?���?Q)O��D���i�*B���P���3�F��7��/PkDYm�ן4�I�����x�	��n-q�4�?Y�+�DD��ǚ#j���W.!i�!#гiB�'��R�d��.���˟�c<�A���.h�ԡ
�g��xּlZ韄����H��	\f$�ܴ�?��?���x�h�yd&��Y�x��"c��i�DY"�i��T�H�I�]A��Sџl�I�\�s��41�,��
��FC�*�x�i�� eQJ�{�4^����������Ϝ�N���4;Vu��M��9��&S�$��%�S�P��`H�Z�����ߛM<�|nZ�b��ܴ�?����?I��Z��'�bG6�,C�DM��X��wO�6��.K��"|:��f��c�P5s�pC�cW�z����p�i�r�'m� �=Z��O��$�O����~7��9��!n(���98b��b"�!�Iʟ�	����Sd�(`ڂ�[SL�Ȭ�0����M;�������x"�'�|Zc�%c�� ��]�͗ 0vs�O��e��Oj���O�ʓz���AfJ�g0>H�Pm��E����ǟ ��'�2�' �'��ɷJ��� �B��$��%.�%zfh�[`�=���@��ݟ�'�4� a>�FS�#E��ڄiQ%X'j=�M�>	��?9H>*O��Z�Xk�,B"u��͑2�&|-x��fͿ>���?	����ĝ��u��@*5Q��K�����͖P�H8ߴ�?IK>y,O���$�D^���yCf�� B&P�c��V�'��\�p�������'�?��Z@Q3�� ��z�KG7@8{��x�P���p".�S�� �g��e�M�Z>)��Ĕ��Mk)O ��	�̦)����������'Č 8�)!��)T�G";@P�j۴��DE�
Y�b?�`�L�Ӧ
Nwe��Ypl���t����	ٟ����?];�}�F�=����"%��2vū��.�6�U�p_�"|���BG	�j؉C*���#�(E�>M�irb�'rb�Rn�zc���Ij?�3J�7��Y�D�4hxP�Δi�<����<���?	��5���c� >-�@�a�/��T� ���ixb�!2��c���	a�i�u	U��.
�����H^�	�n��$��>��̕N��?����?�-O��3�֫G�Pa�X8@^4�`C޺o����>��������f��m�GnjEi�0/�n��Z��|��?���?�*O`�Gk�|:_K��e����.X�9C��ʭ<�'0��'x�ILy�6��)U�d�$a���4N��V�W)�	؟��	��'��Y	� �i�g�l�T㖶h5J9Q&[5~0��o���\�	iyrU�`�7d%�'��P�F�T��+�:i��9	�4�?�����"tx &>��I�?�DK�� 
WHU�0��!U-G7�����v��'P/���A�*1��$��Ωm~y���"+�6͔Z���'�4n.?t��U���X2�J������=�'m����i��l�R��BD�^�ӇdU�,��6��\�p7M�O��D�O~�)�n�	֟�p�iY���DThöDT��J�(_<�MCF�M�����DāI���tmq��`#Ʃ^���amʟ��	ߟdҕE[����?����~2�T(_���	߾P�l�*DF�7��'�rq:�y��'���'�|�QGe��Q2E+�g���銀f{Ӡ��K�;j`A&�T����@&��X�G'�9���H?sv,��Q��7��q+dY�<9��?����dy!�
Үn�Τ*��7r�<��&D�K���&�l�I��%�h�'B���e2�J�0�e�;X�����ڭ��'�R�'ob\���հ���	�5Z��[���dxr�h�`����O�d"���<l�I}"ꈤS\�9�ǋR�<X3��F}y��',"�'��2kТ�;M|�t�Lz*,�@�3�:!sKĖ^D�f�'�'��;.xhc�� �qb�I� �l�H�O�T]�g�ip��'!�	�XC���O|���rc�F5M���A@,J�ꅊ���+%��'>�ɡ��#<�O�L�� ,�K `��v��/Эbߴ���Z�v�D�l�,����O��I�H~�[�[�����F�!l0�ܪ���M�/O:����)��7]��D�e̜9`O��Cpc U,�7-����o�Ɵ���˟t�0�ē�?��ji��O�=X�qx��a@@�ܴY��Ex��I�O�}�У�>A~"	�У���#�ߦ��	����{�:��K<����?A�'ߖ��ᯛV�@0Q���>K]� ��}b����'o"�'m�ƺM�~�i���<1 �����6��O�(���@�����IO�i��2O��D.ع���(�h|�#��>�QǙI��?	���?	,O��*&2��t)g�ۯ5�@H2i��7��]%����� '���'.�ěQ��)1*��7�<&��jr��2��'(��'�S�<�gA����(Q�?�z�Ru��dl�A��$�O��d?��<��Q}��;4��S`��y!Fr1&���M���?1��?��[?���,ʢ�M;���?�cg�
1r<��vg��l�ځP& ��M��&�'��'��	0u \c�xi�#Z�l����$LK��&}�o�"�d�O�˓#�艢&��$�'���!�0#�����W!{�~8p ��,O�O��U��Dx�����wM
� �ˇh�)tF @ �i��	W�v���4���ßh�S���N)V�l��5k
�(ebi��!Q����'���.,�O�x2��LX�st��/.P:y:��M[���(����'��'w���1�D�O,� Sh��>����#�Y�6�&OΦyaeX��|�<A����X`��D�@Y0s�V} ����i�2�'g��Y�06b���	E?1E�^�%I��+��nP�g�|�تT�<���?��{Qp��7[1;�R�y��T�<�6L2�i�"&�=O��d�O�Ok� "I�������!:�l$0��%7��iyr�'�Ҕ�dN6oOJ��a��8�P
v��d�>��v�4��O���4���O���ќ�꽸ע"n)�gn�b-F��E��O���?q��?A/O��#bY�|:��i8�M���@)J����$ �^}b�'g��|r�'f���yb�Dx�dm�dM�D�րˁ�]>j�ꓤ?i���?/Op(�`�	Z�S!Y��axq�P_� :�c�f�Ba�޴�?iH>���?񑏉��?�J��(ӀɩL������ؾED��&�x�6���O�˓!�4�)���4�'W�ԁ�4[��:�i��Z6�H C���T�<On���O���@�O6�O�Ӱ.�ʱ��F�2Ҕ�"	�&��7m�<q�@��${���~Z��������`+Q�,	��^">���J��h�n���O��Bp��O��O���\��؋o��H�`(��u���r�ijމ�Av�\��O������&�D��G^\j�m\P��	���&^�@�{�4?/��ϓ��S�O��]v��	�����|b�t9��K� �T6M�O<�$�O���DJ��؟��IM?Q��	,sh��t��a�����æ!%�������ħ�?���?a�^�-P���*[P���Z�z��'6	)E+�D�O���<���i(�3"ٺ0i���	o�)��X�PHWl�ӟT�'C�'BQ��Y�/ϾM�qE��t�е�$MM���J<Q��?�O>Y���?��B��2���3�AA4�Fq{Bт7l�y9����$�OR���OHʓ1�T8�6�p��BӹD(d��ʈ�a��`��[�8�	ϟL'�<�Iϟ�:�&̟|j�K'C�
ТQ&��-ڶ���D�O��d�OB�Lp��Q�����o�\��aB�[��U�$��R9�6��Ol�Op���O��&>O��'��c�fY�o�|�gG.t��qڴ�?����Ώ>0<%>��I�?�cr6K�l�0M��,���YA�ē�?����������S��A�(f�0hN�<�t�ʶ�K��M-O�$�P+����������e�'��H"�K�Hd" �C�A������4�?��[� ���S�'L�����;!w��r"����oԞbߴ�?���?��'<�'�R��&^V�+��H�.�F%�>X��6�V��;���矄Y��ĉ�����u
�,jw�=�M���?��'L��.O
�'�?��'M�A�0n E$�@W���l�% �}r�
ݸ'�0|;⤋0<yv<Rч���D���=,2�e0bY\���_x��$����8�I)�l`b�Gl��z�f����$�&Z)�l�j���$n�֑դ��9��ū�Ҭ0��BG��Oy2�;�\�,��c��.z��1ZT����(�j߶�4<sQh��t�� �$j��r!��;��,a�cL86=����ݧ�����j�/��S���1A74��#�V#�T��g��i`,��8��Ȅ �?��X���?a�O/��;C���s��a��J:�F!y�� �o�246�8[�C�>},�E~2%
<H�H!����0/S�T��i!�t�g
�,�(u �_�J@1BŻ{� ��q�'V1O.��q�'d�^��H1�ƫ~� ���F�q:���t�;�e������v�<eG�A�&��L�T�-�hO�	���Q@l��$n�x3��ʝI�x��AI���'����b�{����O�˧��!��S���j�.?�.i��I	? Ѹ���?qc��? F�pVk�P�S��W>� 8��#c�9>i��kgᐜ- �"��>i%H��5 ��F�^�gQ?U�U��"V��Y�CB'k����f4}���?����h�&��:*_*�q�F�g(���T�z5!�dБ-H����H����H�ax�e(�^+g�� +�\��X�(GR	�M#���?Q��@��#H2�?���?��Ӽ�ìM�2	�aI�D��Q�6t�&�j� /��AB�=@`�2�/�a�^�P�q��MG��cB��&B���&�GC>�ߴNn�Y���ި������~�,Ǽu��� +�V"�,���� -O8@�����W~�aZ��?ͧ�hO�P���Y+0��
w���7�>4hq"O�5(�H�	8n�""�wTXH$8Oh��_W����'4��(
�|r@�+%���j�
5���j��+Aj���	ğ �I�zXw<��'h�)\Z�ӡ.C��<���EN�R����ٴ=�����M�2K.�J��@x�'�d%��!�)��qRv�ũ��!!ċ�{{B�QQ���_;�
"��v��"?��5w`�,��)�2ʬT�1M�*G�<`�I)�Mp�i��[����J����R���,�"��l
ؤ�ȓq��,ݙ)�q��l(����<�"�i#�Y����,I���)�O<8���"(W���*R%�.ث���O���A�@�:�D�O��Ӷ%kwh�<��\�CF���5L��L�C����H���Po��83B-ʓ@0d"DK6�d��`�ݍ�MS��HL��Z�&�8/��D`-]��P�a'��E-��]���;j���'��	���� bL¸��# �J�P��c����tx��S����TD�#�G�X��hH�8��hO��C妍�`Ŗ%8�<1�a̼  ��0�?	.OPL��FCЦ�����O$�Yp��'��Y&��
����U��0S��'"/H�*@���B�8$�����O�`�����{��!�m��^�}�0jږ��	����bU皭=G� ��e�O+����$�69[�¥e�ԡJ�dz���Oz�m��M�����O��x��Ɍ-�R��tJ�Rk���y��'F�y�	�C�b�͎H�����\�0<� �ɝ|��JD/��l�41q�&�t�QA����ݟ���B�S?����ß��	ߟ�YYw^��z��vk���·�by�Y#tBתc,� T`׸�:T����b_1���O���#j��Uj�p4��y���b?�\:6@�GG�=����46�q�@H�O����-N�!�	J1m�-B�<���Aߦ}��4�?YQ�P!�?�}�'�BeM�#�* YG�Ccv�C��K�:|��A&u,x�q�+[���Ҕ$��y�Ɋ�HO��	�O������i	:kT�j����[�(X�%�V4\Z@����?��?!���d���O�S�l��ɐ��^0�|�ꅛ7���n�0� r%���<��'uf�c%˒�_9��[u��(�����.d�<�e#5Uh���5l C&�&h_���|R���cl:�kc	&R}(�)���0,�RQ�L�a"��/~~D��)�g0�@�N��0>�I>� ���j�Y1/W�A�aB�+�q�>蛖�|b�Ґe`�7��O����"̦A1�FQ=r&��s��.^���d�O,X����O��$b>a8�A�lNl2WLԦ~�������- 5�x��l�
e"4|�'��c�dMsA��=8�Q��� ��CG���tM�.C����Bœ�G&��� Om�8�T�@�+c�Y
w��
65,�7�%�	
75�������O�H���>	����	�����5O����O@�"|
�o�� X�l�C^�e�c�Bl�'Eў��?7�Æ`�\] �n�DjrD+���'Z�`�7-�O����|R5�3�?���t��=��I�+劎��t�$�O`tq�I�8`�h�"�4JH��6���|(V"OF��*���-zl�|�G�a�dAa� �ŋ�򦱣�/�M;��~ij�L��u���`���N�3���tM����	�R��d�ߦ���4�?����F�+/6$rWIQ�+%�=��
�ʘ'"�'6��uA�6|j\�öK09v�`�i>�+���E2 ��՗v/���W�|&� oZ��������b�j��0$@�	ȟL�I�ݍ5L��Cqȟ8^�Hb�Ϛdi��$#�Ţ�錿]�v�Q�l�M̧o��3�m���D�X�=��a��sRl�ɂC0~�A��E(?$m���.;��>ՊAd@*��d�|��*"O�..`@�r#��d�v�m�����J� �O_����	���q&0Pc����+�i�!�D�=m�h��	~&��9��Q�@����HO���O��iJ��KT-�2@�Yx�mbwze�R��9^Y{���?����?�D���D�O��S��X�����C�rR Ѧh$�(�<j�j�i��L1l���ɯZ���p��KKD�hu�:@`�m��RD���(�f��`^�0�I-l.Iq���t%�@y���p&�����R#2�2U�i�������9�ߴ�?�-OD��,�ɣ�8�ѩN!(��+ �����2�O�O,(���1���Q�BC�4���$�Ϧ���^y�N*xn~6��OB��D�U�(�)��$L���аb��,�����O��C'/�Ol�dg>���� d�L!�"$����af��;,x0䪒�3�P�K�w�x�޳y ��r򬀙1z�d((K�? ��u.T�m���#C�6M�(x�b�'3�mr�KݛV�'Vr�� #W*@jՇ�<:����"ܼQY2�'m�',җ�Ԓ|�/�=E��I�,�:��!B%\��xR�vӞ݊F)�%���$ƪ�q�7O�ʓ'�RK�W�p�I{�%��9�rǅ�kҰ��#�nْ�0� Lz"�'*�qe�#����&�ɶ\�(y;%��Z�\�]p�db	()��� �A<բu�uN���I@t��	�9Q����� ��i�.�ħ! 6!��@P�c�Rl�����>'��OZ��p�'�J6��H�OU�TH�h��H7MO����2�[�z���䖵�|�3 � 0�L��ք�$Uaxl0����iu�* ��DrԠ�����i�r�'�҉��0h��'h��'���u�%0�HW�Z��UYǀ!����	�ʪi�L��?q�,F�_��!�|&��9��$W�H��|&���X�c���sK�'0HH6�=#��>�&�8���ѼR���P��#Tz@b�n�MkE�i �H����,O��$)0S��؆��1*(�|Q&;e�bB㉇t�.���U�N�V��'ƃ#���/b����d�O��<	b% ˿<�l ��dh���eR�0�]p� �8���-�b$�ȓ&��1�uԌ/�����_�����M�ƫ�'�1�Jŕ6�هȓX���*���/I�R��C�@WyLh��m/��8sA� �X�uf��Nm���N�`ȚB�G�@5d\֋�l����,�±�C%�6>�H|8W�K&n<��ȓp�>i1 E�9Cf���`K���Ą�{�@��	�5�<@e��G�h݅��u.�r *��D<_���2��FV�<�R��9�ͫQJ�0m�Yzs��T�<���[wZ��Aթy�Ă�N�<����3���k�ǅaҘ�E�F�<Y��݋c�:���%�qȵ�!�C�<�Q��3� �sF�BT���čY�<IbH�P\�����Q�Ԝ��*�~�<9���~$�d�&3SJ���EM|�<���X�d�-�a�M6��e�% O�<!�m�$g����ʅg&%Z�#�K�<��It�-��_�p�d�@q�<�U霮E�p�5Mωv���	�X�<pn�����f]�r��|���ZY�<لA�88����D��87Y\���IT�<��Ĕ�4vI�67 ԙ��G�x�<�lȈM6b���L��Rd�<D�p���N�DhF�QP�0�(۽s��C�	�G)�B�o��Rq�6ɚ"F��B�ɧ�D,��K?}@Q+T�ڥa��B䉸IښIqCFNu��#*S�CZ�C�Ɉ|�@�W����bĔKRC��3Md�7%*�PR����C�ɟ=�� �n�
T�� ! �1V�C�		Gl<!#M5k�B0�cѥ^%�C��sζZ���0/�"L���ӄ.�TB�I'�5�����{�D�y��Q�X�
u�E�M#�������L( �R�
���A	T�s����4;̅ �#%�)�矴p1��.�J8;�
9�|�)�e������s��|rǁ��0�J��UL��0���y2��Y^�F}�L*0Ј�q�r1�cOX�^����W&V�<��;�@��
}>2�`�)������ԟ��Q��]�B��2)���ቸ� ����>)a�\j~"2��=��H�:7� � �^�vB@�"�G�c���O`�h�w��	���)\)��A�ǌ,E�5�� !������;T����S�J3���9�"�P4`L�'H��z�
Mn�45�7R� �"�
t��l�ЌϨH���9ʓ*�����A,]֕��[�-���h�J�NyR�$.�����;�>�b�Ӫwt�Ea�M�u�\!��g�?0.B�xCoI46Z�Rs�	\����*d�Q��K,GaB +TGD�_��L����L=��p.��D���4jL�?�?�$Ae�"%�5�P(=�M9¬=iǘ��#@�$xJ�DH�c܁�`$�'|�r�lO�q�0�&�t{�R��	gK�%�i�a�RPI�_��>�1�*}�� 0�`�0w ���Ĥء� /&��	�t�:H�JMHD�*Jb0�"�
�̸�ygK�����=nU0�d�O���dJ�{v�T�@G���V�P�֦+@Q���#FȘf�B���$:��@��Xyℍ)v*��5�H����*���Ӹ&/B"|�@/(��e�F�e��<�EԴKd ���dN&.Tأ>Q�ٓx�DL�;�ܐ`v�� �KG�y{�l�;RL�]�g��S�L<aem�uI��Ҵ]��(�C��/>V%PU� D*jꖠ�O"lS����C�|�H$���j�]��CI��r!��o��4��Zy"�O� k,O�IHB@�+�|���Gu����WJ�\2##�>X<E�6P8G��!y�L�s���C.� �q!�¤}p'+��~�O�䊖�~�"|+�H�}��肒B�'��I��� �Zꟸ�����H_Q��T�[$t $�³CCT��Y�C� E��M�P��n����'E��X�oT6���r,^<M��Ƒ�EzFG}��^�oG���I8K�~d*3O�X{Luku��+p�0@.?"��'��9�*�{���W������PV� ��+B�p@��s�&]~���RSaY�p\~!Fx��a��I�p|pl�#�ۀL)(��Q4�&��r�W�`��)֍ݛv5���j����6��ʓo7|�nH�"]R�1:,6��f�#Ak2e��Dc����U�Ʊ�0�.CƟ 2ҁډ=�=h��%��D�dLe���U�֑B�PP�ɪkhN(S㭎y杛6AH$#}����u^�)��oΙ)�ү؈/�N)Ey��,{8�-BCiP*���.�	M0N��O�0ܖ����������;���iQnv���<QbW�q�,�� ��u���3��?#ǒ�I�>YC��N:�G�Hlqt`S5K�k��	YމnZ�DƞL�g� B- x;C#��$�9�0(���۟����H�a��ESgiL�:��àǹO
��Ex�AQvC
��ɸ(�t�M�W�U ����[��Ys*0k�~���іw{TY�6ὟX�d���#����;������C��y"�P����:ux\�3�Ӗ<^�л�`,^�4�R�υc8loZ?:���C犴{"`�1�k-Ų�'{`����x&� ��*� �fM�*��G|�S��2��a*��t�ަ�@��DI���Dx�W�+�tri��#�8�b�"�d��h3F@��V8y��r�� �gݍReɧ5���L<1�'D�6����"h5iڮ)�d��sxB�jG �:nFP����OZ�(�`���[�
����)#��(Ըq�"����'%����
7F@OZ�k��f�$�o� �Aa+]�A��������t����}�%M"�Ȁ���t0�#FbB�a�K�l�@�#gF`�\���XH���(P��ēƁ��,Qb?�Bѵj:�D�0�<%	$�'o�OO�hC'*�u�X�D���V�����4"" X��U��*H)�H�:+�nI �&��yB����u��±{����
��n������$`�PR�O���~B���f>%'���?�da�KK��'��,��bT:N���b�pE��SƇՐ:fօ��Q%�0��.A4�ם�U�(�CVG�9�ē_xtt�U*�576H��Ǆ�ܠ��GW7%�Xqg����(O�Č�/]�ܡͻI>>dÖL�8o���۠[:B�lڅH�)Xe��� X[�K&�� ��ץ3@!��`��3��D���}�J���}"iO�R&����ǣ��a&��
��Di��.@lԙć��V@�1��^�U2VdZ��~�Oz�OZT��غK�zP�H�)�6���҅ R�A�1�BP����Wj��3�.\
$	�_#(�a�M<%��O(�	~~�䐙xvT����7�P�!	���	?w�n�+��SPє07߮Js��`���!lע�(ê��V�`��`���䓖~��?�� ���;�̕#:N��G�ᦅRă?���p���O��"�Aq��(�������4@M�bF}dh�$/�S��H�$R�<��9�4e�,R�"��.V�L�q�}���\P�$�D
d)_yr�I�\-��s􆔳q�xa1�G��*"vp�'N�$�
O�D˓w$�����I?��)G�8��P�R�$D9�E�%�ha��AUp�ɡo�)��<�G���~������]+d�J ��U
h;�eEO���:���"��Oֹi�DE)��'h�pY�'�?o�6��p �Wf@A��w}���C��9�S�"��9wX2@ �z��+�Ś*�~���@Y�1Fy�'}f��'g�Lwb��h���� I�%V$q:�icNMEy������Yry2���!2�%�x�����ό�P���c�*�j���[�Z�`4�TI��WrL#g�P�k��\��%W�>��>�"hdr�PX�MR4q��D��y�B��'@bm���S|y�\r��������>di�N���j��H+��LQ��^y���c-lu�'H�Qwr��dP�i���3[�R�ʢ�7F��@�'Nl�He�O�=�'��	@���d�-� C>� ��O���(��(O�n���~�"�63�
�Z[@h��
�q2tV��O
�=�O�^��$V��3R�ȃfة�q���3&J�1�2��2FbͰp�Oh8�Ν|
�ɣ&�v�kt�A�4L�	�y�Q� ��[��0�,O��B��!:��^�q\k��NQy�� J�
��)t"�v����OP��iX�g��}NO8�������< 1��ye���d5hE��O��pU�YIjшF/���U#$X�#�^�k��b� �M�c��7�>�&%] ��O>��m���t@��$�`%��S�0\5�ro� P���I&F�}�0����\4�vg� �y�M¦d*�k�H�J̩�6� �?	b����y"ĝ(j0!���~���$iC�\�+ţ��O*Ш
QӷJO���>��³#�rզ�^>�B'"UW�I�12��eBS�m�j@[r�ɛ}��4X�#�O4��򦝙�)�?�0�)�$��,�����
���)��f�t��ϓ�F�kM1zi�8k2�Xq��=�ua�|1�5��>y�'9��π ��E@�mθ@V�/6����_>EYd�f� �\�dJ1���Q�MQ�)F�㟜yw��#Y
�"�o^E0�5�d��4�O�	�so�S(v����#!?�@J�'��@�/Y7@Z�)A��K�T xփ$kp�t���Oڪ(	E���k�EіM�!ۺU����U�L9Pa��<��e�+hJ5�O2���)�f�VLyiE>Ov�!fʑ��'�H��v썭&�X0�4��=�M<��,C:�C���4& T8򴉁?Tט�O@�rdi���+�t[�La�4&��1G���2g�6:	�e
E��~Y�Zw,ڈi��l���^��:q��1��.�	�}JŐ �K�L`��FX�k8Ɓ�Q�U�4;���K�4��k�X�Z�҄�ZS��6,�GF\�kH��4NA�dܢ�Sd�|2���V� �����Q
�� &�;ծ�'a��U%�%�i�m�(GzZw��@ţZ���ء5�I�R(�rd"�q��0�l���y���:D[܄����S�����O�]��ək�B���''2�;��?˓V8��4M
�����M���v�)Oj��"3��	�)�x��D��?���V(\H`�FJ�\��͓�J�%.�R�&� -�u��O�U[F�U�r�'s$u����N@e��d�ЖE�@Ca���剝�� �%�?��@�2 2�<i��N�% �f&�<�UiЂv��U�'�����Em�����d�T� ��S�gR�`��L�����I,r�<�x"��)6�̕���' T��!|�
�E'��Ԅ�p��O��=�O;�%�'�V�sĄl���dγ2,J�lǿ�����g�IY2/ؼ'�eZ�f�<ɔkʎL���oA48�<�S�A6�򤫟x*�\�d q�P7=���k�OZ�x�1mWE�v��$�Ҝ@�H��F(�.)� R@d*	R.��T.���hBy2/ S?��O��^�g��a��F�k6�0�W�����V;	ڬ���� ��샓�)��h�p��/w8�Ѐ5�2�Pp���NyB�x?���ԟBa"@�*w�h�C$��hLx#�O0��vϝ���Ob�´�֤�?!DMٻ^`�S�cV�|� -s�Lë,���~*��<����!oYF\��F],#�~�뷎T@�m���X�m��������@�gh(�$@��A��eJ�2��t`��hv!�'����:��J�o�*$���]ǟ,B��q�a�/�7�LC�˖X���̍06{�Mr�D�$>l肅�<YH�c��Y��j�$�}��i1�C,;��:�û<٢�XL1`�R���//$Z%�I�]�'��]�u)�6���G��/�dY���΅��D=:���a	k>]H��/�'�bm�
�/u��GЬ{+b��&�6_ �P3�)�N�̸�*��F��.]$��3 @�=���B��*/�|��A� }� ��	D�����S"�a����L�� �$���qc�'���a@f�6q�X��Q(4ɲ�+.O�`�`j����`$�
.�h�D�6L&���E�)~q��
�<�}���ݼ[���1l��t��K��;c�%j�p��V='܁�����#�F1����y�Փ#A�!1�ŃS�Ejq������6O�L���ա3h~�k��X�/�Q��S���"	Q���&�^|\�A�E �U���:��p;E!���@R4�����u��	,���F������gJ����=��O�\ru�
	P��n&�~��u���A�v(������bV�W��-��'�0h{%�9O���T��H��(L2��n����ԅ%`)�FS���'����WeW�<��B���"���R�\�;�vDGx���b��y� ;%LU9�M�@��z��ר��Q�l@u�ɏ��)�s��+�J�]�����n�4�A�-�\}b%�\≼"(���剳 ��q��,�>B��i��m��	�MM��!��'����/�DN�x��V)1m(-��'{"@�D�Tn�'6J�kGQ���A��h(bHR/y�����l'�O��
�>�H�=@*�u�p*�H��ңLL�<��$N�oȾ	k$"�:X����օJ�<�����^S��f��M��`�B�<I��{>ft+Tk�mX�ԣ�|�<�uÚ� 5xp�#	�X�[��Tv�<)� X�c�n]H���J<�$����n�<�Ì�i�m"�̝�
S��; �n�<���2(а"�	^=��S�f�<quc�?'�*��+$.� �Q_�<!4C��A��
�Ä;;�I{"Q_�<a"�1$�HAX�)6}liP��Oc�<1�욿:�:�Sᅚ2=%x�mK�<9���x�>A(�ȍ�<| ;�o@F�<�uǓ�A��}*#��S�0y���@�<�ʙ�^2�00��`Q(���gUS�<�Q��6�����4%�`�Ia�z�<�K��+v��@$��V�\ѲQc�x�<qU���L�����%�%[x�8�s�<� ��tcR$�P���q�l��"O��C4 I�Kd1���lDP�"Ot@z�n��*��0:g�_�%Y"OL�����T�\�Q!w�j�Bd"Ol��!`K�?[Ĥ�6~Ɇ�<�v�a�S4pZ�YD_3߾|�ȓ;fe�Q�S�.pD�y�W��݇�:�z�)P蛱?���Yǅ���чȓ>&�@c#���@�q�_�7P�ȓG���@C��F�)�˖x-�Ԇȓ\$��[��K'�hx��&��	J$���c@��X��1�K�#o��(�,4D�0QR�WC��I3*�3C��02A5D�0����i���)���
zn\Y��2D� r��Ϗu�@�[6["S��/D��℡�+��hÆ�Q�w�-D���En<f�8�ѓ��a���(D� d�>Ʈ��W��6���y�D%D��b��O�ud����/a��£%D�������SD�X��t��#!D�T;�D�^�@��/��$� D����?eL�B��[���*s� D��Y�;A�z�0#E�7I<��9-2D�ԢLU�O�z4!��j�P��+D��xr�Ψ��XT�װEl48��'D��b,��@!P�A�"��[�) D� 9�!ݚL+�)y�f�v<�|���:D�x	��˗��afhò�����D-D�d�!�܉=�.��1�V�+�ZQ�b)D�L��P���h��djR���e$D����ةf��KEGo&���+$D���1�S�6`PSwE=k�X8�rA'D�<[�P0�
�J�S�k�Ft� N&D��0�J�jliJPꄝeE���e�/D����#��Z�:Mk�C�_&��F�0D�42��>-��UC!J$���`5.D�*%�G�8���(Pa���|�+F!D�s%�3��PB��yil1��3D��+�aX'y��a
��I ���G2D�`#`��9B� x� N��d0E�2D�� G.FC�T��=�⩐��-D� �2J���H�HF[��2�*D���%V�IQ��@I[��,D�T*!���_x�,�*T�_.9�q%0D��+�,\�w��l9F.��d��:Ӌ#D��A2݆ 6C4H�7��3��5D���6��;Y��|��Q�	����a-8D�$c�Y3p(������T��p��6D�H�`���Y{^�[&M��!�$��5D�X�JTx���8��܀s��1#�l)D��0Gi(d�8ࠅ'}z�q�׋(D���b�t
���JZ9�Qk A;T� � I=����� i�<�H"OH���F�>d�B!!&�Rg"Ot*�C�,D��)�풻I^��"O���ʘ�5��8��m&R�`b�"O��#�I(-m�a���߮&(�4"O0��D���Y'N׫`�0"O�E@5�M%�^yh��͸35��"O�@������S�
d&:d"Ob���Ѓu� ��fiO	�P��"ON � ������@I�����"Oj�L�F�Zti3��l��s"O�������`�A�!-8d  "O� �m��!�|�AD-�;-�p1��"O�����/�"d�q��?�<��p�24��P3�V���'�-ވ} WB=D���.�<
ٸ4A!�L
���K/D��QۉahE+�I q �a��.�hO?�䇈	H
�҃�4 dy!���RB��)�'$����c��d�Z��5M�<sNh�	�'�h )��1���mL/7��P	�'���:��%u[p	3EE�����'��C���-��QQI�(A��ٳ瓼ēP|y�6�C����b�b�p����ȓ< �d�!ʬ <�*�aW�� �ȓy�^p�6�[F�Z�9��νNʵ�'��}��H$E�V ��M��0��m�Ũ��y�c�)=$2�P��G� N�� �m���y��e����)r�:&�(�y P�0��H�) ���I��P��y���2�J��S�ҏ��@�C /�y���l��]�RM�& Z@�12�yR�G�^�x�Е�zTV�p�yB��I��Lm�1t@<�{�F�%�y�Y�C�|Y@�O�Z|�b��K#�yB#�N[R@�LVP����B��!�y�D��E�%��P�Z`��%���y��-
���$�2Vh�Ӈ�\�y�e���f�&r�@@j
��y�O�	rh`�H�5�JXj��[�y�f����8��`G���7�ѣ�y2
Lؐ@��J�Wzȸ�k�7�yR(ϓ��qED������>YN���'� ��)�ԧ�\�����5D��Y2�C�"#`3�̂�#�z\�Sq�B�k�^�ئHù�cl��
HB�I�JlVR������΀7+�4C�T�X�0@"U,c^M���ST�B�	"�2�҇���[Q0�1����B�	�P\�p$A�+Kn�Ypĝ)�C�I/�``�����+�T]3Tm�IrC�Ʉ���8@�H!KKL�+S��&s�2C��y���I�@�sXF�Ç�e.C䉇sYxS/�?d#������B�I-��P��P�HL�R��W�t��C�p�0��B�:��P1��U��C�I� jr4��!Ҷ|m��m�?V(RB��;u�09�#�d�$�J��J#�fB�	0 h���b�ޒw�*)�&�,~e㞘��	<&S�z���kx� j#��$@�B�	���q��
��fM�y�笅<V˓�hOQ>�"E�1N(����#=�"�As�2D�TP��C$t(ŋQb\��"�1.4D�$`G.O3n��E.%8|R��<D�4�vM)f!#��/mx�u�'D��;B��oR"�	�aM�-����N"D�ē ����I
�;��h��!D�L��a��(ډ���/Ҵ�b&�$D�tka+Վ��!J�(B#wG�����"D����+?,��*&���B&��"%f?D�8����vm�U��[�>tr<"�*D�|A��-L��Z�n� [��<��+6�O����<�B�<^��03-�|y�p�U�g�<i�`^�T�,�!�
�$�z<��ȁH�<�$'@�ʲ��cI��m�v Y��[�<����+4�H��Ã�=`	��86C@�<����"�tH7�֤{���c���R�<�  i9���j�8�Y@FWCE"���"O�D"����I`zL���7!୚b"OTRȁ�'�|��.��*���"OLp�ٲ h�$h���[�@Ib"O���ƇE_=�H����Q#��x��'�2���&R F*�U+�ʁr!.���'1�S�Z&��ڏm�P��'��������И1@�޳e~���hO?uۑΎ�����9�p[�Ht�<QqW�E���5	��(" i�s�<a�i"ʴ�I�e��JXm۶jp�<�VC|d)�a�ԜI�D{�%�e�<��*�E�@�¢zV����c�<�a�ʌC]��
�ψ~}� d�`�<� ?�0rw���~���QeVD�<�`�� +�t�u�C8Xayb'{�<�E�*��p�d��4��DU��\�<��SPZ$�bU/�c#��0��]�<IĆE=4���s���-y�!U�Oe�<���ʥ�j��5��L�G�c��hO1�Za�U�He�,Iv���b�|`��"O��C��ϖ'b��@"��lu"u"Or,��ň�Qm�U@��a��D�"O4`�v����D� ��.u@0"O��MP5hX<H� ^�,_�`�"O��Tl��W�D�)2�ԣl���"O�PGm۔|`>-��Ė@�Y�t"OL�q�E�(,�<ac 㝫Hl��S�8����#���ic��jBt �U=]��C�	7$?b|�ą�r�FdRg��Pw�C�I�l����D�O&�����Jz�C�I$#\ ���L
Ck<t�E�A2Y�C�I�8^�u�E�ϳ	�H�@C��n�C��&|��x��X�i�N�! �!~LC�I*+��3���G�ܤ@�%P=hC�	�&`c�!ޠ�0��CnY�+�=��^�җ%+J"T5�І1gb����L�'��]vvIr�cˡ+�0������Ç�w�u��Ȓ�Q�te�ȓC�ʝ	�`Y�!�	�E�'9����%�eaï�+5Р�c;#�0 ��k�t�&!㤭@�A�^�Յ�8���`��]�=(��b�W$% ݅�U���i��[P��6�]�F.h�ȓU �r���)�\��
+���ȓgu�dR��#z��J���V$l�ȓDHS�+�+-���U��r��d�ȓ�v�s""�>w��7��Og2��ȓ[?�i�ׇ��g�%�'�sǦl�ȓp���gaN!?��	z���ȓ*�j��R�u���� K�p��ozy�J��%�p �`���\����I��9?~%��n\{��0��w{�+T��^NPx��S	|{^��ȓ%vX��C�
����t5
Ąȓ<�f���	]�I΢�i��Z\8܆�
p�(�6�$��P�6x�%�ȓ{;6����LL��@��\	N����ȓ+�J
S�:DupG]c��H�ȓ/�ޭ��ǻ[�qiюw`:���NZ��I��O��	�L6* t��ȓ�h"c��@	`�$	Q<?ʎنȓ���&oͽ0��EQf!n�]��5/03�ї@�DLZ�H'Յ�S�? ��I�b��sm
�˴4��"OX%���P����cH���"�"O��cM �LA��
q�6�"O�Y�`$$)]�X!��ɞ��@�"O��K�K&*����Aw�U�2"O�t�0G;%��U������d"OD���
�+�$x�:��0�"Od���8%��p��a��r�x��V"O�d:�B>5����ݔ���p"O�QTLϷ����]�GL��"O�Ŋ����x�L�l�\�<*�"O�=JR��:r��m�c���TK�u"OT�ᬐy6�h��$Z?!\D�a"O�[�� ������=0�5"On��Vc�&=wJT���'jt̻�"O䥨􏍲bJF�`S`]���rg"OT���,�
F�YP	�;�d�C"O��P���96� r%O�"�zxS"O�Q!q���ĢV�'`[�iQV"O���ŦS�t���a��T��"O�1
&������5:�x��"O֌:#Ɲ&+Ơ�6 �o8�1ru"OJM�wH���	��	eS ��"OdةFB�/
\��& \�DN�)�`"Oep�/�\3:	w�ߵK.�"Oش�$�đ-O�����[?#]: "O���"�_�+?��r���h���d"O��"��,c�fd��Ąu;��x�"O���IO�9�l�(4��O5�d"Od�2��E3)	�@�`�W�M��<g"O����)�4R�"~{�acR"O�)���=x�)�&sF���"O��"N~�f`�OvC��U��y"
A�#�:�(�$�~�e��.
��yR��.S�����R�$��
�"V��y�n�+f�9ۧ�\�!�@��@E	�y���6xf
�S4.��!�pBɶ�y��\3�@E�Ε#�l�+P����y̅.RҰ!�� �ա�l�=�y�o�sm��A�bʭ-vy!%��y�i�%�6��d�B^`� gG	��y�:aP��B�f�46�vuYc�\��y�H�<�|%�q�*0c<	�n�yr� %`�d�#\,-f���K��yb$ï|���i���� a�� '�y�#�l�b�-.�yd(��*0E��'"��H���Tx�fR1�b!
�'}���'�#eY��B'����8�c�'"�I"�OܡC�Te��V8����'~�$��o��V���R4Iɶܮ�s�'$`�%-��VU��4ݨ?��4�	�'��X��0��S�Ӊ7R<i�'��Xs������L��jX 	�'�.`�T.%Y�Kg�M�v�:<��'�.���$ܞ��$b��?W��
�'�L�3��ٟP�@����1=?P((�'ò�YT"�L�*T�s@8YL �'t�u��R�g�؜�VB\�4|j���'� 5d9NF�����9%��ي�'4�0��"A��HW���-}��s	�'$�)ы.;�Lb��L�QF�X�'<U2ri�-=E�$�j |��%I�'�ZAiPo�*Dy�0��ͳz$��)�'���*���74a �
�A�C|�	��� �(4�ɧc�XM��ӄ+�.AcG"O����S m���J�l�
"�� "Ox0�Bڽk�@f��|�ܸ[�"O��孎�KL����5�iҬ=D����&�Z��U��R.7)�mӄ<D���v$ؗv���( lM�`AjUP":D�T��ױe��K����*�R�--D��A@B�&�2,��c��̍Kq�,D�L��"	;5�θ�F= ����1�?D��x��,^ �iB�P>z��ф�?D�ȐЍ˾>^� c��OPq�x$�/D�8�[%'7x� `��~]�U(a�.D�@Cd0Gᠴ���_�>L�5G D�t��O�Kf�ub�1j |��m>D�,����ee���і8_�h��:D�0� � uolj7�Q&N��1�g�4D���	E�%����  P-qI˃�4D�ܒ���%������*���� h=D����%�f�Y�,��@a�;D�\y+ܯiϢ��qe6@ ΅�V�9D����#́�����m�7 ��u��d3D���c@�i�v�S�Q <ڀ	J'l/D�0Zq��=�:�+�.� �H�� D�,�Q���Hu$���j]�� 2�,D�����{4!!�M�I�4�R�)D�
�N�U�1FP����&D��Q0!E�]�<i��	�+�
P� �"D�L��#J���Jݠ	�"��*ٿ�y�j�+Q�������  P|�bb��y�K�1���I�o͵AɘTSb���yRoZ����؆%�i&�!�`��yb��q�����̣�~9zT劃�yB��ht)Be$oV)[�C�!�y���lb4���]�d��T �A�+�yR�\�[�n@q�"�bƬ"�B��y�.ͩr���i�����y�ƎGα{4gǙoO�Y��@F��y
Tp�!A�ټd��tq�к�yҌ�cy�8���B\�( :'�Ӌ�yb��R%���&Rp���&�E��y��?��P�2̄O��C��yr�@�$���[�M��!��1�`���y�¹M@�}X._�����/�yBa��x�V���v}�ԥ��y�G�,H�A�Ӑ}��@�(А�yʖ)j���i�C�b9 ����y�Ꝯ/1�u8�G��X�t	y�J�4�yB�X]��4��,�b��䡖DM>�yR��
�(uRR恆\��PC���yB�,�A�e�Hn��h`�K9D��e��u�pI��
�U@H�`�8D����' H���IS� �zl6D�H���u�"t�D&/����r�3D�`ie��8"(��rj��!�M˷�+D��a�̗6"���J	بT�����'D��Cr�̿{���s�V�����H D� a5iV�u�0��"��8ۆ�?D���E ��32�R�69���A�(D���J�m���p����NC���RA,D�8p��Q�!�t��vn�
C@֭4D�\�1jW�d�,��7�F=EP��	5D�H�d�
k(�j��2���j'�?D� �®B�Z,�8+��C�#ui�/+D��A*�.,�P�����/
��p�'D�� � +v�7c��̉ &��ml��V"Oތ�"/p��� f�<Q:�9"O�r�T����҄U�nI�8�"O��{�Fޝ2�XCׂ�+Թ��"O¸yWʊ4�0��A�#P\��*O�ՈE�R�q�p�XCC'!�z	�'�lJ�#���`*3�U'���'���0��H�z=#�ʄ(T��T�	�'�J�����@^l]�cΏ_C�0	�'�:T�B&�C��{�e��A
�'O��+ea��m���aǈ�	�'����D��7#�P��
�idic�'Ix�0�D͏�Hѡ���'W��Р�'��ʧb� �d��� ϕQ��)�'{�Ը���1
b!]�V�J\ �'\�чK��e�X�F8K�晲�'Ҝ��1�;O�p��U`V2FH�0��'��%��"cH�E��#S�@�X�'��y��X�+��J�G�=RF6�x�'|4������:4H�*N��ر�'�\�g�����v��J����'���PĆ,x�t1�F�X9M@�p(
�'� �sRQ
������K�6d�	�'����"�͉A�Z xV�DX&u	�'p��(�GG�-EN1p���3=�P��'^b�P�,���H2�.�8q"L��'y>L3t�
�͛0@5����'Rd@�I�,v�V�Ig�A�.��[�'�0�k�J59��CƄ!H� �	�'�y�!�,,3�e�F��#V|}�'>ɻ")	�'�1��+",���'�T��c@֦\Th�a�/��C>�([�'v�X�T�V�CA( S�'�C}��'�(���*|��ų���k@��'I����

iI��pN��a�':����i�t*�5k���V�p�'*Xp��ɂ$�Ҕ�AKˤX�4pp�'ґ���T�vPHh�"�<Lȸ�`
�'4V�9Q��<�Fತ��S�"I�	�',��CM��z^�d�#A].U�����'�rcA��p�B�@#	�#]F���'�*�h$%��Ln�mQQc4!�0A��'����`Q�R�>�0B ��0��'���h6�K�ψl r�	p��"�'�*<��)>�Be�ыW2~�>%��'&��ؖ��33:m��`^=z�@�h�'.���ED]������l1���'����V�k��m�p*ɧh�T�B�'�NQ����;$���	.�]�Z��'��1фC�eY䊐V�5��'w|��� �46: 0d��U&|�B�'���Ц��E(x8C���J��Pa�'��PѮ������,n&�@2�'@l�jȒ y�6��$�2N�ȳ�' \yce�Q�Z>x�[����
w��C�<�U�w4(I�խT�R����0l�y�<!�KZ,]<�Sk�*ܸ٠�����y��h�l ���5'ݚ�r�E��yb/؈[���Г�� ���t���y�@�ax^aY�N�%'�u3����y�C�L�$�p�Ѻ����#���y��K9@\`��!٬<�n������y���#�~�P���8>��a6��y2�D�%|��(C-����s�KW+�y
� `�D��,xh%9D.³L�B�'"Of��ϖ��=����lE���"O�5��ŶCZ�x�$�+���"Op 	��+����E(<9�PV"O5��_��c�m�,0� "O��*�\�&�h�-D�"r\��u"OV���N
i�������$
.�^�<!��D((�������~�Μ2�Do�<���ɮ=*I�c�+O���&�a�<T�_�.0��b�RaʺL��\�<9�*Ŵ\/f��WQ��Zp�[@�<�Q	X�)��	�cl��}���ѯ�f�<)1M�
�x�mP �XXb,_�<�BE�=��]+����Z�~A4e�_�<���E,Ȉa�`
�}c�st�<� �M����'Y�@�0;��Yn�<ɓN�,�hb '˔I �ࢴ��i�<Ʌ�����LR!݋j<�#�Ce�<e)R5/�<��3�A�K�:9*��Nz�<�D�ϖB�")��a��eؤ�IZ��B�I�@q��cJߍ���� �&6+�C�o~bpi�-P�C$��h�F�"��C� :8�H���!"�Ա��H�*�LC�ɳC���f��-t�n�����HN\B�	�i���-�}18���KH�2B�	�`ʴ-�����Xy"`&D)�BB�ɹ��(g��%@�4�YS�ý5�(B�ɰ;�+�%_�g���%��iB䉽vj�p�	�����_�<�(C�	)�<0��鉈 P�D�߿&&C�I6e�~u��+'�X ��� ��B��):�0 �;+��}I��E1X®B�	�Sdּ񦌚O͘��%�^�3��B�I�5� آ�[�Ҭ �-�M|B�ɕg�^���G
	�Z|�7(N�;�B�I9{�V,��B�~�:�
B�X��C��
�e�W*�lhjF ]���C䉎mÚ%胊§4���&̏˨C�I.qfFi(�������� 8يC�I	g�X��H�%THء
d��<x-�B�	�ynLѓ���RZ��dD�#��C�	.#l�(��G5p쐍���F0=��C��,k�< ��&vh]��CF�2`�C�	G,� �hG�:�Q�S&�$e=PC�ɺz���h�;^�}�T`�;I&C�I<�~���%˄Gu���E�U	*C�ɧI�>)K"@7ź�4�� 9��B�#!�H<��(ΩC�~��rLURzB�ɯ4qx#&ŐE8��e�t���'[�#	�&�<t��I�I !��F2��	�@dΦ�|ZS(��2�!�$U=86����<�8P!�,!�+Aڐ��!/f�\���̀�{\!�Y�p�Y"��5o�S�E�o�!�䀼-k��Cˁ8k��"PƩw}!�$܂E�:V+�:tT�eP�' 2]!����C'|!���ooHу�G�8J!��\�\a؀�A�5��<&d��o,!�dU\"� �摵�Z�
4"ȵ*!��̟K'��h��ɫ9A�i��\!�$�@8 �����+;$�˖��2F!�ck��9A�VjP��JߎE!�dA5:r��R��7ZlU��cB�!��R�;ǘ��@��FY"���F��!�� ��Z�.bE���v��W1���"O(|u���nM�xZ�"E�U��l#�"O� �p*\�k��+S��Rg2y�"O��θ�@�!
%Q���d"O$�A���#f���~8�ͩ%"O��B�Oc��;�4,`�S"O����c�Q<a@
�|�u�2"Or	]�p3��Z�]7b��"OP���8>�J<��M*H�N�"Op�(ъ��7�h@�ggL��x���"O^y����hF�� �ƀ�lO�i�"O����\7"��K%ʄd7 %�F"OD���$�j��X���+c#L��"O�݂�Y:w��5(���+��°"O`��1�чEH��*R0O�:���"OЕy��շE��)Ë�zY��"O��b�R9avZyC�Z�E���b"O��gh���Jy�ݲx�T@�"O��*�*q��Pq��Sj�@�7"OR�
bhQ?yJ5!���:e��AP�"O��r.ɩ^�D"Q�+tV^�!`"O��h���(�e%S9@f�Ђ7"OJ		��0�)r�ϯM��ʢ"O�0��v��Tz�"�(0��YK�"ObL�J^�`豣T�	�7{$@S&"O��*�$DE��%��L,Ui*���"O��[G�ȸv��rM[�QtTk�"O��Bvϙ=i�L���O)l;,���"Oƥ�@K�72��Ca�һl5�)�4"O��[�O?Md%�ʅ �����<D���É�{Z��Ɂ�I$�4h���6D�����<3<���	-	PJ�K`j4D��A��[����O��H��uk7D�"�Lƈ[mR�Z�� '{X�x�e7D� q��O/*�=Rr	�'8F]�Ƈ3D��UC�&WP�A�X1}x:��0D�xy�d�$7�)��i�o�j(�pg!D����
�!37�=�� Cl$I�� D��c�O�F/��ٗ��fSPJ�	,D��"�#/=�n$@D�Q*v�j�G<D��S�x��Bb
{r�ph%D��"���0.lIs�À�d�X�c��"D��q�藮k����'^1 `F|Z��!D�X@�AֵL�J1���,eG�C�4D�H��gҰA�{�e+��QAK>D�4	ť˾j,�M��%�>	���":D����C���l�8`�Z���K$D��X�OU-P���Ù-rH���4D��ء�]�p͢5ԸP��B�V�$C䉆wD<5i�Ķ
B��	��c��C�	)+�r8:���d1�W��#N!hC�Ɂ+�� �MT�pH�kM/�pB�	�,լ��j��{�|0[vl�3�"O��2qGϙ'`V���H
YP��"O�\��(V7S�fp+��^TP��u"O� a��� ��5�5a��zHV�'"O�x�i��uϴ����JI�pC�"Opxb+�-=�b�I�Q�$�j!"OX�0�
��ʩB���E�h��q"O�Ay2�M�u6�x�BϺG�ؙ�"O �e+��x�ؼ�@/Q�b���P�"O�����а�P�b�pjո"O���A��'R�h��"��CN���"O��h�N�{Q9�j��i,��"O� ��âH�ie��2�hˠ[��yu"O�Xx���,��a�G���t�&"Ox��r���eM��*����3�y�"O��կ�w�欃$@L��\�C"OHq w�['G�@�bO��\�m;�"O����f�a��$�F�@~~�YD"O��"��ߠa��b�g����]k�"O"}��k�7BdP� �:T����"O~0�E�S35�%��	��L��"O6D��LPA�l���m@�
��z�*O��Tޟ8��ZU�5]hx���'��|#�aU�r��z�^�X��IH�',�m�D��-=���	�L�̊�'�2ՠM(+�<Y!v*�Z]t���'�8�2���-bc����{FYC�<��X�"�^��%GX-�h����I�<�p,J�DT��mQ�����%�k�<�TO2v��5
Ŏ�;�蔁r��_�<a& ܣ.bŊbC�
9�0X#�W�<)���H,֑Ȁ"	�0ٓ0��x�<��&�:ƔQ�B�ic�i�p�<���L�V°���;8�&A��n�<1���_�4d���ʹ@�%M�b�<�7 ?��ٕ瑫f�PͲ�X�<y��K�E4��P��T�N=�UB�R�<��A'1� ]����?y��١��Q�<���^�6n��Y��!��+�)�B�ɐO���BI�0p�͙"��k�B�)r�Pe
���?���A/���B�ɽk3��u��3^��X�g�?�B�	$B��2�
M�l�(���M3�B�	+�~Q����5sr6١�]�BC�	9P�B@�w`�7w,1K�o��CB�C�Ɋ(��=k&	���q$��t�
B�I"P����b�/�:L1P� ��C�ɶpv��Y5Ύ��ԌQGE�]F�C�	�L,�"�;w��\�e�D3�!�$K.3��H��*��2�܀�Qc��i�!�^
ToL�8�� �a� 4���L�;!��=�b����ȮU��aӦ
]�P!�ĀͶ4�3Z9M�������!�R�$b@��i�HВ	iu��*@�!��J�/�ax��S�<�dȀ�,[�Py�E�.�F8���1K���T:�y�	#F���EIS�� ��e�<��iD>��$,��5�Qy7��S�<�[�Y�P�s��(n(!�K�<Y��1=� � �jZE�����S�<��H�x�A�$�I.d�z�K�!\Q�<��k}�F�2�-ƀg�=/_GtB�IR%��!�CR�(��&*+\B��+9O,��EGܯ*3��ʇ��� �C�	x�8y�V�`}{���/K��C�I�QJ,��p�F�ע֥V"hC䉪`hx�S�U�M�J"�cBC�	�H�|��T�+Fu[��C*1�C�
U��(P#O<��\:�dυ</C�	�7��ud�:�@W���2�B�I�)l���ɋ�����	k'�C�Iz61.�V���c�N�-�C�ɛ�dx��+P(�r��G�H�C�I4T��<ؖ�D@|s��T/t�vC�	>lT��� �$<R� S�d�LC�4"�$��	�(x�92,O�,4C�)� D���n���q���*R�Tx�"O�������EH�)Ȃ4S#"OLA#T/��Sn`�XB�Q�x��EJ�"O�@j��g�p�H���8��e+�"O�(`ʌ/��M��CB(��C@"O��r5�_�e���-����"OtT+cF�0hQ�0b^�*tj�"ODXC��G� ��Gʭ]����"O�!A��A�0W�X�df��P��y"O:����E�~h����D����q�"O��u�Br̛���k�����"O��ytQ�E�F���b1�x�w"O�9��L�c��B"���,�(1"Op�1�R�\,�Ё�k�a	"O�\���V�|hp��A�%GRt��"O���F�Vaڜ��V�i�`97"OH81b%3��:��
5U-�J&"OZ1Fd�+B,�/��Z�� U"O�A���-`@4�0 �;BԤ�*"O(�jր���0�� �P�T� �"O���Q�U>K��1�#jT�0�"���"O�$)c(��`>0i'f�
 �p�"d"O���P�&:ؾ�3��#/��ط"O�  �i:l�1�Ù^���"O^�����X$�u�	�D܁��"O5�@LKij�|�3I��5��Lӣ"O��s$� )-4�@��3�J��"O�Px����u�XU�щ\�b�b(Y�"OF��PGA�+P�	Yw��;t|@�u"O�EZ񏂚p@�1IĚmh�͸�"O��W�
�I�؛�e�(c���p"O ��!�w	puАoÂG}X�E"O���R��6i�>}�A��� ^`1�'"O8�)�O�*S�A�Bm:gV�t�e"O���c,׉AI��ǐP���"OjT`�D��)��N�78R�a4"OPԂ2�6EL� �aL*N&�h�D"O�pօ��i2�{рI)	����"Oj��s,Н[䈀u�I=@�SE"O���Щ���*1k��֗z6Tu�"Oىċ��0�mE�v�� #"OPTH��h��QbC'|�X�q"O����٘t:�͙怄>T��{T"O�\*��'B��i�!�T�"O&�t� 6�N�K��9�~HCD"O��&�'E��QSq��m��!�"O�<�Q���
x�S �K�и�"O@���`�-Z�8�t�6r#yZ�"O�P�VBY�-/�]�W�	k0I��"O�����:>Ϧq��♪$��&"Ob��[(��tؒ�&cC��rT"O@u���^��d������@��K�"O����g�Jx¬��L P�"Oz�f�B ��x� ��|��"Oh0�	�%G
i�P���0�b��"O��s���mS�LX�4i��t[&"O�0SDf۲m�tt	��[� � ��C"O��R��)PB��(��ː q��K�"O���柠G�t�3#�'V�tR�"OH�ɀ"Y%B@�֗��9"OT9�A�8^Dqca̶>���%"O�๔�T^��i!�I��j�A�"Od�� �ϯ���!b��'�|��s"OD���/��K�,}�� \V a��"O� �x"&��AG���g�]�+��2�"O�95
\�~��$0�',a�̉z�"OPU36k�2�i�ã�:R7�u��"O
����V�S�t*�� �3T2�"OR��#X(�l\�T�Bd2��;S"Oơ� MZ#u(j46BB5*Vd�"O�	�ɘ �D�U��A�-$"O�,�V�T���X�1B��zGz���"O�A�� �s� �&� �"O�	zq�X*+.q�D��' �!D*O�IJb�+}Ҙ�*��ɗW��	�'���y�	��Xd��0���hm\��'u���R�V�d�MധجN˚���'#"��g�]�����n�:N��S�'��%jU��w��	��T�L T5k�'�J�	G�_!"t�T�a�@t�z�+�'��jơ��V&&��GŘk����
�'��-��EG)e�LX���`OB`	�'��1����T��hx�L,\۰q�	�'��y�S�,��@Ir��"Z;D1K	�'��E0�Fm���h�NҔQ����''V@	�*�+@.%P�"�x��L��'� �#�fS�}����%aS�8I�'_��H��?
�Xb�`R�Vy�PX�'����� �-�$�@�%��a�'ϔ\*'�ŜZA�}�t��X�
�'m�XA���JS�a�c�6ic��[�'-�i����'Wo�xR�
�[����'�2��a	�D��0p1�˃a�֐��'k��ai,e�q��?^1T��'W�["!A@U1�`
h0���'�Ћ�Έ6F����*Ŋ`��j�'
L0���[���4�P�P':�`�'>���elñ}Ĺ�ӂ�6T��k�'�^��LH@������.S��A��',|ES`ǌ��AR��Q�L��Q��'z���f�|!��:GL���'�������.r���T/	�mB���'r�J��O�c��	KC�J�l���3�'��	���;#����ڊfc�Q��'�n�R��:[	fp*!�B_q�<��'��cB"�G��T�`.�h
���j�<)'m˹fM�m��FT$� (���k�<Q�b߄~+����-P���ڠ(D�p�2��\��z�N=7�a34""D�����ڪI�$4�4O�S3@�J��#D���0N�fm5�" ���\5�b#D��A��X�T�@)a����<cA@ D�8 ��J�\?�U[�f�#)� ��?D�D��f�.͖P��A��n��E�<D�h0�b[.��P"�*����9D�(�� ��K�Fab�ƭ���m8D���7�V(V�T��'^PD���*O ��JT���h ��)��]h�"O��Ӣ		��`86�TMu�Q��"O�9DԸF/L���K.饌��y�a�6�.�j�b^��$)rl��y�oӘ8Z�:B��#g�ap
�y%ݣg�թ%� ��1:!\��yB#Ƿa���0&�ݭ��X����yr�J�P�d�BQ�
Ê� �yr鍈x�H���4�(e�qe��y2��
�`�B�-�:�rH�W�M��y���.�����9�P�2�D �y
� �̓�o�����g户?+D�G"OĄ�dh����$2<�+S"O��s&gZv��H bL����1�"O�EY:�q�jÝM;��"O����Ŏ���P�P���F0J�"O��y��ԒA 4Q;�CͶ^)6��"O次�7������ B���"OB��q�ʈ�(%�ͩF����a"O�1��b%�"�
�i�4=Tp[�"O�L�E�<� =S��I�c���"O|�c�H�{Ҵ�c�s��B"O`��tb�p����NG�X�\�q�"OFM�ۍm�������qr"O�C��C�BH����ܧ׌}p�"Oԉ� .B���zb�Y5J�H<A�"O�|�t�
1e`�ït^=�s"Oڜ��-��`,� ��I�6Ō "O��ȔG}¸�)#G���)�q"O�m��Bտ�̵�AC^7��@J�"O<�����I�^L��"J=3��A"O(����1^����٪,ܐi�"O(P`j�<~a>��g�����9"O�t��ΞQ� �y�a� Z���1&"O���/� �Ԉ��I��=��s"OBypw�_3��x
W1H�B�*"On4����a�����+�=c�
8�5"ON��d5(D�LG
R�j��U�"O4aJB��MM�# j �&�fM��"OZ��!��v(\I������"O�U	d ۷@�4��B��[��$@"O�5��ۉH�({�AL��-��"O�E��OV)*�8u`�Ԥ<�*Q	4"O�AХ�T37��m����� "OĨRF)�?3䢑�6��f���2�"O�LJ�b>(�(�b�.m�8b"Oh9Ra�#�E�|"���"O`��H�F�&ݡ��Z3^���XS"O��!G�A}<��f��CC����"OJ���✌Siy r$P�Q���e"Ov��R��5 y����R��i�"Ov�H󇎅m�R@��kD V�-�"O��+$-ŒH�,0��L�4א���"OE�U�I5��@s�ǚ��8A"O�}j �>�"�XP��0:�� �"OX�RM�&�)$�:��ͪ�"O���Q`W#Yl��8�D��i��eX%"O4����&c�p��c�2X����"O>� pc؂
�Zd�dƉ �����"O܈!bJ<6���RQi���p�"O:1A"�;�̡����~�ޥ��"O�ႍ:b.|�!�:h�NiyW"O*���29.^4�d/V�B���b�"O<�����2���um�B4Di#�"O�8S�H"f-�# l�"G�A�"O���#l_,H_����!�1Ex��"O�|��ⓝ M�a�bG� s����"O��r�#��p4��@w�"�"O���íTC>��P�O9}C���"O��	��;q��h3�È�_7��yC"O(�a����J�:4?𥑇"O�Cԇ�1Ȑux˜�#D`��"OrX�%*�L%���t�hhЂq"O�AS
&Hs������P�n�a�"O^)'[�j:��i��_$O@r��"O� ������,&H���"�	��M�"ONM"�	�$cc
�p,P�~l�lU"OLt��[)޼�Y7��!Y�@�"O�)�#l֖ �T�CÏ�]�5"O�|�UϊAQ^h(b�5g�X�	"O�IR��,N��A��M�6$S�"O��BQl�r�:��#�"O��b���! ($iREO�/�\5"w"O��� 'FJI��n�:/x�&"O��'K����I"L�W�<:�"O�<9u)��3Q�����	��y+"O�����q")N�TC�;�"O��)A#�n�J$[Q�]u.��`"O��jZ )�f���P1�P�"O´0HU�loށa���XIS"O����٨T�T��Ĩm�!e"O��3d�+p`H�Aa#����A�c"Ol�7��e%d��%� #��y��"Oz���⃻s�S��c���B"OB��8!�tQ ��P�T�¼x"O�41�)_�'}���#m���@i�"O��[���^>z,�w����O��y�
�)v��r��<s~PvK�y��S l0�8�%��8:��P����y�n߀c	���2�:��qp#FG.�y2�Ih��QoЉ�DA���y/^)N&�`]�� ���ǭ�y��D�:<��%�G~�����yZ���ǨڡZhp�`H@�����'�������+�U�C�B�cv,pz�'� ���ƅ1��T��L�]��=��'����t�T��\*�BC�x9�'�����	|Ur5R���+%��`�'�F�d�	�m�w`ҕF{���	�'#B�*��$Qu�E�&"P,���	�'JN�s��B*"Ԉ��f,	�y�ر�'w8ԛ�G֜"N-�"sK��'���*ui�p��ԃ�$eH43�'���ft>Xܛ#JX*Y�Ԫ�'��� 9xn��c3�	d�Y�'j*��qM�7�TX�b�F4�\�;�'}���A���>��hZ(^P�J�'�,d�/U����Hs�u�8
�'�$�2#gC�PfyrB �%ea.=�
�'..D���!e�VP�VIH$c�PX��'��ᚥ(F�nW�P���L[�q��'�R2�(ͼyu�1�$��TԔ��	�'���6-�: Œq�A��2C9����'������T�D�x�� V04�*���'fz% ��?ZyHh�Q�&tа�'#�bHרI����T���ʞ���'�z���"�?y�����L��Y��'� ������O��áM+
R�	8�'N`����(��a��||N���'o��H���q�uI񢕣B�*Q)
�'�J�H��3S�Aa�յ9�h�"
�'��<��ëb����C��7~M����'�~dh�@J����J�*8�!h�'��P� �,Ң���KR�U��'7r�RN�1�N��r���g����'�P@T�- �!:ŦKvzT��'>�����H t��T	f��ب�'J��X �H�vȋ�Aq��q�	�'�f�Hp�B99�er�GDe*D�����  )���->�<���� y":ّ�"O�h�)B2:�A[!�\�el��"Oy7�Q�-T٫�#�/@O�Ӂ"Oƈ�S��d�r�b��Ii�X��"O�s�̃�@�e
!��Y`��Q@"O.p� E�ct~���#jQ|�f"O�(Z�J~�	k.N�y2Q"O�=��V0,�VXrk�7bM>;�"O$9xq#[B�ĂF��NmV�o$D��C	Y�\P�j�.̈�2�8D�гCbC�%��RT��l���3D��9��!��]q6*�H��i5f3D�T	a��sN��K��=���x4L0D�\�W"8_~�1�B��R�@8�C�:D���pOڟ*>�Y�q#*����5D�Ԉ!`�6p��	�@���/^�ۥ�4D��:�kȗVf-1� @��@E�m4D��q��\mjUhݨ[R�7D�TI�эm� �� ���J�&�aԭ"D���5�� �Nxj�%W�3.ճ�&D�X�S�ɿ@�H3�V	&8&1ID�8D���SbI:4@�{s؜R��E��8D���(��v��]�^�+R�+I!�Zz4(��+�%p�p0�7��!�D�e,E��"]<p�6�I� 	�f!�L����� K�y�T�H�&	t�!��o���ʝ���`oT�D!�с2���Ud��Q�8ͪ���]�!�$��il���G ��h����"4!򤍨Z�Y��,��Hx��J��!�d�B1ďV�kr\�RJ^;@�!�d�������K�1�P�3����!�ā�W �@��`	'��`XP�YV�!��e��$	�Z{���⁤�;J!�V�9���Q���88��i\�!��)Q�T��cOE���@�C'o!�ߎ$k�b.(���1t��h!��ƺR��0�<<�i�$�=!�U��m��15��P� �˹�!򄍵	��EK�`*]`�AG`�-k�!�ˤ�����D�U��P�ĵ$�!�Ć2-����N��h�4|���L!�D�R_��2���jØy��둿d�!�dP�.L}���K����!��B�!��<z���U%1g���1(Λ0�!���E�[U��Rh�p�U�<�!�D܁IꪝAVCE3��Х,5!�DZ��9�ǎ-�xI+E�0X-!��ѕ�xD��hl��g΁ ~�!��)b�l����@� 1�#�Y�!򄆤b�>AYAթ@��"C�� �!��ZiD�4Gd̩���Ks!�R<K?ʼx��dR����M!���?M�p�S��bXA�M�i!�DS�}2<���g��A�r��QMD +R!�$ΌX�
p�U��L� ,�/DB!�dȁ9��p�t�֙h-�#��CS(!�$5������܂CPp!RN��!�řn�~����
�&2�5��͌�J!�$Z M�򑲶��y�3��J�!���Sƞ)�&�� ,X:��W!��^��(�Rǩ�:�F�b���="�!��2�,)�L�1�A��#Ԓ\�!�ܗv�Bq��DS�OrE� �j�!�� (�Z�m߿
o��c2@	9^XA"�"O�5  �%Uk>����|UE�""OHA����9�Y�ƁȫG��M[!"OdYP��/+vT�t�	 b�84�"Ozmc�ف],��䡞9d��A"O��*�&��P؂�O�F�лU"O�)$+<YX�=��n��.(m��"Oֈ�CP�<e���T�R�� "O�!8B��%�ݐ1挜q���"O>e�#H�&Us.�f�P*4"O�]�a��~�u��lн"� \�g"O��snR+~�,Y����3D@,�$"O�䳢jJ3:����q�����!"O�`�f��!">�Jt�O�G�Zi�#"O*�ib�3x�` U
9z���"O��Yt�!���t`�qRS"Oi1E��0 bTPc�\R�Q"O$1:�N:U�|�b'���>xR"O�SA�Fk ���e�
tq"O� � �h�v��.F :�Č��"O���GAI�<��xRpC��y&P�"On���(�b�* ��.2� '"O��q������aC7X���"O���Q!�(&5Ye�H�E�(9�"Ox�*��T�]nʕsOQ:O�E`�"OЅJ��:P�-�莢0	�ؖ"O�apfY�� Db�!a��z�"O8l�� Q�� ���X_P��y�"O~�+��Ҵ��4A&�%#L����"O֑z��ԔQ8I#�#^4T@��"O��aiݸ/0�驰�3kJb5�"O�����Y�DVo�O3��"Ohh�'� �'�������N�^��R"O8�颈D� ��}Xᯅ�#��11�"O�����$%Df��H@*
R2d��"O�ж��CL�h��H�Dު �D"O 4!�[�0>P��E��=�	�f"O8�����[����oS�?�����"O$�z3�9!���臎�UX&"O���פRh�"mҝ:���V"O���B� Cr��Uː/�~�V"OR �Ç[�>�aHd�J$RȔ)�"OʅA�fK!TԴt���6
��e	�"O�|�@.��N�H�B��ª1��Ȫ5"O�}H�]�rڄ��F��9+�1Sv"O�}�&/�(}� Y��LA6��R"On�l��_�X(36��'�ȍ1&�%D��q)ѻE�G�āby�1�w�5D��c��?8�|�Q�AX�l��A�g2D��+��Ś;D�La� �j}��P�'%D���! O�q<ιP�I.x>US�*O,�C EP������L��\�"OFaC���GV�M�䊿(iP�2f"ORm{��
V��͜ z~H��%"Ofl
0�̲#�65���^ B"O^�9B%E(�.MqfdN� ����"O�%k�$A+^�8Y��HS�hp�"O,�Ǌ/)G�l0V�ܶu<P�"O��bҨ:}Y���@��*P�"OFA�'V�U����GX�s��H�"O�&#�n�0�p�"��L��"O������A�8��O<C>v=�"O�u�b��dæp��M��:�m��"O�ǃm$�I9�&L::�ʱIE"O� p,�E`��6lc4�I}|��'"O�e DgV���\�#,�fs�|ط"O¸!a
�����-ӀOr��� "O�ܿ;�t<cĦA��ؒ�"O�|��V�&�����ah��Q�"On�07I��^%�ä�N6:!�"O�Ѐ1'ɍ56p�SËGXp8�"O�%s�(�Rp��@ڸ	p"O��y��Q���C�:!��)4"O�a:�-�) Ͷqa���*���0�"O������Xޕɒ%Z1
9����"O�!�b	��E��"�� [��"O x�ŉN�Q=�Q�������"OH�[#�=J�x��Ҧ�mT�dg"O�):b�"wH�ዡdYC�p!"On�j��=fY�c�ޘ�J�"O4���
��
�.d��O�w霼H"O~aY����Q��u�ICظ�Z4"O\e8B@ȃ/s���WC�� �r"OB�[�	��Y�����`Ś=�� #�"O�U�R�
TD0��D"�A�"O�ma�oÄq�x5 ��
�Uz��@"O�R��U�?�A��L%�D��"O*�I0�^�g��`�bc��.&0,R�"O��!����pb��/U�j��'"O�ZW@6h(��������c"ON��Ɵ�s\Jh7�	�xs"O��V�L�pl^|�@lB:p\��*�"ON�#R���a��@�AK[�bƬ:�"O`��@��K��U�+�U\�9��"OR�(S!�
bRlyi��U|����"OF�2��A��B��ܳ
��T"O��9��
��0�ٔ#���ȵ"Oj%���&P�PH��g�@�$"O�c�+_w� #��R��ђr"Of�j�Kӳ%(��
2��Y�~��5"O�|`�B��)��C�@�D��"O�Mip&q#�"�:����"O����N4�yJ�(�7iTr�"OB��� Ǘ tp(�#�l�)v"O���g� pȉq�,����qr"O,�U�ܓL �ЕM��*��xJ"O������e��Q���2�Mje"O�-*���w0dQժ�#,���"O lڡ��T�̡X�	�}�DiC�"O�1�'�S_��T�r`U"O�- %�.-H�׻��a��"O���&�?}�h}����^]�I�4"Oԡ:��_&Ji����Q���%"O��;�(U?I���BA�EBI� "O���F��(�b��1a���+�"O�m�E���6����BJ���t��"OT�z�O�7T0|���Q
G�D:"O��t��IWT�#gBM1,��y�"O���H��<d����[��P��"O�@)�(I|����&T8RR�Ѩ0"O�Q	 �K _�X�cs�'VR<SD"O2�#sbFl6� ��[?J��;�"O&�J�@�%L1C���BJ�M��"Ob�е�
Zy�	S�G\C��ȕ"O� �痏L�P<h a��{/q2�"O�0p���4)r`���h��"�"O��ۧ��_�H�tdӳB�J1��"Ot���_:{B`�2Ƅ]%D���"O� P�{��@�/���SgV�k��U� "O�iyԡ9�����F�/3�V �7"O(��EA�mL����$X-�n̪�"O��b2A�M;�<؇�^V5D��"OD�@�gH y��7 4z��7"O�UˤHÄL`x"K�3'م"O�=�o �@K$��` �"-�&-�"O©�)���
A<�^Ј��&`!���l�����F�Vp4eA�0!��(@����I	�|�2��ݢf!�>����(�~�b10�L:]3!�D�w�Tq�L>�lp�B��!�dS�T3E9 !�:�����$rm!��N�D�(���B�0����5�5{!�$����Y��B�)��I#m!��I��
����	����	3q!�D�Ut��$A+�E(a��;m\!��	����N"��X��ۅzW!�D=�,CNK�pj���5WF!�%1~��+;r���(���DC�f�):t�"�DE�jJ�[��P���(�5!��]�O��L�Ȝ|�4���-�dJ!��%=S�� ��+����,�f�!�D���ձ��TH�m@S�H3I��yE{���'x��QTn��3S�ֆ'���:�'d)����t�*��@)ւ��'ϊ��$!ݣvB=J�E�������'j��#����U���dX���']�8q�έ 8��G
	S�<��.<O��ؠ��'3*Ju1��j�L=e"OF�0��$֚�S7�P>C�qAp"O>�[*�V2֨(p-��<j�\2 O�����DK\z��+���P��%�$(�O��*т��T�R��kף5J* [�
O�7������`��!�CVd@�R���_!B���&囨�P�ʅ
`0">9����'ߪ��2ρ�,�`��i!򤄯<�$<0cB�3�J�� �N�!�C��hA� sq�Pp���e�ў�n~�O5�H�A\�+g�uC��e��!�ʓ\�����T6Eތ��%J�%��d"���s��rP&�
n.� �#�5 f�@�0D� ا� �$H�e�aM�]�,��e2�K�{�O,-�!��;��B��J?�)�'���+��W�&8��aZ'P��P�}2�.LO8eh�dDe��rTM�
^�VS"O4��a"�d�^4�e�Y"��,��P�؇��� 
��Gj�>Z�*�1R,�3ޡ� �<�ƍr���U�����5^�~�X��Y$�M
X>v��N�*��&o5ړ�0<	Ҫ����) ��7Mty��NP��'����L4���Y .Y�q���C�&D�<H�P�ݓ�jճ�NE�W�/�$�<1�4����};��\�x�r
ޛP�zT d"O��`$'��'�a�D����H���]���O�=�O�Mˡ'�oI��XV���p%�a��'�8,q��GJ������5aT0���HO�M� �P#?���3�l��`����"OlԺ���6,�1؄Ih(�"O�!#�C�Ʈ�J�*�f/��Z7"O2��������� �J�Z���	�"O��Z�琤�%��j��x��l[��'3剻j�ĈST#ͩe�F	 Cmդ-R<��$2}�C��y���6b�H�Ɖ���V��ē�hO��� ����	]@��֎�(�lL���'�qO軤m�.C�� �5.̈́a��a���IdX��C��L�P�,�	`�ګ@�v�I�*�O�OPI��P�v�,@kd#	$9�.,�r"Od���L�\hD�r��jL ��"Oq��d��!�e
��Xd|m�P"Or)�7��ST"}�o��d'��3 "O�)Tދ;�(����*VE`"O�\"ТD�YՂ ���Yʈ�@"O��Q��3fT$�ϒ*a���0��?�S�'*�9� !s`p�jVn��	]Ԁ�ȓ"Hm�`@(Ql�� ��~||ȅ�I[�I� �i�*Z���� �O@B䉞M�fh5�P�oa�������e�"<9.O��=q�e^1Z��݀�)�2O�x��Yt�<���?�n�I�T!j�$��p+�r�<�Ռ���I�Tc���z�c�o�A��	����L]�D� �S��6&JC�#6LE��JT
��h�%��"-|,C�I"Ap�k���q�BT;G$װB�*��D��P@�J�'	�T����@�Wp1���$D���"P�E/�1�o�Q!�I��i$D����	ʐ��2�"z�� P^���x�kG�6m>D�fi0D���!P��p=Q�U5&fQЄa��>�1���P;y�!�䈈~�6!�t�$5nx���7�Oz�Fz�O3�$�;FzX��b�9
�����8�!�$�1�4dsp
�#�,�p�I��!��S+r�ȩB�TqU�gm�i�!��|�0��&U�\���[� Dm�Ⴁ�,D�������m�n�*@aɖ:�-�?OFa��dF/�N�Co�84�dRGK�i�!��&��kEΝh.~���C P}�'�ўb?i�w���Is��S*^�>ؖTS��+D����/i�2���W�$sa'D�(A�كA%4i��ț�?�j��P� �On�T��u��׆
K����&��, ��d7�S�T�]�ĻCm�����B �5�y"dߧZ��D�����D�n���y"���1���7'iҀ�]�yb!�sW�` ��d��B�L���yB�7\�L��&nI�r�i�������9�$p�>�'"�I��W�d�7�E�F3�y�'����!�q&��,�!Kvq�}R�'�y�SbJ-�{6�ݷɎ����dt���'2�����#~v�\ &K�7�hc&�-�S��?ٱ`T=:i� Ju󰩡vsX� Gy҃B<W*V�!וtF���%[��y�!���"N g�`���y�J��-�8d�%�M|(uZ%�6�yb���lѢ���B<|���K��hOz��)
�0bR�ä������C Aѳ@�!�d	%}�p� )�*3*=ztoM����`��	���!U�"5}J8x"���D}�C�x��{r�O/C6܀��ľ/;�C��>[�
���
ߔ6�.����@�{��?��I�H�n��1����uOשOm!��y�\4���\�j�v��&O:[!�$a$e4`
�U���:5N��	q�O�=%>�Q�]&oqt칶d��V!�	���-�$"�O"I2�C�@��3��D��<;P�i�ў"~nZ2
Q�MK���?eL�`� ��B�	�F�x���,z)pi{�JD@C�I�7��X���"r�@IQ���^�f�=�	�g�? ,L9p�E�;�R��� �""O����l� o��a�I`��z "O�8����(i��RR� @L�Ń�"O����)9;4˰BV�0U��"O���/U��6D �����F"Ot����X�l'�U1`w����g"Oh1���Ŗ7��I��3k�4=��"OUݡ4� A���81&uZW"ObX�Q(�Hc�� �� e����4"O�qpФJ��.��"��4�b�Q"O�Y;��,P��̱gb�8�h��w"OHy5Eڰy��Y�cG,�H�(*O 
wk�k��ⰌU�<!�c
�'�*My�f�D�ЩH��V�4��x�'@ؓ�U�n�ixF �&9�ы�'�N��Bn�{������ٛ%f�@z�'ĲM�1� +#�BУ�n�
��p��'|�p�3�><�:@&�ʐ|����'��!���p���P%G�3
�@�'����V`:E�ހ�T.��ͼ#	�'G�#wg�vt{dƄ� �N��'�q��"�,����tˋ�xtZD��'���U�A�x�(�Ǐ��!���R�'�~T5$M%PAB�D��#����'=xꄦ�d��f�%K�n���'"��%]�Z��kƇ�Bk	�'��*�%�<\�iF�R3����'���DRg�n,2�kR.,T`P�
�'y��3��ijx}Y�b�V��x
�'~���
�1F��K6=,�]��'�Vq�#)ǎϊ!�WF�=��A�'Ŗ�ے��0�`1�d���8P��k�'��TJeI)Y/]�� ڮ.�f�!�'���K�+X�4�����,"O�i��'
 T@�C�xŊhk�h� Ww���'��Hj�ۦ8�������T&��k�'�"}�5d���n��,��S$9z�'���@��*�b�{'M��R�
`��'X�H�R,���J(��M0sj�q	�'�V��4!�S�q�� ��ѩ�'9>�4�ӳ"~�8�$�/J����'~=���R��xt��M�L��'��u*�m �
�tS4oɻEC`$�'4�Y�JؗJ�����
~NX{�'K���э�!lX賷�[/���p�'�Z�0��[T��G������'���K��<x���%��yU��i
�'=��_�s��}p��^4J�ޜ�	�'{�iqWÃ�{Y�����M#:D9	�'�X Re�c`��ڪ*�0�hW+1D�d ��
$"���`�Y�^��,!D�4���[9�6d�0B��E��S�;D���7���$M@lK6k�waP���6D��HBeQ�(���#&}�:��c.D��a�۫�u�@�nI��+ D�� $����E)eb�j�ڹ١<D���͗&Q�Bic�AR�ߘy�E�9D��3P�O*}�X������ݓb7D��{���N`�틒ȗ��J��5I9D��$��29lz��E���(<ӣE9D�@��+��V
$��#K6���4D�����jL��!�P�(,q�P�<i�@BILj& [%=ڠ�S�^�<���p��й�l��!o�!�(`�<� (	�ȚI��ti�'�>r?���"O��ـȉ7&J�S7M�)& �"O��3׆O!��p��E�K��[3"O����R�p| �Gؙ(R]g"O���a�ahXYCeΓ1@�q��"O��gA�GDļJ��A5��""O�`#�Cܖ+��	�| �Hv"OR�(��8��us��G�
�"�"Or��vEݦN�9��ܢU���:�"O�!B��;g�e�u�B�6���#"O�-�ա��|����t��� s"O��*� �`������kw��(�"Ot҇��M��p��]-GaĤ"O���@�J,D5��I�IJ0!k��Ñ"O���'�Hh��(c�4�!e"OB�#�,S�(���a8_�� ��"O���*�3}:�C���x�l�k�"O���_ � +����X���*�"O"��c�\�_t���@�&��\�"O��j�q��Y�q!T��GA?D����'Ո0��Щ@�Mf^�*�e>D�d�7�/�Z,�sْS�,��0D���f�)��{a��C��x���/D�|�@,ò<�Ś7̘tf�x�'�*D��UiD�+��R����ƐH6,D�x� �Bn[�5qRa6~��p�'D�DP��΁k$���Ք���B ?D���p�
�MR�h�5NE�Ay��	c�=D��Q�N׀J��X�P�@�Z�Q��/D��E!��@yT�&��1"c�����,D��4�"0�R��6;�R�V$D��q�U{��*��nhX�Q�G"D��h��չd>�\�)ʴM��dm.D��seҤ>��E�A��n;���'g+D���ת	=je��"˕'A�|X��&D���L|W�@��fK�RFk%�$� mZkFl�W��↌jd���C�=V��)⢁\t�H
�jǞ���q%��#/��sӱ�r"��<kڹ" 董H-b�-��y��`S�@���-��,�  ��?��uX^����/�Iڸ'xa!ּ;�❉��Z�K2^!Z
�3��L�"醪FO���N�X�r֨A
P���:�iL4v$qO\�ӓ5m�R�[ "��M�sH� &ɠ��=1/f�b�Q��P� �>�y А��D�É����e��B��0!��
�����Z#\�������}:�|�!k�K��%�U�O����O�:����>?��U�Z&T'"�@��(z^B�IG;�%�d��M=X6C�#�F?�9�����J!pv�c̓Hc�Ds�K��ݻ��ϔiyx��o*LO����g��9�ꤩ�%2\1<}Z��P<�j4/�D �����>c����'l����HƮ�ŀ�nɟCn>S�y������sa��� ��/1����@�TI�t�cC�	0]�T�p�	�y�,\�U��*+ƃ8,<p�s�6n��53Ua�W�l(���'�hu��OzN�����*F!\e!!�U���Rf�+f�!�d�M�.�9dD�Fb<��@��B*"-���6M\�)����Hc��1����-$*�S��MYR�C�a4#az¨ɧ/!艫p`�>b�8����K�
<�T�Үb@�w��}�1OH ��E�����w�\ @�D�����<I���- ����O�x�8x��HΏ `���G�Y}����'�*Qz섇�E�ک�w���`�COW�zT�b��~��t �'�v?��@�?2��~�'���q�+��!�t�&i�0�1�'���Ё�Ps.�"�Ua��xN�lJ0Eg,`�^��{IVp�K������%`8���р�D9��I_u-2�b�)%�Lu1������t,�^V2���`1˸'�T���ɯq�|y�.o<\)�3��F%��a��!^�$���)$߀ 
E!�G�>�[ԉӘK2p�"O�M�&l�0"�rx��+d��A���l��+b�4�����0$D�!&�7P�@��P t��ȓ
*��ʥb=d��c�N�����'�"=E�D�P( �luP���87�l��U:�yB��'Mˤ��2�S`�HZ'�I��'�{B�
�MҬ��f�]��Y�UbB��yb�ֹ ��36a��T�:�X�KT��y�I%����B��Z�z̒�e޽�y"&Ua�0Rc�Vi������y2�ݕT��(� �Y�Cp���݌�y��u�ja)։@��Spʖ��yB�F�>��|A7.ٔ(`�RGZ��y�dPy׊|�40B�bA��yBHL� �R���y�n�K�	��y�_�Q���-��D{P��y҇=NQ�2͗f$yg+��y���jF�Qs�!]� q"E�"��y�T�#r�5+��u*�@��Z��y���G�%��&�zvD-P#韊�y�� Kld��ϙ9�,�yB��;�yrd׺g��@��g��7�(�A���y"l�,i�	��II�!� ��i���yҤ�2f[��.ȸTyj1hY��y�G�Y >T�\�@��8'��<�y2�΋U�=F�T"H����vK�7�yb����%�"I"V��DC�-�y⣗B��a9�Z���Ͳ�y���|X�N�(4,�ã���y�]�0�l�$d@
E�:#�1�y� ]_���G� 89RLb� ڗ�y"���#�T@��C϶���#o��yLڧq��1*B�.8��K��y¨�O�6u�DUax�0Pd���y�h�)D�)f�ƧNR�IB ���ybi�e'��1��PB��'�P��y )�x����6Sm ɺ�+̽�y2n�:���A4��O~V�t�o��B��أ���?E�P$�<LT�ȓ�*�P3@�L����.CTADĄȓP`�(@�ނE$���
�,*��E���H%�X�V��$��0|��ȓ[E���!h�9PI޴"0f�2~ d��m�@��T���m/��s��ƮN�t���y��);�T���S#��T�n1�ȓnt
���u��X+�g�R�N���E�δ�J�GC8�g퇈WM��ȓsS��i���Fff�:��,�����
��F�=}�*�*;[̅�ȓ!��A)b �4ON8�̖�"�~p���Ƽb�ޑ ���!�!+.�X�ȓ@z���߼DgZ8��O(���Ԑ #��e��e���� �>���2���+Q2��ZW▉a�0݅�z[)��ΛQɮ�3uFX"���ȓ`�Ȍ��#�] p�f��#����Z2.h�C�	8����Y�~��9�ȓ唤��T�|��9Հ�gǰA��#?&1���y�(aY6/O!OT]�ȓC��9q�C�:����J�����/������S�	����.@�$��L�ȓl��}�ti�2a�W��Cn	�ȓ��@�t�=�ȅwd�ȅ�T 4a��Z�*'@�;�
�	r��܅�S�? �@�#
¶[��� ��Pz�"Op�����.6<(i�����"O�h�S�Vi/z�bd��6|�Tkc"O��t�K�!N%z� _���$a"O�pC�@Y�7"�B/[�T�[�"O��b��K�0�Aqٕ|d\�ST"O^�Ɂ�ox�D+�0cH`�[g"O.dɗJ�i�)���z%�lKT"O���$�*�`���fFO@��"Oh���O�}ՄY*b�Z�tX1�p"O��"�]0H�:]s�j^�q���"O�i�D�J�Tpp̺(��5��"O�t�
X�E�Rg��nۤ4�`"O���/�.&'�(Q��+�2��f"O , � �<`6��bD�\�]�:�*"O	���DB|0�b�s���-�!�"��+AL��x����%лoc!�DYUL48CcJ,�b\[���  ]!���?��R�FV�#��5PoV�VI!�� /_�
X`���`���ِ!�^ &~�0��E	zc8 01��@!��Y�o���ই����z�$�!�4;�~�G���3(*����ښ�!�N��r!�C�q8	4Iԙ6h!�W=��;��к��
�
ϥB!�䔑W4�����P5���G�*6!�T|���#��!|��tH���-!��&U�B�@���##����.C��!� �p����`��`,!+�����!��Y+
|��)4l��Z�`AN�%(�!�$�$����5��%�d��mWp!�L1�$U���x�)�ܢ+g!�B�v+���#Z:^�xB�ڽZ�!�����6}YV�ȅ,V�r4
�"OLL���7!���Kb�9s/����"O���)U�����J�>n�h	P"O�lfI�-W�h2�.T.sºl�5"OB r�xBH�Gn=*.��"O�Y�E�@��d��*+�`�"O��X0(���
��\�re��"OJ���Â\,~�{���V�D���"O�l)�.S{b-։ڳl�~Lr�"O*D�p���{֢u$��0���zu"O6*���x��E�یK��,"O�Q"�:ێ��pb�
,�xI�e"O<+�m���@d�A6Wbꌘ�"O�6'�� �N�
��-��XZ�4D�l{#�*<(ɠsR�Ԁ�-3D�Xؕ��7�����i�C�&- 0D����K]�D�A��ʦ�&(��2D�4�g�ه0�&��VC	PM��@3D�XA��r���I�m�0��%��n3D��R�S�L\N,�P��x��aK%�:D��i#��J��Y%�%r#h)��$7D�������y;"�ױV�]à�+D�0��"nR)�#���v�1R�*D�	R�Z+�T�CF��{\�JR�=D���Q�J#H�&���1�@�yR U&NE,Z |�L��.ۻ�y� ���!�B�i�D�a"��y",��3��[�)�c:Ͱ�ʅ�ybE	�$����3�P:Q֎�s���y2�H�f����]I��l:0�,�y��:=C���f��!>��XY�����y
� \A���ΰw���,M|���"O��a�i˖vz0�D�W;����5"O�	3c���kf��5R��0V"OhZ���-/�Re�d���N���"O�,���S��$�P�6Փ�"O�չEOB*$W�{V��i��"O(�q�_�B s@��>�� E"O�I���3Wf�K��\�0�B0��"O�0�g�L$�A"ǂ�B�Ɲ� "Ob�/[��5���,X�B���"O�E[��w��Ȣ��
�fP�"O��*�d4�Rk)�]��D�5�y�B]�R%�1`���Xr����y��ءj��P����\�.�cA��+�y�#>����bH�X)�����yj��"!$������K�	�`�M��y�eD'���H�L�6wA0�� ���y��֞e~��P��B�`�D�3�`X��y�%X�~���#��b�ֵi�/��yRoڔE�f�	��#]�z��F�]��y�Lq�
`g�ʻV����VH��y�O%,P"[�'��2:�D�P�D9�yr��U�*T3�1��!�P��y�����5�ˈs��(B��F9�y� �"e�L�h��O�ZuɀJɖ�y���|�^=�7�$^:H�fY�y�K>L�)��_�C����@��y��F�IR�)SƬV�e*�=iG㊊�y�`�'CZ2��霾N�z\9VB��y"�^�e$r�+�ű'�YX�J�3�yRh0� ЊB�. c�D��G���yZU��3��TGy�PC� ]P�B��@{�a����HiC�"D�DiRUI�;P�ޔ�CCN/w*C䉓-n̉@MPgM����i�V$C��!����٩@`�:��^J�^C�I�tK��q5o�&>n�p��TeNB��]�bqIR��4.Xh0���
B��&]&ޱ9 ��4����,C�$C�	?N" �q2��-%8QrV!;`�pC�y��Y�g/M4m%�A �V\�C�ɄDS"m�5��g��ub�JF�8H�C䉺*�v�B�FI��:�£ʄ$��C�� tI��|QZtV��>��C�ɐq�<�PVj�!MR6H ��k.�C�I�J������(_/:� ��)a_�C�	��@��7�Y�:�D�*�V
�C�I5����3Gӷ~�R�GfC��6C䉫!S�X�����:&9I�$
���B�	 ���ѩ�+��r�$K��B�ɒK� �����0�.��u-��>��B䉉	͔9z�ĝ�.���3e鉮�hB�IuD��s�҂r�ЛeLD�%�^B�ɲj���0���#섢0�B�I������ �����H܃�C�I� s�
1Z)􌹑��*[�DC䉬r��y[��tt�{�ϡ�zC�	#9� �▢Z�y+Qh���$C䉤>�p��RK<��u��0�C��!rUֹZ�dI�!���3*-<C�I��� �̛�]h��B�L_~��B�	<c�z�yp͆���ܠ�b�qB��$��E�5�ւ^ ��S�C��(O�X��B9���V��- (�C�)� l�c�D@�y��@�SwD|ya"O�`��E�W�N@���N�jU�1��"O
���ީ n�����22��i "O�̩c�I�,|DH҇�L� z܀U"O2�Qr�8��5�wd��~��@�d"OЈɀE�+9H2���|�n)�"Of�I������5J���^g 4�"O��B�鄷ļq3Gg6|Y68R0"OV��`���
�֑8&HO#']"u��"O�5�'C��mX-�v��Oӌq�s"O0�b�h�H�p�'���^���"O����V�@�)�sØ�0����1"O|���P��2`����GR�A�"OԹ���'�1�Gʰ-�hq�"OM�ҫ̏mB(y��P&u0�%E"O������,�*�08���c"O��".�d�f��/n<$���"Ol�I�=\�
]#BF�f��q"OR����/|��Kb�� ��4�4"O|��Ԩ,6TM�D��
:�ȕ��"OfU����|wjE�4 @�u�*��"O����+����5(��F5zaP�JR"O�I2v"G{��d
s�0gj��"O��QA�CSt+�nBaG|��"OPJQL;Z�
�����).�Q�"O��ڶ���:iTd��B9J�k�"Oz�Ҷ�Y�&����0.�4@B"OB������T���-H�s䖜�"O�DH'lP(X�k�L]0=�f-��"O,y���0I���E�՜/A��z"OU�2�Z�|�2��Q�<a) "O��a��%Zx4(���	%:.��E"O�	P��ɓNZ��j� J ���"O���qhåb�6�f/�2Gh		"O:���+�B/0�9��3	J�pe"O&]#ƌR�]��M�!,J���"O���A��m����;
{X��#"OH��Ł�
g�L$���Y(,U����"O��Q�ΐ0w����09��A�"O`[r�?&[x�񂂠�N���"O0��0s�t���U|&`C�"Ov#���0�0h(G�L�FY#"O(��%���^���f�Ѿ'ֈ��f"O��"��on�U�T�N#L�p��"O�ayѦ>v�"=�ʔ�:��"O��H�:i��%�Oq�P�+�"O�����$���3�'m�ؕ "O
|�������0ׇ�:�8�bt"O����S(z� ��@Uu����R"O��Z�hZ�X��%�O m���"O���ŭ�1d?�!�c�X�d��a�"OrA�V�O�hw��� �L�\��PI�"O,B��O�f�4 p��,P��*T"OR����I~)�C��8}�4s"O^�ЁZ<Ҳ��5O����Y�"O:�Q.�oZE�g����%"O���$P�Aw�h{��\:T����"O�x�+L0� i�ˈ�K�F���"On�7Q��0P��1G�P��"O�y(�b:T�<�B���0n%<H��"OL�h�I0D�q�"��[5X�"�"O>�;���hA�#���&ε:"O�`�kOq����N��(��"O�5#�>',�h[V�N�7�)�"O� �PP�(н#̬ ��ϋ&<[�U�C"Oni��/= F��1-K�x���r"O�t�΂��P�&N�j�ɇ"O:��BN?��5S��V)g�$w"O���ӦF }:�D���T�ȣ"O��3#��uҙ�B��x�H�J�"O�����Զ<��Ga�(z��S"O�<JU3G�ƽ{��B7���"O.I&�K�X�]���k��j�"O$�����ԢуR�
0��R"O�M���x&����,�PiC�"O��r�C�-ΒaS#G3~�2<�d"O���#�	rm��C������$"Oj�`�L;;4*q�Fnͷ
���{!"O��ELĞd8� 	3�N�#Tq1@"OBI�DIc����B��W+̬8w"O��+�(�;G&`b�l�%S���C"OB�BDޑ:��i��I�z�����"O���'MҀ-�u��(P>��]K�"O���$J �\��gԔl�P��"On�w���oE�<
�^h�R��a"O:� ��>^4�%:e$J��V�{U"Ov���,
+p��Y���y�B��"Ol܃1CU ;T�x[`��_��5Xu"Of	%���!L6	âA��(�$�R�"O���(~w
\y&���Fj�Z�"O���7퓙'F,��`��rH�kr"O8)� �z%��/Ho>��c"O��ꔪS&T��Y�E�Y6d�C"O����#;6��b��_�i�p8�"O��� nG8v�#ei�2&�p�"O�I���<��[t"�.��V"O4����V���%e+��"O�*r��=f� �,�:葑c�-nz!�X�K�ti�dY
p�jhӔAR�!�ċ&t��ȟ��ہ`�84	!�&@T�	R��Z�@�H�Ư&\�!��B��6�(��, ����n�1�!��X�o%�b@�
�gg�X�!�D���%��XZ����iW�?KHK�'#�̐��ч�� *kެ6�f�S�'�~�0�oM![R!���4R<�Q��'w~���:wޤ�piN%RJ@���' � aSKƦ{��hKa�P�U}��#�'�p�P�!ΣYB����C+SL�#�'/�`�K��d��e��#<o���'�x��f�	S\��&E<Ж<I�'�����>
vt��Ϣ��T��'��6���	��yCd�R�F�Qj	�'Θ�
�Y6#���FѰyN��'(~���A�a�8� .�:}X�1�	�'CP�颇��!�����B0m�����$�.{�>���K�0�r����%Q�X�b�
��?��ɦ%��'�\�K��i4n� 7�!� �ɵs2[%F�)y�H�k��j,�)�'�jH `B�X�b��?F�͓'�%�)�=�|ʆ�.��Q�E��3�P�l�O�Q�"�I�9�y��b՚ބ��&�C��(O8���Ӊ0^�6-�*���Z�M0p�,b�`[�i��(�J���Ā ��}�O?���'�������(�8ȡ����&�����r��	D��(�~��c߳<lt�	.<!��9�W�'>ў�~"�&Ӏ���_5 Ԣ�����W�'_a��"=���ç�b,�dHgK��5(���~��O�?ͣ�H̒Ck�q��ڒj<���m����~�S��}� ��ʲ�\(�S"�5�}*�Nl?a���S=7pL Ig�Q�m:��Y���9����$�S�O���ծ����x1ʎ<
h�c���9���#�͜��#u׮%^B�q���+�/ �I-!� �S'���JP�G��g�OHTGz����T��^��現w&^��v��!���\��(O�>�p��ܡAx�1H�f���|�s��hӞ�3�����\��ʱi�!G�1�ɨ(���Gy��,�'QP�+X?L⤍9�*�?e� 0�SZ(���<�C�'���b>1���O�.v�<Ô�^�9�$p�m8?q��'r��$��f�q�&�|М˷� V�|l��	�5�� �9|��ΓZ>������|�*R-I�p|)��֎��	�"O����q��)���@y�; "O"��e$p��V'M�ž��F"O�� Un^�p"0hZ�Ǖ�
�M� "O2KpES�>���81,X4�J'"O�	*'�U�_{��S��$NB�K@"O�<�3�3L��X��(�̖�q�1"O����JU�`F�2N��Qx�"O� ���x�;���g�pX�"O�i�fm�B�����(Ēgh�3e"O���٢*��Z��50WL�A0"OB��f[�T˪��+0mQ���3"Ov��m��J�H0��
T�QGdp�"O��O����l0�J��H(�r"O^��b̓"w�!��Ʉ=+�e��"O6�b �
i�z�qc6R0�F"O�M��#j]�y�#E�WI��q�"Odl������J3bˉM=�Mɒ"O�9(�,K�P��4#��;�)HA"OV�ZY�_�(�Q�@V�2�9f"OR�[`��eπI�7@ն2􁨀"O.9�(gH��Q�A\�p�"O�8��5{��(��`U}���"O"�!u�t8���%I:E"Ob��RLћh���u��0���"O�y3s��Q�~��@W�\�@"O��`��_0/�h�'EP�3U2=��"O��I��婧I�INV�u"O8�C�$�H�p��:, v|�"O��+���������ƘK�"O�!1��O��@�qIX"�"O��Bs΄��,�[%�B�;v�X�"Oܥ�gl�hhH=��U(U"D"O��is�1dFI��cì-Z0M(�"O0��' E�}[�$�Z ���"O&	�m�5{�DƉo�^<��"OU���-'��r�Aj!@��!�d'vܽ*���W}�$��+Ȣ\�!��p��Bi�0/�|�r��]�!�$�ߴ�ab�Ϛx��
J��o�!���*+���S���-E ��$��f@!�D�A7��R�*�<^�"��E;!���8`%-�F�)�!S^�!�t��(��qή(��J�Mo!�D�9J�!1�/��`p)!&�o2!�dÚJ.�,P�m�3LHءi���5I�!�dD��ƌ��fφl,��%B!!���:I�����-Ƿ�����&�#!!���& �ꐶ>��yj���]3!��?�N]���W� ����i!�S>P��x�-S�AxИc��<x!�d�,F��ţc� =h'n�w��	P!�
|�}�cB.&����(P�~@!�� �!�SGWO���1c�Q�J�5��"O*U��Q��ЁSO�(eP��6"Oh�02#F�=�>U��/�;n���"O�M�⇅�Hv"h��o��-�ƭ	�"OZ��W�7K�h�@L�����u"Ob|3���V8����
��I4"O������ ��Y�J �c�P�"O�{B]�pM�d �h��GJ��0�"O(�"�ҤKR��:�e�1a�2��U"OHI�p�ށ�bR�J�f�NP��"O�s4.Ybd(L�Bi��k|��C"O��k�)'��0�AG6o�<<��"O�q�C�}�ص獚�YrzM��"O�Ԃ%IB.X��RA슥,p|샀"O�5�@ɘUt�e�T#q����"O������"0B@��Ej6�� @"ODLJNW.�5tHϡC�r0(�"OB쒲(���ihсM�F6'+D���a%Z<g
�(���#,A=��=D���5Ȁ�:\�|�q��&��zdI<D�D�C�Ux.^�:��W�Y���6D��0s)���i�Ԏ	�P�H�K��!D�܉b�4p�����;/@ر�;D�0���=O���Ss��ac�)X��9D�)2f[�e�jhr%��X��1�3D�Z``�7n���)ǥ\~v�6�2D�tC#떥7`ʰ�c͂H@z�g�0D����dӬR����A� dh9� 0D����	X�n�6���f�0���- D���3䆅B�ZHQ����ol:��%�:D�����X<�n�(Q�$1�+D��Aa�Bh�����=N�ZC�)D��y��O�jڦ��HO,%*�1d�5D�,�4k�3	2JI�#M��"1 Î5D��;AA��dCt����]�^-���7D��@�)��%:���z\�D6D���E�D�F|�oJ'd7:=K��)D�$�Ъ�d�ԝ�%�ɟ!$�"@)D���f�.�A��Y  �,q%D����) Q��"��E%1��QǇ!D��*� �f�Z����"��-+6?D�p#f�p$�RC��#0́�"D���Վ�-'&Z���Ր`��M[fL+D����&�i�F�#p�E
r�r�3Ǌ*D�4q����E���lm.d𙵬%D�H�"��|,h��cț�@)��s��"D�P*�+�(0բ��dϿ�$d#%�>D������|��hb
�:��2N0D��j�Yy�R� F9�ȕ�/D�c7F�}R¸�p�<��Y��N#D���pƊ/ic6jA�ZPWb"D�,��
�q��R��$~�$���?D�tq1��6�の�����y�1D��C4��G��ۖ��z���T�0D���woS�EŲ}@�<	�TaF,D�8�S��}�@D۵.��q���4D�0����?jG�U)f�ٵa8��h7*3D�`�!��5l�8��ₖ=@<�sÌ&D� 8��˚F��-��$G ��@�D�?D��2r�ؓ5`P�5��n
p\ASN D��
�ɚ�m��������:�@c)?D�� A�4�>	��EL1�4��qL;D�D��V�
8�$�	|((`K�o-D��bGc�+e~��2'gN�P�m*e"+D�� t���g�*Ɲ)�e¬.�����"O��ـ���.I�H@�D�2)�"O��q�L�Ƚp�"�������"O��V'�.Z'��p��,���I�"O� *���q.�\�e �̉�7"O��y�@+�ܩu#�
d�����"O֭����=b�ѣG�"r4u�D"O��J�!�A�fT��@T�X�y*�"OХP�@�&l\�86 ��DF0��u"Ox�i��Mc�p�yd�]:�R"OЅ�ǋ(� M�4�<����"O�Qq�kA=
��3�C�A�A��"O��j��:�z�'đ��j��"O�0#6둸���D�,?`)��"O���S�D� ���&8�r��"O
�rE��(D���@`��R���[`"OLx��C�f\�lu�	�f��T`D"O���d�<�j�*��]����"O ܒ���K4��T��4Mt��"O�����Q�#��8�eǂ�{8���D"O�h�Q�Ƥk`�����+���]n�<�v�lL���c�(f�t���Fs�<�P�рh)���&�Z�l<�"ep�<�Q �;��xr&� xL�qx���m�<��./0�� ��<��t��c�<i�N�<�^|j�@\l��k�<Qe�*75���
�U+���l�<!�nޥ5���u�Ҳ+S��j[@�<i�5l�)���9p�Pa�B|�<qi
HɠX�QA��q��=�R�JB�<ٵ��!�d�"��YR��HbELH�<Id.�� Ğ�{���+ ;*"�$[�<�PO�ņY3 W�<�ѱ@�R�<9����p��P6DV�K��uq$C�s�<����ru��u�F�P&��Y�<ѐ�
K�ԙX�)K��xz�!Yo�<T��%�����>����i�<���^9�჏ z-h��C�a�<����,:M�f�X�s_�q�f�a�<if#��?�Ȉ���i����dƝw�<Q���G�0;�[&=B��SJ[H�<a7g%�4("���h�f���eA�<�S�_�M]��HG̝�$��$ ��Vw�<��PA���PqJ�Y�0<;�^y�<a��A�8@���D#0ְ�`�s�<Y�Jrvpa�O��� ���X�<9�ʝ<`p���g��|��eN�<Fo��Z<�Ca��:���[s�u�<�B.Un��eh�1r���'t�<Q��ϯ�TE�լ��b{���Br�<�a��|�R�M��G��D+�c�U�<�T�2��i�@�����#�N�<9����O��8�D������DL�<��Dԃ�L�%�֕=�tkcC�N�<2�W3!��0����R��4
H�<т�
r��5�Fn�>���pr�ME�<!R���n6`�;*҂	�=P�)HJ�<р���4��O��q/��[�ĕC�<qdhQ1� ��ȡF�Xs��N�<�wm1f� ���^ ;���d�y�<�#j�%�n�[��Cg�l� d�J�<1g%P�{���I�N�4Df!0wg�I�<)�E�"�P�`!�M�LTyb�bVG�<Y�L��k����O�!h߲@:�.�A�<� )�b+S-kF ���@'|�(��"O��B��sdbV���Yx�=#�"Oh �E$��=��\B���D���"OJ�0�@Y���a�\�`��X"OP���*U([w^�"e�Ԙ
�8�#�"O��k'(�x ��g,A9���b�'[JP�����sP�דV�����'kv��Mu�T�bU�����'�x����:��<�"D�M�h�'�$����#3p0�y��ϮF���9�'-Fԉ��M�PNm�b#�70}�؀�'��5��n����iRnܾ¢�J�'x(Ů�;�XUoW�� �'g�9�ƃ��K��t�4�B��E+�'���۶h"��u��d]������'���� ��e=���� 7|�h	�'�d�s  ���   H  `  �  -   w+  �6  �A  XJ  W  5a  yg  �m  /t  sz  ��  ��  9�  |�  ��  �  E�  ��  ʲ  �  R�  ��  2�  ��  2�  ��  �  F�  ��  ��  u  Z � 7  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P�����hO?�ٳ�.J�j����XG@�ʂ�����5�O�k�`ܱ$ڀ�S6K���~���"ObL`�NӘx@�"iU�)��|ʒ�'
��+/�HM��휡*D�H1�Ͼ]x|C�	$To^�C2O
"����+8����� �tbX�Aԯ�'(Ԭ�� m��'����'\�_ͺ��I�$�Ry0BGP�m��K& �Ƹi��'��s�\i�sm�/,1�A���h�d$��o�o�������i�գ'�'v�4�yT&�'���U�����#��������c�f�<aP�'4�ΐ�A4@x�$�)(�Z��R�	�����l�@��2c���`���F�=	�y�gl��ʧ)��ջ7aҏ4�@�����)�&h�	$�HO?�S0/$o�񺖏�P��l�i�<����럜����fw �:VGNAtvl󤍿>��4��>�2M��-8����C^3����J��������s��l#&ǚ�tg����>�`��*O⤣�I\�,���u+��e����fmj�(�?Q��Ʌ�f���C�i#a���P�	�)�!��F9`��ʆl��h��0�7+Ԥ�!�۔l�<򢅄�j�&	ZQ�� q[���|Z�}
� H�+����M��8��l!c"O�5����2��ۆl+Fv�`�A]���Iy�80h��}��m����1Q(v��K؟�K�#�0euh0����$4��=�� (�IF�����ʌ6J؅���'D�w#�0pͼ�ɓ�Y)A��`�H���Z�<۷�R���0q	
�p�L!�!"D��2o�6u���hgO�9%QT��T�>D�lI�I?�$����/7lX��<D��j�&m{�@貍ŽP)T�䉥�����>�ɦ��(N�]p7LH�MR���D%�	����q�S7�$H��h�!B�C��?�
e���)�X8�"�@�	,�7-3�	�<E�ܴz��5�S 
(��'hE": lGzR�|r�'��P6�X�J�F��鹲�	*��ȓM>乻'�H�W�I��n\&.��I�	S�񟤤OX�	R�W��9A��(t.���A���C䉘%�2�@&`ɂN����'C�M�
�A����Ob�#���e��4�8Zs�d�a�'
�'=�����>�z������-�jh���:,O0Q�Îگh P�a��c;�SU�'�S��y*��~�2��(e��� �F�D�6�=E����p9ԩ�Kpv�㖜Fр��'����S�L����:6���A����0�7D�r!�ea�"+Q�z���A'��d"��1�)§a���b�n�@ŉ��P;$���In��w��|JP�L^F���b� ��<�J<����5}d��I8�}(�'ܨX�C�	�T�15�@�=&�i�gW�AS`C�I���
��4�j���`I0D&C�I� >x�6�Q#R�b\p�H�)_�C�IQdLr�"��-=����$S�Y)�C�	H�����U<�<h�Iˀ,&�C�ɰQ9�,��R�'G�4:���<t��C�H�W��_�A)���x�����'��>�	�Ru*!i��V�4`��L;<RB�ɒ/J4���L�H����e��-�R���O࣏}roZqw�y���F�<��q�
���;�O P�@��&p�bI��#�p�u��2�S�'U�h�b���b�8"���	�NA�?���~j�C�9:�p��6T$8KPԊ7J�}�<ٴ�S�7�@0��MU5'����ǯRp�<��Ίs\؉�7a��4�Ř"��o?�	��qC�L�8��{4&�-�����O���d@ӑ�N,�1;��*DE����<!�b<}[�f�I@�aܮV4&�)�)� èO��q��i�4v�\H�S�jy6�C�pQ�HG{*�]��FH�j����ޮ`��h�|��'5|"=�����u��ud�+d?�|b�%�=a�{2E\�8r�e��Z��2ꌟ�y2�6eH�a-H�\�`)������'oў���q��F��a����t�#j0�����&�y�$ ���1C�hQ�Q�
��=�P�)��8�6DW-q���i�q2�,���ɷ^�b���j}E0ŉЧφsD���	y���I^��[�/;�� �%̣t a~BL�>!� Y�pA�y����-0o�|�4�EF�<�LR�H[�諣&J3t����{�'m�?�*cL�"Bʡ1s����pEB��;D��Ri�y{�	0���̔�� L:O�=�!i�6�LsB�ּ<eD0�5��n�'�2����3D�0I2EM3�`�� �����nX��O�>�v@b��]����Y��#�(Vޟ G{��i�z�>� j�\�ꅻ�\=G��O���� �FA�w;�-	�^�A��|��V�d��ɇ:ܑaUb)^jv�U,�8ӨB�-9�н�R�]�d��Z���I'rB�"8Ӗ)")К��xơ�'̨B�I�>T�H�$:c���Ą�BG�#=!��T?Q"�K[�2����ȥ$M����>D�����,Q����%Ⱦ$�N��cJ ?q��i�����H��s��0�ZH�b�>D���Ѓ0iY0�A���6�(hJf�.D���2�ޝgWB�2%�u����M-D�pk+�$|v��`l�Q���2��+D�� d��0F�����A-AX́ے�6D�x6�E�0�F����87
���%�?D�0�:,rz�	���5���!D�p3��ؐG8jQrI	�X �Up  D��r�LA�'?��`�]Ɛ`q��c�@��I�|�!`C�T_�4�f��*"~�C�ɗF�\1rCZDإ"���()�C�I� �`r�얍�8��hՃ"MУ<1��T>x�#E��1�dO݇U�JH��:D��qu͘Wŀ�b���% �M��,D��1�Ao���M&}��x6�*D�t����NL�{!��
�q"2�&D����!�{�r����)d��9c�%D��J3��?�2l��mQ8J�\H� #D�$b���7tP��w��h6>D���o��{���2�np��=D���b [�QZ���~��[��%D����%�O���p�@��fՐ��(D��2�d\$z�XP�w�X+L��l �L'D�� �N4RF�r�Wbr��� &D�Њ��%(��*@JSG�\��a.D� �#� (���G� c\p���*D�Q��^2I������Q-�92ր;D����Vl��aO�&Ŋ@�SJ$D�<���Q�b+�� ϗ�6���"�.D�����Q�t1/X l�����-D�ۄ����H��	�q��M��(!D��0�@��"��0���	c�����?D��dC!mb�<8��@�"�tM�f�*D����I�n�H�7eݶ~Xl��T�)D�8�R���.pl��ׅGdQ��2D�|ж��b4M�0�����A#D��2���8:��Ȩ֪%/_ 	��)#D�̉"o�/���3��8r��k�6D�<D�:��(+�+	i������5D����e�
~$�18�OYB��PGG6D�h8�$p���H��h�$3D�hIb��?H���ʖf5l��m1Uc3D���v I�(;�<����3��yh�H.D���쎥 4@:!@�;�.8i�!)D�A!�p�Y�ТٵҲ� "-!�d�_�����MfM�|0�PW!�Dͮ
�<)��m�6��s�c�>�!�D�Q5�V�l�^4������!�����i� lE6�
����!�䖀pt-�4�R5')����ʀN!�d\��4ɚ'y� ���OL!��]�N���Z�DёE�8��E�`!򄊔M���XK�u��p@��E!��o:��3'� � ���i��ڣ3>!��ʚ0t��5�װq��%��Eک?!򤌡6ZЄ��i� >(8x5%U�g�!���XiV��S� ��ۧwq!�� �a Q��,�%���N�+��@�"OX�Ic�]�q,�M�@N9x�$`Hq"O@��$�6W��1����T�x}9v"O4�@�f� j1��B�@���97"ODe
��]�M
��R0(�4i��t�'cb�'���' b�'��'x��'nr��p�X2@�@m����/
B���'���'�"�'�r�'�R�'}��'�>e��մw$r��G�+|�p�٢�'(R�'P��'1B�'(��'�B�'SX�S�B�!�6�ڻ�lRF�'�R�'���'���'��'�R�'Ɋ�['k��=	H5#W�M�G<8T8S�'D��'�b�'m2�'d��'��'�B�P��˚!���h%��bP9z��'���'�b�'��'��'B�'����`E�^��+R�WWd�S��'�b�'�b�'w�'���'\B�'�:�E%�4AR�q��EB=zX:#�'y��'���'��'��'��'`UC���00 f�F�h!
��G�'���'�B�'p��'b�'���'=<	���)K�D	�� �wĄ�'u��'�'��'���'���'{:3bg@;UG�)�mX
y�꼒��'I��'���'���'q��'�r�'GJ���k��AȜt@�Ye�]{t�'�R�'��'0b�'�b�'o��'����b떈�<7��@��(%�'���'��'U��'m��d�P�d�O$�	S�?��A��ڊYJ̊��By�'*�)�3?Ѳiv����%�
�T�;�����.\`b$��������?��<1�i�� �#�$sra�J�La#bo���DF&T����5O����qGĒ��\�s��ɋg��p���Ɠ	l��vh�<o�b����\y��S�@k�2$C�+��}�V"�gd���4xCzl�<a��$�a��F2S� �cP*Epъmr�j-2�!o��M�'��)�S�"���e`���֏-j��D��fջo�DY0�Dg�x�vBJn`���vK�E���d�'K���W$�; $�qNM2Z���'D�Ix�ɛ�M� [̓,o�A�(�V�6daB�U�X�v�Ê2g�>��im�7-k���'n�E��r�Vy�$m�`;����Op��5镋g�\x#���b�P`���O�`��̭^K ��'� #_oQ��<�(O��s��k�	^�r��
�����p��e���ߴOA|x�'9�6M&�i>�qwfƮN��� -�#T���}���4<���'@n�q�����dԁA��$�v�:3T�r�U�Y�Js(Q��@Um%��|J-OR����hdɘ�}�9���av������ڴb\z��<	��t'��4��� �>?���eޠ0���I���/lӐ�r��?u��#0L��Ĥ��]ʕ�A"k�$�NL(�cF��'^�u"�xbBa2}�/?i0��"������k2�y�F�:�?!*O�˓��~,�����y򬖢N���hT,H]�AV�1�y�Lp���s�tRشzכ��'� ��&�N=x�H�#���\�����L�uD��˙'�Rn�5k�0�aEE)�����8I��p�$0c�N�w;�l{W��P��ϓ�?q/O@�S�O (-�7��A=6����q�8Iӎy�awӺqb�����ڴ��_n���&±H�������N躥R�'o��7�MC��i�҂�6u����']R���@E�7�f`�X�X��h���m�B|q��i>�'m��A�&�l!�G��(z&��=�yr�|�lgӔ4x��d�|�Q��VD ��G�{�z�:���S~��>9��i�H7w�\%>���2��|Qw��wRу��Δ-�n )���� ]� �O����"@�q�a�!@��t���s#H2�lӆj��5B��-d92���+]�^���%�*I�J�Õ$MwR�rnؐ/2Z}37�	; q�Q�6C�w��aA��1���R���.5R��G�I�\����0:��� ��{J6�s���)�!�1N�?r�8�@E��i��A�����AZB<0v��6qlAx�K�%F��4Ʀ�U{p�w��qR}"Eg+B+�]z���f�V��Ƣ�,DX����ݢ]���]B�˧b�rI0�Srb�R�����ۄ.�����2���
�@�aH@$�@�I؟�$�D�	؟@+�R.V^,s�
�Pv�K�B͵x���	̟��I���	��Iߟ��#���M��ꜹ:�ce�'b�4��1�X\8�I؟��	J�	Xyb�۪��$���gֽb&$cᗋO�>(��OZ�d�O�d�<�[J8�xL|갊�7������'m�pA�-ԛ��'�'%�	�+j�c�̚���t� "@��5y�%�`y�����O*˓�P� U����'9���̡�B-+��H�I�������"D�Ob�^*��Dx��֌�!���)j����ֽ
�(���i6�I	,�e+�4D[�Sԟ�S���B��*�-y��9�cL�eΤQ�4��$E�,7�b?�w�	:(�i��;�@�35`kӒ)BT��ŦY����I�?5�H<��&����d��2�i�����2L�$�if �������22m�LW\QQDũ3���(��^�MC��?)�i���˵�xb�'���O�Ii5�@+rmq��J ��Ke�$E;�1O.���O���Ռ~G��#"���|A�aD�RAb\o���4��h{	nZȟ����������	��D�rk��`��a,�(>�*�����>qBML�<���?q���?���?I��-�����5�6tF��:t�h���J2���'5�'P�C�~R.O��d�L�? �PŞ:�ʰ�aƀ�o��Li��<���?)���?����iCa\
umڄ*L�M��X!t.�DJY4~���4�?y��?	��?�.O6��P���iA^m�w&A�(�lD+T���耮O����Ox�d�O���E�9rnZ����I�~�|��@� .}�#)K�@�P}��4�?���?�)O~���	4��I�O:�I=[g�ٓ�2n���HWG�.j�>6�O����O��� 5��oZ���	ߟ��ӝt�p�"�48l����<5|ZU�ݴ�?y)O��HTZ�i�O���|n�-�.X�B�R�@���U&�s��6��Oj��Җx�F)l����Iϟd���?}�Ɍ�DQ�9B|��!�A8uXӯO��dԦ/���:�4���O�Hj�)��@��{��g�~$�۴#p����i���'���O��T�'���'��LK���Q-Ĭ �وrLXׯn����V��O����<�'��'�?Q�K��%����\�1	��9k���'�R�'�=i�m�R���O8���O6�����a��*#�( �!m��,h��iI�'������)�OX���O�DYѧ¼5���
3d�c���I%���y��0��L��4�?���?���3��C?q'�5<�%���$��zF͟C}R#N�y��'�B�'��'��q�MzӃ�0���*��E1��M��M����?Y��?��V?�'b��$�d�6*�4?-�$������у�'�����	韘�	˟L�/F�M#w ŷ^T
��B�E�d<vm�<`j���'U��'��'��	֟�TCy>բ2�J� 	�4�QlP�6��F��M{��?Y��?i��?	�B�Hn�F�'eb*��( �IQo�y��)��[6Pu�7-�O����Ol��?Ѵ!�|����~2f�79�\�;!,I �Ւf��!�M����?��?���q�6�'��'���L�!5�Fyȕ�I:�ո��W#�z7��O���?�Dk��|z��?�D\�|n����I�	C"H���3kPQ�J7m�<�2��5��V��~����5��T�M�0
O���ڦp�p"t�sӠ���AFx��C,~ ��C�g���b�M��Mc�Z�z�6��u�4�?����'h�Kq�XS��%~�@*Z��ŷiYn-j���⟸Q�&1�l�i��J��yD$�:�MC���?���^q��1�x�'=2�O������2㚱�H��p�js��B�1O:���O��d[��mk���D?p�I���/�Ao����2!����?�������@¿ �^l{��Ne���'j}�#ޱ��'7�'=�T��	0�X<5�$(Zw����Ċ2@ðe@�"Y��ē�?��������\r�$�0- AO5ᑃ�rs>H����OL���O ����=�&]w�:n�y��@`.j@[���	ǟ�$���'<"$ҬOL��*϶c�����ŠFH1s5U���Iɟ��ky��D�{�����jT!ֿ`3t��7���h�\�P�UϦ���F�Ijy�C����'rt������Q��T�φ #���ܴ�?����d��l��X%>���?�-�4 R3!œW$��!2BV+����m���v�i�cǞk� #�@Ԑf"X�n~y%�  �6MAn���'���l(?���%�РZ����~��UȈ榱�'g�ڌ��iռgf���dۧ5��Y[� 5G��f�ݝ
�6M�O����O��IS�if�AC��3�8�C�Iη^6����ih$�����Sӟ�V�
v�����=~��f���M����?	��2RR!�#���O����XuZ4�q)�#Q^8(횞G2�c�tJ�!2��П��Iݟ�i����ƌ2��K���l�"�M���/�E	����O�OkLє��p�#+�/��w��8�	�O�,b����͟d��|y���*.p�R���
�!��}��p!�"�	�'��'��A��D�%�$U���:K��I�nʔ��'U�'T"Z�|���L ����>	�1��Iʽ50`�Ҳ�[1�ē�?����<���Bh�HO r��0@E:214��7�ҥ����OZ�$�O,�+�8�p��4�\^YP`���<oJ�,�7	�sG(6-�O��d�<1*Of �?�t��P��� �DQ Ŝ;qx��o�ݟ��IByB��O�������P���c�&�s�o�buK�b�b�I`ybZ�O�S�@�p�r&��iBN�Z���%��6��<I��)Uݛ�ί~����㝟@�5�J<O��	pw³N@N%*��r��6�VLGx��D�U�\`�甒2B��K'�M�S	\Z�'G��'��ć=��O�p����
LR }�ae�28�DJscSئUH�C#�S�O��O��t�����.wH��Ui�&#�6��O �d�O�)0bR�Iҟ��r?1gMЮ���h� ���a���K�[h��<����?Y��A�RI�oɆYVЕK*�=uQK�i�r��uaDOD���O��Okl_k8�eqv�5i p�c⮔��	8=y�c���I����ISy",��m�p��@��ą	����v �d�O*�� �D�<��ރWǶ`���HQ�d�x0�ނ.�xM�<y���?�����d��4j1ϧqpi�'��<Ynm�S���Hb  �'�r�'��'��I@l�I����M]Z!�#nߜxH�u�'���'��\��� @J���'C���<x�򕂣�l䘳��i��|rS����3�)� ��y#���:�<�v��kܤ�E�iQ��'��	�d���J|2��z"�M�.���a/�i��$4|v�'�I�]��"<�O�Fb��
�8�v�X��϶"�p��4��ĉ�8r*mZ���I�O4��[Q~B��5w�h|�HW%�a@(�+�M�.O�,1��)��e��Q[�c�F��H��=\L6흜'Ͼmo��$��ן����ē�?�����2#��/��nD�6���O>����}��!�D��'�*t����?^,�ߴ�?����?� ��!��'\�'c��;<�Ɂ�A"X9�/G%0�O�Ĳb��O����OR���'�sa�\���j{X$�Oɦ���*U��!�H<���?AK>�1T�yJ��*hA�x�aD�J��`�'�b��y��'�"�'"�ɣ�lŻ$�Gl�fm+`i�0i;|�;p"W���?��������^">Q؈y#�4v3�q��AV:y�0�$�Ol���O��s��ٙ00��0����%Dȩi�H��5���U�$�I��,%� �'o��ɮO����
����8���>1�b�ᄵiZB�'"��'l��98��x�i`��'X1xL ;�^1˧�`���jӀ��9��<�'�Kh��vQ��Ř�>��DB�w3X m��(��Gy���xS��"���6Q�F�*p����Oґ@~"<�BHE��dyr%���O�������s-Լc46�� �?vQ�6-�<���y}���~����R���#V��\�v�����;c޼Xh"�v��d�O`8���;�i>O��xr�ߜ2����s�ִ$jݰ`�i��L�#�xӦ�D�O*��ퟔ'�\�I�s,�,�q�Ԑ7Gl`Z�jהr��%��4o9��Ϙ'r�2S?LE# �N�~F
�җ-۩w�6��O����OJ�3 �C��?a�'i�-h��H�?�(��4��e���}��Z1��'���'���If���!冔�'�,9b��Z
6�O���Be��L��A�i�=W����v1;A�3Y������>���Q�<�,O`�D�O�����h���)����!@A�x=�9��5F�*�%���	�&���I񟸲En��8鴄A7"��ӕ���uV��Ry�';��'K�I���xB�On���Ř���V���]����̟�'����̟lF|��0�GmZ\�ԧ��6t�Q��d�3����OD���O��?2�����C$c^�y"��N�$@n^�5�7��O��Oh���O��$��O��'g|$Q�'�<X�@ �dрZp4�޴�?�����c1B%&>�	�?eQ��'@�]���׃ �F$`�����?A��Q�@����S��e��^wֹ�0Ήz��:��	��M�)O����FѦ�ج�P�d�4�'��<F�N�H�ڷ��=���4�?!�W��T����S�'o�H�p���G���POې{�n�:�pm۴�?����?A��b�'��@Z�xe��򢤆�~�4�Ъķ9��6�-G�$3������/�G��ӑ��<0j��Ĩ���M��?��>2Z�b�x��'"�Or �J������gi���B�i��'�$���  �i�O����O����	̯9�`��bZ�!y� ��Ҧ��	@�D��K<	���?�I>��}<衠+��f�5���:N����'q��
�'��	Ɵ�I�$�'
D���%L=
-Xu����pj�J� )��O���On�O���O*P@bhH!}�uS���$Al8�b��\�����<����?I���D�z9*��'JX����eO>p%�%�PU7<ʞ1�'|��'��'}��'�t ���'l|)�c���{"\���%O�|�;�n�>!��?���Ć(>0y$>U��
�#�4�ӁR�'.�c$˥�M+�����?!��
�ϓ��I�Ş������F�R!�b6��O��ľ<q�	�L�Ob"�O՞DA� F=y��`�uв#0�%�#���OD�$Q:w��?�T?-���	N�-�1�	)�.a��c��D�~LC�i�8ꧦ?!��L��	�K��-�K!u�8�Q�̀|��6��Ob�d�#Cx��7����z��Ԛ'ʏ-N����r���^���H9]MB7m�O��d�O$���h�	ɟ̳�-E0�H�d%�{��x����=�MS`��<�L>E�d�'�tL`�FӍ! L1K��+4�fQS�lӖ�d�O��$�ym�ʓ��	�O��	W�9qgE�X5hY��J;[��b���%>u0����Y	�˝�LJ�������6�Āձ���Â��?YAͭ�zQpp@�&pM
0�c�U{���ْi\ J�x3u�2���j��Ӱ(�2��gIʓ,wDPh����V�k#�Զ`�̌����lK�`*`�ֺ<�b�j�L�� /��)u��8«#��B!̄yG�6;� (0&h�;Y����AK�j����(�r���Ku+��V	�$�t,Y#u�P�$NG#C�Ppr /|�+mߟjv�re�_F��O.}��O��dh>���,h[�0s���86Z\n2f 
�!#���2��8��6O����	�F (�H�]d�4���m0��*A�Dh+�Z�_ib@Z�抟c#�-�w�*s�t��<�G��`��hy�C�&rr0����X����K�ؘ'��{CC�<-4��oQ*NT�쫰fJ�O��=ͧg囶m��>�f��CkMR�좐+�&��^�Pz����Mϧ�?y,�z�(d�O�\�pkY�Xˎ�2'�H5G�f����OV��J�D�X�筛�Ab䲫O�l�� ��X�b�[$�8��-��ꗒ>��nݷ4PY֍�$�Q?�e�51�<���ћi����$}��"�?i��h����Q�o��	Y���8��%�_,!��a>-����ą�x���	�HOf,�L��P�fL�() �i#��Ҧ��Iҟ��ɦ%��|YS�Pݟ�����,�iޝR"<#���Q��8#���!CeW2&�U�󤂰*�$0"�/Å:6��|�H<y�)�$����fFBii����-p��i�D�Z��k�&;�<�nW�}A���O9te��d�[*� x@�\Z��� '���?Q�OI�A����퉌D��gk��OU6`Z�C��j��B�I�H�85H�Mv�ey��x�J��({��4���D�<��n�5���!�΋ZB`@v"��$Ux��pB���?q��?������O�Dq>e��)�n 
4���O\�T�@���z�����+��IL��h�����	d�JX�H�&�6���?'�M��皩~�N��6�+x{�����}�'�N�C��!:?�a�K^�fJ(�CD��?�ԳiXf7m�O0˓�?��2���5���%��mH��X0Cֻ�y¨�HH$���9/�t���'?�7�O��gO�-�q_?�I�a�g��7gL��,Stu�e�I埈yta��p�I�|UGR�q{5ã.Z�D"]��4)��cN֒V�
�KfkK.~�	b�V0���Dy���a��P3mO�Llz�x�iSV�A�B�2]���$i&
呡�H$\v��6ɔuP�̻M��0EM�O����<�v�Q�`D����BM6MI"i����G̓�?�ϓ\��$""Q�]����$�G���Ex�i>�شcA ��@�L@�8�q�J��hE��2������*<�m��Ir�ToގY���Ml�T�BN�%�YfH� X���'��Se Q󾌒�LC�X��T>�O����A�?�~(��ŉV�L�XM��)e��*Ěɐ.�W*ΥE�$���p�<X�P�_+T0AP ꉵ���?V��D_Ӧi��4�?�����Ж`�ȱ�G���FΘ' r�'�0A����\~J�
���!}���o:�����&~:����Q	Nn�<��݁
��e�I��x��f{*�ȴ����Iџ��I�uG�kw�4��H�T�)�g�z���$AB(=1� �+��,��U��E���)�]��-���<�U�T5D,X���-��T�`�]ׄ��P�iu��D ��(9�+�Q�X1k�S�]��m�,�M��^�X���S�gyB�'XJ���H�%b
�x�n�Ȱ�O^�C�V�o� $����H�&�Sƞ�����������<A�ݚ	��5C��;p�$�'E�2A�T���8�?1��?����n�OX�x>�*��.(��`w��*���C��b�H��Q�Sf���	\P�x�/J.���[���+'If��գG7�us¯[�Q��zb�['|\� A��t�M�Ռ��
�v�$�P��삝X��і
�4XE�"�&���x؟V�	Rm�������El@4�0>�L>�E��+b���E.	w�\����Ab̓V�F�|k�,�6m�O���s $W��d���
�bA�&v��D�O��-�O�de>!
t�S"z�$K��N,��b�-��Cw�L�8�Y�(R�<T:I�B���C	Q��3���j��E�n\&��ANE�]b8<�q+��5�&8{�H�!s8���6 ��+�B���.�I�*ټ����1�O�Ac���Tq���hT�`�����2O2�d�O�"|�g�1�Y Ф�	���NQI�'�ў�S��M�珍U�.H�@�`����jǻ�?�,O����f����	��ؖO�D@7�'����DH�B��4���ο#��`8�'��/�BI6h:HEߦ�j�n>�M�O���,?H��%�(kp���sl�v(�'�"dz0AԼN&6M�jMP�l.��@5/Ɨ�����+U��2'�H���-�ᆘ�m��X�Oh�[��'L7mԦ���G�'9xT�ѫ��]8(�bO�5@���<�����<I��.Yl �샞~�zͺ���hO�i�i�'��Y��*ţD���$\"P�fH'�{�V��Od�D�-c���0���O��D�O����m�T�g2�@��E��{�ݡ`FT_�>�y%��.=ܠ�N��(�c>1���<F��6oF��!mČ D��`�+�V�h"BH�-��lA���(09�r�IU�?�N�H�'zq`Rl�<P��� 2G ,��v*w���'��9
��|�����'7\� ��(D%�">բ� ��y�ˋ�oʜ�DMֻ8��\3eAH���dES�����'w�	c��l�@H������ӮC�~���+N�,�Iԟ��I���Xw��'���p!:w��$�|x�Aڀ%LTh�*S�
�G�Ctj��$R2j�.0 ���}����mD�	oVX�����p�p��V*�2*������v��.�Y�ēO��e� �k$鋬Js�U=��`��tmZݟT�'�B���� ���ʈQ��xZRJ�|La|��|b�К^YҦ��?�X*�_���'L7-�O2�f��p�i"2�'��i%��T<"�N�q@��!�'҂˿$���'���>Kt|3!H/�=���S�V�R�
Å"DP�(�Y-����Ǔ�ҥq�A�v�� ;Dh�#��� �=��гF�i��U#�4`��'�]J�dZ���'�r͍c~�HC 
[�\��k�ÕV���'���'�ҝ��|"ȁZ��I�Cn @hQr��x�'~Ӻ�"�Dͨ
8��2�&R�ZE�6O������EP���	s���\�3Pb̂�sc\��'#j> [�iW6=�2�' 8��Q`�u���1�μD#ĥ��f����]g��lS�F�j<㐪,���ЬD���=*(�B%CԐNJ�C3N_S{�����h�S�M��9�Ǌ;Q�H�0g��3@D�'�8����Zd�6+3ҧ����Z;�u�FGJm,R`����x�4mӲ�!C:}�4����*�0<aa�	g:��
Ē��mz�#HAm��`ߴ�?���?aūQ[�l����?���?�Ѿ��B�&�V ��s��6vl� h��_'5 �!����@�$`B�?c>�O$����Mc�5B J8 ��Y�(�� L�� ��!aD@�a��,�q�ROQ��M��[�
/�f	�0*�V��Un��M;�[�:�z�S�gy"�'��YS���Fqs�E�N�,O�Q  �~踰c%�	%�|�w������	��~R[��Y���P����N^���@�e)4D��{@l׬Xd�c�Eݧ"��d��1D���]���	��6R�����9D�+pA�2\��sW�M)ܾ8�D�3D����1���Õ_6h�;�bK !�DO�=,�8�I�[TT	Q��1!򤕜 �^�[��$]Ϝ���ꁓA!�$�9ZvH�5Gv��$���D��!�d��!�x���T27�k2N�n�!�Dӈ^o> �)ޢ7�����:�!�$;s3�A	�<������p{!򤒞9�|�qd`V�D_�0�4	�7B!�D-�$ѣk�Z�~8i�b\�a�!�dS1p"-��̝�t��9X�L��?|!��B�:\��	S�C��thd�CPy!��KU?t)b�U%	�Tp�X]!�ξP�P��ra��Q������5,!�$�;w1�L����-���o�?N$!���4x�o��r�0��P�U!�
+u�^������`�]�tLġy�!�_���iB!~�AIFMNK!���?1��iꚮv�h��ϋ=
G!��!zYH�I�Bς�1��!^1!�D��ld��6e����i���$0�!�D�mF>I����<��`s�ڞ�!�$u��A[������@��Q}�!��G�N �@�G�f�m�g��<!�$88�*Ļ�&L<8��'���!��ΉzD![ OpMf�����?`9!�$M�5���Bէ�F��-�a��.x!�$�"�8�x�`�Dh��D[��!�Y2f.��!�O0U|���9�!�����H�A�8nf�h&� /hT!�ʁkۮe
��%[u���*U!�$,H��FM��
��Ap�	�</�!��Jbk��Q�D1,�H�'	��e��T#��}�S��yb���#Eؔâ�r�&���N�6x��9V���O���E�w���oɥK��jS>OtLss��0�p>!��4(`�­�B	���<A����AV,�>ɵ%�0A��ɠx�tY�x,!�M�K�BP��'�H���o)Z\������'���?ٹbF
;���Е��*̉�U�3�q1
p�w�<}�$3���b�))��IE#A	3f��D�k�`�λ��Fx��T���y*�m��!m��H����f �8 �,��.A�]R��L����&�2~����}�;I�0=�&m��8lě`J��o�fP�'��Sg�	q����EEB	�H���$��/Z�1���Ǘ�H��FJ�IY�����#*�|s�T�Z줥��=��0�����7myZF��W���!t��-��	��%t>�r��M�'9`@� ˲�yGc����b�Z[��T ֈ¯���X��QP,��#�G"(���O���f)�}y�Oaތ��F77gX	��,�%Yz|��D���½�˭.�αfaA�+rt�+2.ԫq�`@b�����hC=n����
!d&��S�㋁|6��RR��>)BC�e�� �Q1�ɒ�	��a�a�C �8;�5C,Ș�&�]��Q9 ���s�0pr&ŋ���y�Ǚ�TЂm�"�+$�%#GX���$��db�(�<!��s""� [Q�(�t�ӎ!���K�0$3�����*׼�Y�k�0x�A6K�9K�@�Ӯap���@(�p��!U-��B&I�c"�䐇�Z�68pP�
M$Ґe8"�I.9�tj�g���q�G$]^@�qg׆t����6�dӎ�����Hy~̛�����T.�uw�
�\�6��U�X^���b"Uc�a�l	Z*��t�0�a��Y'vyr��A�
�R���a�287&���y��Of	a)O��"TiQ
����I&'a�屷�� %!��q�)7\�X��KKZ	Pʏ9w�B��U0������A�l�2�W������Z�� �\2���N	ZUOP��\��8!`E�#P	C%Dy-��$XB�[<���:�M�.Lر�t�A��>Œ���<�ƀ;��I��9O$�H�˼4+��ʦbW�C�~@�B�O��I��[���Ovd9����?I"
u�U��,ωa��T�� >��ߴN�x�ސx�Z\9�'}������W T��=�w�N�\M0�Z�H��Y�z�C�j86�\y���O�aR�̀_;��*�Ē#w������#3X��GVi���
�գ}��$��t��S��36�E:�d���� �Z<�s�Ϲ�nw�ФN�Qk@I1#�p`�$��1���F1q�Hz~1Z����
��D1c(pa̓c����P'��H9�L��	zf�^͟t�柴Co�բ��'v�Ԋ �>������f[Q@OgCX9�G�Y�lh�)q�i�Q�����1~���'�
���<�Vj�5�����!t�dᅈ�?Y�(��[��>AU)P��^�d0+�B-�uJ��F�bma��5h��nZ�!�^Is�OĀ���yR�I�i$�q�����( �+��36�P%8t��2Q���O
�thA �?�cdX�.�x�B�	dφ$�򉐣O�8����'f�P�3�JZ:���yj��
���g�T@C��+ ���{L�z&L߻�ph�
��%Yx���?%B����6�M��,�8� ��!@�������<���+>J��9��R�nL�5�\8�����2�P0kU:OȔ����i!:7*&-Jܚ�c<(A��c(0K���!���dà$���p�C1`�9��K�h��N��̐}tv�&���Xź�Vb��ɓ���#@�*R��</�vK$��ȑ��	��y���,�a��P���(�*O��M��g�7����n�"3E��%�$#G%�6An���3[��-�j�* ��0Z��Ծ6�c����%FsX1:�`��!� ��`ܡ73Jy#���C��!�çaN�\B��Æ�d��q��J�')<��M%�~�L�di>mJ�A�X�*PH��Ӈu�y��G���RءRl��nYZÆ�
����)�=jE��'៷$8X�"K��^�d�3^Z�n.V,���C�1w���T���k���i7�d�,0g�� ��_;,�M���ʸ{��O�(��V{�)ro�@�jYX$� n��հ2C�0�V�̓a�)��^u,̑'�H�,�'�Tё�<qv��X�J���A�1]i@��o�9Q���H�E����wӢݳ�%��;�.�QQl�6?m��ߴ~,$�#ӷb�f�L@��W�I�?�Jp[a�S0� 8��͋�tF�ya�$�1�^�+�e��5���$Ck>�8c0VTF��`��(T�>���`�w'��2�G�.����&����ã}�ܜz@Cۄ^q.��6"@�c�̜�&�H0$�m˕�� �-P�#O̝�"�X0d*lɑ�_{�IP?I�OT���,��G��Àl	��P�>9��DX�Y���GI;81�?Ѥd��v���9Š�[24��V��'��$7�SBū� (7�%c��X�\����l(�M�V�$��ɕ��J�`���M+% C*y���sL�#%,՛�-�+	��~Zg�4}ҋZ�#h � �� 0���v-�cn��>	�̈�t��	A�`Iá�<Aa@�	��Y�-��x�H�'`�'
��˓�~RGЄ��	�,a�ŉA����aSc�:�,��`�&2ܢ̢#'O{M@�b���Nf�d=y���iR���@�Kt?��O�Ɉ�b��gkp݊� ��y�1�g�lyr#�"4��8�'�Z��dN���ԓpR9L�J�B��%�ԍڴ�>�SB:�~2�?1+â,3��"3��9G����2S?1"��a�΢<���(~d�R&�Y�Ë�R<:�s��Č/��]��4k~�<�O�:�qů�<�[wGʬS7#B	V�1 0!OdV�䛎}�5jy�G�DZ�!՞Ӡ�p�а�2N��HOe#%ð�h���*	s+�EzSJ_Yq��@*h r�z�
�ȶ��<!efU���gyEH����W�vc���tф��ڌ[ �>�T(��x⟠��#�#I�̱a�I b0{g����Ė�g� ��O����)�0+��0��^4҈pS2(���䖙]u������Oĸ(�'B���.Qz3�䀧�=XCE�O��=�O���Y���u�
*Ό���lS+|����֌d&�O��1+���~b�Ɇp��!+-O�Qs"��`
�iX��V�x콉��å��d���yCOgy�D�77����'R�zŶpyANг6�p����]zb<�cˁ�Wd<iGg�МS�C_�g��'��IL~�^��HB���D�ȳ��	�b<Ha3�z�F��6͏7s�v��?�dd�%Fa���� GVaٳ��?	��'���/�Sz��T�Ha�b"ZF������W (qJ��o���s���OƜ�������PH9Y�lH�jP�{��p��������%���<�'O
:p�L�	{?qI~*��>7+�9�吂<��e� 
�zb�,����^xܭ������He� ��$=U0�6�+)U��AZ��R����'��d~ӰŘQ۟�M�p���jU桋�%֬!�ȪJH�s�D�ƫ=U��4εM!��:��Q4,<��Q�)I1��}�L������g�? �@�CB�;��P���_o��c)�>,4�M�y������
y�a��J�QQ���'�d�t%CP*�R��b���oy2�'$�����)�V����Ǖ��b`����^D	�FٴUߔe�4�f�9��U�@�LEy��_�d���y'DQ//:��I�")�����Л�?�"�"�y��H/Hw�YJ��%?)�a�M�גıeEN�r�����	U±O���tJ�v�Z]Iǆ5y1�P��x�CA�<q�`���~�*�s K־7��K�T�� ��y+�I8�\��ӷi�p蘳ꗢP�^I�
9{hD3��[k�-���@_����ND0��4���b�IP�u�M�U��w��uq�#J�<`Zѧ�6X]�Ax�&M7G���ɇ ��U��l�э	���'���k^�Ry�)h�ɫz�`�"ǁ9��9�IdJ�3v�??y��Y'}�lyZ��It����F�g�t�3ǆ�%m,ѓ�����hWg���M�1?����qoK�̩Ƨ�F�뉣����c�K!���J�KW�tk~����$3�"��O"�ɑ���xi���'�`����J�2s���"�:rV���N���8��T8��+>�aıs0���"\�x�.y�G��5�
M)aI]{��Ċs��xY����R�$�+O��S�'%�		8V`|�v!]x����4.ϟsA�˓4�����Ø|�B
��3�2ʓF�L�-��2f�-��H�d�"�h ��ty�(x?���?���� �Y���y��17��CŪ�����˸IQ�8w��,��PP�z�����X< ���Ŋ(��7�S��@yB)��l0��Ȥ�e�3N�6<b��P�I,���b0�'����o��G�x˓5��H@qH�PnfP饌CG��h.O@�	p�	�b��r7�Z�?9��V��$�B��'N�����͡	�Z4𵊒Tp�|����O��D�U#+(ؖ'�d�������~y����W7D���{EGF�78剚]���=�?頉O�?>ģ<����D<[I�f�̡ѠJ�P�Ό�'��hO�i�8Fp.�X��&`�2�ģ��f���U}~h ��$���:�[��z40���3}�|dQ�&Q�7��56�'�ў�l��˓�H��ab����A�tY�4�@	���O( �	H�?9Se�Ti��k�Y����꒐��I�fN�(3�h�}��IL?QbΡ<����X�j5q��'�,�����A�X��H��C��j�Еo�l����,
�Z4܊&>
\k�n�6�ا�'�b��sj�%�$3m�6A�N!�+Ot�2���eZ�9��X���Xr�( e)�#׊D�k�`�Ј0��<)A؎}p� @�O�FX���ITP� D����>v��<���d�D�1 P4Y�L�a��$�#��0H�3�
�1�.�:�����
z^ @��8si��ب*�@ D/��ԟH�إ�؞c�����gY�X�tӣ�ɿ.���
�C��}G����ߒ
���'��7�B�A��򲮍�s^��SvJ?�(%0Nok�y:+Oq���Q�4��!��' �.>.!*��"��8���m�����b� (P瘓J��)�sޥ"U��;L�����Y8l|��
�å<	�O+'a��;�#�/W)HT���s�'�h8��(ED"�Q��_�0^|msa��3��Dɢ?��y��u>=@H!§2Zܽ䏃/I��(r�<3ǒ�)���~8����/�b7�1w$���;`Ԅ�(!��h��}�4��C�FLĨ�2B�`]��S�P��S�G��� "����U�vi+��z�'�R�RÇM�dńZ�	(����Я��w����B�t��`��ZK}��>1I�d|�iڱ�� h���1��W �0��(��],���xҁA|}���w�4R`�^fD��
@6#J �2V��0'�x2�Z`�6�Ey�C�*G��r�K�	��:a��y��W<Ty���;;�T5�e�Ԝ8�8��x��I36L̋w��h�f!�'�x�`�Ow����5 T�X3
�T�Q��OT0*s]XTӨ�*�Vҳ"ON����3P:��0q�E+0�^�Z�"O$�05*�5�V����F�;�p���"O�AR�($�����eU�CHt���"O|����V-\�I���Dt�"O�0��蛿�`���:Κh4"O0��!/�5�0�S�NA E�@�:�"O��*�C�sh�A2͊����!�"O����Bñn�����Н����u"O����E�s������0Y����"O���꒥_Q�|@�*�m�~�3'"O��Scˤt}�H(���:E{%jb"O�r��!&ƴJ�	A�g
�R�"O��'k^�=�L���84��x�"O��u���W},�0��15Xx�"O���ņ��(RLx���O�G&Hٸp"On��iX�.�t����+��If"OV��O�x�h4�s.�?@�l�#p"O� D�׍��'D8v���I+n �E"O����̻?�		�Aɿ)��"O�t��B�iJ��q�O�&,2!7"O�1AOǌ��ԛߴ:<E�S"O
d1"�I7�B3C���E	v�Ð"O� �wIF 8z�� ��"����e"O� �A9,V�;���Y�z���"O��Ƀ�L�@q�]	�h]B����"O�iX�C�p.t�Re�,t�mp�"O�!y��^�;�м���
b�,�%"O��J�M��Hk�%C����P"O��D䝋eK�X�$�V9  lY�"O6ȸ�AQ1"��p��Y�F����G"OB)Z�������7b����q"O�hT���z�
��0"m-�yY"O��jF���1f���U{%6�X@"O�Ya5+��1DQ3 �Lmp	V"O��
�xK�|c�ɔw��ܙ`"O4l����p���3gH�M4��c"O��ǥ�7�5��$;MI6q��"O\�&ǌ,�>5�c�^&�vA�"Ox���	�i��Q��Iϰk��!�"Oꅂr���U�6Xrw��Z�,� T"O��!��,uF�q���H/��y`�"O���$fT0Θ�sǑ������"O���B�E{p@	�F�2b�@�9�"O<l��@�9A[�\���@"O�%Ȳ�
jT5S �NƠ<{"O�Q(��"��HQ�Q&c�<Ik�"OS� ōg�<a�m�@�H{g"O����(�Y֮�*Dpr"O@|�����5�b�]�<��XS"OL���AQ="JQ+7호*� �w"On����ȅ��M�W,� �,��"O"���o��	����EK!��ixP"OH��+0<:\�nx�Y�"O�HQ��,(����k��a�XY�"O��cA�	9:e�e/�/��؂"OĹ�gB	;
B*=��Mߘ`�Hx��"O�����#_Q#��
�1S"A�w"O���1�=4�,c.νH5��"O��:0`�,C0 P�,��F?0"OZ5�@��:�(���k;r��	R"O���TЏ��-R��ɉN�X)�"O*u³&�=yZDc-/f��L�"O�`c�>( ��4�Ο}���K�"O���&�cs�z�"�p���Q�"OTl
�d�.2���'��
 �eS2"O�T�U�$@*�D	&�#�����"OA��4z(�(��3 �zJ�"O���ũ��V��p#C�z���j�"Or<���$Ƙ�8 ������R"O2��cOM)>�4����7��h%"O��XV�O41����$d\v7�%�g"O$�jbǭ��!�u��$^�aa�"O�����
?tՓ���cwȂ�"O<������	��ؑbW�8�B�#�"Oh�ghE+~3,|���X /��Q�"OT�#C���V5�9 v�-6�*=3!"O�m��ȓ<7�HS�n�"5�2"O4I�5,R��l*-��,�R�"O敲te�16��XʳaP�OtdZ�"O��W�>,FԒ�酤Uvy�"OV�@�F����q�.޲e�>��E"O� �}oD�����꒷>�<�2�"Oİ�aM�vh� 
tk��^�ҳ�#4����H��� �H��P�����3<D�����U�0�D%�(`P6���:D� `��H	/���s@(S�6��5���hO?�Ď_�q�Ĩ��P"zD��'-ў"~��I<r^t�&�,���As�Ǽ�y��W�v��H���F4  p���-�2�y�KE�Q�D�kOe��`�bM҆�y�06| T��.X�Dse�p>�H<Q3���U,��8��P<H�8袷e^^�<iTl��=��BfH<v�0�"A�p�<i���ex逓�QH���n~r�'~�"F/D�<��8	Bɕ+h S�'��yJD�!}�ĩ�Bo�?uc����'� �{��'lDH;R�ը\�v��'tj��/;��
�k�,i$���'��h���e�F�C�@��w��%
�'���2	\=�~h
�n��f��i	�'Վ��4�j�^48D��1��]	�'��SQh�I֔�"�`d��'3�$�ׅ	H��A2�
���)�')8iy��D1���b���6A��a�2PIDJ�%Jv�*0i�m���ȓb��1�L�/l�4B�#[ �)�ȓ Ǆ���&���Ӏ��pt��J�0L�!DE�K�����"�5��5��H�I�T)L *0kV��k��ȓ36�K@�Q�M(�X��M�C8���*��YZ"�Qsh��@�g GB�Ԇ�I^�D��q�`��צM�T�¡R�����!�$;IL�Y�6ᅉP���U)Y�n���
OK��3#r!X�-U�((0�JP;�y�B@��t��䁺Y���8��C��y⎆4cت���h�M{m� j�,�y���[�c�`�oȭʐ�ӎ�y"C��Vmsv�½a�5bqd���yrk�#8�A��B�)W f�[�HL9�y2S�v����i��\�:P1�Ś�y�$C%4��!�Ql�[�n��$#�yr�S9AK* Ȗ#0^��,ی�yr��+4��M�}C��R�	���yZ�lU匮�>8�r����QC�'[� ��
!4�z���kuD���'��-�p��VkXa	a*�#q�,9�'=��1���� '��h�0���{�'t�ӮZA�ܲ�K/d�0ѳ�'ą���	ipH����I�['Y�.OV�=E���
.�<���K�d@�I����yB$>��PR�ųHRI�Ԣآ�yr.�KW�e�a�Bu�Xr����y��&D���.�7?lrܛ����y�
l*�cD�=!V����y�J�-
�T�f�(/۠eCE����y)Cs�nM�c/��'��C4i@��y��/m�4@�.�=��EY�yb�(pDj��J�]��	tǞ�y��u�zUٓA�S���s��1�yB"�����[ք� �΁��!���p>��'��R22Mr80�Ɇ�2T���0wI!��qB���a�z��ұ� VL!���3i2�p��̣O	PqC╷�PyBB�;��T��$ߨz��K@@���yb��"�@�ӋI�o��c'�y
� �P�E�׬L��Ib��ЏL�fha�"O@cU��I�b�ӉT�7V��;V"O��0� �2��}�4KB�MH^�@�"O|ES�a�0��C*�?L9ȱ�c"O|j7��84|�p��B�}2�`���x��'�
Y;A��:}�H�oĲ\>т�'����D�� 0�e��_8bp"�C�'��ݸ��������O�Z�tH���hO?]ɂ�[�2���V�B���jd�Fm�<�d�� `Uy�`��w� �-�B�<��bN
1���dI�ȼ)�KX�<�� O )}� �Q�w�@�9�dS�<�BN�!rrz��C@"}�I���X�<)`��{��"�L�HI9�RT�<)�F��/�6�J^���)Y�@Ke�<��ǨL)�Ĳg�D��t؀�"�e�<A4#X�Z^zaLUx��d����j�<!��ޣG2 HYBeTfPUC~�<����VI8�ɑ/L�q��j���C�<�rI�"�)T���&�0�A�~̓�hO1�����'� �lIr�;?\^�!"O�H�(�r��3� �9Xz<�"O�I � �i�ta���]�8���5"O�M*4Î�K��@�B>o�r��"O��c`��3| x��!Q4`�"�b�"O�X27Q��XR`C(A��U��"O�y��MN;~r�����p�nň�"OZ@�CG�!���%�
5�YӖQ�\��	�r96��q��>�qCE�f�"B�2�n�4�?b�BХÊ7�B�	�:y���"�$Xq,���G��B�I�|!SV-���0]�kOy�<鳏�/����^?"���cs`�]�<�a�2ˬ0�Pb]�c��a$�X�<�u�ڀ{?����9~Vmq��z�<���ߞ�T�21��4S[�Q�Vʇw�<�ak�r�c��Z�9pYc�M�w�<9��, v�=r���1G���X�<�sѷP!,PP�	�_�=���V�<���X�|!��O�!��,�LOk�<�IK��p;�$P�y2�Ir�<iPA֊���t)�o��A��GX�<1P���4��a�#h�uR5�T�P�<��IW�U#��
�K+nuyX^PB�ə[�z-�C*ά#���`����;�<B�ɤ�ؔ��#��^�1̎�B�	� @D�!�E��4��$�1mE�B�	�e�P�2 l��]H����
�
�B�	&���A��5��H��#ʇ}�B�	1)��	��-*���"�����B�+�JY��P.>�4B�G��Y��B�	�=�f-b��-�\XɤDS��B��8��	��9�$�8�j�JƌB�	�S��0XC ��s[T�A��ڰJ�dB䉿LrQ8��Ĺ(0�} ���6;�JB�P�P<���E�l��'�2yFDB䉡\c�,*����i�KڠZ�B��<����Sd��)�	W6��C�I�C�P���Lڛ[@�13RE�`�B�Ɏ`�IS'$6��'Y�$4C�� ���i'n�ؘ��f˩!�hC�IB2��ڗ�X���ۦIT(O\C�����sIǊ-Z��DJ�"zS8C�I�~��i���b:�t���?.16C�)� �Ӧ��<r�LD0�ܘ.�B"O0��e��o8pYcc#�D;��"O�d`�U�w���1����'�� �"O���і3&q4�M�9"͉ "O�� Qb� fS9(�A�/c�v ��"O^�A1j�
8��V֊D��	h4"O�œ�ʁ�O�~�S1a']���8Q"Oh����օL�:���\�ٳ"O��p���4����:�>���"O��s�F����%j�/Yxp��"O�Q�t,��0_0�sF��[P�h�"O(���D>j�����F�	'Z]"OP����2��I�C	K��2�"O���Ě'�2��&���p�s"O��H��T%%�3q+�?<Vt�D"Oΐ �%�n�*�s�雽&.>��4"O�l�c��!�|�@�H�e6��4"Od9�̜�P-��$�Y�:I����"O^xS&%ў�΍y�c��(Y���"O�L;�֭: �I����t9L�S�"O�aѴ/ؔV �b@T W*83�"Oz� �	�|Ȉe��5K�h�"O�tAe�ȴo���ʒl/
�R�"O>=C��Q 4�R���C �&��e"O�\�D���a�!�p��y�aM�-�1��9
�(�d��yr�M�YؤŇ6
�r��yM�$&��g�LD"��f�׽�y¦��Nb����Jh��I'���yB��C?0�A���*R��G��y�J�5@�ht�7�(L�T�/�yB�Z"S�"�r�$��.�h�ɁFA��yL�"LW@��cO({�L�sfh��y��Ky�9��1F}HKaH'�yb�47"�B��Ҳ?}0)�N :�yb����qo�:�У�HW��y2�%��y�M	�z�� �Q�yq����Ԃ6wQ��B'aM�y�F��Oz����F�;9�4A�K��y�I�oΚ,p"�µ����ţ�y
E�.�0n�9���D�ʶ�y���qU�� v�ܭ�h([�,��y�B�UF�|���
�3ʆ�R�K��yR,�2c6xز�݌�@Y"t	� �y�'d`Z�1D�c�'蟠�y�e��%j�E�W��0ʎ4���;�y�F� IWb�����y�9��L�y��H�V��`�ᒔow�H���9�y��B"r���K�Ɠ�`�(���y���2y���֊���V=9����y�"�j6������)9��ō�y��0�5�� 5�N����[��y򯇜0b8�A�D=3[")BJ��y��܌��L��lՎ(?�,�f�-�y"&B�\�ʁ��������1�y2����HF"܂��Y%�	(�y��%@F�x"5�>�Ҥ��O��yM�!$��-z��*�i@�i?�y�3X�0!��H�0 \1MU��yh�0��i+ޕ*���{R��y�ǉ�o������3���lF��y�#ԫ/��eS��)��!�����yҨ�&��)@� 	V{qn�y��^�$W^k�aR�X'�E�e�'�y
� E��a��Y�hԨ6��-�P��"O��,��_B���	�	%�dE�"OF�8�b���E� ���$����T"O�*D��4H��`���S�zmY�"O�a��)=Z^@�2��u���a�"O*���O�2l1V�8rE/M4�T�"O�9�4�Ųs�Vd��ڳD&L�HV"O�ȢA��?��l(��
-6i�`�@"O:|R�B�g�
X��Ɔ�QR�Q!g"OnI�β2Q��s���3$�d�V"O� (J�|��ip%������ "O	!�+��l-�A��J9v9�a�"O^!��>;_���G�~�b�"O��0v&q�����/4"�4�"O^)k���\�T G��`p��"Ol02���}�RM�'/�	8�hS"O*�� ���n�'nM�%� 0�"OT	 _Ƽ���M�b�"l��"O��s疛Ps�*�B�)C7�{�"OĘ"�E8<@����FF#H��"O00*S�âBl<���˿T"LL��"O 	�hR), ��g�PA�qx�"O,����! �ڑ��I��U�u"O0�!��^�#������a"O���(��-`ٰX����!�!�BrFr1���o�l�+��S3c�!�D��XͲ����NT%Q�"�?~�!��
	��� %\5%\PY�:*o!��%zೄ�T�~`����T�WV!�$�(ci����JX�,`�Գ.q!�D�?*/L��͂�0&12�fh!�9.^,``�8)J��Sj�<�!�d� N��!��挄4>��Ӈ	�)S�!��Ձ21�x����>]76�˒�P~!��:�I�2�N@��Z�)0�!��kĲPq�k\8_H�a3�
2�!�dDC�58LC,@d(c���5u!򤅷O�:-b���on��ϙ��!��ϰ�"ؐ�� %E���/³!�Ć6h����􁁳�p�0F��-w!��gWz@hff���J�;���0
d!�d] {p͑r͉+�"�X6�2<{!�$�w�"��7���ִi��S3�!��N�{�.<�`�	Y�0A�f��O+!��T9IN����-��8���!�$�}��Q��h�h],�8�O���!�DS�9w���ӛ>�j<15(_c�!��gH�a{ O�
���a��!�$��HHDl{�o���z+���&�!�Ğ�$��Yb%ß�D���uE�j�!���d6$����ߺ�)�N�&z�!�;����ϽuZj�P�l�>!��ڹ?���H�?����l�5�!�$�G������B�t�`�����&�!�d��r�лo�N�dm!g)�X}!�D�7UQ:��r[<f�n�{dFV�u!���0�Jm�F�D^��}���./k!�䂽r��T#�
�K��]���fN!���W0��X �ڠRtC<�!���9��j��	�Cϖ(բ��,-!�ĊA��ؕ�18͒�0Ԃ�HC!��-8pT���߫e�44�� Ջ5F!�D��b�Ԋ�,9H�:u.�R`!�DR �f����Rd����LXA!�� p	'N��pe�x���7�|���"Ob�j�K�>&V@T ��P�(�2��"O\ثW�_0�����L$"J�"O��2�n
�_����scY%o�^��"O�AQp�Q@Y�0�6�_L^���c"O6hJ�̞	%^)��U�EDhܪ�"O��r�R����H����%�|�#�"ON�3J�@1�q�@�>�v��T"OHKt�<X�͛�@W9�R2A"O(�S4 ���1��C���޻�!��'w>����c܆uÀ&�7�!�DF*e���#qHB_� �ԯ��]�!�-o��E�B��8^�&|p����,�!�D�6kV�тq쏊�
��"��.�!���8v���/H�8������S�n�!�$��j6ɨ�n�+56R!�tf�"�!�d�7*�c�bԪ&*Lh[�d\8i�!��Ɗ���#�nQ8�� !"����7���zšūrFxh!̔�z"X��ȓDu�q����4BH�`U��9/�B���!(���'Cqr^�;"�:�l�ȓ^�̊F��"��냉�-`J��w�xc�)Q�[�pK���(����b��0�b��*��{a��l����ȓw`�Q"F!Wk2�P#��iz���ȓL��,v� ((t��$��pk�H��&��@�MU#}/�aI�6[�LA�ȓp�V06�O�2��L�d"/u���B
� Y�Ʊ8��G[l��
�'���Ī_�d6��V�AA��1�
�'���谀K;��K�"=8�2�'f�3�F����`b�O�7����'�\�2��n9��)1���$�bX��'i�a2g�0&�V�x0��2 ��$��'킔�eAޒ�T�  ��K$�Ъ
�''��p�\2L]�s�GRA�ƙ�	�']�S��'WT��b�C�0Q~]
�'G|p�-O�%�2ى���6+�p��	�'��1�b����B�U��W��@�<i���3yH��a�-�M�$�b@"LU�<Q�$��� �Ɂ��;&����M�<�r��2)����b�n�^��P��B�<a�.ܫ=�v��Tc��PT�	Sc�x�<��֬Nx�=ئk�������q�<ywͅ�wz�(0��0i����b�<���1Cd���Q%k[�����Z�<�'�U��캳F�v�~%Z�	�R�<�� Kj=�,*�H� j�A�ѨS�<�r-��W�h���b��_h�B0C�O�<��$�%c� E�Af�;� 5�q�Rd�<1U��$^<��G�5�"��c	b�<u�5
�W��1V�T��K]�<�Gm����r)D*N�����C�`�<��a[��K7����pN[�<�4��78q`�cB�
 �;"�^S�<��,��@�.����q����
P�<�'�6M�����\{�YrI�N�<If�	d��̡2듆%�>D�`#�q�<gCB!f)P`��=dZ��@�g�<aa,�����Ǚ��" ���c�<t���8�ȠH�,�|�����I�x�<i5��d��a��
�@4��p�x�<�F 2m���c���jZYb��UH�<YAf�?W�D���ëbI��ҥ�N�<� 6*sh��
4�!��,["(px "ObɣS�P�Z��,�w�L�R�I3"Op0�L�|04*�n���8��5"O�=ô�٥-,^�e�@��ڝ��"O�`���V�%�~QP��&�UXc"O��24C�
p|����E�j�|�"O����X�$$m��.	fպ!ۖ"O�*p�ϻb*$�����(�C"O����FG
T2Ys6.�3����3"O.ke���|B3n�,wj-�w"O�M+��3����ˍ�-aZ�c�"O�UIp��<�L���䅏GD���P"O0Y�g/ y�0�`���o=�e�"OL��A�cGȐ+1b
�(ބ� "Ö;�MI�M�Ș�`�-�Ȱ�'B�1ї��/�Jݱ`�~�h�'_>�:�J!R�q��8rR��'���S'/*8i���X�y�ҕ��'%��3 O'X�|�PJE��6a�'��Q0ㅴ���p��؞J�A�'��A0�K9L��)W♢C4!��'h6��@B�3!->�b&L�!=RH�0�'�������*��sD��g]X
�'j�r�مT�$��c"D�K d	�'�<��� �O(�|xC��Y&�Z	�'NR8XR"N�dw�)S":M�ɛ	�'kR��M޵]�,�%��EذY��'Q�)�7MZ, ���1��кJ���	�'dZd#e)M�mν�cc�Io�,R�' h�#g��F���f�PT �@�'��x����L~�܀��c|��[�'~�	�G��6\��R'(n;$t��'rH�K�q��傖�O%89�d�'�[�'æ�r'e�. (�'��Ւր�(hT�0���ġs�dJ�'�8t懍79�w�^�n�z���'F8I�*�i����苒_�(��$�i{t������&C�f �ȓz�0%bP/�r�4��"�֍a�݆ȓP��� d�{.�e��a�w-�x�ȓ�dQ��ˌ�Nc���FĜ|�4X�ȓa �j�%�L�[Vo��_�Zم�I�l$je��1�D�
�+H��ȓ�� Bf�<)Ǡh��ҩT�t��x�����(o>��Gc�o�0���	��}��źe�H��"��"ft@��ȓ)C%x�f۴k/p�-�H,Y��;`�p��G�S!�Y �EđjW�p�ʓy*��1h��=��Qy1�?_�C�	��Ƭ7��[�ոOE++�>C�ɠ39l���*A��b�F+#�C�I�#��Sr��~I���J�1��B�Id	��hw��(�ꐸ����S%�B�		1�J��'lŰ0��S  R�lz�B���X ��G5< �3a��/x�hB��D�衪�������BV6B�	1����Ёi0�(�w��B�I`TT��!f`vL���  �B䉾ZT]cg���U͞�r�R�~6�B�	�u~u�eM� ^���apkދ�2B�	�|	.5�W��Q"���3��Z�4C��Y�a宕�c�^}B�+�޺X�'F��Ѱ��sZ�H����<B�'�4S�B��T�����89���� *L1%���@� C�X��"O2��\�P�R}⁅μ^l|�3�"O�����Ȉ'��"�B�>�M�#"O�p��n��#�zQ7��Ft�T"O�k���8];�#�IK,o{.���"O��h�g�&�JɁR�R�j���"OT����D�n�"�#�a�rG��	0"O� ���B]r��dN�!< h�"�"O�Jr,L���ؠ�*1t���"O���%3�69��/{8	X�"O��{WL��j��;�iًE�8A�"O�`���kEuQB[�.�)"O�S�&��8��<��8�"O�MI���1*0t��r�A��X�ke"O����@͈}�R�vNNx�5B�"ON<� پx\��, �5n�@�"O
)x��M+-�1���TzY��"O<$Y���)���)J:Q��dJ�"O0�"c��Su` ;��_;os��"O���`̌�M�n1٤��SfTѣ�"O܁c؟"w�$sR�éLP�@{4"O�D����Ai�M R�_�@"ژ�!"O�ݙ�H�*t������V��"O��DV�,N �	���/�:�"O̅
�/�����jS���'bZ!�$L.w����1�~Ts�&Y�VI!�D��|�vę��ͩV�,]P�/��m !�D�(	��i�yqf���4 �!�Dţf� �����.C>	�2c�<e�!��N�b� D�+�t ��V�Z�!�$_( D�s��2O|zu㏴@!�E"v.�i���,�Ė�4�!�d�0l��8@gL�1Cފ�J�W�:�!��j��<q,f�~�r���5i�!��E�	Rj�I!/Rn���TMR�2�!�k����G���P�&C6DM!�C")����+��B��ȇ_�?�!�$��_������+)���"�(�!�_0,�l�3u٤T��`�?(!��PXh4��(cs&�vh'G!�$�*Ƅ��
��;=�� ��"�!��.2� �V�z8B}���#M�!�ͮR$`9b'�0 D�h*�F�
GS!򄛏d���q(��$)*�[⥏�a5!�d@Do�\��\.����CN�xO!�$C1�hdB�Ɲ� \*���-D�c7���}���P� 26�{��!D�Xb�n֗(��|ih�P�"5B$D�x�!Q/j�NЈ��\{���
$D����U@ʞ�I����
���s�!D�tkV�۸��P�)�3���s��+D�$aA��iT��UEH�k�HW�$D�̠�Fh��@ ��Ȝ'J0,"�e?D���Ad�ZR���lHD��E��J9D� � ��Bit��"*b*�AZC�*D��
��CT�԰5+O����<D���핡V��Q�2wE���d�<D���$��FϮU��J�9���3�L;D���o9u7����ǅ>_~�)9D�hCҨ�T��ɁG�U!t=h6n5D��P�`[����ɢo�?Pl��vm>D��U"Z���(���x���r�;D���e�ĺ�.a8V��"<��y�&�5D�TH�&Ͼ?�t+֪�]����B�0D�� F���0�P��E�t��4"Od1�78@����	D��x�E"O�5�t���:��ѵj�;����"O�u�3�I&(�+�(��]F 2"O���a�L��$��A�d��yp"O��ڣN�$��\��jJ�+����#"O��G/��d�pu�i�%�.A"O�x@�+�8
�2�h�/�(B� U"O�L#�!�&.i���th��9"p��"O@a@�܁*�*�𡖽a����"Od�1���@�$13፻[����"Od��e$Q�W�e;c�Sn����b"OVTb6��K�2�G�D��� �"OP�Ѐg�UUz�+@'�P�*Db"O��%�_���1s$T��<!��"OX�J�Ő����:�"M��fuK"O��&�$��]s���F���7"O���3���1F�����qR��S5"O���		WN�,�d��@F�	�"O`Ű�È
-¹Yt	�28���"O�ȑ��%���S�\�N-:踶"OV쑠��2,��h�E��v+B��"O6L��n��Y!ʄ[�8(r�4D��W�_�O��l�1�P���X��3D��a��W�Nv���ꂏ]���th2D�,���M�|�HQ���X����0D����r��c����= ���� -D�pc���+�z�b'n�� RByB�I D����a�%
tpV�-a�.��'>D��a)����i֢X�0� ��;D�����Po�M�@e�]�l\�d-D����KE�o�2Hq�!ոX�2�[� (D��
T�_��d��ϳJD�%D�lrW���&�&l���! ,#D�p�C HQ��g�J(0�p+�.D���4�Z�{͘b�$̐��xhb�,D�4X�� cO��z���32	�$N,D�X�����jp�
�\Tѷ�)D� Z��]�VU"�K�$fjd��(D�8�j�r}��2a�n�^h�D�;D�x�4J��Z��2`'Z�Z�:|�`�>D��H�c�YZ!BG�%B�nt8D�9D���f�$'{:\���ӁR� �7D�$��f�Ԗ9��R����s�0D��`���5��S_�Z�q�m�!��[�e���#Ѧ�{���D:C!�$H�
	�(�d�u	\�С�T�H�!�D�y�$	�e�&�z��$��3�!򄟬S�4�ca(h��<��K�?"�!�dR1&���z�K�$i� E+FMW"O!��#L Zu�A��,I+v��u�!�d�1��,�%-P��u��h���!��;�*��0�W�@��Iz��ũ7�!�DB#b�T�%�@�EO*�x�I��h�!�d&9�8�&�jt�X��X�B�!��
�$�B"E]d�����p�!��T�m�kF�:S�u�Eǒ�M�!��>
����=��[P��	�!�D�:|S<�g0YV��6��'N0!���>�,����/$�g"O��س#W�eʒ��d̊�ca��
�"O�h�j�0m?%(ʎnP�u��"Ot ����Z5[�	�td�)P�"O�a�q�	:�♊�k�"\�\2�"O� ��ɕ(�F�h�V�٤q�.�ic"O���	�L���ν3C�xJ�"O<iŪԽh7���P&ޢh>�m36"O�t���Q��9�se�I�U#""O��0���2�@@�t���I�驅"O�c�"��tp`b�U& �p�"O�6�Re�����=J�c�"OH���ň^��C��T�JѾU$"O���2ؼ,}���bP/g�~���"Op0˅�)�*];�l��S�aS�"O>�(_Q�����[  vD-��"O`L	��hz*��`�ӹHD-9"Ob�!�D; r`M�bA�y*fP��"O�,#e�
s�p´�W�P!<�i�"O��*0�0�>�3����,��%"O�8���_w�tÂ>w�:�zs"O�luo��c��UX��ԋ��=U"O�̑g���L����"H�Dtz�"O85*W�G,@�U*ŉ.���"O����g�!]5x]I��ԓH�4�Pr"ON�����-X��4�����u1�"O�QSq�_��)���QJ��$z�"O.0!��V2|ܤ���sD� 
"OF8z$�M�u���ԅT���F%f!򄞴p2�j_HT��C��Α�!�D1%�٣R�ƱL@L���>>�!��1|qr!��*Y�-����Ǩlc!��85�p�!�b�F� b7!�I@vѪs��[n��"�
[&l)!�DZ ��{���JG�d�i9{j!�dPG�ip�� z(�\0#��]!�����S�N&܂�e�A=!�$ʅ��hu ću�����EO�K,��фN�ȥK��4���&�خ�yҢ-R�2�.9wR4tJ昇�y"�:Tuh�(`�+��UxԤ���y�+H�h�d�ّhS�vٮpIi
�yrM �$�\Y�X�q2�Y)���y���_W~���8o'��NX��yr��F�|E	�,Au�ꨘ B̹�y�!�#xU�U�$��t��XC'G��y� R	B	hS)ZW�ʐ�����y���Nd�pĔL��a�ɗ�yr�ν+�6���k\��A���yR��o�.�є���~B4��O��y�OD�5�:�1��T��Q���(�yr�݃~z��I� H�Mg�(Y�nF�y�O[;ZԈ�ro
�<}�l���F��yB�'$P�"eH�/7,lY���y�'˕'� 8��X�#�%d"��y�I��:?�q�$� ���)���yB�,
�N�BbhD�lf��r�Ė�y���a,��gF`���&���y�!�Hu�u@�iʊVf���*D*�y2�[��������S�X��b���y�A�.�ܽ��,�J�FXX��W7�yH�*���+%��E!���$Q��y��$�Ɛ��]N�V���E%�y���KN^P� �G��� ӥ�yre�z��e��8%���)ł�yr���,9��
rܢC�bb-� �y�
�4m��D@G�1�!�y�ǵ~R�AJ�eX)�vB,��yb!LU�r)� c
; ��	K�ʁ�y
� ����!�}�dԊ!D,I�}h�"Ot�!֧ �`���(�M�1"O��P�\(<��ʰ"��hy�"O�hJ��Z�	���� -H�(�y&"O��r�A�(���ɲ�Q�q�~�
�"O�!uoH)EJ�Q' Y>n8�"1"O܌YU���l0q����W����"O�P�7	��|�a���Y�:O��R�"O��X�∴�5{�,�{T|ȁ�"O2�qG�H>�Z�cL�����Q"O�{v�:Y	 ��$M��YВ"O0��C�9z��[��Y���R�"Ob i�]�`B�k�Y
"O.�CX6'ϔ�҂�P'[��ZW"O����d��!��A�08t���"O$C�ȃ�������ٲSŘ�Q�"Oe�Z���$�t�N�M���"O���AEUrۖ\����
�إ�"O���Ck](�&�E=��Y��"O��7-�#I���R%�	mq`Ł�"OV)q��L�f�޵1������9�y����n�	���N��qq�ქ�y�Ҫ.J�Xq� C�M���J��yB��XI�mXg�+�´jW/��y��}�@s�D-?�Lq�K] �y"��7J%'C��K��;VD���y�-�/���ka�V8\xtj9�y���Gf��#�5��"ȟ��y��Հ<�xR�9J���Q��,�y⍟MԀ�J�xi����*��yG�_��p���K`(t�qP� �y��E�Hl9x&CJ�Q��)��ހ�yrN��0!��%LL�p�;�#��yb,I�5�u8�۾z�*Ո�˄��y2aǓ-�r�
��P�<d���L_��yR	�&|�h���0���qԎ��y���;<t��r���X�
���yb�DV6��b��$V#ԨRj@.�y��E�"춼a����T��4h5mD?�y"�]�r�r|C���Ex��x�+�<�yf\�=24�ԧL�?
�(r5JO�y��X5[j媑a�3�"aK���y�̃{m"��� ,׶0:��y���g�r�bNH�Y�,��đ��yj�2m��,Y&b]�QO��i�^��yBk�!8oz�bm�B&(P� * +�y�&�B��PP=Qg���$��y��F�q0ꕻ7��p��Ȕ�y����۔Iz<p0�N���y�H<d��P��I$�sA�
�yr��赺4̛�w�r�/ �y��ֳ;��!��/ʣT��i$��yb�C>~�LAb�1>���2���yҭT2zA�3��)0�(1��P��yBș,]�U��?+�zQ��ߥ�yF()Ԟ�p4#Z�xI$�ss�Ս�y�H#c���w����⏋,�y��[T�ے�lT��A��:�y�����3$jS�]��M"�ݗ�y�G>��
G�T�P��1����y�nլ��\qUE�-R,> ��Բ�y­�4	p&ؙ2�X�E��B)�yBe��%;�܋:G((�@\��yRaV�MRL��	F8��aZIZ��y
� H�S�-I�}	p��6�w��D"Oa�f��<���:R�N�us"O�Uj��:@|�e��d@�7���9�"OQ�C%��Ih�IGdU/ ���J""O^�PWg�7���j�a��,�� "OL���kLV
XA��X2M�4�R"O�{�c &+z��؀eM<r��U"Oby�K�(TC�Ή�3��	#"Od�p�	 J���+�J͈*���z�"O��E�S�g~���:Gjn�sV"Od<����Z�dt�c*�sT�T��"O�`��E	�,���/�sJ�D)"O��S1�
��`�+�.�����"OfpA2�}C�L��i�5��|�Gi#D�H��j��m8l��s��36���F�4D�����{��)�3�A�ȡʂ�0D�\� ,õ!iP!���F�i���&-<D��NR佳�fA;.�4��!:D��:��,e�~���ߤ|�4�g6D�|Z'B��,X��t�?:�|�#�3D�h`���^����σ�H�`��q�0D� ڑm�_ֲ3��#9�l�$D"D�|��O�h*��p+_�e�8e�6#+D�ԫ�i�TH��x%a�<��qA*D��
t	Ԉ��l����m����FE(D��9W��&2��]b�� |w����%D�dI0ʃ�[�¹�EV�TDh� �"D�<[�G��v��]�d!�N��U���<D������;X��%��P�P/����:D��⧈ݥKf�H8�eu��$�E�:D� �"��U���I`)L�":X+p`9D���r�#[3>��F|�X�n7D��
'nӒ4�l�����:2\�!s�H!D���D�M��~��SH�9`�n��4�9D�D�p�K�hd��⠄��^��z@�#D� rG,�G����D	Wd��p�%D��
��Y -E�5�G�@�"%I&�>D����@��`$��
�}�P�1��)D���Tk�N��k�H��Q���&D����IG��S7'��-�@�?D�	E*�1*���)Pr���>D������@=��a<gX�
�=D���D��;������0"�pӪ<D�Lx!��/
�0b�ӱ[�Ҥ��:D�� ��Ͼ ��� 3��?��I�1.D��aC�D�&|3�E��^�����$7D��QJ��^��%j�>V-P�+�� D���A�� �( �RLT*0�BI��C+D��ɠ�ħjQ��!�S n�Q[��(D�䩠*���Xrw�.S��c'D�@ɶ���1��\���U>C�(jFg D���!@��]�3T,������e�<Y���u���S@�-dP��M�c�<�vl�;\���#IĦz���OUa�<r( �e@�2��	�v��4k0b�f�<��&Q hY� �L���U;$�Lj�<��V3<T�"
���p�dj�<���Ƒ,f��sHԟ;�<��A�<9�e�5�dx��Ֆ.o0���`�<	%$�]+���s	�'�r�`���\�<��7P��� ��G\��y�h�l�<��'E�oZ)�F,+[9��Hk�<	qˁ%�ܱ�]
$���2�Xg�<��bD9m�d�u�T/{�(�׉�`�<� �i%��?I��y6L����,R�"Ov���u�.\C�k7 ˼���"O��f�O��y�%�^t�1"O`���6<_@�pm[�-����"Ox ��Z����AV$�fI��"OpL�k��3�l�#!F]fRY�"O��h���=&A ��<[,{C"O�h�u`�`�,q�OO%a*�h�"Of�,�U�f�޷=���2�!��T�,a �G�m~�LB�%�!�D��8�4���L~��!�K$W !��yC� �嬒�B��dk�k4/�!�c��у�� ����Q
�:N�!�$
*2.dHf	$ �N-rtI�|L!�D������F�w�� �0( m�!�䜠:�^]��h�>B��řu�_��!�d�)f,Z���M<� Q���!�	�BX�X��따F���T��w�!�d�>;vL�тEXx������c�!�$@�"�P��&�!o^����� ^!򤘃b����[������*q�!�DI'��M�%G�Q�*A����i�!�d��"�-҇��E�x`	�l�!�$X30$t]f�;#���)&&�!�
�Q;�Hpq+Ԙn�P�"G�0N�!�	Y�\��h���@��&f��]=!��`i�q�b��\Ӕlç��+-!�D3C���� t٘�	@�O!�DI [:�{��*	���z���!�D[+qX�i���l���f��<�!���9m�d�E�IV@f��b�4/!����Q���^-$����K�J!�Ҙ4y�����$:�,�*��>x�!�$M�	�hXk�nҾ�|�8%K��!�dƔ钴8�b]��0Ui�B!w�!��-�	�хG��8�d� u~!�D@�@��Yj�DT�0��I:2�]�d!�B�J�$y�'
�j���P5��
�'�f�s��H�m�%���h~�!
�'�ؘe��8^��"#c��X ��
�'�"�qa/Y�<>���iIA��E	�'"�y�,��f("��ݵOת@X
�'��"!�Y�阒��M���B
�'Epx4�7o����b�M�K����	�'�4H�ɍ	�Vm�Q��IiH� 	�'�@Ck��J��@�MɃ9�F�{�'t���[�,�p ��&%9�}��'�<p��*ÂyxFP���_��I�'�|���m�oB�&NG4Z��P�';Խi�/Ǽi`mP�lճV~����'=��3�͚$�8��f�V7b�K�'GD5��X���������FDX��'� �	�̚�^&L@��E?�	��'��X�+�LA8)����Jٸ�a�'�֥5i�%}���0эҙH��C�'c4�a�f�u��`�n�8�\)	�'�X��b�hj��ȁA�"(e0�	�'��h¯ۡ�,��1�������'�t�jT)�� 9!я���U��'�H�Ǟ�DHz�QM��z�X
�'�H\�6_�~)NQ'f;��	R
�'����g�5Ą�J��x�Ҭ	�'y��H���S��x~Q��'KR�)�(΅4�ryBӡ�ktJ�3D�� B���/�(<�X�$CWкi�0"O�S�>hd��:"��l��u"O�����]i�:��W�ıHb��ʑ"OR�*�&R7u٦�['��kPp�Qv"O�H�aͲ%m�¤�_x@�q�"O��z��Nے���IR
�A�"O�Y��<L�ZeF<+`H��"O��H����DB�a@����"O:�����k P��}1�U"O�!�s�a�X s/�-F]�e+"O���bE�M�h��c]8LU��"OD�b��;4,@�㚅+��0"O��(�Ǘ����S��>h.����"OnA�ƍ��Dhp��@K6b(F�z�"O� #�!ש%��\s��2�@�d"O��i �;n�$�`�S+S�h���"Ox�Y&��=}v�C��z\��93"O���1k]�\o �he�I�_]@ K�"O� ��W9R�X@���V.TVa�"O*):�E�4$�G��-0�F<��"O�!Q�/Km��93��G�|P��"O����,���dhUB��#A��c�"Oxx
�'&ݰ�ad���F*@ؑb"Oj��E$
|�B��{4��f"Ot��i�mU�h�d	�f��M�"O.d�S��`�T� ���r��"Ot��aȑVQ4�*��L�����"O��C���9R0<铖"�|<9W"O���VF��6���Š���ڥ"Oll�)5Qa�|(�N�/n���j�"OH�Eh�m�$�vqҡ�"O��!JeJ0���G&H��"OdzsOé��Ђ�C�2�};�"Ỏs��M�ؽ�� ���$��"O��@lX)ua�� 3E�I�"OR�QR�	w���!�B����"O�MA3F֊� ӡ��#�A"Oԍ $$X�ޖ�[�q0ֹ��"OR�`a̝~O�e�B�(:T"O�X��E�.��AE��F���"O�Ma��֙N��A�/�4M�~u�"O`|#֍�1����L��q2y�"O�k��q׌�LH�de��q"O��B��I�3h�����k����"O0�A k�`�b�G�|�|�U"O�����Tb<C#��D��w"O���J҄2�(�Ibl��73L��"O�����.' 4� fB$?0��b"O��(U=S20���^`=
1"O�8�1�	 7D �����)s)X�b"OҝP�ȭE�`K��ߦ.��Uz�"Ol��k��8!�t�u��t�L�s""O�P��B)��-KCb]�%̼{�"O��Kb������i��̮*'��jW"O<�����
��a�F��"O��+R�Z~R :� �?ꐘ�"OR�"!]�'瘹���*1�����"OP� �!"��.R�G�r�c"Oh�+�h��sb��m�A���`"Oda�㭜�G#�t�R�H��ةK�"O ֍^�$dStd�=H�ءȁ"O���Т
OA�-@���[���z�"O޼����1.r�+T��<�f8�"O�9���֙%�x�Rq匵{�\5C$"O� ʐ� ��(f�tI�%}>���"O��y�)ػv"h����a�jԃ�"O|��^6md��2E���3����"O0��Bj��Mg�4�F�a�J�I�"OZ��#�d�� ��@a�H��"O���Ue@8��9j��:$|T��"O�����v�:Q
�:v_ 0�W"OTႃGQ�=1����(NN��"Oj�{��%w�R�� E8b�P9�2"O�Ab�aK�v�Q��C�E��X33"Oന6NλZ����I��'��̓�"O�q�εDY �&$t(�q�"O&M���T$c�^���	�<~�M��"Or�x�aV��	���xlY�u"O�4��+��}���Dd5)d��"O�L�R��#
.tc��9X��D"Oq��Q��XE���f�X�V"O4�jω2&�á�$�hC�"O<�҄���X�p&�ȺA^�li�"O �*��I"R�e�����+�X��s"O|,B'Lë2�̹�4�D�t�x�q6"O���4����U�%�C"O�4@��Q0CXؔ	B�D1[>�E��"O�"��וXH�	���,T24���"OX��+��0����t��!,��8"O���`T�_�<����֎���)�"Ot����C�"�֍W�#�@�"�"O �rCɦO�L�r���,4��i"�"O�C��&L�5��L����)�"O�13�+ް$@@0���z� ��"Om��陆!�v�a$f\.�"�P"O�-xQO����kI�y�l8qE"O�0�##	>���B�,M_���"O(�R�k�w0���4A�4:]Z""Or�s��2vB
���O� +e�ܣ3"OͲ� �2\�� �l� =@2"O �Id����]� �ۢܳ@"Ol04�ۇ{)��;2����H�t"O 1Zw+�&Nj4�CH:�4j"O �x �- f@�@��*B؉��"O.���)R4�d��x��}0�"O*�s�&D�,�H}��c2!�D���"ONLbD%M.>��!bL���j�"O�Li�N�A/j�I� ���V\)�"OU8U���os���V {ϪP�`"O�0`Vg��hS��	�ډKj>]BS"O$�)$���2U�n����y
�"O���D�[0�� 5;5b��S"O���$X�|D�6,�P�4�"OC��/2�0�qd�5GjR"O�<A���D@rA�P�_4f&�)�"O�p�c��7P��t��"sj�-�0"O�̃�/ζ^b����fV9T��a�"Of�P�[�>�M��K�<Gp�!G"O�l����1�ps#L�	" -�E"O�m��D��A�6�$X���"O�E�eς:���m��U��,�4"O�!҆�t�El��c��m���<l�!�ׂG�Ьآ��2���aՠ��b�!��Ռ?S���m�7M�mC���;2�!�DO-}dA�1b�
pQar�Ԧ�!�d��~I(Y�pB؜I+��Q2&]!򤙿{��I��Ιͬ���l�9|c!�̔p�^e�@�L�v�
��I(!�� D�!7g"tp� <u��M
!"O��)DBΔk$���E=%߂1�"O��f˞ z�x�D	�h��Y�"O���bҦmo�U��i`��*�"O$  I�E�����aѦF"���"OJ|y��b������
� �2"O�����o�><��H�9 �  ��"OXu����)�!񦧄�~��P�"O���f ��A@Le-�S"O$ѓ�K�;`�e���#R�#�"O�H���&jTYp���tZ.A�"O�#�O�\�x@�I�k�>H�"O1�C�R�A� �!1hӭh�$t�"O���F���l-��*)͚��"O�Yjg3?ydLX֤Q�0�@AqD"O^=���/D���K'mV��A�"O�U���$�(hӁm�	4id"OlT���+vm�U���	YT4�K�"O�ě$��DT�y�,�	J,���"O�̲���0`R�UK$��3��q�"Op�8V�Ɲ=Mz�Rţ�	$J�d"O:� TLʎ��4jcB��=!,<C�"Ot�uI�|a�) F��7#"z�3�"O�Yt�O>j4�"յ:�E�"O�u2Ѕ��@�5��)X��s"O��
W#՛Ov�0��,͖^�nM��"O����\,,��XX�+ӝ ��u�g"O^e�CҲ`�P��P�����1�"O DA��O>I�� �/w���x "Ox��4��-P#Xt8��u����"O�BSn6_n�r�&�hQYw"O�	��)���!G�+l�"O^	� )v,4�7��><EeA�"OvŲ�)�-V~ �Q<���G"ON����z��B�C�TA�a�b"O���e]�$�P
�o�9°���"O��s�d�/FK����_�]�bQ��"Od�ڂ G7a�p�����$)BF�#"O>�bDH�'M�����ں+$A��"O )rR�֣Ku>�p@�1]πjc"O�e��f�-wrB��![t�:<��"Oh���/l�:�" ���yd�0V"OJ쀱鏍O�����ŉ%c�-H�"O �ڄş�7u.$g�	'V�-��"O.)s����6L���в "OFy��kQ]p8lH"��W�D9��"O��0�ǟ�,6@�6 ۏ@�v5j�"O�9A$CϺ}�B�� I&t�l�"O�x&#��;�dܲF�=�d��"O��)�*J�xa�����c�����"Ob� �h�kz��&\!K����"O:-�q�L�r��;�Q<;F�u"O�u"�d�YP��@���7E�Kw"O8�x0逰V��P��ȋ?+?Vaӕ"OڕX@�X�/��$zv��Eæ"O�@�Gn]�3��5 � ="O4�9��ʉKʸ��w/��Vبx2&"O,�KU��x�la���%t`��@"OਥmI=%~�\���D?��� �"O��r�f�&V	�w�	;;�j�P�"O°X釓
�t�%dO�|�Q+�"OD���t���e�����}z4"O�e)`ʊ#Q���g�\r&-�"O0���'�a2mi7��fR��"O� ���ȀvA�}bj��R��@�"OXip���1�hԌ!���"OTT�
�X�Л�I�(��y�"O�e�@��T�
��!�^-��l��"O��`4��B�Jm�1M�_��\�"O|ڗ�C�^��!�́�R~���"O.@`w۫s���X�lųjf�)��"OJҤA^�y���5�ǰ!�ʝ�@"O`�@)5�Lԋ���?��b"OH}ٵ䚨h�RDq��7��8C�"O��#�`��D���/$a��H�c"Od����
���O��Mʔ��f"O�@�e�2fu��ǉ�'��$�F"O,�AE@�V�B7⏙k�rD+%"O�i�� �`\2a I
Z�:��"O�ub4&T7��4�v���0���*u"Oz���g
�]�$1��ԉ3?f�b�"OX���)"��=�cV�64��2c"OPY�c߿lͨ�2�l�5G(L��"Oj��w��Nd�Yc�)#9-�	�$�i�ў�w���Ot�B���,��-rRI��\m�=q!"O���Vm�*s��aň��O?��0"O�h@�R��8]�7'_��x�p"OD�(��p��CF��^:��O�]����ҋ<H�S��w���H&�y2�ݖ;(299gC�o��A��y�bQ�<G6բUCӹ7���׀��y�ERT��ܫRG#@C )RV���yr K��&(���Ժ'�dx�-A�Oh��dוob�l#��J4��8�kѯ_!�dM�a���aD_<�4`F�$!�"s�(@� C��q3o�+���a)��z�d�`���y��2��O2���:���k1�fB�p��ӡ�$aӄ|Y E����g�K�#��%�WOv09�솄F�*�ceoF�7j(��I+��蟬��F�ԣ�b5���ߋ]�"mj�"O�X�K\�*���"�ق]�4��"O���<}V41�����I��2b�I�G�	Y�1;ĥ�~Ǯ�4f�y��T-��C��Z�'?����,A�ў"~�k�a(�iU6�2�H��EN���ȓ@ U�����X0��xr��lQ �&���O<����^)\��e���	!�͂����I�!��٢f�,�G���U �YitfȜV��O�t��	w��)�E�=E4Hځ�BC��/)����r���TĚ��O�D��p?�V�!l�]��mćL�p����~�<I�m����7�?|(��.�w����'g� ��ŉ7+�.1pO�A��c��9OZ�q�J�+�Z��N�	xg޹at�'��'��-�u/G.r��| �K>��a��'pp�X@D� e�8ҷ(�1��uSO>�,O"7m*�' �᠅E����SGW�B��ȓ{�| �	��m`����D�vE�'X��hO�.?��̂ѡƸqX���k�
%JB�	�npx�t�H6d[�5�7oQ2-[h���8ғ:˚LXNS�!��5����Q =�ȓL@(�;���� ��X:\Ȥ��z��P#EN1(� �I�i��Ņ�~S ��`D 9�&1�!S{t؄ȓ9`�Y�F����5i�*�� ���Dy"�
�����Nk|>��W�!��>�K��*\�K������&�Y;�(��3�S�g�? M)�TP��]�㨋��:@)��'qO��F���Zn^q1Ve�L��qa�INX��Ț*6��x!MM�?��᧨/�O��O4[c�ͮ|�Lܚ�e�
�>]�"Of�R�\�E��\��e��c�d��"O��SiF���-����o�8� �"O��p��5h�苵LX-jU8@��"O ��ň*pG�98u�aD�@�"O���sL�%V��Iu	a����"OL�ҧ.H7R�6����q��"�Şw��������v�)�=��O�j�Z�D��vグJ��
 �f��	Y�Ih�P��qBQ���#! C�ɂs��%ۓm�x�,��ףʤ&�"<q.O�=3I�$;��XbS��$P$�Ii���Z�<��`�$n
�,[@"�C�N�pw� r�<A��]���uJ�w�v X$F�l���ɶ9�9GGLA��%��PC��?�ɱ2�W�S7��r�º�B䉬U��g��*/,`x�BS�����d���Dk��4A�i�DfE/n,��b 'D�+�+Uj���j�l�|�ЉU$D�X�j!�8�pVF²c�����x��P�)"�q�E,ғKu��r�/�p=��dL	Y�L]� J�1q�Q�@�''�!��]�V�@�͛KS�0H�ሶ>ܱO��Ez�O!�d��n�dI[�g�C���ᑪN�!�$ɹ���Ka�σ)�Ȑj�-}�!��:�6dx�\�P�sM��!�$q������>�`�"k��(J�$D����/��#��K�wVXYre8O�����܊ך`��NO�B0�0��_�!��ɋd���R�̙�i!�U��'Rўb?m�RCH*�,��`ԫ!{���� D�TX���]*�|�6���:D�����
Ʈ��r�ĳY�����4�O��r�x�bAʡkxu�1Ó*Q�����?�S�T���x	Z�
-
���qˋ#�y���z1���ۜd8���CL�y"IT"[05 � уM��;El٣�y� :m�89�ӯ<f2<h�MO��yrJ� �8���@ʹ,�@��6�Th��.�Ds�>��'�rp'��o_6��2��%;.����'�a�A`�CC����L8��3�}��'��1�4w#��s/�7#�P�1����v�<�'��-�b �R�$)�P�ƭĘIӫ5�S��?���R:�Tc&o�&f�@���gUqX�DyZM�<�х�()}Y��ʖ� �C�	-K���0]L��S%A$�B��EdL�dm 1��A��+S�kS�B�	47��|9�ǌRJ�}ئ�ώ�P�=��'7�y�ւ�:����D4�B��y�UXC��oE�"��;��EzR�'`ȉZ�엛	,Ia�aJ��E��'��Ȼ��>e�DI���  � �'�u���ɍeҜp�Q� �wYx�ۈ��9�1�c�cI�.P���ƻ:*�ȇȓb	���Q�4�z���� ~�t���H	AgHƢL���K�.Δ}Up�>9����$�ًC��@��I-]a��6����0>�C4�2l�7o�m������[Ц�G{���ij28�e��h�A���Y;]%d��	�'�(]�3�I|�6�i��V7d��	�'{���E�i_�9���ĸU^���$ �� 00��턇+���q#Q��h� g"O��ȵl
$ ��p�AEvn&�C"O��q�Uq���9#a܁ _��P�"O�y���nԬ�c�)mQ���"O��'%}*H3�:���p�"O�yI�@ϸ�ڗ��	�e:@"O���&94��qp�#���d"OܴK��]�oĤ�*�]'~V�"3"O~l`vOB�~*����=9�p�"OФ�#.¥H�6��E#Yd.r���"OdqA@����A��+C:G���"Oz]Pf���C����X�>,>D��"O��	��՞G.�McP3}H9�"OB�9si�:�nl ��Jm�p "O6̳�B] z��iC6����<(`"O6���>C�Q@�Uc8Cf"O���K�n��T�s�&g��SS"O�,��=>3l1�!_߮�"O�!x���. T��^j�rݺ�"O�l��~�tx2�ꓶ ���Ӏ"O�Ł�e<rV�y��5��Ԡs"O��ђ��=K�Q���Y6�*�b"Oi�瀨k�n��@һgЦy7"OQJ�J4�vP *�.R�r�2d"ON( e%�43��h��(��w��A3�"O�=�c�]�>�:d���؉d4�%��"Oʕ�ÁǚB���ş7)B6y��"O��fϡ^�� �dS�@�Da"O��Q��Dtxu�P�W4���A"O��"o>O�t� W��!��\�"O�e)�	�mH4��D�7n���x5"O���Ak^@'P�AS�!�����"O(	�ю����A3��I�bA�B"OJ�x�lQ�,���Ae��6tC�"O��X1���h�������y�"O��{s�G������e�L��w"O�Hc&�݌f�v��iϴ u�m��"O�iyh��H�ʠ����40Yp9��"O�1:���>D4$���ժ!@>��"Oxb��=T[�؁�	9.M�"O���iV9B���SL�H�b�"O4��Gܔq��Ep��ӑ<C��T"O�p�!�G�r 2G��ZG�:�"O����*�W��z��kI�(�0"O�]�pD����dK��+%*O@��0�_X�X����GΩ�	�'܄��+��k��9��jEj���	�'Ү|j�#A3E�� �LW1ly
\ �'򂑋Q��4o��:��C�YH�j�'s�����"V�6A���X�,x�'�pɰA��a��X��v!f �y���>��|Z�
�q����d�R��y�Nx�Bh�e��yҤA�҆Ƴ�yb�����)�)�<f#��3O��y�%o��X�lF�kq��iӧ݇�y�Ǚ.��%����:3�
싑�M%�y��˖#:NLj"�,���h�(\;�y�Ƽ�����
|��� W��%�y�Q�s�z���h�p����F���y��X{$�#P�~S�!ۄm��y�E¦����`�3��HsT�D��y2�*h���P��&-جq��^�y���Tŉ��ʽRR\��S���y���V��(['b�!=��!F���y
� ~�p� �a�"ՙE� ^��`"O�lZ!��SD:��AD��"O*a��
.��� DjK���"O�0��&�q�xys��ې+��t"O��I�x�v�;��;���E"OJ�k�l��@�*A�PM��"O�uk��I�!P�Sc�ҏ>��i�"O���!a�)��y�h��V�I �"O�:��;8.ڤ	����?u���"O>Ȩ#ÔYH�i`sf7/�B�%"O���3ؠP$�arF�� a�y@@"O�͂�I]�v���v�F.@�� "O�1�R ��T����u�X:y40@�"O�d�E�].|���/D�X���"O0�Pr�)<*�kQ��+Xʌ��"O�!EfJU�H"�/[�VNP�"O�� ��ުBL ��NK,vᮕ@"O� ��16}��żFpB��"O��(q�^�~>�d��FN���x������@	h�zR�қl>"�H���3O�\��%ۼ�>��)�6x�Tj�-A8X�����i+I��eG��nPB��9z��ȗg]�^Xց��"2���<)j˸x�����)��Oj��%i�	-ҹ���S�
TJ�', �%��CGXj��r�(p���CZ��$��d�tu�S��y�T@���t'R�Dېq;�����yrB�)e����ɢq�&�K�+��yrFܼ&�ZWm�G�d��ɭK����V+�/T2���bO(��d�!1�HbV�C/O�� b
d�)@r�P:%I��R#C3"�B�I.^A�-7L�-鰬r��K�v��|рN�X��d�N�$X/�e�|�%Н1t�U`G� 4y��B�<qeKR��ළ]7l�nlb����V3���e؈xP�U�f�F� D��'��-����*DŰ���o�D�&�B�'�h��N�_�x���K�J�����^�1��	�lܠ)�d���0<��G���d��疷3h�rl�_��pSacֺ$�l̑s�hb�1@�!�ob�A����<�|��v�C<a�"J�`�ȱ	E� ɖ,�T��V�%�  �R ���r�#s*�����ʺS4G��fḰr��=�:@��@Y�<�F��Fؑ*b��L�ț��?�
10���??H Y��'_��@{�g?1�#�;;�< p/\�!T��R��R�<���!}؂$k��K�
VxP,Y�<����3%��:!�ÖO"\�=!4�I(5�H��ڡ\�(pt��D������(3**����8;`}3�l�=8�*�hE�!�|䛣�x��Lx����9��Ȩ4�$AP��͗r@qO"��˹!��Q��A�,0(���M��h
+`�ҁH�,K���=R�E���y�OP;-������� S�(�Ƀ��Mc��P:{�0�p5@j�p��?���~�'�.�QĂ�y�^e�W(U B�\ͺ
�'B:y4��X����N��R�,�P7�s�h�Ea�}���>��?�I��FP�%B�5�Й�D��2cF���g��@�G���4*��4�P,!�H:ӆ�8bÃ4�Lc�� 2�'#�1J��A��,f! �h�w�g"
�(��Z4�%J�� ƘO�b7	��l�d���e�8��S�Id�<)F�9VJ��3��&Q0Ċ@ ̧f~Ԥu��>W�za���	�`�''���g~�
��}��9�aiF�CpBy!$�Z,�y�!��58�p��[OۖP3�LF4�c㈃a#�u�4�I�R;1O�y��y�oκ����m��}�'�&�0=�kR?s�L����xu��0�����%p��6{�X�p��܊��'�^Ą�2,`�����J�y��7�xb�|��P6�l ��&@h�5�|�2f��N�:��v�K�*5�5*�M�|^�B�I?ϒ	S��P���^ `���p,�2Q���a@����ԟRɪK?�S���3��\�6xT�N=SSL����%�eȉ/��x��8�� �M��[��t�ҫ�5�T��=��. �	�F$ %1E �'\�x�]t�8��� KR�C���A�J 
D	[�$���'D
�%P��Qg�)ib����2{O���I3�JUv#ۖ��Oll����d���;�����S�? �M�U&Yv�Nd��� l$��bp"O@��!�ԩc���+ՉG}v,�ks�+�H�2�4������BD̐ye��Yj,ə��ҚD6e��Ѧ��p,s-�܉��+�<�'�X"=E��
�$q�݂0�6��QS�
�	�y2n_ \�5�RB�~�j8j�����'��{"��69��}ȓbZ�^9th�!��y2�2u� 8��?_��� h���y�(��k���K+VwP�{�#���y��"__�Q3!��{�ޅ�fF�:�y��S�54��(G�2"�<������y�ۚR�h�G/��&�b��J �y�CV�p��d[��J�l܂�[b� ��y�'Z=��ѡC�4Z�4i�o�y�-[q>�|J�%�=�T��a"��y"��XȔU��#:���;A��%�y2��3X��YPX(	�����Q��y�ě�8�E�'EؗZ��g�^��y�3�`�����NL�Y�gMH�y"�Ғ~�jQ���1V0D�	��y�ᒏZ��+�� 5V|���ǁ�yb/��@!Rbh�#�"�NǠ�y2��8X�-34O֤�n H'fά�y�M�	��ЙD!�.;��T�+���yR�r�܃�M�
;�R鐓m	��y��F�[ŉ�AS��0��ؠ�y�KH.y���F.�'v��Ҧը�y�ʨ<�F`�QbѾE��X�����yrk�#�|p:�� 4lHܢ�'X��y� X
�ʼ�5i�g�:�B�#]�yR�[=w���D���Q����R��yrᜦG��8xv��P����Vā�yRW�2�lX �ޚ<�ҀV����y Q�R�T����2-״]�T���y�·�$��1Y��<L��A�Հ�yB�D�@@VD���Z�>��h��M�&�yR���HM���.�d	�⃊�y�.X3^GB<3�O�!�KX�j9��ʓr B�XQ�@�0Eи"P�B�t(C䉏 ^���G�<}��! .��4C䉸`<0(r� ]5����v��k#C�ɵ>��	��D�)-��Y4J׿C�ɴo�.́��rT�y�h�39C�I�q�*�ї$Y i�@��.�8V�B�	�4�6�H�,�}�l��-��x(B䉥pD�ѱQ��&P9���r�B��ui ��dB �����/�:��C�I:(�0�{�Iȑr�5RaƐ��C�	�V j�*����&f�
JC�� �hł'��`��싣�C�~C�	,���@ܡ+%pM�bJf9$C�	�[���c�h4�(�&�@��B�,\o.	�4�Zm�l_�EPC�Ɋ.�5��ۚv*u���܁p��B䉝Q���Y��̬7z�Rq
5��B�I�(�@��m��v�����&�8zΰB䉐���Ċ	|�<��E,� -�B�;�J����6\[��#ǃ���C�I�,q�$CF��}��[*)erB�	�6����M�>{xY�,הRIC䉽|L��S�N[s��SH��B�	�	��x�cMZ��d��jQj�C�I�h�|�	�\��D\`%��eC�I1O����0U�<","��H�	Q*C�)� �x�S��W��Q�7AםuH���%"O.<�gO>��ey� Дv_RŐ�"OH�0���\#����HGB5X��"O���Y��^]X�F�%.8��s"OI��燙@SX����1�H�p"OxI���=_P�`cZR�|Y�4"O�Jf��|�X�B��J��`�pD"OP�y�\	��B�K?Jþ�u"O�$��%Z;V��U�2\��h��yR�S�^
Q�1jA,_<��c���y�̆�b��``2aFH�������?�y�`8zh��;� Z�=м��CЀ�y�϶C�l0�ըߌ?!����A��y���d*���S)B�+�"��)�yrk�<����v J .��8�hȌ�yB��*6y(�*�	E1%��KC$�yb��;ަ�@�?�ёP�9�yRmӦt�	�"�7Vi�0�@ �y��	
x����(zi�1�҆ ;�yRc {���a�Xf�Ĳ��y�喃uj�Ai��G8����+�,�yRB�) �X	 fMp�b��5�y��Ȳ6z����W�,��  #f�%�y2����ʩ1s*&/�,�r.�y2�R���v��0��X�"c��y�D�� k�ؑ0D�;�yiWn�4�y�6DE�h��X�4x�����y����J��åM)�T� ��۶�y2	�}$\+�K�r���+��P��yr�ݘv��P�I�%m����.T.�y�#ܫ0�]K����$��N�6�y�߹.N�C`�	��P�a ��yr��L���b��9�x���y�E
"��`{��IX��ͭ�y/�:4Q� �D�����.�y2�$[B �ca��L3�I��y2�� j� 5p��D�Z-�Z���y�D�@��F�'��a�ŪX�y���	^�H���G��B�Z��Z��y�/ kx���!T�x�V�ڔ�(�y�o��g��d{!�G�"��A��m��y�I��J���5'I! [�,�A
Y��ydV�L��(2F @#V>|a�Z��yB/G�+��M]�fX(|�0�N��yr��Er ���QPz)�B��y�]2�2e;��-_��A0D�yR�3�أ���/q��u�O-�y"cM�4/����`�e��׷�y����XX�G�i��8�����y�+�k.��Ӗ	��,$��A�y2 
�{0���7F�W`@!��U��y"iK�0i����&�`a���y�b3g�����F�gSH�Z�k�?�yBcSQ%ȡ����P���񔦜��y"NU�^Jm�E���E��i�M���y@�?:N�	�bNC�EM8�@��'�yB�ǁsV��Piޤ1�PC��"�y��D:;nM�u�M�+B��2�#T��yB�Vh
Y%@�'s����E�:�y������2G�ĆH�	�U��y��$}���q��g�j��FI��y�#(Jr�@���]	d��H���yR�ÎU�BѨtOH�ag
�aF�Y��yR��SF����Tg#��{�o\:�y
� ��x%�8FW�]{u��c�@1"O��G��55��2�鈄n�U�a"O��d�ݮw��2�����'"OBTB4�,��@�r�B�r�"O�)�$	[�^���0n��~n��"O
0�R�Ța�����o���{�"O:`ڡ�
�W0$�j�L�u����`"O��B��JN���O��"O %� 	46��1瘁X�"O6P���0<H�����za"��4"O4,���.9���Ӷ
�QP���v"O��d"�0�]��c� �XA�`"O%�0���
�c#�R v`�M�d"O~��g�C�E��ي��N4	nZQˤ"O�`�A�S|�I6Cɴ-A�G"O�0�Ҍ��|�&������0�l��"OT]��>V$�U➗_9N��"O��l�U�����AT�T�x��"O��"�>(p%`����KF"ON�c��Q
������>��|t"O|���k�.:p1W�T�ty�
�"O �c0��"<b�$p��Oa��A+t"O�Ј���
��  iS%c�̹�"O���e� -�̐�U	��x5�X�"OʝyQ^�AE!�8B�h�"O����c��]���L�h""O�u���Q;l��R�`8'Ģ�C�"O��1�K���1�/Ɉ'/�ex�"O����a%Z��3��C�f:�"O�I�ee��ڈA��\
)dDx�"Oư���I�m�$�{�`Z{MB�A"O�0�AL�/�	� ų|"��%"O�t��'W"p��O���<��b"O���%�Z)�Q%MC��b�"O��h�OI�>����ΜU (��"OtM�G
�3���0���*�t�"O( X��Ӓ\��i�c`�4d\�ӡ"OH SUKU�9�\��O��2���p"O��Ap�O8��\�sN�дJG"O�8�Z�n����������bP"Oΐ�7��&4�z(!&K$w�p��p"O�I��BC�C} ��ݦ6�¹Cb"O�]R#�Ӌm��pS�5{�~�	�"O��s���m(�8���M�uJ "O�|�C Hen]�H]�_�l��"O��P���u!����S"OJS�
D#I����	�j�|�
�"ON�JkH�?'�KǈY5_��9�q"OJ���L��l<̘��̄�O7D)��"OԀ9�(k�� ��H�(@a"Ox�2�%>�L,��#ϣ,bJ1�u"O@SS�?d�#��7#�����"O�u�$�H��Qz��٘�|H�W"O����yF�=K���s&"O~�3V%ξ!݀�Ʌ
_�G�0�p�"O0%@v*��N�+8��8�)�e�<I�Cv ��ٷ焀M���BG�\�<�lۇJ�^��a@M��Ҵ#��s�<�2X47�U�P� �u���Rb�w�<�Y'[�4`2�� (V���a��r�<�ADC�%@��!߁H䠰)�E�<� %��.GVA@#�D-�=Y�CK�<y�M�?����nܛ#ȵ��*_~�<y�J�C��-9�-E'�,-�Rd�G�<� �LaG����X�`-Z;���C"O�\iV.׿X6�(UjF�Q�J��'N��i4hg�*�"�*#Z �`�'5Z�ɕ���T�`8�l�@�Q�'����'NR�h�rL��a=����'�����,/hEc��c�V���'��u�ca����є'Y�Cx�|;�'�<�R%@?l���X� 2]nū
�'~�M�3`�7unH8&.�+9\��'��ٸ�c� ���?L̸��'��A4ǝ���@�O1i|I�'�-٧� i�~�!�*C-c�$5��'��]�g�й>�5�G�^�B;�}h�'ix��Ѕ�\��%�W���B����'>�-"'�n�Hy+�V0��*
�'��H���O�tu���Ե3h�#	�'��<��!� x��	�P$�
]�(���'�r=��@�1��*woFn@�'�2�s�T1A�j}����$1�����'�ҭ����]%DH婄I.�'lh����ٗNH����Y'}���c�'æa�V]�Wx6��7� q.��'�Eɱ�i6�@R-H�=m�<2�'F�5��G!9T�+q�(.�h��'��0��J�+�N��`�Q1��'64�--�в�N(i� ���M\|�<!'ʆ�h���)���8Ʋ�[�KB�<A��� ��U#� �"?���qD��l�<�b��f̚��E�tHy��u�<��*1�0S&��*�첢,�u�<iA��B�6xsr*C�0���_s�<)��M�d�ڜత�L?r��"��m�<��(�P��,q�+�	<������v�<ybᅸU�z1�u�=d�Lr��m�<q�BU�OK2Ÿ�aUV�l�S�Sf�<� �N&]-���0��C�0���g�<Q&��1�L�O�2(�!)bbWa�<�Ԃ�q48b'�S-@��U�@�TX�<Aª�=n2��z��K�3!�	[�<A�bR3V�a��^�3�8�(���]�<uO�\�l��	W�tjt�XDa�R�<��K��^��EjC-heR�����Q�<��>cʾ�j'�]1?�`� �^I�<�5������&�^j�4��cL�<��L���8��!�̒�@��!eO�<��k7eA��H�"Hy���ZI�<��-�Zv�Cg&��?�t��UB�<�v)A�4�P(ƭ��I��Rt�K�<�*�'�X��F	{9�,:3�K�<q��ۇd�h�
��U�l4�D���N�<)��H�L�j���#�J �NA�<�ŉ�?Ӱ�P>N��Ñ
�C�<�⎝_c���
,xeK�OPq�<�4�R/2r8�6�L�w�8�0��l�<uM�d�t�H�M/k��] 0�k�<�saƙ~��J�'�CRHT�iX�<9����qkЍk.���MS�<iP��?��D{ao��Lj�=�+�M�<y+��o��:�#M/�:9c� N�<9���s�Tz�B�p���נNQ�<�$a߰e�*Q+f���~����u� `�<����T�B�����/7�`�E�^�<1aԻ*�|�����hӊ��%LT�<��oɹ?���3�P$``�q`�R�<� �I%رJ��C2)-vV k�"O�A��`�$ �V�w�I�~&�"O\�)��;a�!����	�(a"O:D���@"�@R�H;n�h��"Ox-{�"��`w�M�$!R!��0�"O���Nk�@��1 ͸i��0"O�<	f�.B�n-�0�~pt�b"O��X#j��V����� _�<	�g"O@3����@�0cI�1N딘��"O����ĸk�h��i��ղa0�"OLir홋]k��ˁ���n��8��"OΥ��Я]�����D�N�z�"O>m�A�	Gtb͛�m��\j�mp"O�� �Q���i��+Y��R5"O���d+�#nt����8���"O*��!�Y�Ni�u	�/%�H�d"O��G�_zP�iY+�<`b�"O~d�B�����
2hZQ^躁"OJM+a'��6���V#$Y<Es6"O�0�O�oԅ"J�4@[����"Oj�C�
.K��`
�7���"O΁�Fi�}#������{�"O:}�°=��X0s�"�0�"O^��6�� F�0����a3U"OrD+э�-2���h�왩r�f`)2"O�y��`�@U蚂\;*5�d"O4TX���7/�,��ҡk*��A"O����N�:� ���(9'�<�K�"O"d�È֒JS¹�&�ؑz�,�S"O��S�CF_����π �T�0�"O��郜sR��� �=��+�"O�@�u��h>��v��13��a*"O�M��➆�D�W�M��T��"O&u��W�,2�]�9���p�"O�� �*X�$���7D�C�Xy�"O��Q������K#C��2a�=9"O=P��I^����	S_g�-�`"OL}�@���~W��b(��]I�:4"OD��T�OU��z���^��0�"OtA��f�(H)�Q�ϮnvDt��"O�d�d EP��  T1Q֚H��"O������a���&Γ/�T���"O�d#���y[L�Qr�n���)�"O�U0#՛xt�#�!i�q@�"OLa!�$Թ��d2pC��(�4��"O,P��H$��j��S�4���"Ot4�5`Y(�p�Λ>���	 "On$��n�&���BDm��jbЇȓ M�Et��6��U�S�03�L�ȓNÄX*���,bŚ��bᗰ �v��ȓ�m�!�N�@�A�I�:E�!�>D����`ސ���_���e*�">�:��F�D�(N������*~��K���(���'��yZڴ~�đ蟌ꄙ?Y��M3���4�jt2�Ǟ=eެ���MS~rH�O�]�=E��F
�>�̤cs!C;t�,S�ķ�y��O0��=E�d*@7Z���� �j؂�!Ag���M�V1�S�Ov�t�fc�!m��%��n��au�I��0|J��F�i����>Jj��$Gd�Z3�<�{~⫞<ZL��b�V�CL�0A�ύ��$���b?M;�.X�C��9H�'Me6pE��<����Z��`�Ƈ�NĠH��ȁ�{Ժ��.�S�OP�Q֭����Mj�杋��*��� SDU 7W&-A@��h��,�s�\Oy��O��)�'t���څ�J���ǧK�9K:l���~r�O��S�π p]�Џ����`�px���"�u?ɏ���3\���@�.b�t�l�q?���5�S�O*,5��@ r\�(�1+/c:@p���%�@M*T���g`���Dۯ6��4��?ړ|~�0r[�#F2[)½S��׽i��O��Gz����*MT����:�9P�Ξ1�����(O�>�J�D��h��!�\�P��f�>ph�����?�>h!�6_�.$���Ft�L|Dy��$�'(����0`)@�1x̸q��LD�~��<���'|�b>��C
@���`"��#��2�??�T�'F(� �Q~q��R��V�A!J����k�&zqU��H�mtΓ�dm����BH C� Kˌ�0`�P+�"O��9 �qy���R�^201V-�7"O@�H��X�W�ܝK��[�(�"O�(r��!&�9a�F1K{Hl2T"O�ZP�T-\���vN�2�Z�ٖ"Ov1����r],�E-���TP�"OJ��S�,�~E�7*F�Yv�4 "OJ)d�M�9j��h��DXzT��"O�,A�Û(A�d;A�PR�#�"O� 0�KY6�rŦ�O4��r"OQ�Dm�
�m�Q ��'�`��"O8�����j~��qNӄ-�����"OBH���6��	P6G��k�*�*�"O��Y��H�S*ܘjB��?��c"O����vU��
�\�^��Q"O��x�(��=�ʹ$)؍T�B�i�"Om���v��Ũ$XK�e��"OJ���L�P(�`�6ȉ�D�|!І"O�h�C�K"�Dƍ�xx��W"O�!��-�=>�x+��3e���7"OHh�E��v �-�B�R,K^�p"O�Ii cV��(<a -�(=���@�"O��a�d5DY���^���"O |��kJ-!0l�M��(���"O���r��+�X�T�	L|�Zc"O��X*[�W/����کzd�h"6"O8�ˢKH+v�4�/��A4��C"OTH�7���.ľ@k�d�%g%����"OzD�u�-^ٶ�@���,oH)�#"O�l+��"R�@{"c�}Y����"O�R�9:x()xT#�\�LS�"ODZ5
��BOB`Y��,\�̩b"O�t�fS66�9�HO�
��u"ORR�M�F��`s�\�wO\���"O���!�C�zF��i�"_�J����"O08�f�G��<Q��,���$"O�yd��è�:����&�(b"O&h:�J9huZ#	|h��k�"O4��k(r<z���©d0��J�"ON�� �<.x����&�$i"O��iu��l�V4��㎥F�&x�"O�z%���r*ne�(�r`I�"O�d��0Q�&�yWe�*?p���
�'��U�&
�C?v8�R�B~�l��'�a��-�~H����F�'�< �'�����O8P�8x;䍀�$�8���'�d��!%),�}Z��Й	V��K�'�2�X��ȧO���B��̝��'B(��C�F�,^" #L��(�I	�'�Z雇G�R;0�)Bc[�tx��*�' I��L�2�eH�EϬl��)	�'�����S>PRr�)bCI%^���'-ȁa�C�g`�k��VTD�
��� �T�E�$��)�ì��~�(V"O8�J����-dҵ넯Bjr)��"O4��%d��<�H�k*z.�(;�"OV�;��H��$� Qz|)
W"O���f���]��u
w��2Qk�l)�"O�Y��FZ#eW���@��4=g�H�"O@yRU,(3���0Gl�`�a"O�\�b`X}"��o�QNI�"O �`e��9�P��	r�F��"O8x�f�&V�J1�d�ȩ9��3"OJ�JB%o���2 ��s!��Qt"Ob��l�?P�����d�
��9`"O��S���n�i�$Ҵ��	c�"O�a���:?��A�(�[-��,�y"&K�l����gOo��p��y򦐘` �ٚ��C�g�j�r����y�ŉ��8rF$ֽb�Јn�-�y2̄:�0퀄.S!0���P�y�l�\ڌ;&]@�8	�vkś�y��]1FX������;�Խ���y�hS8pd���f��(Ժ�)U���y�hNT��sG&E% (^�j��H��y�oX�fxP���
�0	"�LŇ�y�% �T��yT�W�^�2��B����yb�L3>�3b�Б(���y�I�?�yG�Y,��,����@��/�y�ȟ2�rd8��H��X-�O�y�4}��	P�$�!$�fy!�#-�N�2m1J�d�!��$B!�R N���dM��<R��T�5!�V�>'2-��lިG�8d�RdZ*!� �]s�&вOʂYX��(C!��vRLy#�՟'��`��6!���AV|���
K�F����äU�!�X:I�$T�2�;��aR����!��Өq��p�B'W��x�(��ׇ�!�D�!{u�cӁ�(q���!��"t �	p��1�7��!�!���
���H�t���3��K*`!�Ԏ\"(QUB��<i��	M�RM!�$G�;
1�7�=n
�IDC
�\J!�dS�J����n�\j��bwT!�$#I�|9u��gK��bOD�c!��Km"�6B��Q�܁���+d�!��^��IsDK��o�v�+�Nݺ!򤐔(�,غ�D
�+n)i7�#!��_�mjRd{v��'X
a욮$!�D�y:p���D�ZՄ�	3��!o�!�ę�;�5�a���($!ꎾC�!��Q2�����X����!��w�0mY�Gg�`���	�B�!�$/x+zTY7EA�w T��V�!�ȕ�̔�j�W�-�H+@q!��H�n�
T,�#���.�!�ڎn� A��/H
'�d�cw헨;�!���N�@BUf�49��1P���0*�!�$_>ZgX�(8z�
�g�� St!�$�y�:u��/�9��59AU�&@!�Dӱ8���5��C�TE#�AҩE)!�E3�4�r�T�@��̀�܎{�!�䋯q,b8��-V�rQ*F�ŠB�!�L�F�{�Γ����r��.rV!�D�$�ܱ1��ΉR�	s�ȪO!�$^�>�$ԃ�*��C�\�H�*6n!�� ̡����J�%�T�>K��A�W"Ob@�U�F)#F|9��r	8%�0"O�!`�*=
~Dc���4U_ά �"O�h�iد hȐ��@Z�V>x�"ORY�7ϐ�W��@Ԯ�0d�dp"O�iR1d ��u����g����"OX��ML�j�4���X;c,@AE"Of]��O��ϥd�]��`�PCϱ�yB'�Y��I6�4PЄD<�y��:�����.]�kU\K�Ϭ�yB):z�\���as�����A��y�MΒ@�=#�\�f�qJ��y]C��@�T7�εq�Z�y"m��k ���E����-Ч
O	�y2(����ٱI�jtYw9�y��#Z�����4��Գec ��yһ�n1!!,�1h���8�@U�xk�B�t�6�d��'� ;�6aI�B�	�5�^��6�?EJ��i� B�	:�6DICH��vMk�a*�@C�In��1�u�Z8)��+1��̀C�0ⰽ�u�R<4�x��T>C�I�<���q	D���Ѣ�/�C�	P�Mz�g^�~�4��&!L-2��B��(I^,5;��<d�H,��>[��B�	�Y�~X:�$�\��ꇽS��B��$X}�$�3�k�t��l�urB�I�pn��(�,��H�)�W��e��B�ɵ%��@u�3_���s�ܘWw�B�I�}�0�5ʃ�^��Su�6dH�B�	�ظh)�MZ�f�f�C/@�"��ȓ|r�뵈J�#sN�hP�ެ8����ȓ"���P ,��%h���NҨ~lZŅ�op�I*,��`��� �L�ȓ�xl�3B�Tp�� @ē8����L#����<������W2L���]7*� #K�|԰�i�Q�A�i��D���P��C����Ǘ�l�:	��� x�7 �(|IH	�쌬?�4؅ȓQe|��M�:���eÃ!'d���S�b��_?R��sp��?g�݄ȓ�m��o#��1�ջZ�j��5ұ#6O��/�,��t�5a
��ȓ��H���5�4�HA�S�'����/���k��X�)E�I,b`켅ȓ��������U��8�	�E��P`1�M���F�F��!�T�ȓE�Dhq�m�//ߌ4���)L�����q�X ĩ@�iTZd�˃(r���ȓKk� ���ړZ�عx�$��>�H	��1�X�@��Y�>���ȕ`D�L�xC�I8n۰u��C�,�rX�qMǚB��!{��c�jԤ0Odz���kAHB�	�m�(<˲h�+҈5��g��B䉦/�:Hyb�N# �R�4�:o?�B��/^�ޅ���Śn�ܭ�0�(�B�I��ܹ��f�8(_�Y�ȋ�obB�I�p�DU�5� �t���K�).*>B�I;,r�14b#UΠ� ��	�R)pB�	!��I�.K%>	R�(�Ƅ�"B���ܸQ�Ń`�X1�D��׮B�I�AO�8@�n�OzB���F�'C�C䉡Qǎzv��9^�Ƙ�C�$J9`C�	.e�ɠ��%�L1p���q�B�)� J�(S'��&0rED��Gbd8�A"O��z� �.8�([�F�Uy�`CB"O����<aHY�@C�y��4�"O��6FìZ9]	�H�!�N��"O�	�Qn<Z��0��g�`"O�9Cq�H�)&�H��svTe�c"O�xJG�;|�>���{��}  "O����!ˠrS��*�
ԗ��̘"OZ���D�,*T��C���	"O�0r
J:2��$��)W(�����"O��Q'�[���1�R���3d"OL q�d֓���[�A]jR�K"Ob`��b,���
��=j�A�"O2Ep5I!w�������tL��"O�=
w��-��!������4�v"O�����.����%e{���
�'m�}#  ���   �  ~  �  1  �'  �1  8  `>  �D  �J  0Q  sW  �]  �c  @j  �p  �v  
}  M�  ��  ӏ  �  X�  ��  �  _�  ��  ��  ��  -�  p�  ��  0�  o�  ��  J�   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6�F{��'n��2i�'��L���LK��!�'NHɗ�@�x����F/�h��'ƚX
��[T�x­V��q�'"�����X���22R;S�����'(<�1���$h"�N�4..�r
�'�4����!A�U��;)�XQ!
�'���{�V��&�I�f%��j�''�D��#ȭD��qUB���8�'��8C0iY�=���(�+��$.,O��C��=�6tJ�$ҋ�^�!"O�%V�E�d��R
�DČ�(�"O��A�a�7��BR�G�9��@r�"Oj��;NA��J�b٤|�H�1e"O�%�->UD��0!��Ј���0�ŞC�}
�J�'YV���[��D�ȓkG�B�ጐ����H<¬a�ȓ4�����
߳!���q��;^.�1�ȓb���b���0���QM7X�h��ȓmDx0�ĭ@-պT�q Ĳ7&�X��	T�'VQ#�@;J�>��6B�p�D�	
�'�Lɪ� ՝%~���X�l9*���'�l�J���0U0P`"��&M����ēقt�gO�Sq�mY��ߟg��ȓD?�P�@�Ցr����c�\���ȓo�X�������?�. ��'�����<)0T�G@!Va���� tm�t�t��� ��[�5��l�"Of��Ѿ� ��b\5i攅q!�>�S�S�y|�"Q�ݺWH�H{#	������6?��b�B����[5|^��´�W�'�ay�C��B�bd E�c1�yd����xJ64�|S"R�)���q��1	|bO�|�c/�F���`�,ܕ|t!��'-��%�x	��5c���1D����:B`*D�̣�nEW��c�`�?0ݘ@C���O������Ɛ�6bP;Fr�D[C��9)��C�	�@�0��qK_#x��Hf��o�Т=i�-Zf�{S�� w4$�#V`�j��Ɠl�1ڐ���j��=(VI�#Z��E3�'L�����+^Hq��MVh�]���_�>�R�<����O�9 �ƮrF ��4G*��,�e"O�<�f��6��q��3Nn��@�Oz��DޓC�����`��D����E�y��{��8�E����@^�h���\�8�!��}��)@m�:j.�(�R�Jġ�I���41n1�j�wL
��C䉱fH�g��#u@�
!"W�\7n��d"�d�+Gk�M�eǥb���f��!��߁�Đs#��#yJ}�Aj9+��>����_�7NQa�K�Miʔ���U�b!!�$�s�h�7%M�uRh�H�h�	C�!�d�u
�\���&OK!�@�Zl�!�d�j�n�x���sc��Z�{.�B�I�~U�-[�L3Ix�p��ք~�8��d6�Ƀ)>usd5YLH�Y��S���C�I�=������.mEv"u P?L8�듅M��O;`����F;�8��È˚Y{x����qa��\�"�%h��?���'�it��z�t�	��X�Ta(���'-�ʆ�y�v�c�I�b5�y��HH-�y"\��`T@B�-j��r$-̦E{J?E�=���C�Z@\��� H�1�0l:�)Cw�<��+�:�h5y���7��RC�Z}ў���˖��F��9M��%�jЬg�XC䉌!�Z���CҰW��A�BL�ljB�Ɉ?t���<E�|A���K�:�4B�	�6|���D�,am|=�-�!�XB�Ir|r�Y�"[����4B�� ;"�B�i�2	�y0ƍЂS�B�IH@���f% �e�$�Z#T+B�?�XI@��Qjd��13���C�I�W����Q:v
F!��m\=H�xB��2�@2�C��0�A$mœ-?�B�	�$W&L��䁝�<h�׬�>c�B�IB+B��6oߞ�:� ��	�+�C��64Q�H��T�s哫(�C�ɽbh�h [��<�sG N�C䉣p��Ef �Wv�p�E֢"�C�IO@!c�,̣0rd��e+U&-b�C�	���킃E�	b8C��P�9�ZB�	97f�sb@LFP$�BB�J�<c�C䉴}�3���
I�ʌ�u�I�B��6L��s��nK��j��Ɠ��B�7C3x<�S����x�����KhB�ɹd\<�X������ ɓlP�6B�	�H!�H��Y�D���%��B䉠!�`m�ҥ˯�(��0���J�B�	�l����GɆ��q�/�,�B�	Y�]+G�8u(��[C&V�d4�B�I�~�~�w�)ʽ��LهxZ�C�)� `��`��7�L��cMG?M�1e"Oz���ܴ5GZ$UTM���9�"O�)��@�}����GL�5��8�"O͛!��7\���Q˄Z��-�$"O"5R+�b���`�ǘh|b��4"O����M/\Q��5iW,��""O��)�`ȉF1�I�%��'K8�f"O<4H&��7 �V<SԡT<uN����"O���g�(5�b���=��{�"Od�!`��t Ϝ٤̨�"O���4C��8��i���[;	��a�J�<93��`w�ɇmD�Ҥ�AJ�E�<IAcĴ1���I�'��o�5U�^J�<YÃ�>G/.=��X8֠! O@b�<�����%؏5��A󋍏;�C�ɚ�쨋3L���bh���J]��B�I	`	B9S�"S,$:��5脅g��B�I�6y�=³�L�Pyt��5(��B�ɖ
��a��@�|�DW(0��8��"OT%�s�F;rE���Q\oT���"O��EK"�"%�����]����"OpAJb+t����!NAD��"O���7d�+vE�EDI�w�X�0"O0C2%�0�>��S� c���'"O���C޵d7|�RbL5SL�H��'ʹp� ��Jr��tB�)�T�1�'S*�bƎ�(	��Ic�C>�'�]E(��W)�d����*���'�Fa��Ḧ5:&4�Pn	~�2$��'���B�L��i| I�Ul[�y_� �'�TaPf�͓~	�Q��n�\t�
�'��%狗^����E��nʴ��'�hd3�����1&@Fm��`r�'l���§W<�ځ���C^5�$��'����Ƥ%sM�D��*ϧz�p��'5�E��gA$�����~Μɓ�'��҈٘�x�F+zz �@�'�"��&+R�s[֭6ĝ>\��'����N1gU���(�Lq��'W�	@S�:?�lX1�Lǧ8Ǝ�i�'�4ZT�Q=6rB���H�&<��A�''K�9N2���C6c�š���n�<A��?}Bf�:&��:]:^��!-�T�<"!��^�l��U�Q�$a��h�<Iׇ�:Jjl����P|d`A�3D��y���y����O�S�Z��p�0D�����+G��%��M�op��d/D���W8����jIrżؐ�.D���k� f��؀��()-�,Pa�.D���Q�*xF��ŮB�Z�r���c?D��3Đ
��\�����w"2��WC<D�����5C@����".�(B�0D�$C6)����U�	2q���-D�<�/+���ڠ�9U��k��.D� x�eQ�,p��3v�W�I��A[UB,D��hR��c��u�{�n%0��(D���LG$A��]Sgc&|sR�H��%D������.�v��U���i�T!D�����T%9\�b�	Օ5�6�
��=D�PP ũe�扑&IӐF�c�<D�<8����I҃
S0��U; .D�8��a�<��G���f������,D�<i񮈌Rbz�QT�̴-�0`m D���fm�sS�7��x�4= 1�8D�� REc� �\�.H��iL�0�Y[�"O�Z�� ܰ���iI�U|�%Yc"O��!�@�T�j)	�'\�uBd��$"O��qӉ��7��Rw&��(�"Oxt��HF8$�ʕ#���P������'��	����i>��	�����l�ɫ,C���%� ���[�JZ?3?��	���	����IƟ4��������@�I�c�P��b�V�Y�LǸ�����	ԟ���ß�����������ɍ,�*����[5z��p�P1Hh=��ȟ ����	����(����I@q�+�mD)��hvā%J:��	�`�I��L���T������	�����MQ�	f�X�jTx,s%�ɻru$���ן��	������h��Οt�I����Irt4@qGBP,�~���K�
:����۟p��ǟ���៨��şH�Iȟ(�I�Ye��`i]B���scϦy�` ��ϟ �Iǟx������П@�I��	(��<��� N^B�pVOѪ'v��	̟��������؟��I��\�I蟸���Y�PpKN��;����C]#��9���<�	̟ �Iҟ�	������I�Y���䝨 �`t����4�X����|���d�I����	埬���0�	<A�
e7k*_�6��2�$Y������Iן�I�����@���p�	6�E+7��(EH�lq#d�C�x����|�	ȟ��	ʟ��	ǟ�{�4�?q�6����C��_T�[&�N-W\ђ6X���\y���OBemZ�'�(9����*�8	�d�B4|ZhEy�2?���i��O�9O"9mZ�L���SS��(A�M�9�v1�ܴ�?���I�v��͓�?�a�ȥTl��$'�Z~R)� ��H*��V�>R�8c�˘'S�^��G�T�BZ�xD�+L�<����4JVh6���)�1O��?5������-=�*U��iH8��D(8Q���kqӒ�R}�����%p�'BLh{rO6`�t�����d��'���yv
}l�y���i>�I64+&	�`>U���C��n��PyҞ|&hӐ��e�7(��t �9U�4�rA�4+��
�OjoZ8�MӘ'����_�3��A�A�td�E�ǷL�j�M�b�0W`H*����|�� I)�H���S�ڭ��� ��8u��7rQ�u2-O�ʓ�?E��'���S@'��!-A�R
os>��'V�7-��: �	��M���Og@]��OJ-(�L�G
K*-��';�6MЦQ�I �Ȥu-*?�#ш�0c�Зfm�PJB�2�q���	��iaN>�.O�	�O��$�OL���O��V+˹D�t�����'�l�q�<�@�i���8�'hr�'>��y+�1,�4s��z�@D���^p���0��(h����	\���?��ӛVy� �
R�3 �/��mܺ}���U����X����#ݾ-^�+͜�u(�4m����3�ӗT��	Bv(B�I-�����V�,l!�DN�G��1�w䂷!Z��(�J��k@�O���D�ȝ;���3@o�hL���a��-B���YCI]�5����gLܝ{?]���S�/482�	w���Y7�Ӡr��%+3N��d��JчOW�K���s�M��L����F�kT�@� bs������^�F����Y.g��{�D��DW�Բ�Ä�q�ֹ"BK�<N�F�
��H�u╠v[��@��/1�H��?���?1O>��;���O�j�(�,vnd��6���u��1y�4�?1��?9��_��;x�zخ�|���E��:�(Xe�Ah"ـq&6��O���,���O�p$�i	F�{F��q�B�T]1,౸ߴ�?���ĺT�0%>��I�?�{B��tF6+� I�#�����M[M>	�'���k��?����?)��{RP!r�D�q,P�!I_!F7-�O����D��,mZ�����O��	R~��/��Y�'�K0=����$�
�M����?P�"�?Y��?��\c`e1r�Y"%��a�C��0)��4(Z�	ۓ�iJB�'	��O��O�7V �R����.jP�Lވ@WJ]oڵ$,5�?	�g��?	ի�-Q%`����� �JA�Iě��'��'�<D���8�Iȟ���g��(�QĒ/!I�ˀbޯ.4��>�F�A̓�?	��?A��I;3nN-APf��Q�zi�ƅ[9��v�'4�"�e5�4���d�O��'n	r4���*��&��n?Խ{�O��)��d�O����OL�c:(�A���kJTH����7�*��V�e'�'j��'��'k��'<�r`��%��P�-��\պ#����'���'�"Z>-�I<Y��O-�)�>od�Ѭ+y����O����Ox��=���OV��R?�j��Xq̵P�A��ke��P��>����?����T�@��$>�8�ߞR�HY�#M��<hC�k�6�M���?(O��d�O^�Ӱ��O��O��<�7!ƞ$u@���k��Z*�5�ߴ�?�*O.�$�?2k��'�?	����1
8�%��h&�����M v�D�'�,��ڟ(���w�	[�I����̪$�>2�^Y꒥��?��	埠u#ڟ\��ɟ<�	�?���ug$�U�L�8Ǚ�Ff����M���?�v'
���(��Ź�&�_��-��B�]y��ײia�zCdq���d�O�����X!&���4qp��D)�"��mpeƕ�7#����4Mr�p(���?����?����򙟜��G�O��*3 ��O��X�g��,�M���?q�Af�m�r�x�O���'�>Ѩ�G�mC�S97��\��y����O���:V��=���d�O��O�? ��D2@}m�Κ�� H�i�B��*��O��O����<��4������nP�!�Ф�)�6�O�x�Q��O�ʓ�?���?	+O�sa�
>Mm�TBa�1V��t[Q�A�x�'���Iԟ���Yy2�'P�n�H| mУ�ǂzlUi�"�q(|(J%�'��ɊSc<UExJ?ax�l)n���U�Qrb�v�*D�(q�
_�x�x��6	O~�(� $�	'=nsp���P���c��'��ВbD7	;�Ȩe��7cf�ux�	T4I���
4���7є-�&�Y��x3�˷v���P��-Wf�9BY*u�h,˷����D�ҥ���U7���G�F�{��!$�k@t��5��snZ+g�� n@�9%c�3eU4\�$L/Oh�L��B�9f?��$Ϻ+���2n��`�@�#����O�a�uI�[@��&��&B$nZ���i�|r�
LJ q�� P]��`�QJ�B��;.����*!'�(a��\���B��xR�y#�"�&��`R&$(����!�ٲ<�}�O��kC�O"�D�O��=�CD J֣�)^H�D���A��b��	sx��h �P�Re"���nԀScHD���$�?�u��T8�.��iQ`)SQ�� c
��7�i&��'R����L���'���'��wEXNr�(SS!=*���Qd�T+�]c��C�{|��|)��AA�|2�ՃR�hy��b�#?ҵ�C�,����Z�mFذ* ��3v^������xr�R4d
����� �<`�o"��a�.�O���Ot�d����qU٩��ՑF��� ."D�0S� ]�U[т6�2���)??QA�I5�Mk�����	��$�3�C6q�L�	ªK�-�a�u.��^$��O,�D�O� �;�?���?�FEZ"v4đ��%Z��E ����M(�[D�V�S}&9I��ꍆ�m2NP��E(s�X���.@�9�Ң��$k[�D����K���`r`/ړ<;V� #�5"�(�˳�U.(!�5
�џڴ ⛆�'F�Iɟ��?A�f^#K�:$��C��آt	c愼�?����?a�L�����c�#t��4x5ٍM;�-�L>�Ӎ���|r?�;=�NI�8����՘P����]遦�k�t�3�KO
��ȓ�|pFF:j3j�b�RV)�ȓ{9*�L�@%`��7OFy�ȓ0J"�ЅfbxQ8C�H� �r	�ȓ1��|@tEQ� 6����1�R���`�lY��lU6j��P���2��]��F�qc ��W�rP�ԌN����ȓ;��9�Q�@��Rc �O�!�,1�ȓ��ڣjú}���Þ>��d�ȓ&�5��ǂF5v@*�J�4��ȓSm�����\o25�3kV��.̈́ȓ8&�=z!'%"*�!ֈLO����ȓ/�Z�Ѕ��+�dY
υ|�<���$�&��e��F�]I�CY����?�1	��Ϛ&�)ɵ�0c�e�ȓ}#�����Q�Yy�m�s�T$��h!h���Ξ�T����G�Os�4\�ȓA��|k�G:�pe�bf��n1�ȓ.�\�2��-X�pH�it	��8�U�pč��,����)PAxY��:�6���I�j2�8Cs��?|���ȓ��b��!0��������ug�I�ȓ���MFy��ң��>�4��ȓ{ �J���y[�m�t��`���ȓN\^T7*�-t0|�d���_t��ȓ�U�/C�f�А�������}�ЫhB��
E;T�_�*цȓ���CA�,W*á,Q�$pzE��\�ؐZ�bŪ9�h<�E"N��d�ȓe��s��)h"���LT�0_r݄��<��!@2\ިň�S6�(��ȓ�0$r�`�+an�P0+�"���"-z�p��� O �#E���f��(��L���	�/k��r��+%꤇ȓo8A�5�������� :������	��(��	�jo6��/�#%�� �C�4(�nC�I��L ˵�?fP���������~B��e�|�y�NU4��q���0=q�"��
F
ҧ� �t#ŏ�%���6ㅊt����"O,����E�aMt�g�ihԱ���)�԰Љ{��$v�����ȵQ���w!��y�aVE�����Ǉ
���ڢ��-�f�R��>��M�B���L (�~}�$�,�Ԛu>�;!$Be5z����soa|���3�<�yWb�_g@�bG��q<lhB�P����rDT ��˖T� $Z$��n8�4yU��
'���D�tN�ȅ�)\98k��D�U�N��U�:k(2��'�`��g�G8x���åB�	bj$��j(<Q�+Y�1`�n)w�l�ĎK
5:���i#Fm&�rƞ1*,8����� v:ر[&� (Q��sF�z�<�0�-��飐l�(e��`ub��k:㞌9��~>yBG�$�F(�Ҟ>A1�  �2�C4�~�S���w�'���B�����ᏸ�&�� ͆���g'�~��f��RlY��I:vθ���6k��Bl><�P�2lJ1=
�"<)�O��-V���.�z��c& }�kJD��D��/߼T��9��IC=����]�lxB���8^Ȱ `�H���1��TxZ��&H E�V�4�)�;W$(a�Ω$���LW>`1�$�ȓuI-�PMR= ��Z��R�0��lX�h!�I�#���ӥ*� �c���o�Y�|,Bu�*�8$���R7V� ��I-�����yeÏ
e1J��gJH�65�(#�'K�7�|�S�T8&��jWK�"��x�@@.� ���#�*5�u��On� ��Z�� #Dj,7��Ti�4��d-0@xF�'��)��ܣ/Y6���'��z��X� Uh��\�=��c�	ލ7��`��B�lN���L�&ɧ�9�n��B%�'W�=3P��Y�����"O4�
��3:a��☀u��HO�p� ��'k6��f>7m׬��:"h=}�.�"kf�jR�CO��	���0>A�l]���D��;el�����	�.xrQ��3,�dI�U�����U�KO���DR�Q[�H!#E*
�jxa���w=�O<�D~����z��ӈm����oPKd��G����m�A�ށn}����eu��k%Ƚ=��
%Α-J��pXR�;�	����A�`w���#$}bF�H$�KDkO%�m�4�^��ȓw�`P�):�z {�A�u�`oZ6L*"�#AZ/$/:	��w�)�����E�	�~I�w
�!P�����i{N 8(O2���I0zf$K�
U4�´!�#����t{µ#���x"i̺T��p怂�W̜�#������'{�)af`�D}��%/�8��|ZS�)N�X�壆#��|%d�3��p@���p?�fHNԁʅ���n�t@�Sdo����'5t��J��~�'5 r���?M�w X�g�H<�%x��ɿi�<���'�8�wO�;������
T���t���C�L���c�9�sGڦ�%��V��B'��X	�s$�0qʉ�c�2Tᠣ#lON8�t�G�j�tu��0}L���ҥ0Bb��A�"8�����.O,\',Y ,�7�=�L�>q�Θ�?O�y��L�WY@X7�p�����U#F�=1�Oe�\d��y���[d$�Y��+ɰ�:W+��c1}�AN�{��X��
ʺnM���(E�>¨Y�����*����lQ�R�'��5�~�O2�韔�λJ⺐�b%�1h��c+A:cԇȓH|F	�⇔I��9�A��t����O��	g?!^w#�S�K���� h[)�$��.lb���`X7����4Ν�T�a{"�JYƸQ�"G6[�؅�Q/N<0������ٮ��h�O��7�K����X�q&��U�	�z��Jf�W�:)�(��͒!)�$�X0 -�\u �m�1��2����<����8FL�7�B�� �\a�炑�#Dd�s��B8^t:V�қ+
�yq��q�d�*��U�#�.�D�7W_p��AVʟ��»k�*���ףbJB�Tjt�#A�S !�D�� 8�� !眚[|�=W��6z����R;��$)yg���g���*f�I�@�����-rSeE
6����d��j�R�c�&�" , �"�ҙ��z��."��H*W�i�(�{EA���� V㙄2�,�?9�&1�*!8�� ���L��o_V�'����v�	�T@t��!2�b8��O�xxǁ�	eݠ�s6�I�]�a�wD��7�H���X o�@I$X���"�@L p?������d�$	R�� ��T>�]>�-��X�|{`a����2SˀC��4���p�LG�-|q	�c˷'�lL1D�(��3��	��$�b�j�[0_۾ʓ���p���� ��.ƴG�L���I44��<pa�Ont���3�p����}k�����F'\:�9�-O������O��IP��s1�UK����R����F�ɸ(����'j��I�COI�TJ��F���o�?\V������?��9#5O� �M�C�I��$rw��2=x��D�}����{��d�W��"���>����<�y2�_�J�`"�S&`��p��,ާ7�������<�ԭӆ;�$��v*/z�^�*�+�x�<�
�)p�+K�#*��z�h�l�<�s�W:�U�bߔE#�Xa�"j�<҄�7T���$H�m^.Ѐ 'Ue�<��b[�Rnx���X�J
��:��|�<�����B�^;`��B4�y�<��)�4%{��D����R��[t�<�-U���"/�3	8؍��AKx�<y�厃/0x�2#푱$�(��`�j�<�N�hk
%��K�6d��T�6L�K�<���c�iC�O|�U�3��a�<Q��R>s�乊rL��i �q
�\�<)�ϒ=:�D��6�1�r�*��r�<�k%�"��a���S.��ڲ��E�<��LO�*S�gL��(��D�<��P�V{uR��fC�u���D�yBKE�P!zh��Q(l���GgU��y"�������F��#��9!��HV���p��9\��h����2�!�ڳT�t�6�q3F��U@ ���C�	(]ʨ�z�E��XP sa_$D��B��,1��Eر�N�=�|;tD�B�B�I#^�T��%\�4H� ��B�	��~�KTn�^k��G��,c^C�3��p��@�)4\�u;��?9��B�ɇ�6�x�ᛯ6]>��r"�9~� B�ɽ�j�	%��y�6ea4��>�C��d_`,X�mD6�*ٱ�ee9rB�I�'5�h���Z� �B��22��B�	�}'N�r$GF�p�0�^�x�C䉮9��A�J��@:�[!'P\C�	�d]��	3M΀m� ��/2�C��=[Zrܨ� ��+de�`�XvC�ɑ�╈�j��)��x���x�TC�I&2�̹z"hN36 !�d/B�d,C�I�~��y��aL1Rc$�i�K��7�HB�	29�Y�,��XU�	����$�C�ɾ��Uk֊$�M�v�9Je�C�j*p��gI�
��d��J�ZB䉶S�Qz$A�1O�"���P�R�B�I>�v�P3�9^�BK�}� B�ɷz;t�3���(B\���G�iw�C�	��QbS!�Bx���c�Fk��C�Ir���9��R�P馄�`+�*
RC䉴k\�,��`
	WF��q�G�
o%�C�~�$A$�^���*[�G��B�	�|4 B��I{�X%[f"ۻ��B�ɹ8���#E�I8� p�X�%��B�ɹBH� $G�x��̞$�B��.`�����mƷoO	���˯6�8C��o��XP�%�E$F�ZU�\��C�I,\��cd8b
�����P�B�	<���H��<!��2mǴ�C�.D����5fM:��C�Hc�E��,D���v�e��
A�3�~���8D�ȨҍN~�����bA�3�f�`��5D�T��YD`���Q%.�5�0D��8a�!	[�Eh)B-bR��UK.D����J��L�9�%�9� �!/D��5k'*����-L4 ��'�-D��a�*�
BLͨ�������/D�� R��R�nGN����@'"�LU+"O\�*���=zI6��5���O�:�8S"OJ�8�B�0(l��AC�7_P�b�"OL%�W.Hf��*��nn.�"OL1�3�Q'0���@茠~����"O����*R_���P_�UgJ�!�"O�|¶��,;X��hF28r
��R"O2�s҄ƃO2�I�GP�<�	B"OD|�6kXP�`Pfu\�B�"Ot�3�ǛE��lb&/�� c��0"O��˳��4�Jb��+H���"O�����C�fȀHx9�#�"O�YE<�\�ᘷv&��"O�	�/
"$p���:��"O�`� �;����c�3��p"OV�����^y6�br-�

*�`"Oy�&7�j��-!,t0W"O �;V�X26R(t�Gq&A��"ODu`qbۡYV�Q%]�6u\�ӓ"O" ��aU;@��gI!ofJ]i�"O(��%��8����fo��PXB"O>�`�T�9V�$c7��	�4a)�"O�D#Ud�>(�n٩b�=����"OJ4 �H�=Z|��`�(h7X��U"O�$��1}S�ً"Y�-�t�Z'"O�P�F���A�^�}��"Or��r�T+#�H��c�^�A�81��"O.T��п
����5�O�ZvB���"O���%�P~�x�6�����d��"O~5y�bRI��!-�>h}�Rc"O֝�GL�Z��V��<��e�4"O��
��+�ԙW
ьXp�LӅ"O�B&f	��M��hX�R�pQF"O1#M]�Z�2����?UO,���"O25�����d���'ƒ_�!"O����O)H,���D�����"Oj�Bt�K�,ް��4D�� �2TR"O�� ׂ+>PQ�g�&I��T��"OB�i$�"�<(��H���5"O�4��#�4q�v �&@�F8D�0!_y:��J�}��!���:D�$b�(���e �20��|;�-D�d��B?����c�؞s��Y�l+D�� $B�k��S��	V�4ka�*D�����	p$�p�套6Lи<Rѭ"D���S20)��z$#דrP� ��4D��A#�c6��X3a�0vMf��"2D�THs�F�Uk������:|�A�J1D���A�/\-�J��\�&a�(�"D�d�ujH-[�*y!�Ǿ.�.�bc�!D�P��@*D���$��y�^����"D��
PK�!��Uɖ.J����4D��0��ǀvC`]JVhT�o���ŭ=D�H���M�77��26��_��\�d!7D�(�ѩ���i�O�xX���5D��۴�P&SuԤ�v&��g/l:��3D��`�ܬ'ؐq`\�Axz3�2D��{TkQ�?Ѡ�:1�ى;Qhh��d.D��04D����h�6�b�Rh@W 0D�%a�_~����U�i�n�Z��;D���	F/%*e��<��({:D�k�&�C��
e�Њ3ޝ�K6D�ĉ�O��JP晹��ybp+5D�:��;8�3��1}��Bu�0D�� x%�@	�G�����&㾅�!"O4BÉ�.^@Ā��ٻn���Y�"O,�k�O�i�P�cr��Z�~u�a"O�<�F�.N�$�٥i��T��X"""O`�"�ʾh��XC�ь4p�i��'�.M�����1 Y��Næ<k.�j�'hj�[*��~�1p��<5l��!�'�(d��#ʖ��������{ˊA�'iP���0JhÇM�q�4E��'�-���H���v�<R-V9��'>2�Ô�OJ�'dB�t�j��'��4!&/�Pj2�
W���nP���
�'��   �$d���J�����	�'*J���,�44�~)����/��
�'�b��Z�ԋYg4�������yR�ۣcbR�5⇗Jyt|�af���yr�@l����d�R"H�"�P��+�yR.�0qq��l�?g^ys����y`\�j��TCPhaC4�9�΃�^!�D�6�r�)]e �B2I����YP�T���8D��{g����fQ��jYzm�p��'���啒h���a
��{�,#�n�X�Ԏb4x��Gz�r1�O]8ؓ�@�w�.\�ȓe��4�V
YX�&tsЎ�0���%���B	�}dD{�nZ�	\,|��[��]:�/ u��+$4l5�T�ȓ��h[D�B*!��$s��:�(��}K�L#�g ��X*e�V=#r	�ȓuj�\���L�*����!z~<��ȓJ��E�$Y�<�'��=`Y��K���*F�*���a*�=�����+s��!����R]N�� ��B�u�<��D�+g�L#FfN!VD޴���n�<�� �A�\A���K�"�rF*Ij�<�̜�s���B"��'+c(�b�M�D���j�N����9�,�e�ľ���=�A�b	�C�F�a��K�;传�ȓD�@ProN�@���"��ďa��5��j����uƍ�	%<�6���m�<�E�b֝�@�	^u�t`V']N�'Eax%Vk�F\��Ɂ�~%�aǖ�y��Ae����E�
�NH���'�y�N72|�Ħ��|0�E��@��yBI��n�����K7w>�ܰc
]��y��-�&-K�M��r�������y��^�{�6ɑ�����A#)C�yҨԺ=' �I ���t�l���E��y�[xni���ڌf&������y�Y�,RTR��R
N�2�dm1��'�ўb>�QpH��"PB���o��t�+'D���b=XD}�d�ˈ�� ��b9D� �&K�w:��0�ˈ��0H��7D�\��NB�H)�K<X��s:D������(���b���i�8��V
7D����,i.^!9��U�
���Y��/D��5%�<��X�7��	f���#�+D� ��BC,l6N}�e��=�^DӶ!)D��0a/�TR�+C�Ð6l  -&D��k�G$Rx�1�Xd�m�C�6D�ta� �-�DE@sn�(�!�bI5D�4�� ��\��"}�ڭ`%�?D��)E�@���cK�>͚�a��<D��a�;W�X�'�ʶ	�½ %0D�� �<�j@]�������'A�"On-�U��Pʂ\k�U���lje"O��$�Y!r%� WDb��s�"O>�zQ��Q��0�m 	YTL��"OlaT.
�2r�Ys�m�4jB��"O�Q�Oۗa�R�8���`0��"O���w��?�dዅ5?q�0:�"OX�����U*9�V���-��:�"O�����M�B$�`J0 M�q6"O���ĢM�;҈���D�Y?]�g"Ox��%V�;`�(�#R�$7t��"O�����R� 0C�A��+�lC�"OHA`��
hB-���4Z�8"%"O��ȀE��)�T�X��
1�>tУ"OZ9qD�<(�� 2�դu�z}�"Ojx8Q��)R������ތa� 9�R"O����	�8iK�a��aܔ3���`2"OrH��	1�.�C�ԟ	�f�Y�"O�Ȁ�l½4`X��4�� K3"O*T���ϗ����"]�l���:"O8`1�ъbݖȘ����k��(�"O�ԙ�� 7��r>aw�1ct"O^8�� UAr�+���3E��z�"O:U��'	�C��e�3)� B��"Om�����P��@yF�ߥ],���"O4���Fa��d�p��9_$P��Q"O��Ha�N$d�bgȟ�#��,�#"O:P����#�>T�D��1�2"O��1U�-5XD�D#�<�Dy;'"O����e˻8�� fb��%��"OB�P�&lF����pۨ�s6"Or(c&��]3�]�`T�=��;d"Ot]j�
F)�FV��_�
� �"O����nX�c
���M]�s�D� �"Oک�@A�-Gِ�"gM<��!�0"Ob,ˀ����j�k��a��y��"O���e�+{VL�ڤ�:p�(��"Op"����A/�P	*A�R��"O�S�T��LIF3h�$ r"O0�@��ظ�n����0�"O�����5X�ʡ� P��Q�V"O)�� p�~�y�N��Ű�"Op-�VBG�2��T��MU?$��s�"O��b��0zJř�+�-2����"Od|1��B�q�R���,^�?"�H "O�Yi,Ml�qG��V�5(�"O̽���k��ܪ�O�1w�^!�"OBT;U��Qw���=?bU�R"O4�r���:t�'-2%����"OĹd�B��ԲÊ�:�5�"O����ᕌ\'nջ4��F�v�t"O�5�%E2Q������M�`��"O�y�D�Ex6��H�8[���"ON�b	ƥ�< FL�L"���"Oz�3�m*ޖ!cK�-& �$"O��G�P7jr� #*��h"��"O>i�c]1�b�s7ˆ2 `�)2"O4�a%,ԌWk$ar�3��q��"Ofha��I�}�H%��h	�(���"O��J�T�B6�hʰ(W zpfQkr"O$9��B'S���'��AdNi��"OjE���'*~�3���7B��3v"O΀2��K?Yx��T�	L�~�ɔ"O��XFf��i�����I���@G"O� ���JK8�nt�$�ۧ(��}�"O�q�"��Nj(�0%�@�,�A`"O<�`#gM�V�D�?���"O,R���/"��XZ��%|�E�"O��Fe_�,Ò�	�%q�ޡ�"O�؀�������D�풢"O��1Eˁc��I��.E=j��%j�"O8 �1���sz�`�)�r���"O��p���9o��1!�L	�x���"OR��A*�[l2T�m�
>�����"O ���,i|�Q�f�>��|#T"O��ѱ(B�Q���d�G8*|`P�"O�|A��̯Yf>��J�,$���"OJ��2�Q�0J6�]=M�ك�'���y�f$02�YY"�ݲ{��В�'a��Z2��F����pDO] ��`�'�D]�p�A�a�)+#��P�ތr�'m�Ha�$�,h6dL@ΥO��'<�8��1�pI�A@�-�P�	�'*Q TD�$l��-ѡg�)]�lP�'B�7��	Ty����L2�d�ȓp��z6j�?j��HP��1Z��|�ȓb{�[7C�o.����EpN<%����lCI"$Bpi{'o>���ȓNF�5�G�\�`K���L�$�����8�QnA�E����� Er`�ȓ~Z�����Tvw�)���͗��9�ȓc1����ۮN0&#�j���ȓnra���q��$�٢}+���ȓ;�̑���,���[��@!U֐ͅ�,~�P��ڶ-����!#!��ȓco��6	I<a��q@,B�z@ͅȓpTQт�܈u6��`k"���SRhQ�t�2&�� ��v��8�ȓV�^@�$��d${e���P�ȓD�N���+OC��z��� S�x�ȓ��X�G�/jhZlzQ+>t�,I�ȓԐ8��E;�b��e��E�F��ȓ,IzZ`މQ�>�)��q�h���k�1��
	�+S^�g���ȓEˮh9��ѱJK� ��ȗ�Ff@�� �"m*WBҰ� dk�j�U��q��AH���U�_�<�����? 0d-��%/hm��!�>-�0��M�%��͇ȓ�[t%J��f��h%b�����	��բOlP�` ��.�j,�ȓB��HZ4n�L�2e��3�ְ�ȓ#�����l�~8 �+7�	������
t�i`�ϒ�椩��؜\zVi��'�Z�J���0LD�N�$I��Ѫ	�'
������A���-Nة	�'p|�2���<Q��äd�*�]��';Ј�vJ�bPV���J��\���'����H?��{�M}��� �'HNI"u�J+*I�H��֠E+
)��'��5A�n؁d���!ÔB��#	�'|e饃V./�Jq͎�h�H�	�'�	JE-5A2̈*q�<a��'^�U�O�4�j�A(�w�@��'#�#��-���� 	۲Xw8TK�'g�� ���p�΍h�׽ad�k�'��3Qؾkp���BOޣZ�Db�'�6 W��4�v!(�"T���)�'�:`+��S~@��xu䊆K|qZ��� , ��F 6�x�iƙ\���"O(�b5+�W��!ɓ|���F"O�x��AnPQ$��h>��"O��R!��5D�AfV;f��)"O��d��`=d�z���*��U�"Ox���G��<"�߅tmx쓃"O��r�8pƐ��j0k^>mk�"O�Ű��EV�)��Zqĥ��"Ov ��,_�n	� 2���8{�)q�"O@;��Z6N2�"g�1Xr�QB"O��r�	);슽�!�W�= �"ODyQ�R�咦EH���qJ2"Ovl�cE�0��\3V�1��,{R"O�Ū�)�0�Q#�b�6@���{�"Oԅ `��$�<=[aa�&U�%�&"O���,ZCa�-ғ� #�"�@�"O$�� ,i��=Av�8�H��F"O�ABl�z� ;�J6i�t��"O�Q���	"�\��Rȟ.p�,���"O�Y��IZ�	1�!݌;�faz��,D��ze��O�hj��TX%#�-D�|ɃaO�!S\��&��5I!p	�R=D�$x�I�z��A� &3�~ȷi<D�x9��c
�LJF�O�e6F�E�9D�<�D'DbUڧ	������#D����FA�RL�,�s�ˌZw*��<D�X����^3@���O6(�#�<D�<a�i͕"��H��M�a-���b9D�d`s`σ6ܚ)BRĞ�x��
�!+D� hS�D�P:�8��b�$D� H@�� ���	0�8;S�#D�lq���%-�j��ҪKj�|��J"D� {O�Rz0���O�g���abc*D�����U��l��La�X�#��=D��k�$���Z��Sf�7�J�� �9D��3ՄL�
��0UF	 !�p=�@�#D���!�^&7y4ЅE�^��Æ6D����ʃJ�޵�!IE#e��e"D�����[�ZRB�1u�5t�f��i D����;5NR�C�"v��v�?D�$��X�p� D���Q�,���S�=D�p*e�I${J��O�j���9��.D�\C"(K�:�بbR�R�^=� '1D�@��mW�cr�u!�	-u�2����/D��� /�zw����ݳ	�P��v).D�`��H*~x�M3�%��S�� w9D�p�A�Ġ	���Bϙk�2D��	6D��$��-V�v�#�.��e4�Ci&D�� ���#��m��i	�:l(HFj(D���E\���F4�^��׬&D�X8UeO�^�.`c���tJ*D����6?4ʼ"��2Y�p��#6D�D��ǝ�	kvxy����0�,L��)4D�t`1˖�[��t�@ ^#~>Ј��,D���A�ֽ�ŢRd�o��!�*D�BBΩO�|`(��P.���o+D����.T�#��]�G.F�f��w�(D��᱈����]q�e�U�\q�+D��rV��z�P�"읛�:x� �+D�("ІDQ*���K��p.���'D�$���ɰ@e��4&�5j�i�d D����c�q=�m�W��S��%C�-:D�0��κr?����*о�*��3D����y�"����k���Um.D�� ���օ��P��%)��!or�b"O�8`��އ\+4���ϐhWXIs�"O�ccfx����^f;�8� "OR�9"̘3Gb�5=^!KA"O�� '$�oi�y6b_�{9�]��"O<�a��^�-}��'ţ!@�DPC"OQ�6�@<in^)c���21�q�"O�l+�f�6I�
���d��1�6}c�"O|���d��Bm�x����7(!�D(�89�@��M���)歀%XA!�d�i"��1NI	L������p�!�d���f�&�ѽ|����,	�!�DW+6%�T�I�I@�l��q�!�D��L�b�.)9~�A!����!�$���Z�\�P!�� �%Ļu�!�H�Z́�U4��K���v !�D�~嶬�-i�|�ߵ!���R/����|� b�� �!�D(ĉp��Z�=Ӗ��G�˶^�!�D#����cѨW �Z#h��m!��!!;��"�G��V��wh�!R!�݇_@ �2�ǋ�*��`!(٩OM!��)N�H���G�Q6�O�5!�ч��\)q�)W0�c�%��%<!�\�=��� /u<�\z5�4$!���}��b�& �M<�<���=!�P	u�h��� D�4��] b�.A0!��
eK�@�R�^�*�>|�#ɋ_.!��$	�Xb����AmH=8b�ĥ6!�$�-�,P�Z�kv&�z�+)!�dǑ8gx��&��-E�ca��<#t!��N�M��CF�x��aa���:Z!���np�� �
�F���6!�dS#~��i��<=B�٪��5u !�$�2��85዗�|	ra��	�!���v��͈'������T	Э5�!�d�;
��u�5igVMS1	�'�!���`F$��k�p�����h@�s�!�E�¬���(+������{�!��@ej-q�$�7<��$�����s�!��S`Cn��+�ƌ2�e��%�!���1#�L��D�R�����c�!�d�+5���d��c��84�{�!򤝡�� bd�<i�Un
!{(!��!Rfp@��O�~�R��S�U}!�,p�3b�<� ��O��ld!���}q��@k^�n6V4��"7J!��t�a;)��=M:_�Ԉ�"O�-�wC��m������C4�u#c"Oܸ�*ǥ��sr��3�L�"O�{�/Ъ+��0�/��G��2"O��sRGʊ=�b|Su@	j�؁I�"O�)3�ՂK5���A��<n��`)5"ON	��٧y ��PE'X�^i"O6=�Eb^�s$�0E�E�R�|��"O�M���v�����Ҡ˲H��"O����3V �(�aǂOĮuYC"O�� p���LI;!K\��y�"O渫&�RN�d�A"�V�~@ �6"O����F�s�.�&��z�
l��"Om����h��I!��(�V"Of����.a�&yb��C�Vo�9�3"OtE��A"��A+��U�TDX�"Ov�Y�d�6_�P�;q�$2�La�"O� ����c��V��yV#��g�5�q"O(�A�%��c®E� �[�`���)W"O��2�A3q�l�� �}�ँP"O�\0�DQ8N�`ț��=S�"��*Od�!�)�2)�\SWE�*_��0��'����Ҏ	���( �f"Y1���'�H�rLT��a�P�O+T�
�'�����W>W�Xh�Q�Atw���
�'���Bf�/9� ��W�<�0*�'Bf��RB(h�<E��@��3�����'p�!"e�4a#��2*�:i��'��U�E���\�b%O�/���`�'�Z ���&�
�%�;p�U�'�,���<*皬�Tf�fJаc	�'Z$����]�\��%��_�̍��'�6hB���&�9�M�)W-P5��'n�ಷO��Y,� ������ �'/ʑ���.U6�P�Μ�I����'��@��D�3>�09 M�0�49��'E�����J��9z��O'2\jЈ�'�f!+�"��er��ׯ&0FY��'Ҩ���2�,���G�3�Jy0�'�%��/�"�u�w" 0��]z�'w���Rөz��'�	�>6���'i>}�H�a+��#*�d3�'�:�!�%W�bV ��(~�V���'�*�!j�N��q�I�d`��'h�)�+^-8��4�SlA�`����'aQ�e��k�JE�Ҫ�;^�ER�'��`�#��,*t�q��#]����
�'�Q#�e�D��]�1��K�x��'�M��oW��<&^�m����	�'����&d�3�`���(Ƚl�xu�'�`D��@P2{0�j�g�Qz��X�'�����B�<�(I�	�;LA����'2�Qy�	>Aha�� 9q���'�����b���r�ǌ/�]A�'�z�qЈ7y��ag��)"��'d���\�.+����_�z\~��
�'?vl�����i:H(�*4w���	�'6`���e�Y"*���j �f��Y�'z�<Z�+K�W!*�;��ǐ�
] �'vfH`f B�������~~�x��'bp�@��(n�
!�(rCNu�
�'�"��S�T	B���0�7oI~t��'jf�y"L1w_���@ I�tt*���'��u�g�  ���� e;�0�'4N��W���3��قe����'���Ƣ�Z$��y���` ��'�$a�&��e��@a�ڈv���'����D6���x�^�r���'�頒��(�T4+��![#pr�'ۮ���R��`����[�r(��'*�P��W[���K$��#N�D�Q�'��X!�*#-�,�Ui�A�r��'�yKV,K�-�`���@4���
�'�l�2q��ƅPuE�_�~Ѳ�'��8h��F8��;��dA(dh�'����2��S��Ǝ��V��ܢ�'e�%�� V M|��ʑ��J��qJ�'C�P��#Pk�M`A#Ըn�E��'v	kb�իq��X!�Ԉk�[�'Ja^q��Li�A+^�����`1D�8�vG]K�b�y��8�tM��:D�� ��XfG�4mtL�$� �9�"O�pZ�����)���߈a���0�"Oy��
�N��L���\�iJ�"Ot�� �s�����5oF�aӢ"O��Z��H2d�`�����>0`D�"O�a�]���d�P�R��@8r�D��!�$Q�+�ą�CC"��"�� =~!�9��a�G�S�b�-�®�+Lh!�$�
.`
��#	0�`=�E#��M�!�D� ��`Ȓ	+#�Uʅ!ێb�!�D�)\���K����Z�D��v���T�!�d�/����פP'�2� �Aw!�VV�$AQ�r�ĄZb,ԔQj!�!<��Ys Z@M��	��]<=Q!�d)������M�o4��	�o.8!�dT�c��)Zg!y*z��Zr5!��֛"���!C�
|��RN��]*!�D@q�<R�h��TY��$.�;2�)�'0V* 5�%c�_�i��5��'�" r �_�:�:� 1L���'z�]��K�*�2��'G#Af�\r�'�Ό[ue�O��傷nX�@��(�'� �8��Y) �L�a�#��5N(��
�'�u��E�Z1��!�-�3ҾD"
�'���eUjcTT�
Z(0�P=�	�'>]�c�.l��0�eh@<.�bA�'~.,���X�Qƚ��DAC"0 ��'5�Q.�zրA�G���A�'�N�+U��3�@�	�*�0o���'��W��\�F(�n\�S؅��'?�hC�3�Hآ�K�4�{�'�F|:%��=3:E�'Sz�hI�'s4Q� F�" �!,�.V�!!�'}���5Ō0tta@c�,$�
�'�Z`H$Ŗ�{�:5Yf��0Y��p�'���B�׼b������7� �'~\q�$)���Z�+P5���'���cO�/7M}Z���C�1;�'q�H��oW�y>�YAL�?�x1�	�'�ΔK���F��a #��
�ha�	�'h��IB(�JzL�Jp�#(
Ic	�'*��1ϊ�2����`���45	�'2�����	�B�2�/�i����'0����.9���
c�d-�C�I�F�
��e�X(�lB�R�$fLB�	";a`���'�A�yp1J�q B�	�!��)��L�V�ܠ��j�>�ZC�Ʌp5���$D�:���E��Z<.C�	�>��P!���
d�c���[%C��o�:�#�->�2$���5�B�I�l����ƕ�tE�\����}�C�	�A�0��UOɺ+���B$	Z+I�nB��4K�fy���݉��Pd��B�B�ɳen=����;'t|pX#�@�S��B�	�(�, �̍*kb� p&]D�C䉆J��ZS�����b�h`�C��wl��.@�
a � �	�x�zC�	�{]�0�e�<b]�����&fC�I�Z��G�ͱ��9�vnY�BHC�I'�r��f/[�C{2�b3�U�2�FC��9�Z��4���o�>-ʖ�֝V>,C�I,qi�\y�V('��	c��e��B�ɤN����C_�)�a��j�6i�xB�ɳb�����)T���KAG�=
âC�)� ��i�܈I�����jE����J�"O�+���J_��14�� a�0\�"O��Z���Qp�ƃ���R`"Oda�Ó>L�f@��\(@*q"O����i-W���HT�A�	4yR"OV�x��mE�}�Ŋҝ"d���6"O�LAvM҂0)����4Z�]��"O�Q�8O����ƓHNN�pq"O�ta��\�!eҽ�p��uE�ѣ""O�p�j��nuL�CPdG~,6���"O�1CwG�+Uւa�@��!�� g"O�m��B������QH�$�x�"O.���hZ��,�Ct��.�`�"O$Ձw���Y��T3��@
i ��s�"Ot��g�K*.B)�����L b(s�"O2E�piK#/8af���1��6"O�a�A�7|u�]#���'*����"O�L�7�
�n���C1H��]|�Q�"On�z�CݤXw����eP+<`z���"O���)N�V�H��M��VQL�I�"OE)�Ƅ��0 CӅ���["OZ5�OYp�`��$�%���Qf"O�)2rƍ8x�A�5FY�y�����"O�1K�ɋ��Tmբ�	w�X:e"Od�[5�żAv̔:D�G�k���A�"O�t{!��.�Хx�o�=�Й04"O<<��Hx�"#�Ξ8���{�"O�_����cO�yO��V]�
!�� ���2r���?D�@�a��2	!�D�	[�P�j��7!ђ"��(�!��E/k�f5"��;5�DkG�Ɖ]M!���9B��eo:p,T�@a�˰eJ!��G����W��d� �S,`�!���J�� ��&Z���`*�4w.!�D��)��y+C�U�RcI0!�ظ���"_�i���)_\�!�dľV@tTѕ�^Ȯ`��A�@�!��P����O��[1�R1�!�π)J0Ʉ�)5�P�Ua_-y�!���S�B��nͨ`��t�v�!��U�E�$���n���,�����ej!�J'��ɇ�6�vHc��4GQ!�D�0��`����4w�<}�F!eG!�D�fHN���%��C�b���<m!�$�SX �b��<�L�Z@.��!�d;*�d�2v(֝i�f��Ύ�!���s#
�"ଏ��&�ajژOi!��4qܨԫ��9�8�zT֓J�!�$;D.�� Q��1Rd�H�χP!�$S"UCRɇ�[�d
(� *54!�dG�2t����K���m��!�$S3Cp�C�E��DP��H�F߁i!�ęn2�!D>`Ar���'d|!�d�-fv	Ç�43�� ����!����E���Àƛ>��4@t �4MU!�DĈg-���[~�ҹ(�n |�!�DӪ{G8��e��J�R��-���!�אoΘm���E�*�2��!A�$�!���:\T@ai���k`L>�!�܍U�r}qeٚ^� �*�D#�!�d�[S,�R�����Z��w"O�XH��M'9�⩊B�K>4��qw"On�w�,Y��yedW�*��"OY�ѯJ(sA�I�B��s�x��G"O� v�#���k�t$�BA�6⨬sF"Oؽ�ᐗUM:PB��/Q�Fİ�"O�q��[�+\�ɵ�ޱ2�\�q5"OF(q�/�8�tt���+	jt�+�"O ]g�@�"��:�gO��Q��"O��Ʉ�O�n`
#a[;K����"O��Ad��,I�D��'߾�"AR#"O�%�T�[1@�rh�'�3Ĥ�ip"O�d)��S���EH�F��ZY�� �"O���'!ϼ.ʾI��Y`@�Aa�"O�a6���w,���DZ!��	A"O�a�S?u�fM:��.9D�`�"O�<h��� 5b.Qa�!B�8�#�"O�
��^�j� ��jݾ_
ɫ�"Oa"�I�
?��PɌ��X���"O̐׍�+b�\�ڐ�c��5lL�y�aۘk����jp�^�Pb�+�yB�J�Js8�Y�BtT�<Zq&���y���R��`���xZ�8�,Z��y�`�� �!� �ܜ�W����y�,?>&����۵#����Feي�y�<��Jݳ"�X`�Ci��yl×BT�	B	��X���[*�yB뚽Ji(3�ߍJ˞�c�I��yB�R�-J���Ց<���l̿�y���M�~��u�[�G>�T`�U��y�jW�ߦ����uO�%��ړ�yG��y,|Q����v�L���O1�y��+4��06%J%kCUyiP��y��ˆ����@-o^���G����yR˄)b��q�"G�-~Wz!�V�K>�y�!�Dx���x0
Y�&V$�y�!��-��g�'�2���R!�y2́�D��Ѓѣ���~q�5�ӧ�y���x�����$ԣ؎M���I��y�#ЎLˈ��Q'�4n����	�'�b��D,Ҥ{H^	��ќ�����'�n��A�O����£��?��D�'��}�A�"��"��:m����'e�� �G��X���gg�P�
�'���c����r&`�c��O<c�����'�t��
�T(h�_<T�@���'�^ SD���W��I4,L8!<4��' ^��b�_F$r�!"����'~5�P��������_m�� �'����DO�>�F}c�i�D��'FX�P�MA&j���"*��j&x�'��Ԑpb��#�"aS�o��Z�'tlA�+�5&W�CRG$l|�{
�'ZHX���T�J���j�?/%*�i�'�����E#=��#_3,G���'!�Њ��T#� �:��%R*HS�'���aU��'���C��P�X���'��"�)���@��w
L���_n�<��L:`��9VZ����O�<�1c�9	�U��-�4/�����K�<��S��4�"QM/ ��S4�m�<I�D̶FY|��-ʬ8o�����S�<�%��5t
Y9�-�����W�N�<I".�0Ggr�H����')D���L�<!2�Q�l�L�!0$�Y���a�<	 Mr0� �d��W�Tb�&�Q�<	$�\[])A�T\.Bd÷KO�<�7���B�I8�c� }�Fi21j�p�<� ����_�Vؾ�0�I 1�^%�"Oj�ۣmўKΥ��SI'إ�"O��u"ڞ�ur%	)��5W"ORXSU�Ŀf9�= d��c���@�"O��h��Q8X(�K�DE�$=�E{v"O�qL�&dĊ�d��# �"O�}����md���h����2T"O��`m�6��Y�cM�8r���""O��:���deFEpp�߳;�`��"O�P�a�e��
��\��m�f"O2�%�	���C�ɂ?\��)5"O�([B�C�g���*сL$��)j�"O�ȩ�O�$2FnG��V���g"O�� V�I�&Q�-#1���%,��BF"Or�2w�$T^���K�]n"`��"OF]+���ea�k�<9P�� "O��c����y9�#J�e*E�s"O �ӠYq9��B�v*���"O�ٓÃD�s�(�*J�� �p"Oȕ� �W�d���+u�`"Obd�'�u6��R!�U�9[`iy!"Ox	���&~ XA�ET�R �"OU��E�:
dچ��s?��"O���(�A����#Ϛ6
@�rV"O��x0�:w�V��qァR8�I+�"O$�HЎ� H����C1h"��q@"O�=�ukD�*[��n�+O{0�)�"O��Id&����m��}v$8�"Oq�w��x�V�赫Baf(�v"O��C��+N��i�$뇯Ho��u"O�,���ޙf�|�#�Ob�e��"O��3�ʻ^hИq�'!$P�*�"O\9Qի!�V,�p��3Dv���"O!�v�ݖs��M�[�9$՞o�!�Z)yBp�k�T�|�r�S"� <M!�䏨x����M
�G��T+R�S(S�!��^�*4h��㌕Q�T<�!�@�!�$�.J>�����i�������K�!򤖠b�6U!��֮\���XŎ::�!��45�>���FA/ :�5�$�P,)�!��Q�=� �;�A�:*4�$�̽H!�ā3�6����?t2-�de��!L!�$	�;��vk��{k��+�G�h!�O�?�`�)T���=��eB�4V!�����z��D;����D�T!�N\i�cS�7���
f9M!�dZ��0$ɀm�� �nT���WJ!��R�f�  ëۆQ����D�y�!�D��61�����3L	�!�D�j|�gaB�h�� ��M�w�!�S�>��a��`��'���!�� j���BȟX��t��dN�S�!�F�-V�!�@C9�x�R�&C�Xc!��˷5��|P�L�<�脒��Y]!��Æy�d��h�<X\ ��#%�@S!��Xٚ�<CO��: �L;k�!��P�s�0�3��G$�M0��3�!�ddH4���Ab� ���(`�!򤟎^ r]Y󎓆]#|=� @�"�!��^"�Xa��_�u��Bqd]3q!�O�/ݠmҦ'q H���>E!�dI�Z~&����@�r"�����	5!�DY�A��8W�FT&Mi���+!�ċ�\�\�`0��<VL0c2mT�9�!�� 2�C�W��҇�F�E�|)�"O��᭜4w.<[Vb�!�H��"OLu��'��F�� .���AW"O`���W�<������ƅaq"O�h5 �> �Nz�'�6,��`�"OVQc�ʾlMƩ
��+t���J�"Ov�3��':Ÿ1��6{�. @"O���3-�1�E�!]|�X�"OV4ۤk�6謑'��ET"OD9ЦE�A���R���� 8�U"Or*&�$�����z����"OD��"��h!Y���}�2=��"O@�Q)I�)�~��G��N�1"OĽC�K�*+�f��GR</�Rxj�"O�h�� �E��\)�eM.3u�)��"O�р�Tk�13a�\VڨC"O�k�e"dd�Q���"O�����"M��pfɄ'O0c3"O��w)L�0�H��S��`/��ct"Op��lA�QKҭX0,Sd�U"O��(�H�� 窌B��e`$"O�kc��b=914��?���a!"O�$	gdX�,"����]J�"O$ Ŷ�������B-=k"�WY�<9��^4~�D Ǖ�Y&*�P,�l�<��4����,2���b�Wj�<i��Y�y���xt�9�,*3K�`�<�3�La�����ĎB����![�<IE�#"�zЉ�]G�u�b��O�<��mK�Q��%�����\a�<�(�\iz�l��<�N�B�d�A�<Q�!uY\h#独_[|��m�}�<)����� �G&;�̻��}�<��o�iG�öhX#a걣D�z�<t�S��.գ�p:�h�$�[�<���
�-�����H ��\O�<I��9l���f��	?S@1�)N�<�(K>�m	�N@+H{�4��F�R�<�5���l�օE�����;�]L�<�@	�)$��#QK� {�F��3��l�<���Ϋ#܉�TB�Nw\H��Kh�<���Z���b� �tex�,�zB�	,\~�m �(�~
��yG�P.��C�	Y�֜9��L/���QңȑAbC�I,qy�`X@�S6U�Mj��Ć{��B��4�%��%\�`�B4�+A�;[�C�I�i;�	��`�?�J��00�C�	a���bnG��F4p�W,~�XC䉧:�i��M�	^�VqB��U?`�C�	%�L0Fm͂NM9!(v�XC�I�� �:�n��+<The����B��{��� ��H��q
����"�.C�	�P̤�K���@L���a��N�C䉚Xżm���_ǞYB/X�T��C��0}☛�oK�5��%�	�~�>C�	�&*�9t']��׬����B�I!l=2��oC� Q��#��@�j��C�I�'טHx�i��|I��m�z� B��:+�Teiԟ{����*q�C����i�a�2m��\ې.JY�"C�	-W>\u����ZFb�a�d_�C�I�N�F�H�LS|[z�j&I�p�C�I�2v�T����5�@� �C䉫rV1�c̄��F��mё<�B�)� ��B��~��	���wU2q "O0�A)�;>&�hR�5QD͐c"O�a���L�/���g^�^���;�"O4�Y5NU1	EFqHq�;k%�ܓ�"O�}ʟ<c��8aO�:��<�"O��#cK�5����$Z
S���"O i�����)d��><��f"O�p �E�P���;��!$0yi�"O�ǮBL�se/7�MJ2"OP��KՐZ8��S�ː)7.�y��"O�X �>ЬX�>t+�K	�'L2��]�s���+��ǋ
^
�
�'+�Pfj�/!�����{hB���'��eA�+� ��96̟8{{X0��'��p�EcA0N�!K��A=t��a�'7l���3���jLpK��{�'�	��lʭ/p�D�ӇGac�L)�'�Ҝ�1�ǚL;�F��6D����	�'ip嫅-����u��=����';z�R����N�m���W!4j��'����Ɓ�.0.�QK�6@�R]h�'T�xa��v�6��c��?j/NE�	�'�@@a!�nX5[T���i�t���'f�8A��oMX��2�]=t����'`0�1Γ�)/V��q(.D\��'�hT�ӫ $6�����
��y�'��<{��H�P�"ɢ5O���S�'tFy�5$ �:ݔ�����i�R�'fT����եI�.t��U�����'��=P���.Pa~��2�Ɍ����'w�1jDi�8o���rI�.iC�'܊��$!L�m�R,��J��y����'��@`��M�u��i��>}Rj!��'_�0r�H,0��K�E�-=�HP�'�ؙpޜ4'����.�4*�mI	�'b�	'A�67��1"�%+�����'��9��&V!���ST�$$�`H��'��HK�J���5+�+�Lr�AX�'��)2s�L4���v�E�XhX�'f2�[d�jh(}8�NQ�7���'"��Q�Kg�LxF�@�DuZ��']���5�ݏ[D��#&+�:>\K�'��]Q��U�D8H�FA�v`\P�'�ēW,J??1�H���;�p�*�'����0�L:wt|{�I�D\���'*R�ǥ#S>���Ȟ�*��'��v.�>;��(� :��)b�'��x���	�f�XM��@�5
�����'��<c�Ǫ~�fH��0?F�h�'�l�Kӭ�":a�*�vX&�3	�'x��S�K�m�Ҥ�U�Kv�T��'�|��ȭK`��9�i��torP��'7� "� 
q;ĭ˄`nN܃�'8�ty5Vb'��0T�M:m�zXk
�''��P�E�0jn@Q3��O���
�'^�d�M�7s"M3���W��t��'qƼ`�aZD �2Ћ�5(�<�'�,��r�N�5��4�h	r��'aXp��v����-Ȁb/���'��X�mQ�ggT]�6@[����:�'���K�~%ջol4�#Z�Y!�D�,��R�W22��1%ϟxM!�dF�DTfJB%�% h$RwO�,c!�Ă�d�xCN�D�64A�X cl!�� ��E�#l@�����?-J�Ab"O����	>`�(9�%�(Dd�p"O^
�[��C`��&)i4"O|!���U�cD�ݚ5f׭!	���"O�L�5�Y�6�D����6S�Jl��"O"L��+H�2x�d�%�$5�6Y��"O��x�j�]O����*F��P��"O����\�~��,J1���*"ON����(��K	�n�� �P"O�j��'T9�8����t賀"O���)ָ�qu�R�g}�8��"O�a��&���ˍ|s�<�$"O>�B MOU(����RhC� D�丧o�7T����v�?q��A=D��y�bQ�9�\��R�U�;�c�9D��{P��9mL�0G��R�	�=D�h��!5�D�p,	2?��=
��9D����`XEyD�;��˚-tU�DD6D�x���"rets��!eҤ�)D�D�e�2�~�+�aLZ��(9�
5D��́{�����G � A��5D�0�2��
!ETap�L�5|��#Ʀ4D��1&����C�#ۡo�F1B�4D�ı�+��\q�d�a�B
4D�$QvH��&`У¯2|C�@d�3D���o�4s�Rw֓�l��A3D�X���qf�T�T�S�άI�2D�L#S���5�
Av� ���i �1D��PK�4M4�+�+ :1��-D��jU���  ���B0]C0�,D��K�i�05�<��3f�@H&	"��5D�<�t�Fu��5K��P�2)�5�3D�
@��3+�ӣ�Օ��ɖ�2D�<jdJ�;(��(S#O'n���w 0D�D�4�S�B^P��C �L��!�:D�L�T�S,	T�pQ�Y�z�:D�@�U�W����2"#C3^�mh$�5D��x�쐹<�"t�'DNDa��u3D�d;g�f�� �̪=����(<D����a'6��3��&]������:D�����˭$˨�3�&ɜ:���7�8D�x%�Րv,b�S�a�8�A�+D��8Ug+)_Ĝ���\�cl(�$*D�����t��Шд9��-�u,*D�t�2�E�L1ӧ�`��Jץ(D�$� o���r<����S���!�(D�`�l@N6Ѳ� �l!��f(D�T�D,Y�OlJ��lާ
�ڱ" &&D��ȡ`�.��`��s� ]��a#D�����"�X���Z?&��S��+D�)�H�kF����!��	��(D����@�hdD�J�Lb��G&D�@[`��r����A6��M�2�.D�DsQM�5�IQ �bt " �+D�`�dK	5g�b|��c��,"�7D�h)q�I9p+�=:AK��C�����*D��2�$�2w�`:unG��(P��&D���̇�NS���NY/E�\�3*D�Ⱥ�'A��${D�]�,��&D���N���9@��S�wt��r&,8D�|�5gӀ��I�V{z(�bB9D����ζ-3�D�d\�6�$�[#�8D�����>	|�07/��{K�{&�4D��F#M��q0C�K�D���&2D�� J�pŦ�po~U�qJ�>i�p��"O�98��2E�Ќ)Ej�
�t�3�"O��ѧ���Ԝ��@,�R`5�"O�b6/�[`�!��;G]�H�U"O���f �fk]��P�8E�e��"O��! �	n@�7dŊb(b���"Oh�ɢ�0r�lň��C����3"O
���jV�t�̑�o?o���"O�d!�C�n�����al@��"O��Qd�+9��!�`8��,#D�4���x)Ҥ�!]$c��}kt�<D��:5�X?y#�U @���/醵YD�8D�`�嫍9r��8�+D�}�z�Q�6D��Q��؄+H��M���1��4D�X�6	�,=}�{w�	`LVq���1D�L*��ق<<1�`�#}��F0D�$˱�G��5!`�9,M$�r%O2D�s4�L�t��p�E%P�����:D�4���3]`yYAH�){y�9SE�5D�0� ��0y��g\�@:��j`�8D��a
S��\;2�>i���R�$6D� q,�aJ��@��J���2D�(q��~Ѣy$�ޡ5D�"V#D��I��1)l!���8����i>D�T� �%S�l�0�Z&d��0��N'D����L܊
�}8Ƃ M�T�0C"D���̅+�*�RG�9"
�,�w�?D�8ۄ�Q6j�f�kC�"�H�bB2D�H2C�'B���O��p�Ɛ���=D��@����Un�[�GLż$s��<D�x	 �ٸ F���A�=�X��o%D��`K�7�I�C�ֽLDj�8�"D��ڑ�
2R�D�@��3:0B,"D����B�K;,�����'r����"D�h��-D�`*I�iS�hS���5 D�p���$s&�r�!?P��˂%?D�Pk�/Q�}��x�A��J<ꍻ&�>D�dр�j6T�c��]^ �k�H"D�`�qh�;C���J &f� -�ac D�P�dƝW䉳�Ϋ
n ���:D�Ȼ�o�'E	t�A�����!��>D� x��_�}y���bh�J,���¤=D�0�$	�/,��H�	�%v%���:D��ʴзO��K�@ S�ѕC7D��#$�N�I�b�ؒ���yh���t�!D��!��
̮}�g�����4c��>D��f�݌q>Ĭ��8����7D�0H�%M>0r
hx։ȃt?�e2D���a�#d?�!�i�,x�U�"D�@[�@�2^� e;�J�[��\�� .D�ثR%E\��@n
���" 0D��+pcٽG~��ˇ�
����.D�`�gJ�?�җ�5���F�!D��*&��f?�(�u)E;)�(u��2D�x(���f�z�Xe��2G5�Ȃ��3D�#�D�M��,����fx���c2D�t���Y	Ll:8�E�ߞ�~Ȑ2a0D�1Q�	E�J�2���5�!�R/:D�PӇ޻d�($0��:��(�P8D�|ٵ�O$�lѱJ ����Wd8D��*�*�+�<��G/I	iihr�N8D�����M2 ����a�8�D����+D��
�h��BO���2�^�OA
� �6D�XY��ފxhu�[�MТ g*O� �ũ�G���lK;rP
y��"O�8y��Ė9J�0�t�ߍlU�\�"O��	B��~���*�\�0�"O`�a@��Ƹqr�$Tlqh�Q"O,�0B��3HiR�\�Yo~	 �"OH�b�)-5�4U���+0���t"O�("@�V�8�����
�u��"Oh�2�K�<42��K¿.�b��G"O�Sҫ��]by2��,�tAG"O.L��c]�6���h�R?z=FUT"O�1����1���%�+. 48� "O���dL�3&�&�@��8Bᴁ�"OJA�f��'���ۖ!���8"O��AA�&>ld!�$�Q�]ƪ��"O�%iEC��&�9���>�hA"OR�;�fZ5Oj�R�
?���"Ob��P�W����%j>A�6��V"O.*	ɎJ>���T�"!R�"O�
$F!$U�� S��(,
F"OhD�g/[h�q	�n�nT��"O�b�@��O.��z�D�e9r���"O��3��V.d�iҦ"�R���"OZ�3�m��ڬS�	$�"$J�"O �QiͅA�.D��,��"�"Ofl�Сx(0u"��rQ!@"O�$2I��$�Ԭ2L��+g���"O���(��F���aK�z���"Oq�蕂r�4��gl0Q�2]ɗ"O�@�%��5�d�A��eƸP�B"OZ=9���:Q��J.b�pM01"O��q�+�N����M�r}�@R�"O``�^��>1�Bٞ*r䤁""OXi�V�פp�ܥSv\f,)�"O.   K�>\�k� B�'ª,"O u�� ��E#�E�ab�\La:�"O8�'l�22�	� ��%L޴#�"O��x�k�5:U�1s�N�;/��K�"O��i%c^�hY�#��K�`��"Oڕ�f%�	gє"C��(���"O��;��(^R�`P�`;�D�T"Oޱ��烰 �b��V�
�\��g"OnҢ�N9E�r���\�"�>p[""O��e	�+����4�>�"���"O���'�f#��ia��[Йʅ"O�q�0.ߌIR�-SHV�/��!v"O���E�Xrcf��6�j���"O�0�QgX�0�ջ�e�BlI*�"O�ԣ���>.T��DS-��i�"O�8Y��V,,�Hȃ╹x�t䱖"O�e��Ƅ���m����(�� "O�M��V�V�&���E�?6�:B"O�E�se�("��E���ōYtPh�"Or�(�C�#Μe�B�y��%i�"O
8�"EV06�؀{�g	1�r�z0"O6�ʗbɚwW�*S,�(�\Њ"O �p�!�0&�!�ؒµI�"Oe�	���l�t��"s�Z���"O�� �c]�؈F7M��H��"O�$����O���3�o��x���"O���L��jf�x"3UR�ye"OhHB"d@��2���qrl;�"O4�ƫ՞�j �����50�"O�$aq���T�t�,xR�h�"OE` �!i�j�1e"�1{�p�"O� Z8���W�/&�ҡ2+��$"O$���̧y;XX(�T�r ��"Ov �&Lh2��r1�ʢ4�|�R"O�9�s��Ss@��/�=��9��"O�`�&�!.t��"��R�Q��@Pc"O,��A��!�G4�r0Z0"O��ᆤ��}!80�%�C �Ի�"O�`���O�͐nF8Kt&���"O���dI��j��U�۫(hȑc�"O,Q���� p������$j\���"OP4��8z����e@@<1"O��[N#�����ޠ^��"O�0��Ν�x��[t�h��(IA"O�:��<"h���%$ʲ); "O��T��$�u��b��@8h�"OD�ac��_L|��4(�=f!B\��"O�"�'�k���R�ė��PU"O>�3��E]
05�۷b��- "O��x1�[5xT�,!�T
��Ĳr"O��6�G�T��'Б@�Ĭٳ"O�Ik��YE�t-� �ϒ��%Ҧ"O�� C%�j�0��&��/�q�'"Od<;�\$&��E�𡀌/�<���"O��֣F?8����Q��1��0�"Oz�CC�BVh�!5
ÍoT��2"O��)���qx����P��P�"O����i�y��e�UlK�Dɫ�'�Ā�j�w&�Qk0���i#>���'���+$�ȣT��H�ڪYX�A*�'� ��G�T�����X��ܓ�'v@� �h Mqj�q�޳%="�9
ߓ��'\�H��lʐ��ƐΨ��'ղ�z#O>:��er�(B)�
���'na��b�FJDۗ�W4^5��'�ȁQ��W���:�k��$�$�s	�'(�%#+Ūi.��i�ϒ
)�&����y�+	3�.�3MI�I2���c���0>ѲN֕q��T��.[�`Uu@_�<�'.~Z�0�7�-n��2�Xp�<q2m�9e����A,X�� J�i�<a⠇�Wp�
��P w��ABF�`�<���̪D8P�¤S�*�Q�JLR�<)�U".Ina@g(@<n�($� ϑQ�<�"�A�\�J�ju#��>XqX�O�<�@%�)uǨ9�5�®z8̓�-�N�<y�@AAi���m|"�k��A�<�� g�~lide�=��k���~�<�!�3b�La�C<m��e�@�y�<Qr�S%��`Q�C6G&���d�'�ax��R0�e;���v� %�F#ݬ�yBߟ7����Ќ
s�^�r�Q��y����5J2��w"S�r%���Ê�y�ǂ��hh�C�daʑz`�X��yR��L����lP+ �P��J���yBM�.��x���p�ȠY�`̘�y"�V�
��zV*Řg��x5@_��y�|b�)�V��#Pd��@-'�0m�� �]�<�f��ys�̱��G*:v��umZe�<��K�/p��Q# �"E��A�.�^�<��5q�<ā�KQy�(���W�<1ROT�%tBD�\���0�/HR�<9Bǆ%m�`��@��M��T�Bh�Q�<�J_���AǞ���t0�X�Ē>yc
(�S��NV;����$�M12Ѐ�aGD]aR�O� �8�F��9BR,2CA[�;h���"O0�[T����6�2��<~S�G��}}b͔\�dr����
�%�m#�i\�6�]�D	>D�,��$N�xA�$\�q����c1O`"="a�2%�h��׃Xa(�zV�b�<9�'�:a 0���s+�<b7�`�<Y%����A�ZZy�e.GE�<9w,�4=��A5��'�h�[�f�~�<�4C�~����Y,�֡�w�{�<I��>sD��gC�&Kb��E�`�<�Ɍ�E�G�! L8q%�RX�<�h�CV$����M�j�Xt�JI�<Q�N&Z�N�!���ߊrq�TB�<�Ն�,t:@9���!J��Qg�G�<I�l�@"�)�a̜;ԊM
� �D�<���q��e�� �'5�0�͕u�<)�)��+�Oƕ�<#$��k�<1&l�y�F`S�.�0"��bi�}�<��I��62�aQjƴn�j� ��L`�<��)}�L��U ����X�<�dL�*$;��A��&$�:Q��K�<i�<Q� ���!Z��܀c+MI�<Y1"MGOR�@%��P��@b-�E�<��I�9�0c�рUr��XH$�ȓOeL�h�ܬSxٳ��H�����0L���Ɋ�&d����x�X�ȓ�2p��J�H8�)�	Y���ȓ�(��AOE�(�B�Bv�Cϊ%�ȓ)�A�J�CD�Z��+,>1�ȓ$������{!�0:4#��I$80�ȓt��Rq��
<z!2w���<u��0�� ����n�%$�65�ȓn$�8�nϿ\i�}�&l�l�p)�ȓD:d��˶O@��F� ����ȓ9�`�Kq�ҧ*fF$��.N3G��ȓT�
�s0��,|.`[3ȕ2ց��`����Z�.'X�5�aW���ȓL!��ˇ���C|��B4�_56Px��E��@�#�!a��-�Tg�%Qj|�ȓ	���hY5v��q啝My�Ʉȓ8��E�d�6�z}itb�IV��ȓHJ�K�oч$�8L�B�T��A�ȓ}P���g�<�b��u� �!�r��ȓwl����+2�J�8n�.bԝ�ȓnq�m�2:\X�:�o� X�1���0q�w��DFR>az$��c��e&��3D'9ف�|e� �ȓ"�v�רhru����S���ȓ[|����GN�!�8 �M�
9������f�ɱ���ʒԩ�B1u�@�ȓ:�̐c�G� Cִ�a�Я����ȓ*�f=!��ޜF66카�p�깅ȓY��Qb��'"�����N�dYJ4�ȓ<,$1Qs����!�Մ�5 �z|�ȓb����	�){b�x�������ȓ�֥g!�$�I�Dɟ�=G���J�P���l��s�F��qkۺb���� �S@nײlR��cgc��o��ȓ7��;6�ɩ-����k�'d�D�ȓD2T��c������9<|������"&�?xP0hpNFX�ȓhvx̳gfЪM��H4�Y�����-�.!�d�wH��SU�
C�X��B��a��j�P���:P�UC@����S�? qy�Z�\���J�78�xK@"O��[r!S�s��0�Ԩ�,OF�)�"O���q�F& �XH[�2�5�"OU��!I��鈢�-K �0�1"O�u� .C1��EА"B��p��"O6!b�/f�>-R��ؤ�9�"O~�жK�����Y!�~�D�@"OnI���A�:̘����l}R�"O��(�h��4L���c�^�"r���"O�Ar#	�+fY r��W@����"O�� +'�����*��@��'�̔Y�j��k3�4��ʰ\�<�C�'i�T��Aֺ9��$���N�P��'�0	�nj�ٷ�Cr�IB	�'u���#�Z"IA|%17
.9S�a�'�R�bb炽c�t��̂ \k����'a�aa��C=&�q��M�
@�Hq�'Tq�1J$0-�1M<��9Q�'x\�H���
~�~uZpf�}����'�@�T!�9�Z�r'���p�9��'�*(�R)��a�:E:��B�z\�@8�'~RDeN�!b�a���k�bЁ
�'0x%�a�ԣ�p��1N�#p��U�	�'�F�%n��W��D*���4 	�'7ʬ�wN�-)f���ⓠ+Y����'���.�����#�>5��p�'b�)�!Ƅ6^"M@����>�`��
�'9��pQQj |r3#ϩ/��	�'ǀABq��-�� �u8(�h���'�nԋW��N:�XzU� ?"c*]{�'���"*}����Kt|$�
�'ڠX��f��m��x��%P��dH�'N�0�E�0#p�``ܳ6��
�'���%(F�������M��1r
�'���2�S�2���� !5b�i	�'�tP(di�$�)H��_=/\���'��%��yCf���$K!�'����B�u�D��FJ�kF��
�'��)sA���?������<LT��'JB���NB�;׸${"i�5F#N:�'�6�y6M��<1�a��*9�ɒ	�'�,��r�,�����&= �"�b�'�@����`
�rb[!pqXJ�'��.X��j���:#����'�x�GL�IA��#׍߿i�1!
�'z����NO�VL!0v!,]��1c	�'�ڜ�'�/T*Nm�V�F�M�^��'�H�p#δ#�4��@�V�F~n!��'�*��ao�/�n� 0m�<w����'����b&"+�1!DOK!��B�'���eL:RcFU��H|$�z
�'8�L0��\X��D�Bk��u��c
�'te	��X�~���Fִk��
�{��Ӌ6x�8	PˊCh8��Lò� � ֏�yHȄ�*����K�"K.��D�_�&N>܄�Y��:��H%}c����b���n��刚�"%mH4̘>|br��ȓ�d�;�OE����aT!��oU ܉V(��v����V I�'6�,�ȓq���K�&� E4AKGA�#1ν�ȓx�N(�؜#��]y���??��A��'@.�@�O�T��P���?�P̳�' h�I5z�ؙ����/���`�'��Y�g�Ǣq�|媖�Ѵ	�A�
��� PԑsP����#,�$H��ڦ"OR���N@�U���h��Q��d�"Ox���N�L��)"e�vwd}k�"Ozܺ�葼[n8U%�@)bP�J"O|\*#�Z�8��"C��/����"O�A�0n
� U���3$�;IvV�7"O�e����]�z��1#C�U���W"O\��R �#��JF�pr�"O�TFZ;}PTY`#�p�HQ(c"O<���9�b� �)D��h�"O���ŊV�w��A�5�z��@��"O��䕲�I�n9��h2a"O���lS��Fp�1·3@ ؐ`"O�q�W���0�f0�sm���"���"Od�8 kR�3_�@3����ĵI�"Op5B�|�Z�Rt��,Q��|��"O��ca�ޤ'~�%��N�nT�"O�\��\�5���8�Û�b�j�bS"O$)���šZՄ��D *M��|�a"O�񦊂����	Q��a���"O���NC+"v��L�i�D�a�'���q4&�1���2 U�ܣg\N�X0#��*;�&�Q�b:D�L��dئwM(��BI͙.nX5�/�<��ˊ%4d��y够��0��I	�n��i�l	^\Ľk�B�*s!�DKc��!v��P�,{���-'b��&��c�XpŎI2F �Rb���}oA�U��I!��ğֈ[p����p?)���<M^�	ae�Zй����e��@5�S<ur����n.4�Pۓb�|IˤF�A��|���:�°E|B��h���`e���|lk��R�7����S�Pܔ����:T"� 6m��yML��%���F��db'Q�g�N�	.�JD��'u$BF(Djg����a���4��'GS��L���䃇-"�}�	�'6A���O�d��V�Y�#��t鑁�	l�Tz�A/k��] �����	�2�|QN>�6�Gc����e^#D���%�NX��`g�K	�j�P� F����a ++�t�&��$#�A 
{
ؙ�7jC�yr���w�n��(�*7D*V��6�(O�asC/Ѐt�`5�7@.>V8j�m75�h�LA1KFP"�/�_����K;��DA���}��$h�T˶$U*M�^@���N���I����oLB��T���<���0q��%m�DӖ��L�XH�����yw(�3-Y
a1p�6EM�²$��y���>Dzx8�H-~1(�)��dPx$�ӄƆ!] ���V�5��		��F�>Dxp ����K*nx#I^�yG�ܠ-�UP4%��B.�|*RG��p>y�)H�G6t�y��E&=:�ܛхѨv|&1�� F<�HI�cʾV�"G��2:j��y�(��g둄C�~i�3�E
U��=��*
U ܓ$�M�_�2,&��"D���e =I����*�%,���u�S<��p Ҝj���P�8�O��j�(_�\D�)6G٠2�HD	�g	,g���5��gx�9Z��wq��*���1^@�1' 3�HH�7��dc���v^LC��U~�X�
O�5���5I�x��oвNg\Y�i�8C|qD�$I�%�Ć�y��)��$��M�h�ԯ3MoNq��ɝ3?MLS�k�:~����ISL��|b���0<��τ-M��tB�ES:n�-\q�6�@�\6D �B&�����XW	�(���8�@�#.bx�H�Lw�*�r�h���'QI`�I��~@��	# ]�E��<��O�0;S总���I��
 
�.m!a��07l��Hݝ=� ��(��\�y��U�Mf�Q)�$��[0�,E�$
V5�T�:|O|�Jq�ב8
4ę1d�J6���Ŗ� p	��@�H��1$��XZh�Γ:8�١$LH6��5���d�^�&�V��o�U"	p��S��4$/ޅ"��8�f%�.g�L��kL4�h�H��#iT^�z�N�D?yf�FV[ a�jV2uG(D��战b?zQ児�C�h�"b#�4�ٴ���2�""?�f�W �ݫ!�p=ĈIu�ݣm=��GˋIc5��E�"����@@�A~����ёkZ�=�]�O
�KtJ�Lj��{2
̌=�4@ɐm#ZP�������$��n�����.{��S��F�M�D���Љ)
:񒷎J?Sej̡f�ܥO.��F��WB���M�nL�m�$B_ip�Z% $\OnArҊ�{I	�� A&W'!��Ѡ�4t��(p��n`YB�
Q� ��GH� ��X�f֤'�N\z��ُ�X�T��~(p��'�������b*�ف�nͮ"{���6C̉H�l�Jb����B���n9ּ�O-c!���qL�&|ʘ�V�K�b�rf���0�Y�s���LH���)[A.#?��Hh}�ѻ��)�EI��xZ�ʈV�2=���;%���2w�K0P'���39�@�s��/w�4k��
	U�>%��iz�Z>]���
�.P:�Hr�M:-�y�'W�e��	�>f�Y��R/��QB2%+�\<����n�:�ڑ���ry����:�tl���� 5!��;�D���Ǘ 0�z
� ~�Xa�/��Y8�b�8Xj�$�Ə�rah^!+���u �O.p�pA�A.��}`Bb;^j��Ă�vX���dF�S�X��5�I�%6�!W�'^��$��o�l�j�.x=�-� ��%2�T艆��Q�f��]�[eJs)�i�~�"��z9�%��$�%��5YZ�����<��Aq2�H�.��MA���
t��B��Ȇ&��Jwe�w1�:�䔷&�h�c�n�,���Ү)fEFmcҌ�;���"��,.���"քT�$�~�;�}L���Jr�
��$��=�q冗����
mM:}K�
,��ٱ �)A�X��D�6d1���"X����A&\v@�q�e��,�4��-zJ|��5X���m�Q@ͿO~��x�@O;)��i���������	F
������o� I1��>M{��H�@�:*�����%rZ̔jg�O�k���!�4���'��a)@���d�0}K��L.&�y��"ͣ ��S��7%���QB�z-�<*X$�5�Ĺi����O����L�i��4s�	�@�ȑ*�Ym��y�N�A�Ν24�E}�(���D�'�/g�0��ʘ3�=�0)w��	TĚM�ӆx^�����B��?� �����+%F����$�"�MIS�|�W)�E�Ogʉ�씁 � �ЀN�:���u��8a�L �^@����0{׮,��}���?���5#)�"Z��� ⊍� 떽h愃�A�f�<�Т	��>!+�	I�$n&=��&.��
�O�@Z��e�q��'w��򨂳F�����"Uh���'u��痢� Hv$P�����P�U{t!��7#ڕ�@*]�Cb@�E�:dߤM��ɄQ�T5� ���0L;�hq�b�9?>(���B'!�65���0Vĉ�O�$�pC�g,���06��q���1�l��פ�EPb������B��-->Y��,�n��ţ�
h-c���e�L�k.�xB���t0�(7hǙѤ�a#E���xb-S ��}�C�����:�n��x�l��/^G(<�e��7��iB�쀢M�"��&��J8����i�r�G#���` �)2ژv(.;J~��ȓ[��0ą�9wđrR�_�{h �ȓqǶ�A&#� 
��Ѷ3z�D���1A#þ���q���@]��f��=����)]�y1"K�.NA4�ȓ%��,��O�8�J�!͇���ȓw쑉�i YǢ��2��XZ����l���%(ڲf/"@�e`E�N�U�ȓ7l<���d��okjL�� =L�u�ȓhh��%ȗb�t�{d+�aR�a�ȓ
M^�ώ�s�;ԦW�0�(�ȓᕧ��lD�Q�v��D��"O�i��OB�F��U�b�=�d�b"On�ٱ�Y3(�U���\/>q h�"O���险GLb �uBT,a~lб�"Op����@?b��
qaԚU$X�"O&A(�42ذ�έ���"O�ɶ�G(i$d�8$m�&y�r�"O�) Añ\����QL�K3"O(�[!hI9VZ��8��s�N)��"O���d(ġ^Ŕ����B�FI{�"O���&�#y�,����6|����"OHM�UCؔx��*��*S�>�x"O,�CTO�	�&���녾���B�"Odm���0v�����,�H�>y�"O<y h� *��<#�
Y�pX�j5"O�|Z׎iȱG��v�6U��"O&�����Eg��1 R�Im40�0"O�̒Q�K�E�RT��Y�ظ@�"O\�B#��C����+�1O�ͺs"O�+!O�LJ����_!^�𑃣"O�X�+��QR�៲g�"qX "O�iEe�QsP��Co��}�fe��"OJ��b/Ⱦ{vn�"��Uo�Rt�P"ONA��o�){kP�"A�|�RE��"O|�"�Sm_��硑=^�d��e"O�%C��ڤx����5�9�,��"O� j��%FE�#�X��"F��,�ӷ"O���옺N�@8)'�O?$��5"OnuX�(�萩c�f�*%��"O 9���\g��r�qL�is"O�|Ѵ�t�6�Ȕ��)�b�"O���6O]:8�pS�\�<|�6"O����B+����׌X66R� "O��a�(/b)Q*I�84P<�"O�*���Jk,��A�Z�aA�"O���L�6t���X�� �P�~�HR"OnC"��#^�8��h�39����S"OZX*rƑ�7��ǉ�&�F�P"O�;b��=�z�F�.
B�a""O����s
$� �d��^��p"O��p`�ͯJ��P���)��V"O��:wI�4\vSe/�:�B�AF"O�� A �323�8-�'�h�8`"O`t���i�@���-�y�j�ۓ"OP�j�A�x� ]Z7��GF�3"O[��R�+��
�
��t%0���"O�%�t�|�.c�J˼/.�mr7"O���d�\$�H ��i\#��h�*O��:&̗�(0N�`�*/Q�k
�'
�����ʉ����v�ŀgG��Z	�'g�ã��@8ݱ��[���a�'�
�2��2e�<�K���^7���'ޠ9�mP&c�Ƒ���9L��؉�'eZ�s �M~Q�٨S���s
 |�
�'4�i�4,ވ���r���$J�Q�'�qÅ���(�ɟ;2�r�'/���#�I�9���\���p��'}�]&�+C�l�Ңy��P
�'�DЉc�����s�
w�Q�'�,�`���L,	S!`L��j4��'/������/k��{v�ĊpՂ�'��|:�XF�y� :P0�B�'`�Ƀ���n��0��Y�|��'tV@bEֳ_�M�S�B*U�
Q�'�(��®ʅ��D����F`th��'op@���ɱ~��4�"�(8 1 �'�>�
�%�"�|�g��	dT	���-ٔg��j �wϊ�[����'R���%��Cb\5{��7Kg.��'&�h釬�<q�TZD�@�p��
�'�����.�9�Č��"Q�olȡ�
�'@�S��]KpCB�s$�Ii
�'����K�U^�*K�<T�T�	�'���R写"c��F .���		�'�J,rg�S���l��'�\��	�'��ai �A6#�.�z怸�楡�' ���#5q�<Igb��E��'�f��t�U>br��6E�]+BLh�'EK��7H��&�9�Ll`�'�FE���4�h$�p(װ �\�2
�'�>���5VM!�^� ��@	�'̾����XRm¶�3�`S	�'����ӇD'@-()Q��i��'0x,9��,8���@���0X�Ds�'���p��/`���7dW!BVҸ��'��qE#�1#Ct�#g'�9�ഛ�'> �#4'�(�0Ѓđ�<<x�'H�T%C/o�*%���Y|�Ɣ�	�'O�Br��MR�ʁE x�����'vzA��BĔ%B�3���x\�y���� ��(-�&��&��I�� c"O�����(�R5��9,��#�"O6�:vo�5u����v���+CZȣ�"O6ų�@7Ro�����.OFX��"O���k�:T�ȁ��U�U <��"O�� �ņ&$+$i1�B\[�p"�"Ob���ɩb�8�R�ᄉtAxH`�"O<���a�L��ψ�l��7"OUCS��G�ȵ
'M�6uL�|�D"O6E�B1�zբK�+����"Oh5�7�{��Y��
�`S"�r"O%h�%�P�p�"�#����� "O���t	�t^L]�r��.E3Ԝ��"O�d(�b؆;��h ��$^D���"O�l��H_��4�a#M!l�5"OP8�)��D/���R�W� p|��"O��R,�L�)���Ư<&�#"Oʠ
�)�/\�N�3!'D�3�"O��Y�i�2���K��܍P�pq"OJ|�V�Ҽ h,C���S*Z<"�"O��"���"l �S�!��%�p!"OlQ�(�4]���QH�8/
ё�"O6�����РЀN��8
v@"q"OD�a�G�
l1��u�ߌ$�^��7"O~T�4jI�|��p��֊M��3!"O��S���C�LJ��)U��4X�"O���/~��Lb��t��H��"O�e�j���mB�)S
G����"O^,q���U���z����&f�2�"OƘ²*
!/fƑ�"_�Mpa��"O�[�b� H4��眆J���q"O�}"�͕�oD�xp�eڗ)�4ʣ"O��0����g���swn�c'��CD"O���f�ؐ2�Xʱ�T�`s�T��"OR���G�����Hs�P|����"O�(���K<@`%8x	xW"O��������b��M��M��"O�ӡ$��<��]:v�N</wt�K�"O����3+`�b��JsP�R"O�@���\�  �'a׶|h{g"O|���$��?�R��/����s"O,�c�J�=Wa��+�ș� բ��t"O��6'�2v�@a:�үt�,9�"O>�:%ӱ-ST8I�b���(,��"Ot̓&C�t,p}��1&kL%3�"O�l��˒�*�"���ϙ&w��"O�i�"�+OX�QZU�Wwb�@�"O������S[ntQ��ߪ<���"O��Q5l��Lw��vF�.G�"���"OZ���)�M?�m;g�ٛX\�Y�"O��AV�W�p9N�p��,T̨!"O�%+���R6�	�,IQ�`e+"OZ�B�Ĉ0crH!���+�HJ%"O�%���	���1 A�Dv�K�"O�0"�c8r�TѤI�"2:DI��"O~!�W�?q��ŦN:_>�<�'"Ol$#af�=�u�ڈ�*ѓ�%D���cD f
�S���Nب`#D��:��E�e?��i"J�@�H����#D��wf��%8��H�]�?e r4n4D�����40���kZ $�:h���/D����dL# פ%�`�E�lCv.+D�(#��
`�p#��>1&�yw�&D����*aR��� ����!�E�'D�� FY�#�&v����pH�>w�6�� "Ob��6�2��2E��B ��E"O��A
J�>�Z��c6 X�X`"Oe��T�S�P�Jd��);4(���"O�,�Fc���n�S�B� -��*�"O���tK��+Pz�3 ?.P�j""O�l+CɁ	V�n�X�N�$:;"Ot2i>e*���L�A>.�f"O�`vMQ\ک���q��	�"Oz�k�e!��L#����P�H�"O���!�\^3*����ĥz�i��"O���N�1��}K��0�\I"O%Q�͕1jY�ICf��Xl|�c�"O����,ִK���a��?an���"O@!����'2b^%W�Z�[`�� �"O^5ɀm�&������|]A "O�5��Y��}���X�dEb�"O0=�����.��w"�~1���F"O$�X5B�ɡceR�8�4��rm_�<񒡛� I�Iu�Y9��ET�^�<�A"zj�x"� RD���,|�<Yp�D,xj��c� �S�@V�<��	�!{n8ZA�áG�hm;#�Q�<�oñ"z���CRK~��ӀH�<�V���T����ӠA����0H�I�<1�*H?r�D�t��8��ʤ,KG�<A#g.>��)��@�L|B�	s�K�<!�KP�m���i��1�\� �^�<)��n��<�6�1p�d�At�Rg�<9"FFr�:�7�.h�&8���Z�<��A�D���+ .�O~�0�m�<q�l��T�h+�2��I� �l�<Y�(߰J��,Q�g�(6��p�%d�<A�S	.y��(N�'�X�t��{�<	F���X!����P���,�o�<CS>&�|��Cb&�Qfk�b�<Y�AҶB���K��З{��<��"QR�<�w OQH���Ӎ%�n�PUȕE�<��& O���P�[>:���dn�<9��%�p�0&C)'=��QA�n�<��K�!�xd����]Z@�����r�<�&$�!s�TR��Ec��.��Ć�2,D���P�[��"W(�&)���ȓvk��I�KώV�J1��Wzp��ȓ7�X��N̢E|n�P���S�̭�ȓ���a#dɧ;C"eP���|���ȓ��]1&)HWDi t�I�v���:�D�A����k�ӑH|�х�wfTA�ՋB�l*���!)�x݅ȓm��h7G�6r`�<���A�+����2���4�]
4�$����*0=X���*���8E�X���Q!,�\��ȓA+\�xa�o����Em�Մȓ <T��t�V#{:�uj_�*	�ȓK^�$�#��7�b`0W��4N��̈́�>��E�1���	�P��Ӱ?�D��sh���H�b�1��˝�P��kYFEy��^��8B$���J��ȓS$�}Ѵ��j^�[�O����ɇ�	��� �B"UF�z�e�=hl�ȓWg�A`v���#���Z�O�Cz�܄ȓ^�`!�TG�zx��wnR������X�H����5�8�Y���!1=���arrx�S0�"T"��!%�䐆�S�? z�"!�ŭ|t�ӗ�W!H]|��"O�<j�NC6"��d�"L�4VM�Q�"O��R��]��]h�N(|<�e¶"O��JP�N,,~��RC��'�U�"O�pS��n���q���F�F�г"O�	��J(r-@ѠS�˕P��0�P"O<Hk�L�8*A���嘩_�\@ $"O��LC&�@�cÐ�Yv@x�"O<�9A*°8	D��Cc�\3�"OIP�W���u,ۊ_3l�ڢ"O�ث��$,H�!�E����"O�A����gply ���?z�I�t"O�	�E��5�6��g�U	gJ��E"O�51A@
������l#�|"O�yIB�Бc��<25�Xi~1�"O��K���B\�mY���i+�!"O��g�4ex����,C�=��r6"O�M�v�P�E�%�%�)uI)�"O�4{�M�2^�������e#�	j�"ObA�t��;����Ę"&�(g"O��rS��S.D���_�efuX�"O�,�d�ۘ�M����E"O(�x鎷#~��c��:��cf"O$	0&!�8�����E�y�P�s "O�u)U�.]:Vy���:�8�S�"OP�jׅ�H�aǃ�9f����"OP�شh�д#��	�8QR"O�L��� ��S���0T����"Oj����V����3�:|�LCw"O�Y�D�)/@����L�Sh�I�"OH\��%4k�L�3ɀ�6��#�"Or���I�S�h��di����6"O��*��Bk�4I���V�{���"O$�ۃ� )"�3&�B0[���yB"�3?��V���dX�t��� �y�MR<!� ����BD(W�z�~���1e�aĭZj*�0Jt��8{��ȓ;`�P���PT�B�H+�Շȓd��a�򀋶g��i"��,MFd�ȓX��-�3�ͣS�80�^/A3���ȓ}|�cK0�=DN�+itՄȓ�\<j#6t�� ��9霰��N�
�JL�F)
��v`�:ܶY�ȓb5~h���<-~�I��=:{va��Zԕ+@T0<�qÏ<P���t[��YRI��8�Y#�;�.Q��vp�k�,تc�@�u��8�%�ȓw"��f	�PE�I���)�Ƶ��.}�m�S�"���CC(_L��D
���! �PND���ӦfZ�ȓC��ER��_,<��;N�>B4�ȓUK�8
�a���PQ�Gt0��ȓ,��H��@QK"�������ȓXVn���ݟN ȀA��$]���`^5������<�����)Q�܆ȓ|[��%GO��� �Z��ȓ�T,�7��
x���'M>C/�I��Y��ఴC� `����[�� �ȓ`��ps���9���bN{�p��C�\y���P}�с�����ȓM��9e�ֿwY�P�"��\u��	8+z
a���)�$P��NO?v��5
"�%��=E���"�|r�O0=D�Oq��X�'H�e���2��N�*���eS��;��^��
�A�,��;�XRrT?��S
/ {����Q�^]�}�Wƛ;���
���1�����y�b��� n�(@i# 3Ө�ej-Ö���8� �&b@��A���la�V�(�(�2���q��
>&Ab��A��O�(��w���k
�'dtz|��(�1�t�B. �HbTiKV�'��ˡoG/� �4f�v>I2d6^5�\�� ����&$BTe�EÎP �Q���h#��s��L�9�DP�u���7>�Xc�X)g~��lD%[fj�r�ε6��z��7꧁u7�A�l2�M `�/zh-inkB �6#���|5����V�d�ç����7@
Ř�'��!q��B�!	�	I�}K�i}�'�n>Y�&'�"
b� %f�$b�|ٹw�Օis�()� F�PcTH*v��{v^�	*�W�fQ+W�g<�=�g�um,�x�NV�q�p�s�#�{'�4X��M>U;�⚟l�.`ɞN:�M���5/���Β����贳iz��F���Z�}ax�
���^�������y㠠��g�t�qӋ6?���qO���������7%�n�7��
lD!�d�A`U2R#�4e��!:d��Fb!�$�1A������]�������QL!�K4W
��K^g۰���EGF!�I����"0��1D�0��WȜ.7!�QG��U
�h�L�68�Fˍ !�ğ���4�N���\�qdH�q�!��K.&���
M2:��Zi�/�!�D����9��q�R���9R�n�<y$Dv4�P��,���'[j�<YW^m�85��.�&��)P�<�*��W�j�0���h��tA���M�<1��S!RL9� e�+:������J�<�P�F2hx����&y*Z%�"�{�<�c�I/?��@�%T�Q蜫B�]A�<�D�z �9"샦&���8$O\A�<�q�M� �()Z:_��p%�y�<���TD9�d� Dw�`8%v�<�f�
p7���4��sGXّӮ}�<���߭^�d��Gh�l �c�|�<��Z,e�R8�cG�b[#�_�<aVʯ���ڣI�*���TOZ�<� ��������8c��bV�<���ɼ(+(��I�ꤱ��j�<���^��}��.�1
���9dj�e�<I �W� �,�@���<@l1���a�<1���))���G�H�L���BIw�<�7"���(rA���4��<Y�# q�<!�`�7�X��%H&9E��P+�m�<!�"�)/
�5���
 P5�8p�m�b�<�NP��D������&�T(s�<)碘���� �Oĩg�ha��$Qm�<w�
77��hsT� 	��UyņNj�<I!�J�D�Ьۥ/Y�w:��u�O�<)���'R<�y��1cY�`H�I@u�<�D#�L�Y;��/@&��h��x�<�� O�YJ.�r�AU)E��MXS��s�<��&��=4�i��� 𔰻�.Up�<I�B�hYHm��Ϲi^~����*T�`"�3	"��UHܞ�`�P�H2D��I�荛,���jc�؃L�$���l%D�Q�GҵGb�d��Z�"�21J7D���3萿R�h���j�@����ZC�I�;�`q�`�R,rA�\�W$Y��B䉑:��HS։��.�pl b�~i�B�I?���S��A�i�p�y��	�dB��G��Q'ߎ$'�Iklۜx\�B�I22oB|�(�$;��A��똃QQLB�~���Dدΐc�V4T�,B�I�k3�A8 bS�b�be��.�z<^C�3=:��! �a	�M���zC�	-22J5�ëG�5��mS�lB=M�B䉒IP�)ڐ2rh�P�h[NB�)� �!�0(P3�^-����W�6�;e"Oƙk���V�4H�HR7xW�%t"O<q�4H�/k�r�AG�0L�� "O��b
�$�
��f�h��z�"O,�æ�_�*����G�E"k���S�"O�,Q4�ьpP���ԅG���홶"O���i_����(��X+'�M!�"O��ɐ��==��E�aC�TP��"O�\Y��jM�q`J�8Z�x��"O���و6Vu�U��%o�Z�b"O�AS��*0d��)��BDӅ"O��E�I�(��p�[���)�2"O�$��n�"ʺ��ʘ~��z�"Or��-�0h��s�@J5��h�"O��Rb�]3e@�ʗ�,�Z�"�"O i�cOó%��]aG���t�H0�d"O�8R@�/��I�MK�V��|��ȓ+��9�%���4=�l!K� h؇ȓ/�f�⡂(F������eΆ4�ȓ,oX�j�Q�"����D�~�`��ȓ	e�Ӟ-D���'	q���-\���l��l�������z�[��ek�m��NV�rf$8Aa���ȓH)��s���^����A(Z.Da�ȓs%&uv�O�z� �R�ӧ��H�ȓ�^M���J$�;����-B���ȓy���GÛ3�8�Ѧ�dy4��,��I�!B�� Q�^jj=�ȓ9����H�l����QA�P�ȓ鞰�S���,Ք���K�+|	�ȓ]�C`� �t�D���<!�Q��i��4P� Q�?v�Pjԫ�=jΔ��<��'�ݠYd��& ��?>��ȓR�b�"w
ѣ`�Z���F�0L!X��ȓd�ѱ�%AD����/D��T�ȓM�Zk�d�u��a�@�����f0D�Lj��ނC�� RPN  <:���,D�H��d��Q�S�z�J]b��&D�Lp�-�A�Y؉pE*N\�dB�	�K����b��o�Ib��
9�nB�I�.�	���X��i�@�ǜQM�B�I6��k�n޶BЉP����}�JB�	�Z��U�T��h�1��4&0�B�ɸ'�|���J�"���CpA\�f��C䉡A����+x��&g��D�f"OP�aӈWk�j!쌰#Î���"O|d��j�
T*�#�?|��-��"O�qy-˔K�tt	ש��&|`��"O����BŵgW�Tk�gD�it��E"O�=hti��o��r�fa�@��"O�ep��R�i��p��h��1��4@3"O�Uk��ʠ"����hU�,��S�"Ol��DE�*#*J��MX������"O�ظ�j��v���H0�Ϲy� }�V"OZ1����ܫ�j��v(���"OB<�T��B`�X�ui� �H �"O��������Y�EH�6�d �0"O���U�Q�� �F����W"O�BN����� ɦU�%"O����aZ�v��ͣ�oJ�]�Й;�"Olbb��7_Ț`���Y�Sh�� "O
�`!IX- 0�2s'�W^v��U"OL 9Ӈ͟������%R-�W�^�<�� D���Q#�2P`ب2��S�<� ��'�.#�:���υA�m��"O��B+�8A��ɑ+K�E�"O5�����U�`���-�,�
g"OlA�V�Ua�rV�6�d�r"O6��  ,f�e��ҝ}(m��"Opd���X�ބ;!fK7w���"O������k�u�cۍP��у"OŘGj]�/��պtE�0^�.�[�"O��3&EY`4Qx ��x �Ȩ�"O�۵
�c�mucK�P^p��V"O�	W ϔq���G�x.6ɫ "Ol�c��"uKdn�+5��e�3"OTxҡ�0k`���X�{�`	�"O6�t�Bw~H��S�O%��6"O�A"�n�5g��0b�#�ĩ��"O>���n�"rN�t��`�e���S�"O��2J�ԫ���jǸ}�$"O�<��17�����j�����"O�p�L1#@58��c�t\3w"O� ��R;#fv8!%�* u)�"Ot8��GO4.htQ5C2���8�"O
���BD�,���)�F�g��e�a"O���b�	$�i�DGE.^p�R�"O;b"Υ7=Vh�AlқhBl)"OH��#U��r6+�!F � �"O�$��b?��\:rh�8*%�V"O��;ąO�J�����䗨(�"O����O�����ԅ��"O�a��W�M�����c���"O"X3C ?m���r-ř=N��"O��I��F:J�Q��K�Z�j�"�"OH��"��]/M��ꗍT�J��&"O@�s�,������*L,~�z�0"O<�"��;�6)� +P�H��Q "O�X4��)��8�#T�aa�"O�uеE��V�"v�J3G�T��"OD���g�]:�=H
Y#l���p"O�ii�HY�J=��`�1(�-#"O�aa쑷^jȅz�f�x��â"O��J�T�n�f(�Y� �h��"OZ�Ì�-V'�$
�
FT�p���"O*�`�U!ZE~���Jv�x"O�bj�9/��B����g=�%Z�"O�@�CD��jL���ߣ!��"O� )b�O+K_��KLؠHB"O��2�Hoƍ��$H�r���*u"Op�`�K�o�L`Ѧ�������"OB�� �4@��X�f�O�/~�#"O��c�$�.pY�j�<Q\�1"O��;��N=�\9�I��*;J�V"O�]��kW�`ꔥ�)̋v7X]�A"O0m��cŨ�����
�Y���"O�a0 �J�47���d+��h����W"O�1�"ᗿtX�a��E�(����"O�Iqѡ*yp��+_�8�]9s"O��jb�
�e��t���F�t�"O����E�!��r�Է��X�"O�%���� ��\[KY����0 "OR����ݍ~4�H�ǈ���"O���g�F�UE���fV#Z�� t"O$�u� xň�A υ�u�F"O��s4��g%��⠀Ɵi|%�d"Ov��Gn]�!D441v��г"O` �pIQ��H�Ua�,o��$�S"O� ���Q@W�#4�=�d-J$h���I"O���؎`����wiW���0�"O�l��B�j5��(�RCB(}�"O��#��/a7�88b��8�:M��"Or%YG���LPQ�T�B�N�Za"O�z�C�!d�sG�2:���0"O�E7�ŭ6�R �4m�b�ɩ�"O�����&YQq�)g��"O�̡�n*`�Ġ&(�d T�#Q"O.��QDZ�$J�#��R�/Q*�0"Ov-�U�$w�$	�O�:�5��"O�=A���<����>j����6"O�D`L/~���,��%4bh�f"O)+���#3�xXŌC��i�"O����ӯv�FE:$�ǟ$��M�"O�d*��̢&괁�ɕ\����%"O����S�,��x�O�5�$䫆"ON<KѨ�."b�P	�-F3s4�`$"O�IY�n��A�Æ.�1�"O8hj��[�fv.�cXm�fQ�"On�a�[Ί���`}I;4Ɋ��yaՊi�\�zeO�K�N��#��:�y��UBY�][Ń\F&��c��yBƅ;z�&@��7����a#�y�A�&>�`��f��0ɤ�R���yB@���0�ř!�����M	��yH�: `  ��   ;    &  |   O,  �6  �?  ^J  S  bY  �_   f  Cl  �r  �x    R�  ��  ّ  !�  ~�  ͤ  �  S�  ��  �  -�  ��  t�  P�  ��  ��  �  j�  ��  � {  İ���	����Zv)C�'ll\�0BL[H<yVCQ��F��e�P(������C�<��	��e��A��+O��$���X@�<�v�C��p�TJ��izsf�a�<�&	�P����w�&H�ؐ���e�<�0i�������^z��B�V�<��(��Fz,Q��!\:�\U�N�R�<yӅ�I~��3��,}��٣�JVy�<a㇊)nt��;G�ʏ���b��Kv�<i�B�r�8��L	�W6�}�=T��zf���R]��0/�6őf?D�haV���  ʔ ݿ���1D��[�
(m����@!\	{�� 7�.D��`ƭ�}`|��a˚t���Q3)-D�[2�ߌ=�v!����ɳ� 8D�t���O�u|D�Z��Y�P�1c��7D�LÐmֱlGfPb��U̮L,�0C�I�[mH=�W�٠d��C�l�&9�dC�IMM^� a!1�>�Ie�?`'�B�	5Jy�]��tn`���JF}��B�	�v�6��V�+#*t�c2H�`��B�ɦr9\�{��*v�h��⡍��vC�I�v��ɐ�ƙ$�P(˅��=EItC�I��9��ǟ l�����&2lC�IO��P��(����'�lZ@C�I�aS����k��p,rI�3%�`B䉅%���Gk�S�X�z'.�#�C䉙U���@
��K�V�j6.����B�I6\�qi��-d@��4�\�Y�B�|�d���a϶l	Ҭ����_��C䉈-�I�����NL�,�ب�E�8D�l�C�*&�n�h��Ώh�YS�j!D�h�$�$!��0*$�b�p��� D��3�X(q~T�אFbv��K!D�ȩrMY>n��ڵ��$V�$�P�5D�l;'N��d�MJ�6[EHS�%D�����£j|)��f�}�� �L?D�,q�
ۨP>&@���S�b��K� !D��`�AJK[�D�!�Y��dZ��Oj4���wyl��p̂
��: GǄ��̇�I\�'؆�Ȣ��{]؈� j]	����Q��/���
���?����&�>6EZD�O��=���bRjI�u�V�R�Ӂ�Ukܓ���H�(���#;���D�ŏv�nqjw�i�ў"~nZ�a��q��e6�-�0�	`"=qǓp5J);tGO3�,e+G��(�ц�s��Hx�V>��RӠ��bʎm��݌���G�9��@�׮T�xDb�S� ߞ,�B�őE�Ψ��f��=�Ó �6�+��^ HZV�2��[���'7ў���I�|]������,��4�Қf�<9&�h���Ϙ'ZLL)�@Khv���$�
D��	�'�ў�}
���'o�����'q���b��K�<ɓ�G;�$K���~G����^�'9ўʧG_�d@Xi�¤0���;���!��	V�O��=B!��.j8�x�Y�6���+*��hO��G;���6'uD4q�g�##�Q��D{*�,�W���P�F�`��	s_Xt���=�S��y�/˽*R�k��M.z��,�΍ �M�O<��O?7�L�R���;U�Z+�|���%ȣ9!���nw ���,k���i�F*Q��F{*��ZbȀ�<b�h����$2=r�ѧ"OH���,��*�~5�M*��B��b>��!�P6�8��`ƕ9��ɋ�"D�� dC�@Cx����䂘?n��j�O���=�Gˍo�hlAGN�10w��)ӎ��<Ɉ��S5}��L��@�d�l�V�ڸ?�C�Ii\�D�ҦR#d�0���C��*�~E�E�	��Q�-�*z�#>���d�~*R��wB�k�-63"ɸD���<I
��[��TR���:�(9#e�y�����Vr�r�#@`��t`�deV]�?�	�q�,�5'�	5ȍj@�Z�������YL��1O��R��'<E{�G3%�89JS"OQ(#�''+�����j�R�r7��l?a�{B�T-L��֝�v}��R��7�Rɛ�Y���B����������GO��m����	٠z�V�>Ɋ��O(чmF��j���-����e��IG�O�؂'	��l���#_�h�~P
�'��=
F+�ٕ�W����O��	f�S�OFXi3'O1��yZЊ�36�����M���E9;��h2	�� �m��CM�<����0~5�h�݂\|i���K�lD{"GW�Yh�A�~��qQ�N�����<ɐ�'Fa�dJ;'Ն4B���T����Š��O�~!�@m�p���ΌgOt]�'�k�'��xBd��tA��y�7eXMb�(O�=�O�*w�5WK�u�1@N���Ұi�!���8xb�1'̎qQ��g���O!�d�R�$Y"閑FY�}ZA �(�!�Ě�R��$�XbR1"���!�D�-B>���ŰQ� ��3~!���Q������b��!k!�����lӢ�EU�ْ�B�ip���E{��th��L���-#U�z�$5C�"O���G��/;oHE��-��Jv�l3�'Cў"~"'d�c��H��!�,/.��2���ybfүt��+e!�TjB�߷�y@�&�<��	ׂ�lqÆ���0>)H>�rC�{ȼ�	���5Y��K�~�<�����i\(����ڡ%SNѸ�gP�'��Hp���H5�5�����)� �:wQ4!�d�-��D���(Tvu��
/)&�����O��W� �G��irQ��[�s�"O�\z3ě�1�Z(ёȐ�cX�D�U�O���D�;%�<�hv��QL�A����{�!�gm��3B̄��B�+�!�X ���g�1/D��g��?�L6�>�~2R�dT�l>BF�i����6"�?��̋ac�"�� 3�^�a�a���S���
� �
�� �F(A��enZ�P�v�O��'���MC�c>8�,���$O<Nm����H�'��D8?.��a92`n�/�%x��J -K0l!��I�},���i���n�|�� �	;D	�ά2��D�sk��L�H��A~�j]� ��q1�Ysr!���:I��(�a���a&%�Phr(�v(�u�A���`���?E��'y�Xc!Ο�]@�k�e�!=|��),O����I7��j� U�NI�<3�&�=U2�O�NU�g�p�EZS��6�1��GP�{X���I~}r7Oޝ��D��.�Eۑ�ʖ Y� q�A>�h��lT ��-R�o݂(�f"<lO��4��]\�� ֍{���5�-D��8$GǑ���w��*j_b��0��~�S�o:.���O�'W��1D�P�Q��B��#U�9��C?bl��"!����X"H�"~*V傼qp�(SGت&�0h��=�Pxb�iҶM�g-�-F�`���,L+���P�-ְՅ�I�V�}���^�F6���O�8�VC䉽j�����4TV�h0 D�=OHC�)� @	V-֣ t> ���])��p"O�=6�^9P�h�B�!dJ�k%"O�0¤
v�@C T��((�"Ozz��_�� �N�G�LI8���i�O���j��]�$n��p�u�&��2m,}��Oh�����~�	�o����
/傉Ba.(���'����D%���?�̽�V�4s9f�R��/1���	b��H�ׇܝG��e�t/SX{�,s�<��5�<�D��O�&8�$�̢~����'�a~B/C-te�EHJ�)l��fj�	��=��yb.�J�pq�W-�9z`����y�%M� 
Ɋ�]={���iaN��y�f�,?�9
�'o�A�@V��y���E��Rk�$y�ȲӠ
0�yB�*pt�m#Q��=f���c	]��Mc�}�4O?7�A�!td�r�jӄ# ,�І&� W!��ڟB\�C1�θF��P���YP�LJ�'瑞��GC� ��#R
��L�$$�0�"LO21�4_�$��'e��	El�*����ήv�qh�'�
,X�-�:�\��%EC1g�"����d�l��6§'�
�P�Ƃ�=�R��f��d!��FzR�'��������N����܋y�Ltp� �	�<��'��(W�6@b��(��?�μ�6��t(<�B�F�9�l�W$9�Nl"PN��?�L<��}���=V�9���h�P��󯙓Kǡ�djӶ;�@0�\�+�R\`5��"O�	jB�[�(�B��fؗ[MT(���'��Ol�S��e�TmbAK�2HB BU"O`��A잟a9��2���e:�iA�.�S��y���zYƀ�`M\N��	a�J��y���,�İ#�N�_��<��iW��yriXP��zפT�[�n̙0N�?�y2�ё����j��M�*e ���y��U%Z�@��ÎN������#�y�g�5
�����M N؍s"���yr.P�5*�r� ܸ[\�T!����y�*�(�xq��*Ob\��m_!�y"�ϠI��)���Y�E���w��"�yR,V�\]��NYE�����U��y"䊱w2�*`�'�x��@Ӗ�y2H�`
*D*T�([�򘢖�U�y��X|d��B��J�����+C��y�̖Xp�O��Mp��c�Q��yb�5NV�U%�|]�-)��D�y#�	搈��8���pPꋯ�y�+(����������܉�y�aU .�B@q��Ե
��2%D���yB��>��i��ن+��������y�K�~�r�����<%�t�%K]9�yr΢!��yE��&Cv��dFO�y��
��H�$@�7��JDc��y`�>�@5�I�
%F�!��yg�D" pBp��T�1��$��yB����±(��J��8��y�"�7M���DC�;��"R���y���bO\�FI0�d��A��yBߓ/]��Ð��x�Y�@B�	5I0Ȣ�b��x�� *u�hC�?2J���3�!g֤ �v&=k|RC�ɏm�� f�»�8ͩVO��+�C�	�N����F���5}2��;�C�v�z1Ȣ3��T#��NV[�C�	�c���P妔�h���p��V<�C�7ꀴy��)I��А�d���XC�)� �����~�B�q�Ə,�.�3"O����``�$��P�"O���CR6l�j��[6wy5Q�"O�$(a�����`G�w��`�"Oȡ���N��u���ZZ�d���'c2]�|��۟����`��؟��I
Q��IR�1�� �c���f��I���	����ß���ݟ�����`��%ym h�3��P(蔮GU_�h���x���d���������\��՟\��-G�p0�D��
�T�BƁH+q�,�I˟p�I˟���ş���㟤�	�8�I�!l�� �ȡ#?
a���=��T��֟p�	џ���㟸���<�Iӟ���` ��KǢ�p��x��!e4$��۟|�IП|������˟|���d��&Ai�03��S�D�Q:f��%�6�I����ٟd������t�������%(m����)ۀ�S��	 \������ �	�� ��ƟD��ş��Ο��I� �� W�T�����(xe�	�����ϟ����������	ӟ��I�r$a	�mډ`��4�L��+����� ����$����8��Ο����X�	K �``L�:]��5!�@�C�(���ß<�	ԟ���џd�����	ʟ ��64QT� �oF�7*�t	�&W�D�T����l��֟ ���d��������ɋ#����o�6��%ы@`G���I����0������	�M�!�i���'n�% R����r����/��	"�����IK�It�����4�Q��J^0���b�i�E�HE�qf�<y��i �|����^Ŧ=�w.J�y�`���-ҫ`������@����IQ_��m��<�)���H�fX:+�ԝ�'QNa��-����=�@'�7������O���h���D�(0��⃦�<%��!4��զ��"��U�'@���w����B�=t[��uhW9r�.=�Pg{��o��<ɭO1��b�*r�b手S�yӡ"�q��EصA:Y�J�	=�l J�Յ^JԥG{�O/R��$�D�pGJ�K>��[elQ��yRR��$�Xٴ#RU�<�% B��,+�/��`�T����Y���'��"��V@Ө�I`}��ѕ6�š��A��#��?���F=-�6�1ҍ�V�1�ƴaRJ|�y���a�J���'��k�"�9��"8�X�.O�˓�?E��'o���X�g��!s�M7�<�ٛ'8,7�F�qf���Mˉ�O�ΐ"��M�&|��Թ.����'i�6�¦��	p԰nJ~B�)��z0(L=\�����
�P���2)�/��i��i>�'��O������D�W�����lN�*�xa��O^inZ�9>�b�t�s�!��̨6�ҿL"`�*p%C=/�=�O~`nZ�M�'��O��4�'�,=Z��T!� 	Q�ܲР{�ܘP�FQ#�O�������d]w$��'g����� �8�0�����H��I#����d�<)I>��i�rI��'�\�J �Arx+A�"wj T٘'�~7m.�i>�	1�MS�i���
��ʡ"H9��Y�VEҺ����a�i�R�h߬HZ�@=;l6��O��ķ���_c4-Aׅ�I��I��بf� �)�'\�T�����P� r�)�MB��ζ��[���H��G�5?A�iF�'�����/p��Dn�4{���:O�қ�h�:��ײL[�6�v���D�tQ$i���G&`Vl��q��6�P�k��(8Ō|2v��K�f~�O����QA�F�Ȃ=���̀B_����d��$� s�4&*���<�/��H���֝y���r6ߖ��p𑚟x�OulZ��M�'�OB���}��y�j�4�D֭�XL`�a�M�2�(!�O�����k�ޘ'9��!���j���
�{��@�/OH�$�<�|�'��6m�3BL	�/�.$�`�0*�7N|&@����T��4�����'Ӣ6m,�Be3�Ē�0}>q���4O�TmZ��A�E����Γ�?���w�Ȥ�`~b��bЕ@U�j�IXCi�y�Q���	��͟���џl�O$���E�0`�4$\�B`���s!tӂ�� F��	۟��&��Iӟ<a������p��U	fgS%3��4��	 ?7�������4����䟺]B�X�	�enF�Cc���,¸��s�x��Cǅ�^��}#!�V�'YR�'4P�X��.����H��!��3�'��b��M3��SD��n8�����m�D	E���I�r�>��i�7mp���'�l<3��QqXQh'!��r��D�'��-ql3�N	0��$��8��M|ݹ�����6n�2���`��+5ט�3B��O����O����O�"|�ߴ�?���]�CUҘ����1VPꅛD͛��?�u�i��5�'��O��'�剑q��a����szX9�"�&O|�Ɂ�M�P�iׄ7�V�&^6-/?Y'�5`JR.Z�2�`H���
<�G�ӭkpČ�H>�/O:�$�O��$�O6���Ov݃$f߭͞�C�f������<ᇻi� �'�r�'��O���F+2�d����Q�7����h���I��M�2�i����&�럶�	ƯHmr�2$�K�J��g��O��(
/k^Hʓ|��3�Jý�u�+��<��
i�����%���&e�g���$�O����O��<a��i墘'(*)��H�I	� ���T�;�ĩ[ �'�\6M!�4� ��'8�7-��Űܴ*��i�/ɦ\>�[��M�2�2u�N�M��'_2�Q6@�l���_�M����?Q�_� ��v�+c�nq�EMR�-H�i��:O����O��d�O��$�O��d22�4&~08�S1*b0U�����$%NXΓ�?��2J�����y��'�R�|2�T>��$Aɸ@�z�A�V�T�J�į>�D�iJ�7��8uht�n�Z�I�3�k?��q���I��E+VJʓ%�~0P�FT.��E{B�'��Iß`p�ڒ_<h@���!/�܃��x�(%��4�]�<����sȑ:J�ѳe&XU�i2���x~2m�>1��i�7-p�d'>���^�(1p@J�,4��A�o� &�HP�ue�/i8�r�*?��'c�dh:\wU֒Ob�
�NA�sf~�8��X'��٤�<������
ߴf@<9���M� y�ē�>�*u�$ S~��~����s��ڴd�:�;�bW&����c�;M�h���i�RlV�%��&<O�W���`����M��ɣJ��	3v��o��S�	[/|��c���	oy2�u�hxz�Ċ�h���еn������4W��Q�<��t%p��A�8h��â��	r�X@���!n�M�'�i>m�S쟠pǻ*�&<O�J�l3z�"hi�G�Dthp=O"1�)�#H��#n$��|����\�T��u�D�'��8}-R����$<���զmS�?才`�`�I֠[��A;:x���	Z�I����pش�y�T����
�R�f�I���q��%m�d+EhF�$ ��q�c��9��Ӻ{Zw� �1�d�Q���D"��8o�2ۢC�h�}����?����?���h�f����>��3�B�>��7�M6_iv�D�例�C%u������McI>�缳U�A,_���g�[�d���"����<���i�6MS���t,L��uΓ�?aO�:���5�K,\ފ1�pjY�%&|��g@%��N>�/O����O���O����O^}2w�3�=���.K��t�T�<�չi�viC�'���'��O���J�����Y8�0@1`!#��	��Mã�ip�� �'l���D��O�����'Gv�+��{\�;/Od!���ޚD����?����?���?	�W?=���R!��m"� ׂ�?����?�Ѝ�>ҶmZ��?I��ip��\�!i�N�٪���]�-��zY	�(�I7&�O��+�$�٦m(2An���u`��Ƅ ۴_Ť�"�nN�2B�bŢ=z.ia��ұ�Mk�'���������"e�O�rA��E)��Cx�	J MY4S��p㢢D,I�9���i�@�Iwy�P�"~Z�m�06��dƝ�,c����M̓51�F��.�������%�\"˛xB��ʉ�d � ���<��O oZ��M;��Q�����4�y2�'�����Y'&�+צ�,E���4M�*?��}�B�rlў�Qy��'��L�����|b�0�1��*u$�8��':�'6�f71OJ�����������F��F�҈0�2se���حO�o��MS�'��O��Ԏɠ6��0�Z;"��`v��$���#�>I��b�OB�i;�����$, ��B"R�;�9)��!Y���?	���?��S��Ύ��M#+O��m�I�*	#��m���s��΄~]z̑d)r���	��M����4�ڹ�'2�7���uAԱ��Ǒv8�xŏ0ADMn��M3����M��'���U4.��q�a�?~��#\�29jQ��8�5/~�h����O ʓ�h���JС{4P��í1�li��ʦ�:$)/��?&?M����c�䐨b��`��B@�!S��?FJ�V�z�r�	P}�O����'b��J"�i��h\S��OM�HIulj���5d�DJ�y�Ԣ=�'�?�#�ی08!�HA�(b$!1���<�)Ol�O�m�E�c�hs��'�06�'����ް�?�L>�'Y�tyشD%��5O �l���,�i�pq��Ԉ!�|��?�5�ܔmi�����l~��O����б�fa�I>k_�@
�$D�{H� �"�9Ӆ~y�^���)��<)�#�=�գ��ϼ?\ɛT�X�<��i�2���O@n�@��|2��@,@�����fEO��3gOJ�<��i��6��OH�Q�!t�:�ퟄ2G͝'XsW%ֿ7��!�Rn��(Z	�盬B
�'����$�'���'�R�'x��t�F���u�
�zn�i��T�2ܴsV �ϓ�?Y���䧣y���?B%���&��9Y_�!�1@����M�g�i!��D(������)��X�2(U(�*��@`��d�߀z�2˓FĄ����u�
<�Ŀ<Ѣ���Ja�pS#
>.�Np��ې�?���?����?�'����e��h���Ǻ��U�Ѐ�A�c��pSش���|:�P��4w���j�dt�!����&��4&\Vz�9kf�ԑ\B�7�v����+g���E�`y4��'��$�k�!��e��ux�!���
b,�0Pnx����\y�T�"~���N�R�{�	s�#��p�j��F�M0��DE��U'�0��S�8�$��!�5�<���C�<��O��mZ�M��SG��+�4�y��'&�ᘴΖ6_�Z(��V�B"hDp�-�z�����l�v�^Ќ#>�㢔�h��8��K_4p����z�<aV�ʠW@���?j`=���f��Re��4�
1�C�קi	&��6k�&[
v��(�/H&�:��D�r����a��3]�|�E�L-Xd`�,Z� ��bgx2#�-p`Qh���5��ƦA;t<� �@��8r���EI�,���H�-C��� _x4 $C�(���H�c�vq������)�Iן��I�?�Hքǯz��U1Õ?z��QK�'C�ē�?���jq��A���?�����IW�S��<��NG6g�d�`q	�3��n����"mc�4�?Q���?q����)� Z<�w��E�x-�2�F7��='�i���'�*hr��'���'���	U/�(�p�Cb�**U�ע���l�ao�Ǧ�	�<�I�?��H<a�j�D�:�ȖJ������I����i��l���'�"�'�b?A�	�c�!ݙ��<�T[=J`�}��킢�MK��?������c�xB�'B"�O��9`�J�/�؄2�g��=[�Kc�i��'����BqL�'�?�T`A�a� �k 5O��q���� � 0 ��{���"O<���☶V��ƉNIv�Щ��'��y�S�=|8����e�*P���,�J��PF�\q<�0*?�88+. ILШܸ�z�b!fmq�cc�� �2ع�(Y2,/�@@�lQ�WD�i���śSv.��0�	�n嚄���Y�e@���0 ��|_�U��O��|*�,��$A=�`AR�� q�na+KFe��'/BFڛ���'���FL=iC�E�Y*���5��D�)�	E$����8N�T��㉰p��ĐQ��"Z���[�'�y1ƢNt`Ҁ���f8|�Ǔ;H�Y�	ٟp��ğ(ըT�b�st�X�(1J���Cy�'V�O>i�Bg�O'"�"LڬC�D�u�1��i�4KV�![!'g��$	�B�������)c�6�n�p�IZ���#:��腚XR�a�t�˄U\��<4�"�'�<�!����Q��AqΉl\a��~�.����dBD�"<�!%�Y2
�����>Ɂ��+Qb�*�+N��0qݴx�B�L�S#�Ep�i��^<�4���5h�h���V"WKݥO�ـ��'�R������f�4f\٘a��:����#E��'��'����՚Ψ�B�с2���F�i>͸��䌙1vf���A�7Wܒq�f/�7��m쟼����d�2��2-����ş��Iҟ�cre@`Qbg�	�ԧe岄3�6$�����\r =xUCV�'h��kl$̓�)�?h�֕��	�+8�Ҵr�@��L��ʥlP�X���.	{�'i���5YN�+���2i�
��Wز�#��iK7�O���a,�Oq���ݟ\�R B�>,A�	6'�x�{�)�h<y��X�7,��'��'%�мj�H�L~B�)ғ��I�<� ��%����fO����
��w�Z�I��@��ϟt�	�T�_w�"�'����?_�QB�ǜ/�x����H<V��F���G�щ1G	<EV�l��I�I�D� #��J���� �Zqv�Z��	��F���o}��b�۷��qE{�eB�V�2�h�U qG�L�#�.~�Z��I!���h�(�$�<1���'�
f�͹f���c�a�� ��`���S�-�Ɋ�?����靸SpL\�<����8�?�-O2ԡ7k�ۺk���?IH1��	��МVp���!���?��M4��Y���?I�O���'eY6v� �gW�"�6���'����U�S�G�pቲ ��p<!�Hڬ|�����GV����޴�$$h6�#2������8M�ч�I8����˦m�	�б�t��*�B�4MA����d�Ɵ��ퟠ�Iɟ�$?'���S�O&3��8��Z3MR�1��;� �4G�1��CSOK"�s�BE7b���Γ���Ūd��5nɟ<�	h��لY/� �g���cG޾jLph�v�^/$�'f|y���RFj=+�F�<�Of���,�P�I�r��fF��f�'��`S�n����OY�OA���� 2<l��reM#27�M�I�,{���O6toZ���'��'�"5b"�V�j+20h����x�<�����<�4�WX@(�IS�H?@:��@�^�<�����$Q赂 E��(��Q���Zx�HnZ����ʟ�14�ɺ+���	ß��	ޟ�1@|��T�O�8���	/�<"�"X�b���Č�6�ZX�Q�|��ҮT6B�`.�Ld���N���Ic���<! �L�e8�>�O�$iV<�����ȝ?VԵ p�RЦ1�/O�������?����?!�mH�p�S��!6��59��(��x�� �Jc�!�c�";f�q�A�����K�'h�Vy"�ēN���m��
�,�..d���';J�I����?����?!����O8�S���HC��1rQN�K *�[��� )G�h�jDc�b��H(N�(m �`�-��1Ep2ӠΛ�>2�L�RdW���=��	8_���pJ��w����`%�Z5���� �MSs�xB�'�b�d�%2�h�A	�<dC�͛�e|�!���/��i��0I�R�����o�1O�'*�'� ��i�%fR���QQG�,6�R�"O
EAd*�(^<���^�u�R	V"O:1ł�{�~0!�k�#�R���"O
 ��˅0���ieŜ�u�~Ig"O,�Z$��4Ĥ�+��ڶ`���"O8 ��K��9�>�行Q��*'"Om�f&Cd��i�֫�K��K�"O��I��[�;���0��)&Vx�f"O |�`����R��� fМ��1D�� �9;A$CJP���cԭtvX4��"O Pcȉ:&��3#�4Nd̀�f"O�|AU��	{����McPL{e"O�����~q��B!r¸4C"O�hiGf��6B}�%F�*�@-��"O@�ʇD�?)iP����.�$��"O0=���f�0�B��W$4@���"O� Y$ЊhK��rE ��KV�s"O|�P��I�dE�Zc!EJD�T"OX,��%KR�P�RG��UѬ=��"O
Q�R�ң=B��6
7l�d�#"O$��@��6�m1�/�(/�5iR"O��)2��3G��4"�k��@RTI$"O�p����0�dmbQkH;8pc"O��YF,ݗp���EO�b>x!"OF��	��$��<��B-���'"O��r�$E���;7��t���ht"On��a`J/ .�X�MB2�i�"On�;Pj�%_��дO�)�1"O��Pt��A�Z@��D�Z򚝛 "O�t��FA�4��|Ȕ�O�	y�\��"Of��#��
תP�ٿqK��"O�a"�&W9>��4�d�"u����V"O�ՊE�V!{
���l�M;n�;C"O&8��H�\�� m�p#V��!"O����Q�!��q�NԒ1����G"O:i�p%I<u*X�s���4�pL����Oג�Q�v�l]B�K���öN��YF�aS��D8�M��[�����w7�$Y�����a���:����N����l�N{�e���+�P�*�G���\"=Y�
H�}t���d���(T����l}�$����	��7z�� ���O�)BT�_��py��.2�����']v���#�t?"��]�0N�Ej�47�z%ن���I��m��F~R�] }nD(6k_�Q���	��L��~"�P�{���d]'��E+�&��hO&��7��>z��ə7)H�K8y��d�8?s����6r�n�����R��9j�O�5Rvi!��֫]�-��IV�Hۙw��a��
q�R5I�O��ż-
�{"�Y�"^�2��3^PT�y�R>˓m�����9���T�I�;.��Gz����ie��<Kl	��,�=��ć�P򶼛�Nq���x��1|`��8X���"x�f'��mo���M͌y���*Xw�|�و��K��A/��RV�0d<����?i�=�g��5Jj����Ѹ'=�!B;Ob�rA\F�\���Q��ð Fɟ�b0)�N�����L�b�rE,�~"h%���I���Kr��R�T,�#�FI~qO�Q�#����~rrO���ed��~Q��$O�gw�IiQ��p<q�/���О46��5!R�2�vo�1d��c([��WP~��tI�ъ#�L�)��	5OJ>g�4L(���O�'v~œV.ϴ�#-���&ҩO��r#*�9��$��L�F���Z���Vf�r?Q��D$`*�r��-=F��Ţ�Ob����:{"��ADӰoT�1�i<b4[cG�w��i�e��c�F�ڍ��+,X��*M�[5�����3�ڰ�	8��seڱ�F�5�p�f�j�cދ6�`6)��y�4�eV�&�џ��s�	�1g&!�@T
F�Գ2߹FY�6��D�H�<gd�m|�y�B�ܔ5E��5�ug�x`��(��Z?9N����!9�i�3Y<0P'�(� ��w�H`Pp����ݐl���d�(����C,h���Z�c��14� �Z1/��Q-�$1}��'#B�F�@��3�.	$����0�U��?a3
�0뢴��aݟ>�ɢ6���A�nM�v8<��׏FT&p��n:�?;��R�Nă8��@�P�
�����'mD=����H����%�*;��P��$�:bh���ۚ8^PJ�ᑴT�!��[q�'��$3?A�j�/�8��0r`��K�+T�&����C���<I%���(V�أRn��fd�%xZ<d�T�1�^���'����i��WJ���D�z��A��)�N��<s��HO\AA*^�w�H萀R�8��X����A"jg�	yůĔR
�|��#�O%�'%R�'��6�ʹ.�^�)5��"y���Ja�'n0*e��j=�H�e,Vo:��s�4��SR�W8	6����Eײ3�&�F~��		�L��t
_�
�f�,�%DȜ���Y?�3KG� y. @��$�hO�8���SH$��K��R��Z��r螃{/>DG����h�xl���6���T�I�_�hȀB������B�f~h�%�� ��O�Rt�t��Q�3
I3��6�IW�$�@ ���� ��s�P�� �ƉD�lI$�鉶@�tѻS��''�P�@�J�d�8�V�2uG'o��܈B@Q����=!��?��*��{8x�q�V4B���@��lsP�Y�q\ތ!G�_����s�~ӊ0i3�ۻqd���d(O�V�����	�R�p��&�W	X�\I	�*2�P(��*bz�R��޵D��l7J�~�r��D�+,S��c�_�,���e�ưm��6MP_�')�� z"oR/��� M:�6���lw��L���5�p<I��$;<�����I�09r�C&�F?���=	�J�_�b傔���*�ȓ/��ɤQ�SR��s~	�#�
s��#=ipd�-��(��ѯy?�b�Y}2�F	]�h���^(+�U���9��On���V+,_���jL�z\�A4�'ԥ7!�<;r���D`��H`޴b&��cO��=(���<IL>�E~"A�,"TH�`�Ơ2����+�~�J�&��r��\-w0^@��Q6�hOQ�Vm�$G��Xu���)!�a�P� -U�L��	:i�����I�r��D�@Ǖ�_y���򤟋jd���	=�~��w�`����>���J���+5~E:��� �u�ޑY> @��ثHj^�HD�p� �=�pl�/H�t}�"��W��F+�T?16�
 J�[0��<�\I��#��'F&�REP�0�&�K�it|���'�!����/Gm>�ht�\'cbJ�A�Vΐ�`D\	��D�>����9<�"��l �!��]8�e׏�7�>MK&
L)(N�O�� W�37ax=
���5H7X���P�C!�Yh�'W��!�$J�p��P��"z�]�3Ѡxo�Eo�,���'q�#}�'�\|��b^��x�g�;%�|��'W�u*�F�F$%�s� _F� ޴� �
�����.��D�=8�\}p� ՆN��a)b
��a{�!@lŌA3˄���/�1-S
�
#�Z�&#T���=D���pK�m�̸���(+��yE�'��`�^P���	��>IP��<a}6���л��p�q-:D����'����v�Z5G{`P����;8;`q�4 �z�IW��~RM
�>Z�P�4$�a������y���-5��ɩ�É:��;��G�M��.�yv9S�j)|O����Ì�g�p�0V#ʕ^J��iW�'FjE��Cٴrm
l�ɿliJ$�C'|?�8�Eb�7 C䉡P���Z4�J�aV� ���Ӱh[�т_���~�H"/���c��f��l���̫XP�%��%���<�	ٹ1��ͅ|�F�RB�-Z�jG�1�~�$S�w��D&7;:.��CO)l�P-���Yd�'O"P ��=]�y٥�5(�p�O�$�'рw��RR L/+��ݪ2�IK�zS`�	e����6�͍jӆ��{i� V���)���6#ћf'!SD�8�E��%�� �b,J%��O�c�/�%g���ta�7�>�O,8�1���K���c�i� h�Ȱ��	 $�*A��h��kϩX�r @���0��?	�`D+�Pa���x#����0�F���0�p<�e��6n"�?-HB��C��1h�Z@����`�~b)H%L|�!s��!p��)F:z��R k�'yX�bA�P�����]��A+�O���/�?~���P1G##hԘ���0>~���*U�T0 4�V�I�����m(j��*D�t `"�ݨT���U�B4PD!���.D�D���F��O�t+e�Őn� �)A�Ńqt��hqbK�6Z�RR�R�Z��_�V����5�1����m��	���m�9%3$]gCa\џDP�>�]].|9X�c^/8{>�sph�$7�����ʇ�U����Ɂm��X�w�
U����X���7����}B�=}��_?���7y�P(P�Z�:��B�?֖��aJ�q��#=QG+mX �Bg)�?+K��2!e�؟�l�69Ԫ� d��T�HuYA	fꞢ>�G��, �j�Cq�D�E��b��֟��sIW��ީp �=MV�p1�z�.���)�U�aҧ�يW�Xa��	�����)��yw(]��ϟTY�����̹G�x�Ǧ�9�aQ�'�j�+EO�e����۶���;Q������D(�j �N[Q���IC�V)ā�]q����
Ǔt��-c�:� }���.=WX�+VbX(:��Tʷ�'���I�< |���B�4q6|��D��Q�"9�Í�(�C�W�x�>�R&A�ȟ��ζ>	�DU�H�������X	j��� ���R�d�ڟ�Q3��/M��Ш�� �o���Q*��OFԜ뗨��M��%�Jd������?�(`}R&��/�T�蓠�>� �^
M��A�DN�I�`��Z?�Q�rj�Lp@�Xp�a�v'�F�''�@����uZ��U9K��=�w��m,�I�E�ܕ��IճZ��S�l<�a��[{��F.�>}����b�S8v`!�	Ǔ${�Px�>ﬅIT'g��+�
��JK�@���'K!�����Ā������?af動p	���hҖ�¬�&�?Y�dx�%ғH��`0aۯ,�VP͏� �2=���� R̛d,=5P��r���0,�tດ(ͬi�2�R�}�Ɍ)2�P�H�	�@�	��D �vb`D 0�Q?-�u��OJ/��F�H��8�c��.U�H�䭍 �~2�I{�t��CR7�~ҋW7��s���$S��L�'HǛ�xt�u�LW��L0��'t�[��Owў��ֆ"��U"�G�Jl���Ҫ9�`l*�Q%b������j���O뎀�����8C^�%hQ�-ȋ ��Ǒ��tY�� O��8&@���5`�#���#�%ځw :�
�)yC6<�#���y�K�3�p��'	����!�Ψ�qFƠm���ÓJ�rt��KF�!#<����I�>g���Y�
�:p�!+ްQ���q�ȯp��đ�[M��q���HD0�(���+N	���@���ɓ9�q���Y�����VE��d@�np XPI���iHf��;&��E.D�*(���MI,�r��ԠJ]��C���I�z�Ж�
?���D�x�:����ۻMR����b�!d��	=M^�l�6��V� q��֣= �� _�Z8#��H�|J��WA�	򡤅#RZ^@��÷$������|�G�z��=A7J5���;z%��3�p<A`(\l��đR���c���Is��L��(7?�~RH#�es���'L��0u�Āx{dip`-B-b̑��9?f�Fz2G�}249���V��I�u��?�?�%G�#GvY8�CL�tGn�q�7F��=s�e��S~D�HM>q�m���D�Jq�?a�qa���ӟ<Zq�Él�n ���<Z�Y��nӮq:��- P���CKۃp���{��'@� R�4=	�X�ړ+C0�tA�Vģ"j �x�̽�غ��z�SHգ$n�ˑ)(ړQ7�q�-�>�X���"��<q+�.X�]]nY!��ţ��)�Ӂ��D:���_&�Hb#Ҕ��aX�����)��IQ�wTy�n�*|���c�H�)yҔq���IE�I�8xF�$I'�U{"��E3��ܳe�Y��刂�hO�I�Af��E<���dW�>֢h;��O���ł��L���^
S��Z�_�h�>�Rh�7kV0q(V�:�L�a��<�R6.`�FE*y,�h�j�<qW��<�\h�,�
ɚ����Nl�<A�kݯj
�se5��4��h�l�<��EˑoC,�rXMe~Y����@�<a��S�'�(�QB�5N�#gEe�<�7�͎���a&E%�N�  �Ja�<��E!*�Nu�E/ƘS:P8��TV�<х,Z�pQ��ϐ[�r�����S�<Iӈ8D��Ke�
%� �+CP�<��GS�y��c#��@!���5(�H�<��C�,v@�0`�S�yX�:��G�<yS�U)�S��ǂ:�ҕ�D�<��,C%'Ԡ���u�x���U�<�w�Y# �RtjE;S1�%� l�S�<i�GK7��YPj_6gu��AdeQ�<�6��1���AB[3c�&T鵮HG�<9��N�`y�wL�2��TD�<1r��%���e/[�0q8|���P�<ٶn
	�쫑��.W����t�<��Ȟm��!t��n{�����L�<�3g[1'�6��_�A�0P��̜F�<���� �0-*�^8�h#HE�<	�O��8T�L�P�:�@�[�<QB̝:�Ƚ�6�Q�U�( �E!Hn�<q3c��!�b͊�d�.4\f�i�_h�<�PJB�y��@��T�	2��6��c�<	4W��Y�P�/IQ�y1Vdc�<��Z��K�4� �*�
���B�Ʌ+�����
�����ͬ�B䉼*��E��`֜E!����1�B䉴D�h�����6��P�Q(�vq�B��;nd̑�)��v䊌Kb$�:)�B��3X�+pG�!�h(k�A�E^�B�I*)H��?lfXt��fT�(z*C�)k��k6��>�4R��ųq�
C�	:^L�T�5#�j�@a �B6m6�B��=����/YJM�FCF'��B�	6A�<�s�j��D�����V��B�I9?�U��ځ
������=|�B�5w{�y@�+� ��Xak��C�ɴ+�v�
u/x;85�'�W"C�I�(�#��A{,��$,C �B�)� ����F.٢��Rh޳�.L�W"O\<!��35��6�Y��N��"O�Ŏ��;P6]i���4�d�"O�@�=�f�����Gϲ��"O�1E�ޘw�H���d��h��"O��ّ��\`v�3r��hu�c"OTU)�̂�&Ѩ`��.\1Y�M#@"O�@y��T$p�b<���1��P"Ox�8�*P�h��.S�/� ��"On���@������U?A�A0%"O���	1�h�'+��3����"O>$`dn���x��	���)q"O4yy�����rb����q"O%@u�ݰt�)�1�Q�n���["O�Q0Ɣ�~��"T�D@�n� �"O��ї�]�hd�}�� :���k�"O�Lr��}�ru��h�Pk����"O�T �0���"H�Q ��"Oܑ{�"�!-J�l�&!�P`�"O���#!L!@��p��kQ�J��b&"O�P��G�逷�צ0��I�"O�H��/ڑnb�� X�g�6�8V"O��eM�f@���CL�$"�N��"O����g߅C��h�c�ݖ5����a"O~DrI��g \�M.c�16"O��b�$_'2ܬe��&E+.�,���"OKB�k}F�h���:�R�ܫ�y¥ �|:��Ђ.h s� G<�y⁎�M=�X�1��l��ٲfֵ�yr@D;@�Y����dTE�5�V��y�e�>]��%��)�Z�D�AD��yM�<G 0sI�G_,��2�S��y�|�h(���
o�&QHs��y2/�� ��9qeJ_ 7��uPr'�;�y�ZG}�]�dc�1_��Q/���yR�+и�D��/CZ� ¬B&��<�����D�q�T�%A]đ�6�A�7)!���Uw8���ۑ*S0 0��ؚk!�$��q�(!��A.iݘ����D�/!��V5JWn�0�mQ�Ä4��n	� �!�h|D�xqh��l��kN�f�!�d5�9�d �%()�h����5�!�ĝ?���j��Q�3k2�ƨ�wh!���x���U�N7^E�pYq��N!�D66*�p�.N�e@0����{%!���Z)j�M؆[?l)���0!���k�ތ
�@��A/�	J�L�G�!� �5r@��L��pz��	^�!��Ю|����N�q�lHS�đY�!�3$`�0C
F�)�F���-M�}?!��pn���
ө�b����y*!�DF$���8A�� &��QB�lZ�z!�Y!(��S��(X�Z�ac�(;s!�d�;}"��C"�:V�츻�Ȫ1e!���@�ЈQ�խr�1�BIT�WZ!�X�#
v	h!'�9٬l�&��~�!��xv�k @K�gp�\���Y��!����8��,�&X�%1SI�I�!�D
`��+�oM! �%�e��K�!�d�D�x��cA�>4P�D��i!�ė*j�L�
��H����՝Od!�D�C������o���;R)�ub!��<�,�3$f�'�R��?-�!���&�Ċ�#�L�����6{���)�'�� ����C��1�a�e]�PQ"OZ�	�f��w�ȅ���	e\XmZU"O�D[�G-픬��#Y9%�Vu�"OX�����lⲽ���L u�K�"O`�NǒT�B�@��)T��A"O���r���.�hr��" R.��"O��2���)�@kńhAt=k"O��#����~�`����A9�"OH��W�0Y/,E���2�4�k"O�L;Ӣ�%zR(�@�j�n���"O��&�ϋ*���Q��&U���c"O�d�3,ږI� �:0��;bG��ȁ"O��̆'���A�-'Bn�{g"O,}�E�]�:0��Y	4%n*"O��8�!�lޔ�����bf,H0"O�I�ӵ�y�+Q>N��k�"OF��  �8C�tȤkΥ3ۚq*"O�<*���R�����i�'{s�sB"O�#���n�&%C��M�3���h�"O�����R�j9��
���*�z@0�"Oxi���Lr~H�'ǈR���[g"Ol�s�'U�V(;�kΩ&P�̪�"OP)Y��#��"������:d"O�{6��,3�l��nA�q�=��"O`�B2��g�m�f4Hw�,  "O��@r�15<��rOP�t�ʄ�E"O��+W�X"V>�$r%�
[L�8��"Oll(6LW(*l�4��SW�3&"O���v���6*�˰��"uMth2"O���4oȕx��·���J#"O�aB�K�)lN��&��0R�"O�H���[�G����c�Ԩ6-�`JW"O�թ�ƻ;�����c���s�"O��4AZ�L�ܲF�
-9^9v"Ot�����>A�sB��<�`u�f�'�'@�Ϩ��H��F���~��'	䱹���&grlр� S�	D�É��+�S�d!�eh�I�`��x><9�;�y��߆G�|� 1杍s�t�WA�y���"n�\��:p���$A���yB�ݨ�*E[AǕpP����'�ўb>��ŷ/M�`Gǆ<����?D��;��
����2Ԛ���������91�>9�
ŴH���s`�AҠC�	�&bD	s���*a�i(N��^!�B䉲9��2e��S�<���Iæ"<����?� A$X�l��))�C�1|�bHa�)D�����,u�\�y���.�
�;DC%D���֝�����W&a7*�kE+$D�T�H�1V\�	B����Qak!D�\�ȇ��>ᡃn�L9օ�`*D����&ЂTؘ�H��J�kq�$D����KV*����KjϞ���!D�p��یN�L%�DJ-3�v|�q*D��	�!>f<��J�JxIJ'D��+q�D(A
,� D�H���C0D���ȉ:OD6EƋY��D��1D���u�W��*IuZ�$�z'g.D��)��ЈlT��W�T�(��F+D���`n�Wl����C�~�И��)D��3U��
�/J�V�|��D@�S4!��}\��	K�N�N�d�ؤG#!���C�]"� m[�a£ε~��S���V��Rl���X�J\!_8�xw"O� �@a��´3c�س��s���{�"Ov'D˙nWڠAI��l���Bg"O������.�p� ɑ��L$x6"O��(�c�$X-��)��y�E��"O��0��
}@����ґ!��e�"O�H�*�6%Z<IDAK^�""O��+�ʂ�!,|-X¦ł^dҕ"O�[�RF8̢���
�б�"O���R�]�3�蠢6d��;��Q��"O ����\��i(��2DƦ��"O*QyRlL�2����QBG]�0���"O���Ԩ@.k���:!��hG$�"O���g��y�x��.1A�H��"O� ����P� ����R�d�̺r"O���tM�b̒4��C
��"Ot���b��R��5��N�#�܉��"OLER7 ¿d4��@u�ڙL�fU�"O��Z�_2g�l$�ǎ�=v�P5Q"OFQ`�kʽs�4�2ǎ�{�`�K�"O�DiumI7@�ʝr��q�-� "O�,(�ɀ
n�N0�W�����Z�"O�1r��,��	 '	�u�Ԍ��"O���8�����E#u����"O�d�I��`sT����H��"O8�{�Oٌ�:DYS%KP��P�b"OV��D��HC�<���\y��H��"O��QB(�:��8�P�I4�u��'��<�ȓ�L�<8�"%[���	�'���H�*��*Ix�M$x��$P
�';� ���&�`���E'#f��	�'���6H�������2�F�R�'� `�ĥѹ
�.qX4��d̫�'ό\ ��71X�D-P��<��'���3�W�'��2ɟY�Z���'Ǭ�����2�Vt�b�!���j�'ʼ�����ѹanߜP��a�'�^�եZ�^��P��ɀRV�B�'���9�.�H�d�1 <#��
�'��!�Ձ�w��؉`ķ39*T��'����-��$֚�R�C_)�̐�'$����\%� �g��"�����'�X� � �RԔ[b�H:�x��'5�Y2��@��)*������
�'8�3B�� f�����\�8 ĨA�'|ެ8㉙>{�2A+g�F�.}�'�: �c�_�d����F��!�I�'C���R�2[0�uVL�H�ZR
�'�B�0% � /<��S�-H�ܤ@	�'�<HE�I9iZ�Ф��"�48)	�'�:@2b��1R��d@$���z�'�J����B�"GrAc�
1����	�'���K�� +�t}x��`�䔋�'EN$��nV�_��q�I�(BP���'dS-������C"� �X�<�T���J���͎�\��8�5jLp�<�E�S�,`�E!�9�N"���q�<�@`L�Oތ�V�۽Y��u	T��o�<	u�y�܅�B��I��+��T�<�)G�y�f��$
�)���KG*]O�<�S�ژG}�1���mh@1"���<�S�]��,l�e$�K�hAc��{�<q��°JQ��Al@-,����gHw�<)�ʺlw��1c�:r<��H�W�<Y��,o!d��3�ˇf��%��W�<� �Y��`��|F���kN9|��Y�"O4���&��1���JC�Ұ\�&u�s"O�y�ׁ*3D�i!��[��첅"O6�{��@9��L���tr��y�
R�p�He�g �ⲩ�#�y�#ߕIj` C35�ٰ`
��y��T�3�^T���+fm`�'�C��y2�A�Z�~��cD�j����f�%�y�AA�.��9W���XTz�h��$�y��AMqΠj3�H���F,J&�yb
۹y�Ƭ2��Ա*��8�hD�y�lq� `�[ ��ܪ3b?�y��h�x�`I��,�l!�DS�y�%Z�'�r4�癑|����y��V,u�L؀���tr����C��y���/-��Yz7�T*��B
[�i�'�ޔ��I�8bf9#�(S�P����
�'\ i��۟hh�T(�J�[����	�'`̥Ck%l��I��ѺD^��	�'�\tz'�G�i09/
-b�'(d�2�U,!���Z��+n�y�
�'��%H�ۦ�j!'*�)8pl�
�'G�W�X�y*6��� 5���
�'�H9���
`ȑ3s�ʒ�V���'%��I���2T�T�qRȑ�k\�+�'u�E*#	���9��U�~TH�'.DY���z; ���+ediy	�'G\�b'�&x��	�ׯ�4�`8��'�n��L�~�x��K
.9ΐ�
�'q܄B�^�ZҤ�HF
;�v ��'`H�9a
�>@]�0A@f��2�'Bp0�eJݼ6D�փV�qی�R�'�I2"��g�d��꒫m���'�H����V���4�ކN<�r�'����G���A���4\0x	�'����UM� 9
�+��8��h��'iܕ�@�	6����H�� ��'z�M�Gi۱sd�`G��-��'/(�f߱Cq�:�KOpq��'�셺��Qu}DX�����}�8��'�bt�MA���i���(t�b�j�';te�Mg؜ Zj��8�'���*��U�|����O>[=tIy�'��5*� 
��4}A�O�
<X���':�|�L����Q�z�V�K
�'
t�:D8,1$d:@�A�D�
�'���D
<,�z���1e���k
�'_(4����{��h����4^�h
�'e�(��*3h2����0g��0��'���-Ŗ-��Y��'M̜�)�'�P�hDIA��4�arJ�(V�l��
�'�E��,��@��I��a@�I����	�'������Po
24l��X� 
�'%l�˄�ɚa�lUb)��F\�qh	�':��N!s�J���)�P�y	�'��\c�GC�0݉��L� ڸ�j	�'�J��G� �4u��*��x�@�'���1A�,)�b����P���'`��[�Na�"��!��%4����'_p�3l#*��c�LŇ}�XP	�'|�����[�n��qZ�FIsX��'�������*��A�DD�g��u�
�'�i$��$�uP���IP�`j�'a�Y��4�$a�n�*C�z��� �M� ��4Ftr����lp	�q"O&� ᦁ*/T$�9焁 O�ma�"O�@��N��"�I"���+�Z�x "O����H��v�"H[$H��/�*�X�"OdY�Ӡ"VX��g��M9!"O�L��.D�yl<sC��/c���jV"O���iɣ
����bEH�'���s@"O�"��LDh�ǁ �?����$"O~��$�K�k�Ƚ9����hc�I#"O����n�2���#�/����"O���-_�ʈa���-�V�@q"O4IH!�mBZ�0����t�I�"O>x����#gb��0bg�27�N=��"O��a�4�Z�����Sn���W"Oֹ��J $w9���rc�! ���"O�X���e92M�=r�P�
"O�|�VcB���5) 3��W"O�xjg�Hk��a�'ύ8ݔXȓ"O�<{���N�<QQ.M5fz���"O����g�k^u�p�χ|��"O�P������sj܍y��P��"OH}Gh��h�����f��pv"O �Z�M)y��LJc���'�Q�"OzpH2L�UI:h�f!Z�'�:L��"O�1#)�&Sr�hs�/I�m��`�"OL�눈+n�L�/L8��᫰"O�pS��(#�r�`��I�m}�M��"O%a�k^ļ�s�C�Sg��s"O�P	߯r�� t�M�m�f]�4"O��h5#�=b��ҁR�U���y�"O�L���ūcbla�q�
x�^�"O��
E+�-�2@B�c�a��A:�"O6p3DLdQ�E3�bM���5�"O`�)�iY2Ya��/%s�4��"OV9K#O�Er��z�G�R���`"O����ĄGi��E�;{F�(""O����q�J!�1�4ڀ��"OfH��Ā���Ă���>'��y@"O�<[��)Y.$�� F�����"O�A�vƈ&b����d�QsC2-z$"Oh����~���B��ղG�P�"O
������5��Z#�Y�"O�|뵄F���L�L(i�piz�"O8U�bU3�x�0��,=�|��p"OB��K�z��-� 3E�2Ib"OT��Dc�%7Yd!b���L�L�r"O	��	܇"��u@��G�'�fA`G"O�J�n�9#��U -�~��*�"Or`����������"s��ڧ"O�q�l�./P�y�F��	7N�;�"O���	ߙ ��$���2UNa�"O����ð;���@פ�"d9�`@"O(�xP$�%PD��`���Y�"O��1�D�$Ģ����h��!�"O����!���cT��Z�ӣ"Ol푴�Q�.�Ȃ/��h���q"O�1�V�J2��B!Y'�z9�"O�qK\�*����ت7�
�"O�-+�Su��S�'FO��9�d"OT�;�l=\�ݐci|?�4s"O�=���q=�����iO���"O���BI��
���\(e��s"O��)�%R�I*z��2���TH9�"O^�S5/�}��a��՚/��ŉ`"O� ��+�zv�a0�8C�����"O�����-E��� �R;FȈ��"O�!yԌ@�L` laIP�3�� Bd"O4Aq�Cb5H�{s�2�$���"OvՈrm�I�:u�2'!�N��"O��@ �$�Vm�����=�н��"O��$�WR}2�1
 :��I�"O.��@cfd����C@�t�#b"O�5�_�sG���nZ�j9Vp�"O�4�6��y*8�'�'42Z�Q�"O�@�䅥D]2�����x� �"Oz����<��L�o��H��"O�px�,�ES��  �q�D�hA"O�Y@V͋.d'،Y�A�x��4!�"O�Ւ0*�
�AxІ�-6H\�T"O�8�!Ú>Z��9�@�C�ȹ�"O�,y��F=h�6$eF�.O�����"O��CFI�)8}с�	�H0r!"O���c%��M����I��t0�B"O5(��Q�F�TU�deAw61Z6"O��3�ÿh�|١�_�c�l�@f"O��8�b&�����T1F���"O` �2f�++��(�O U+: ��"O�-xv  Rpr"GL9)"��	1"OF���j�~��w%��:w"O$ �ÔZt�Y�q�ҿC�`��"O�����[:?�p8�-@p-P��G"OhAbF�4pd� �ؼ/q^�"O<aj�	I�*mQQ�+VX""O��9G�߸7� TO3(�x:�"O���宅�|"��`�#�1`�P�W"Oʐ����~��ܛ���q�q�5"O�,�T'H�<�	VZ��L!g"O|U�ӨPR�a(��U��Y��"O����)m���g'J�0Ԛ�ʳ"O�-K�V�Z94�S'�M#9���"O��I�ǁ^�)R�F ,��A��"O�(L��Y85P�Uج�A�"O ����T(��j�O� ��rQ"Opr@�W�"�E�%0'<��"O����(-��D�:*,�"O��!U�N�J��Yx�*D�0�MrC"O�4�"�V2M%Di��Y,:(�"Oʍs �ƨ<Kv<p�E��M�X�&"O|���*%-� mæ� �4T[�"O�\
��S'T�B���Kz{�� "O�E�d���1��0�� 	�~4�"Op�+��D xŐ 
��E a��"O��(�nϒVK�<����/�	��"O��Ae�-��!#�N?)*b���"O0�;�|rs�Ş](<D��"O�0����.
Iڜ#��=�6P!�"O�t��ы*3��p惍��>��"O0� 	��cZ�Y����' ��!"OԈ��n֜`z(�&���)�>��w"O��Q���CYV��A`ӛS�~5+W"O(�� D�8}b̽���s����"O����ǋ}���ሐ�R�<���"Ob��h6L���3V4��s"O�ع"jʠg�+s�ɛgl<<0W"O���@^'�� X���%`d�<*�"O�i0�*��	;�0��ς9K��"�"Od����A�0��zqD�
@-H��t"O4<�����0�8&�Kx�`g"O� )�m�).o�k���)b��J�"O8�𷮝�_�D����M?�����"O���2�� :�k��>0�;"OF}j�cQ�sƈ*U��.G(^p;V"O$��
_�D�,�i�	$XD)�"ObEHSB�X�tT��'��[ �Y�#"O&t`�!2s~�UDN��x�B"O��ۅʄ(|ؤ0�B��_�Br�"O8q�&@-\�����a�*�� "O�``Cadd���f+
'>ntm��"OX	#�`ɿ���K�+��bD�y�"OfX��CʕQf��b`؍07:���*O�g�G�a�p�@��|�HXr�'|L튣
�#$�jP2>�:u�
�'
�D��k�&l�Aq�H2^$ 
�'��8��IO*�Vp�C	�� w�4�	�'��UC��,�ZU�ah���1��'J�`�숺*5TeSV֦�L��'�$}C��ȃf�ұB��zUp���'醘k����q�)�AS1	�fD�'-��Yf	
�9 
U8���U�	��'"ΜYpѓN�nՈ��0y�4�
�'.���Q��/�\|��띌�d��	�'�D�3V�Z�Fb�Y3��R,�`xh�'t� Cƭ�����Wi����E`�'��ABo7&0z���>��D�'8�s`�G&"�%�c�ǘP(��'j.��j�G��]�"�V�cL��'�hU�%j��w������F�W͡�'0�T�'��F�F�cQ��KJ>!1�'�:�x�k��W��Xf
˱Aw��[�'��E�#NގD28�iE�#ha��k�'p��h�>Mt�bp��dx� �'	�У���Z�|$sǩ��S,�p
�'�|�Eœ:�"D�'�	�'L*5A��2��M3̈�J��8�'Y��/� &$���d��=pHMb
�'�̡���Jк�A�B�%f��ܢ	�'s�}��S(B�Y #� ]��m��'��s!��B�LE"c�C�ff��	�'pbA8�@M�o.~�9�A�\^���'˰��%�Q'S�>���A��lP0 ��'$D9����5mtl�P#�kW�-��'�.�b�
N2.����0L�a�8mc�'�����"��l��G?`��k
�'"Ľ1�÷<m� �d��7����'ulUa搔4Z�P+�j�J�M��'�Z0
���.�q;�D� 9PTi��'���8�l��E�� bD
ے*��T�'���c�
�� #�C�>lՊ���'c�E�B�%���Ѥ��']��a��'�H����U�D�D�ta
�j8]R�'^h�B�I�o@2x��̓�ey���'�>�k�`����Z����O_�5s�'F�hp	�oS`��g�?W�ػ�'�V��e��6�>\�D��.X����'��Q���#���p��Ę#bzE��'B�%b��۰S�fp�đ1�<��'���B'H�[n��hSf�ِ�'p��*w��Zv��H�[�wΈ���'PX���7*ΰ��R�O� �|	�'�d�pL
���X��,!,�����'$�aS�ܖ��$@B�r��,a�'dQIg��>`y`fˋ�b�	��� `����@������U,Dt �"O�pZ��Օ ���zЦJ:��9��"O��Aan�	, �2�A��FT�v"O��dLOb8E��W�0���P�"O�l�!dT�n�ЁE�N�Ns���"O��S"�ÂV�t��0�@M
f Z�"O�eS
붨贈ؙm�dU P"O������y�#�7�d�q7"O�ԡ5HW&aN!+��c��B�"OE �a�!/u�	��.F�<�"OA��ȏ5��9��[�M����3"O*c�
3X��O3W��,�v"ObP���Y W���b���g�N=�E"Or����`�x��W�A�ꍹ�"O:`���wM�����T�p8�hT"O�lI�T#8OĹ�,f\HKc"OR��a ٱ3���;B��uJQ��"O�%Z���{�h�!�~,��"O
(��.�h`��U"HZ�"O*9"&�7��G'��QMN=�ᢛx�<!d*�f���d 9eѲ���Vx�<1#�A_  �l�"AR��w�<ɕ��9=N���Z_*e�Ix�<Y�MM ��( cH�=`|��Iu�<�Ch��K� \����}�m���Cr�<�AW,nK��k�4��<�5�Yr�<�a��Ձv��:�������k�<��&����sk�m�İ�r�O�<�F�s6���E�ƪ�h�9�N�<�B���`��M@�"�xQ�TI�<ɵ�'_�5Q"Bd���V��G�<� ��:�"�P��+D���)@�j�<�M��oL�Pwc�)\�����a�c�<�B/@�II�	ᷧ���[4��d�<�C�Z_��;el�3w��}{���Y�<y�j�'��Բq�5Z ΀�ԧGU�<�e�_�<2
��7n�]����jT�<�s�P�x��������P��f�<I�gQ�,� �㕩]�d8��`�<1A��8[�1aH��q�4�c�O�\�<y`��4rr2]C�����6�SW�<�Q&�.Q�m�&�3S��h�&K�<���ϚkԽ�'LU�;p��[V'Vo�<Q����"%z'��(-#X�r��g�<�`�̻R�����/�$i��(!��O�<�f*�6�؃,�Sv,Ya�M�<I�=\�j!��`@�Ar	��bK�<1�ŕ�*��o�O�h�h�O�<���*<
xB�Tn�]0��G�<Q���h�؝��-�?�:y� ��\�<�1��� ���U�IDz��f��R�<q�eV��SDD?,Z%�vM�O�<�h�u1�m:2C�"?m���ɄH�<y�*I�
Z�5D�=�0U�	�H�<AF�ԚJ������?]�IQD�E�<i��D�d� ֫ё)��E��E�<��ET�%t��>d,9!!QC�<�v��xZE���!��K��v�<�
i��ipM�jV<ӵ�Qo�<�����l4ՎI�]&f�p��P�<��fL.�p��3�E�Z��Afn�V�<I�`Җ:T�1 �� 5�8���VQ�<	�E�:5ʜ@��Q��)ÎG�<�vi�;1���Ka�X��S�f�~�<� ts%I��&��uK���]��"O�,���4d-Q��Q�'��<��"O(�0�X�P^Ҹ�cU�G�<	�"O��#5�:Nl4S�Ĕx����1"Oέ�v�\B%B�hf��]��%"O�� K� �ա��D�~�p�"O�aFK�+EX]�nŠ�8�ZA"OpqBlM�x�0����ޖ9���Ӷ"O�qhe�C�6z�d��S��$t��"OTm.)[�t�8".Ʒ$U`�"O����`\�o��WLA�X�*�(�"O��W�6l�pmۢ(۟򪰰�"O��U�\,gE����T'n�P���"O��*�ɄP��6�E(�ΩA�"Oұh�%!�$3f�<�8�T"O$��)%`օ£���B�v"O45q0��2Ui�u�<���"OD�h�c[@TÆ�_<y��ݳ�"O�iKFʞ�"�H(
���q��S�"O`���ݺG�J���E�7<�����"OZ�k�����Y抎P�%�"OF�2���KԈ9jpÇ�N��)0"OD	��W>��z����[�b��e"O Y�cC�-w� 4҇�Vx�J0"OD�Y��K/J7HyD�쌤s�"OƵP���P��@SB�:�f��"O8�*P�`�w��18�Vi @"OƔ�	�W�|�a��=�Ѝi�"O|x�aͅ	�`53&�H?@�(�k�"O���c�� T�~][���>��Q�5"O�P�T�7&BȌ;i�c�RX*d"OY	�D0RM�aRfϬ/�X8�"OP��A�@i���A�o�\@U"O�]�XA��ӲK�9Wm�HB"OHE�FjT�N$¨ӢJG�&�B=�"O�$�!��u�.�;�ĺ݆Ts�"O��4`W�7?���>.��`�e"On]��ߠU���Ǡ�7�(���"O\J�oG�2���+��@;���Ȗ"O�)��k[G����A�(R��xʦ"O��y�ݙ@�ڤ���$Q`�"O$�x���`�9re�	f<� �"OD�� �*�p��U�JQW�d�"O�)�s+��&u�\3�!	�S9��"O25tL��Jb>К%�8�19"O
���h�s��R�a��$��"O0�[Ui[�[�D�J$/�)IIp� �"OBd3��Y�ceP���m̎>8��ұ"O� 4���$��`j� ҉�6"Of��g	��&i��R��%�$��"O�5�L�g�LN^Hy�"O�UsF!�7���c��-Dr8�"O����M֚.f�!��W�B1D<(�"Ol��C�) � Po�4&�"O��T
��l�R A��?T� "O�}�����W1���iM�m	��	#"O�� qA˃|z(����c�=��"O(5Z�i)X�B�˕JP��K�"O2L�V$�Q�X�h��O�'?Ƹ�"Op�Uc��]�4�`�ܱ�=I#"O�t:t�ߠ+��҆�Z
tB!�A"O�uY���@Y��E1gPr�a"OTA"���^�!t
[8;Jh��"O�yˁ-H��*�rj�.e�XP��"O� B��3%bl6-�rΘ��Z5�t"O��H�gҳ��b�Ƌ��α�"O�H�ukR4$t赓gf���٣%"O�m�ub��J 4aa�υ5�xq�"O�m�Q�y e�P�%D���9�"OT��C�"�p8���Vm��"O��B�'��>I	!��uG���a"OL<��jW9I�|��i	K.X(yb"O�y؁#�5G� ��&.\=��D"OFD�Q��V��y�$�>(>�E"O�E*��� c3��C�b�!�b���"O��鑈�� !8P�˜i��;$"O�P�A]�=�|њG�־|b	�1"O@�(�*ƚ!��ݱ�E�Y�i�"OH���Ơ<5����$bt�R"O�0�wH�%Y�����ȃ%#� S"O Ժqf�7o�Hy"���#@���"O,@��m���>�`늧{8�Xc"O ��c�	%3��Tˑ��31t!�"O=q�$�AK����"4��0@"O�D���B�3�dq!h�<T�U"O�Z���$fF�P�&5&d3�"Ol���[H��� s$���r"O$��kD�0ԸQ�C�-:1aC"O���)�9k���$MD�XP�"O0,��
�c�f���C�7"��9�"OVL0�.�NŖDD��-�52'"O�<E���&��rn�"l���"O�Ւeg	&V�>�+v(>ir��f"O� ���)'�{�8Y 
�� �.D�D�V��Qo��'�#��@�-D� ��g
=x�P�YT�޿FI�9PwF+D�\�͐Gw���Ff܎m�`h'D�p��j���E���YUYR����&D��(����4y^X��&�"C0bU!�o%D� �5�=��R�j��Q�#D�@��̖>��rv�="���!D��H�DS��<)��<J���s�!D��� l#���ٷk����:D���k�-6��R"kN:j�,t	w�,D�(�Ԃ�0h)��Q�K�j�p��+)D�����
�d��`�1�ɽ	��!�g�)D�8P!�3<H\<�ЯF�AF�iY&(5D����(*/�[v�I*Ulz���3D����	�a�ȥ�gJ�'�>=�"c7D� ��ḃHOF%3�č[�c�3D��Q�T0�=Q�hA/P
�s0�>D�|C �ݏn�f	B�)�2u;�\U�)D������,�΀K�zmր�")D�Tb�Eb|�#i{]��O'D�|� � �J�l[�
�)\/����J0D�|��*���8��BOJ�^��`��N/D��A7�H�?w|0�r%ʨO�� Pc�.D��j �_9�j�h�*ZIt�|�tA(D���ra�d��sCu��	��$D��Q��1 ��v�����''D�[L	=p2����/W<��RK?D�xI3�ȸa.Hq���[<��(!D����o�J�r��U�J��Ω:P�=D�ܘ���i[T����!|u���+ D��:q�	 $�z��T�D�B	��	?D��C�ǜ8�}S�(rĀɫ�"D�85 �;L���9��4
��Ѳk"D�<s$/R�e�؄f�XXO��Y��<D�� �! d��D	�ep���5���ٶ"O<<5��E?�e�0�ʯ�z�h5"O ��`.L3t(ꔮƇ��ᒗ"O�JkC�*3\��gA�V�)�"O*̳�hЦG�P(ї�D'��5��"O ��˲)K4��+i�!�f"OR�j�hI�T9Fى�$�D"��'"O�� �Ƒn��3&��g鼹�"O }�wH�!fO��!��Ƅ84�P�"Ol��(S����t��[4 �5�y�J\�:(�1"JӘ(��u��L���yběK�v���@1����)W��y����J�b�֑>����E��y���H��(�ecK��T��#㏓�yR*�?B�U.l�:A�ăyB�Z
�'z�KC	#sp(�S���;�a�	�'n�y�dF��Ȧ��F(�-:.2i�
�'�zD{a��5�|e`F���2E4	�	�'S����MB�
��� .|p	�'���i
&/�L����ԼI�ya
�'����e��Z�����4@�.a!
�'pZ̊��#@���s���>0�(
�'�V5�&��:ɡq�N �4�b
�'l�9`�H����a�*z�Ё	�'C���$�=�b8��n[� �h��'��!�Ƨغ8����كl�<���'�V'�K�|0e"�4b�1��'�� ��~=2��d�ߴ+����'^��A��,iڜ���R�lLk�'�b,���ʳ?�,ڕ�L�"�d��'�j�Y%Ãz��HvNc��	�'��X�C!�E��Y.˟%6\�
�'�>�S��O�k��r�Bj:��	�'[ �YF�X�NĘ#�P�a�11�'FH�J��	>�^���� <\�n|0�'�T��D���%��3l�p�Ҳ�}�<����|@:��&�
,R��@���{�<1щۜ;UР���0`ۨ�#Q`~�<��IR6SIh�+۱Y�H�#3a	D�<A��R�at��sCj���m�ύ~�<��D�*c�[�F�-"��d�P�<�tG�
�ld�����I*4Ȃl\I�<q���:�d���Z�`Z��b�E�<�ѭXCڄ4��NF�P|l낎�j�<Ӏ#,������+Nu�%Ӑ^g�<��H
d��Y���)CL���EY�<���	+T�b�1��N�7^�����J�<YTc̐.�� �9��BPF�M�<S�צ&k��Fl�K%pHACǇL�<y�G@�&��RoѤ@ʭ�cK�K�<	@��Y�$X4�["WD<����R�<��U71+\�14�H�O����u�<��_bC %�97�v� 0�0ړ�0<	���E�6��2�j�2A�p�<Y��.a=�}봢��w`�5��j�o�<13��$�"ȋ$��)�$�{U`�U�<YSCH�&��y��97v"A�ǥ�G�<��j�v�:L�4�V6b��-aQ�F�<	��B~r�Y�e�^0~p0��c�_D�<i` V/��!���ٲmp�4�Ney��)ʧE�:��'ID�Q��8�DL�8���},�KfA��"(�y�� ^숰��<�fT{C 3<��ћG��<>�����\P�*�:¢�_|t��#�"O� b��G�.�Z��¼�"O l;gLQ�g�޽F愁�P��"O�Pb0�ёn�f��c\� @4G"O:aSs�A�W�PH'�I�N:�A�b"On�h�D�<�Ƀ�!1}4ܓ�"O:�!F�R �B�� X�$'�x	v"O~1(�,խ2�� A"�[/6*���"O^��ԩ�y0�&J'[PԘ�"Olh��F�99�؀A�L�w� |�&"O�X�E��hFH��wn�7@�":�R� ��`�S�Ob���wFAa�G��@B����'N����%O;1�V�*5�#4-\�	�'��ujP����k��]�3o�9	�'���Q<v����Ô5)3(5k�'�u�`۸G�$zG�;U@���'��0��~���d[�h	�'����T9r��pA�cAC꒍��'�2L��#C�_��ͱ�S�<� DJ	�'ц|�E�u��L�� 8W6�#	�'��"6�-O�K�m��f�e��'���`G�;��hJ"A	z�٘�'��9�&꛻2���h�X�	��'m&�� BĿ���Jc��;�'�<@��L�N���I�&E�~i\��)O��$�<�K~�=97)��5�v�c ���$'y3t��V�<�Š:+�*xJ��Ȟl�gR�<����e�U0���QZ�pp��J�<�5i� �H�Ѳ"Y�a�jl(���J�<���D�b���YT&^�-6L�ca�P�<�� �F������;R�]���V�<!��E�; |�%�@�����}yB�)ʧ>����G !O��1&�*�N9��6窰���X?��sc� ����� kMФ�'/�V�x�ϙ�4h��ȓtP|�bQ[�4��HZ��׶D����ȓj ��2̸U�x{��ӛ1���ȓj�ܝ�5��		� s�/⸆�6lt�s��N�)�q�<I3*I�ȓ;��h�G,�$D�\�)�IQQ���ȓp��CG��Gm����;ZODɅ�*ci�DM�1��E�HιR�ʔ�ȓm��3�F� ' H����3r��T��c1bY�%�ËC�"u*嗰(��?a���~:��̭-���D�#'�",*#��uh<ɡ� \��b��O�@�4(�2Gܕ�ybH��f��32C,d���X�g9D��zfGL Tu���P�W�W�ĔK+8D��B�LB��O�?[�l1W�4D�Lyp�P��D�/��c�0j� 3D��Bdŋ�q��+u�Ђr�Fu)f�/D��i@�7B����')R�E92u
��.D����I?k�<�C�ѭD�(peb7D�(y�uL �ABP{��u�8D���㉐%�"9ꀫ5*5��#��;D��b^/)��c�/�
E~�Je�7D�,����?rjmȀc~dy�;D�%�
0��ղsi�*\Ұ�!�8D�h�Cϋ�D<|�b@
�,���k2l9D�`kGH�2 ��ہ'Y���R�;D��	T�)B�B�3�$VU\���E(6D����`��Xa��U=�DR��2D�<� ��D��`Z�ESb������*D�Ыc�Y��J�"	�R�й��K�<yƦ�W.�����8��A;ǩH�<� Zx��ݒPJ��'���:T
��G��h�� 9�S�O�Na �Z�]�$�R#��6ݰ�')jy�u�+\����cbK?�8eh�'&*1P�F�*q��yك�#"�,
�'N��ِ`å%�� ���B�����'6��p�%�(��F&�v�b
�'��| �,N�GThS/��u.���	�'t
Ĥ�/4���C�̲mr��I>i�����G��bc�
V5�@CB&M!�Ā�]�8��}hY��!�u!���~�d����� 4"�
!���L�LE4�����+!�DݮVb����*M'9�`0�2�H[�!�d/n_d���W�q�(�H �ȟL�!� �]2)��C�7"�|�ہ$N<l�!�dJ?D������ȵ0�)��!�$݂|�z��ƳT�R��,����'@b���R�	��zS��^U)�'�l�kva[(.(���� 
�����'��I�p�D�}��-�6�� �^���'��p��ߤd?��c��6a8�{�'��� �M3(�*(p6�H&`��'|���F(�%J�^����ȮZ7&�j�'Gb!2iY4�t���烓W�<8��'�
�$�)����u�C_h�Q��'�"(��aD�@y�M2�]@���'��Tɥ�P�YF�$C����O�A�'����2��=�@�ĊޏF����'�*Q�����`�{��Ê?Z�у�'�� IC�<I�|(��^`9b�b�'�rlS� �0	Cܖ_C��2�'zR}�eb��H^�`xe.�W~���'�̃�f{;tIPթ�K(j,9�'`�-�@e	�c��N�q��q2���"H�F��X���o^����[�<�EiP������Sќl{�J�U�<�@`ġ}F�@�Ǿ(�������v�<�F.�B�"���Gڐ�"�H�<�B�Q�-�ȡ"�U8Ѡ���\�<Ab��BQ�o]=��W�<A&��<Y����p�Љy�Dk�<Y�)��S�L��P	<|�]f�< �]%Z�D�zpˀ@�^�����b�<i�g�(Kbrp�R#ݍi�z� $-�Y�<�un�Kђ�!�F@dF��t�EV�<A��Ơ]��`#FU<9�z��E�~�<!s傟) �������1AB]|�<Q����b%X��dF�-�R���]�<)eFT.�89+�섲B �d��_Q�<�ċF�d�:��q�T�p"�5�`+AG�<y�C��Z�v܊�*�|DSP�Rn�<S��0�(I�*�_�ݮ�	�!򄔹*��S���
=�l��`�01Q!�D?�V�i��4�(X��+�!�d�D<Є�9A��%y�a�
t!���0i�s�"�0&� t1D�V/	U!��H���R�; |L�r�
 v!��ڂc�1�0`�2��ů�?:!�d��Dd�÷ �hy����v�!��L;z����ؔu<���K�2y�!�$�!=�P�+vi��M^���a���Y�!�D�Z�`��J�eS�@T �X!��.j�J쒔? E��٦�:!򄉲>�d4)g�$'��Yd���]�!�� b ���mo���17xh�"O*�J6��~��ـdVc���"O"��Bf�2l�i�M�7	MI "O��ҕ�Ҫ0_�,(�e��0Bt�ht"O<T	�A�A�^}�#oUk>�y"O^�3��W�a�\���� O	�!�"O�E�v割fD@Ō8p�<M�A"O,e�GZ\z a7?�Ju� "O��Y�KϾ;���J��V��@�4"O��b��ˉf��3��L����h"ObɱRg6~�~y�%^�+v�� �"OԽc�+�5C�d5�3Ɗ_WD�
u"O&5*q%���TM+FDیLWp8c�"O`��'�+|����C^'8�n�"OV��+RI��RT��9�x��"O&�����
Tk� 
gB��0A8�"Oޝ[a����a�Z�x H�"Ohm�wGP!X4I��1O���Ig"O����k�B40e�n=���"O0Y�w�V�����e#!o#p���"OL�:A��*�i�N�3zФ"ODT� ��;R!�%��h��"OvXB�#�8�tRP��69o<�1"O�X�b��nX<�x@��m�\lpS"O�ɢш�H~�����S�ă"OdyBW�D���m��M�+�|�R"O�@w��.8ξ��U�q�����"O&�c�a�%ZX�Z����-�b0�$"O$X�db�!b�\}i��ȣsjv�iF"O��3�pT��2�-D�nj:d�"O��c�� ���aJU��"Oȍ:��B�'k44"c.�"L,�	�"O.�pRIB�Z�*)S�M:J���S"O�c1�	&8���#/�a��"OxYK���c��"���o���B0"OX	�pn4T0R�c��+�~�8T"O���]�h�&�)��!���"O,U��oK�v��cd�Z?+8�"OP�A"Ú	 pU홱�G�)6�]��u����5�Y�RbB��� ��K�@�����,P6��B��`��j��+&p��/���Aa���R�Dx��͎!�&@�ȓ}���+]iRP@a���;*���r"O��G/�3R�F��w��*�5z�"O�I��ɠ:�"�F�"��A��"Oހ䏖�$%9�� ��+���7"OXq�VaǾ6^|�yB-ָ�m� "O2�[��U97G���*�0kt9�P"O]c��-Vt��gF ,��Ö"O���LҦ/m��3t��4�;"O$ધϜ�3������A]�l���"O�͓R�3���#'g�@ö"O��╉_,.����"�no2��"O�Y��).��%���2�N�H1"O*iӣ!�/d����O���I95"O�F6?̴M�dl z�@�j�y�<�3L��ڰ��&h��-#��y�<q��J�;Lx�i�(S��k�<��_��]���[�q,�i�D�^A�<Q�� e�X���G�!d�4<��	�|�<Q�Q� �8�@�O���^�<1�M���q��)�hDA��@Y�<�B��d��s��& ���R�<�d��Osұ!�#�Se�T�*�M�<� �H7�_� ���CW�	8H��l:�"Oг�d�S�<@A4F�E[*���"O���T*2���!��[�&K����"O����Φ[#
�Q���9L5����"O�a0N2�P4�_�dTL\Y�"O�a�4���%R�h��H��.��"O>�HƂ�?�srΞ*(�r�;"O���!� 4x��#F��%"O<�OՑL欘y4��"q�q�"O��AC����dn�^D��"O�\BChM��IA��U���X��"O��@BJ�pǎaX�
Y:{�y'"O���!�& hX���I��K��8�"OP�r5�D�muD�è
f���P"O���P!Zi�ah��"� ��"O��`ǈ}<V�PQgï*i��"O�����h� E�Ŋ�-�T�""O���aWo3�4r��^�Vz�Y�7"O^�k���_\�I��e�9h= �Z�"O�Re ߄1��O��Pb�"OF�a'��S��Y␂�4����"O,@�G��-s��S��,hkH�v"OZL�a]��PS���"�<jw"OJ-[766+��4��(�ā
�"O�Dh�*\�I0��tY�!T���G"O.��vω<u9`1rG獭k5ƽ:�"OJ�$nF?R�>D;��8nH.��"OƤp�T�4�(�5~��(�$"O��X��ʒ}�J�9�g�dv6LE"O�"%�Za"�hg�S�\���G"O"�y!A��D�P|æ��cN��"O� �,�{��h2�U�bЩ�T"Oj�Bm�w�Ι��]�!T�"OF�`�ϒ((؞��%dK%4h`e"O��S��H@�BD�v%.8�"OJ�'-Ab$@�Ȃ�j<���"O0d��.4*X��錉\}�Is"O>��%��\�m�HY&l`"O�}C��U�iI��fδt�a�"Of�h0I;J;��H�R��50�"O|2��DA@�S�g���ȔK�"O��*���D��B��^�`��Y�"OtM��-�*i+d0	W)%u8��0u"O�g���>�Z�����)!�Q�D"O���'��Xrzb# �]�ɸ#"O���퍿xW�����*\�(l�F"OƜ���/�R���!;�$�"O�9��@�1X��w�X�dH�"OTa�ۏ-�D5��F�Ѣ`9�"O�Yp��8�~@�P�Y�H�N�B"O��掝�P�V��-J��@84"O�Y��I�gZ��K��[*,�-y�"OIȥ�?�:eS��Q�n�<�
v"O�u�4M�4+^�\��Z�T��܂T"O�tB��ܐl�`1#h��Pm�i�q"OTK#i�"M���蚶*y�Y�"O�T(�b�fX�X���SHfx�g"O"d���Ït�b �`�I�W7�I�"O��(A��%D� [�j@R��B�"O�(%�y��xC��_O4E��"O����L,x ������;\���Q"Op��!���:��LY琇BK�=�"O`��A�m׆A�U�ǹ18Ĵ+D"O*M���o�v�J�OLN�[w"O� �!�Ê��M�J�zg�ӹ��"O<Af'�p	ʁX3��IDN|ȗ"ON|��ϭS^� �&��@92A�"OlT��lg�H@�%͓$lH[�"O�]H#�
;�tP��$�!*��"V"O|��EH-VP��*�#Øx�"�w"O>�j���W5ʉ��"B���a�"O��2A���f�	'V�J��"O�UpѠI
�YR�<18��"OҐ8��7f�,Й�ĲwL"���"O�8��� ����O��vΨm�&"O(�q'��1��� $n[+���A2"OؑP��(?�ޠ#�영z�V��3"O�����i�� ��"8a�"O��csi��H�pt)V``x��"O�x�'E/_Fdi��$8^�\�%"Or��ū���uQ�L;˴�z�"O�D3 Õ�N�����Њ�f�ڣ"O��pף�,�<|�\}�@��P"ON��D��e����J�7_xʤۇ"OE�'�#h��k�	 �HYT1#T"OfpZSa[�jĊ�"�7T>2]�"O�A��f� /R���A�5U^S�"O�-06�8�T����^?����"O^hrAd�5X��:I�`,� Y"O:���(�j��`���:y�P�Ae"O����N�;S�x�H���e�4�j "OD�`Dh��C�"H���H�+��"T"O@XK#�ަ�Ґ��(Q��Be�"OJPB��O'b��1�d�p(�5��"OD՛�'�DAR��e̻)0L�F"O\�b 7ט����݌H�8��"Ol��G��M�0)���+.&��"O䠉0*ڰS"9�1��PBDz�"O�,;��S��L��*@-�<;�"On�1�[30S<)��H��*����"O�9U
]0l
���gW)&��5�P"O�#�	�Z�t��s�Z.\!2�(b"O���𨎋\@D��Δ]zD�V"O��
�Y(M dTi7�"d��V"O"�[Q���	s�n�"7Jl�h�"O�8����)|�Z1+�흋|/�q(�"O0�QN�n,HaY7l��y:v��"Op($�Q�(>ny�ʘ�X7VD C"OzD����6a��$hX��0,h"O���<W��A  *V�XI2"OP$��j�+�ea 	I�h� ��"O�}��c_�jaT�Q�@��$�6"O(����?7��h��Ο��,]� "Oٴb�3#�
%�� �>����u"O��g�l2j+���F�p�ҥ"O�y��6f0R�{P�*�����"O�t: �Q=� ��ō�0��["O�X@�0k"j t�]��q�"Obx
dDJ8JdM
����"O����ֳ	N�S@Mۀ?����4"Op{w���B�j<�Af�"�Y�"Od���
�(i�\���f��v�ZD�4"O�����Ԭȹ�*�! �,�Xb"O��JvD��[R�|�WOS�J��A�"O��ʞ��̌�F����8��g"O\�ʂ�i�b×h�	�pY:S"O��3)N�I�ب�UG[*=|آ�"O�Ue��YQ�\����`N�#A!�� 0D�$��� ��`�R�5��8d"O�q�Э\!xD։����=���ȕ"O�aB���[k��A�,K��"�"O 蘄�W
E��K�i�D�
�"O�=�aY��z��`(Ψ1���"O�D3���	+.�hb2j���"Oׂ6,��y� �o��(E"O*�˷5�P���Np~4��"O-:S/	�>4S0�ӑ~���"OPl�V)Tb���b�S������"Oz�W��78QP�I�O�M���Cd"Oz`H�B�(ѐ� 04�\��DV��G{��iJ�g���g�Z�{_e'�Ɖa`Q��D{*���ê�i�"�"�&ƒ;r�"O�����E(�~��P$șF�p$ "O9�W?VY�v���DLz "Of�����<Tv�,a֪
;!��`�"O0	��j�0q04h��_\�V"OBt9�f�:0�����I�d��3"O�x��̅I�|Q)Sh֢9(C"O���G��-)���ǋ�lDE�P"O��ѣ��#,�xm�"�Bs"O�9�ǘVg8-�C�ܨ	�܄�w"O|лsk_�4��k+�,<��"O���ăRҘ�;�Jj�|�@�"OZ���'��7���1�)����g"O��[U
QfUr9H�mɈO��bA"O8C��33&P2s�v�=�"O����h4@�
a1ע����"O(�Ŧĥd����B�%��10g"O�d`S�ͩ�=��
g�i�F"O^�� ;�� Yj`bi�"O���ua��r-n5be�O�SN-s"O6���o�6(T����J�>�@("O�D÷M;���d$3�ZE�#"Oڜ#��"r����BN��8�`�"ODZ�.V�Rڈ{�F�Zu`�r"O$�3�ŷ`W���&�!l�Cp"O�m�s(K�A�Ջg�V8Y<�bQ"O��:nD>Gl �؁�Q��"Of��C�D�h���#�qKʝ�"OȼAU��l��-����E?��Z�"O�����jXZ�	�T�Ҡ �"O���0�T�d-�B��V*Eb�"O�	[tCˎH��Q?P`|2A"O���'@ӊD>���ܭ�*�Q"OT�;҉@1qyb��Te �f�8`"O����6LL5�6��3���2"O�\��f��\x�-��O�,	�<HG"O�*�jM�++\Pq�M6c� MY�"O����<�m@c�J�6�&���"O�%Z���	+�zr�����"ON%�u��eYꈊ�,��|�Z�;C"O������mntaR7���7��� P"Oh\�f�6�Nl��KV!Ev^��"OҀ��l#<D�8C���'[,X�$"O�dk�k/괹P�bF��`�"O�A�p�Ҵ_���E��*4� "O((b��D��%bBh�i���w"O���RY�s��d+�M�3B���H�"O	J��T�pd�l@;��XK�"ODi��@M�3�MâM��C*~��"O��#��/cK��G-�y�d)4"OB�u�ʪP��e`��R�ܕ`2"O� ~H��ƞ<v��٤�@�EC�P[�"O�}J�CD�H
"	�U� .�4)a"O��*�C��W�� H�E������=��{�m՗�������x�����H���yҋA�V�r$[��?x����2!��y�m�<�	��ES9tRz���ی�y�c�-11�MI��}ex��Ȥ9�B�ɰS��Q���Q�:�XƆ��	�B�ɪ��4m�r� �6)F�F�B�4A��2�Ϗ���ہOXk$B䉟5k~�r@8U�|zu�x�(B�I�EU�dQv'�b`097l��1��C�I0`����B��#L��1����pC�7A�0L�$��:��K[�i���4D��[�#D$6Ҥ�a�EP����3D��J�O�9L1l�!�j�!�u�c�1D�<�.A�~��� ��^�Z8c#e%D�Lc#aC�V�S��y;28K�n(D��Y⡚�Zh"��.���$�8D�P�#�],4����8^I�E���<D��C��L�P	���\$D���A�'D��0,�B������ڴX���3"�8D��k�� L`V�xb�F��M)6D�x�N�Q�Ys�$�%*z��I�m3lOj�̐�'M(�xQ�b�A5�]8�	0D�{'��)2D��w�]!9�]C�-D���A��W��U�Q�T�d�0�a/D�0����_�Lp� T�7����(8D�`#��E�`��9�#B�mF�1P�+D��u&H3o6�p�VJ6\��)4D�l;5�Z�����ӧ��鵤3D�p���X�	a�ms��J,����1D�x�ե��a�P���g[�v��<A�`1D�ۇ�57��$��,�(q /D��R�LI9|��Y����
JZ����E!D�4aa$�+�|�¢�X���Lr�� D�XH�BחX�D��u(׏�R����*D����M
%�AA���Hx>��"-*D�\hX�[�8�2B�6�ؓ5D��� ��tt��Q���i��[�2D�l)��$�ѳ`�H��@�k6D�<"q+�(Kr�! 	�,���Y�5D�A�ǔ \{��ۤ�4%�iJ �'D��:��W4	�:��1A -�p���0D���O�"/]j���G��D'���aH,D���"�����<��/Mjj�,�$�)D�@a�)V$J�ҙ+�h��s��d��E(D�Xc4��*Q���StFL7�ź�L0D��#e��#-�V�hD�_�Td%�Ǣ.D����Ԡ>�S�O8+�lİ�-D� {	3G[xMS�F�(�0�+��&D��pB�Y�'j^(�ǨQ�Z^�-�"�#D��K�/ޫ<�z�BD�vݸ!�@N.D��I!�Z#�
��pw�M!�9D���@)�{,uۑ	�V��)�J*D��е�ķM1���*�k�$b$H=D�h���S�=��U*U��<�` ⅊.D�d����_��j�E�*L@�j)D�������)���y0�D�je8ao$D��bA�!���)O�O�H�A��"D��`4"����aw�ۛr�2���!D�YU��<K���`�Y	��5P4F D��Kq�ݖy ����SR�2�9D���W�	,M�]R��0F�Q� "D�� ��in]�B��!. ���ʶ"O�8;�Aʀ��5��/�/����s"O�8�F(�#!)�3�v�`"O^�R��T�f�6Mbb�'k�4���"O����L�[N���kQ�b�T��"OV��wkY;g���79�J���"OX	�ȶz� ����7vFī�"O��)ӊ�1X��R��۲\TY�"Ot}�v�ڴ5[�HY��Ĺ5��{v"O$��E�C2#^����+���3"O0Lp�#�5<��Tb .��V��1�"O�a�g C�/X���b*����F"O�i�h0��v��~�g"O�8� ���!j�CC�Z��sw"O���(۾3��(N�9����R"OR-����!-�@��U�Q.<�uC "O.���"�&d��A��T+x�A"O �۲��N��B*O�)
l`""Ob�"�	:ABt�;w�@�:��*"�'5��ä��nh)���O�|	�����EzD��g��5KEe�	�'�f�Ѐi��,��X��Ҩ@�q#�'8���3MA�}�Bt ��_�:�����'x��*�큼�6��CѯDZ�9�	�'�(���"��A'�k��>����'���da��j��F�0����'D�� )�*p6����ͼW����'(���"���+�l`�'����LL�7�Y:խũ��0��'M�Q�q�Q�?K@��ĊX����
�'YD��i��RIh�R���hHT�
�'�v89��ɓ6��hf!��PV Ax�'���.��	�LeI�P̼��'�$���J2�)�E_,{u 4 �'���	�!�u��ٛԏ4>X��'�rI��K��p�$K��5�H���'�P��~|�1d�(бS
�';�H�,Ưg"��#��%=����'�����T�{������;*��[	�'r�1�2S�l� z���|܂I��'Or K�*�u�� hsi^�~�P���'��Z'��*9�L
��_-r�Ԅ8�'���EI�(dӴ�8GF�d���'Ema���"k)��8��)�\���'J"`4k݌g�z�&�ԣJe���'��!j)�
V+�̑���qFPh	�'C���S���T�q�?O��	�'M���N4�Y���"xV�I�'-l�h*Y�I�$��G>*��U��'�Dt�R��wy�����r��9�'��X��A,�J�S���lԶU��'x��)�F����cF�:(�B�
�'��M�D�G�=3L�[�*�>!�
�'�V�p�"
0Ѽ�R�� �D��'����@�@���@���(�DTK�'��Eb�FЀ0����&IM�����'������!	��Z7gL���[�'�j��#-A�v��ˆ'F�}�	�'��Iu1c�����R�|°O`�{�aӭL�R͐�cV�6Y�v�'��O,3L�E4�e
c]U�訊"O�ؤH� :jH1bJ�1�t]���d.�S�'O��5����#Rmz书��$YB�t�ȓk��$stI���j#�Z�hר)���ZuX��^hF䣷#o$0�9��
mb!�� �|�d�)svx�(�
?S��Ũ ŉGH<Y�m���ë�*6�)JBQ�������(d�hPEnҦ
�V���ǚ�{�!�֣FSd�"A�@�4�چc�7�qOLiGzJ~�Сܨ3�\�J�\�>��=jV��Q�<IWΟ)�Dt��Z�[:�)�R�'N��񄄮3ˮ�ZФ�F�ޅ*q��H!�d�	���ƯH+`~v�ɵ�Q�p�攠	�'��hZ�L�Ĉ��B+_�^A
ד#|qO������A��5X�Ł$�dx�"O��R��0i��X�A���B�byAP�$�a���'g�Z���i�
/�ܡ�!�ͻz�t�ȓU��Aj�i�H�*�K%S;L�eEyR�1Oܹa���0\r%��� @�歘"O�a��+�#�\ k��	�f1��b�6�Px"�+�n�3FA-L�Y&�B��p=I��$I�LQ2�k�/v�ia
�'3v!��Z�3�哱�H$���2IS�yqO�dEzJ~�4��X�e���پ[0Dġ���C�<����A�]�'	?���Tz�'CB���B�i�f��e���O�ZH�r��c!��e<:HS�OԷZ��C�Aj�Y�'g�R��Kz�@�o�-�X$�	��ҋ{��Q�@�(r��/,��7NА�y�MUR�pVT 8`L��J�}���E{J~�S�M�z~L�#Ԧ,7� P��JZ�<��&�c\�D���(;���+EO
I�'�ayb�-3"D��!|y���ݧ��?�T@�2]Y�iP��[ n��I&�@��!���?4�"�K�"ZizSWH�mp xEG�s�R!Fy��"[kx"|��00����Fh2�Elx�2�#�Dj�'����1�rް�CA$�4B�� ��O���>�)�';p$��)܏1��!���.�" $�,��O�-�qOq�~�Q0��-=�4��Ő _`h�ßxb)���=1"#�Z�*F��??䤁	ĭ� %qO��&`;�3}��Yوp˓%�
pB��+��J���x3<��2�W�!��t2��0��#�Aq؟�ف�	���"t��3��q��4<OđF���w�!�׎ݩT�DU�.�^���ȓc)�,�焝n��,Ba�<'������O2��� ҨN�JA�׭\�+����'��2p�Z)���3�)��).*�P�'u\A�	,]��v��	+���'~��e�^�j��TH����x��'t�|�W ����:T(�8}и��'���[
K��-�r�	P���'��x��\�%��iY����Rd��'��ѣt��NHD\�A���x���k�'"A�X%:�����;pu�9y�'Gz�K4�S&=?�t��'�"E��{�'N�يV�[,}�h��L9W����'���;MȂ�j�Ɂ
cN!#	�'2@��	k�HY2�jۂ�f]��'���!t�T�.,���7.�=���+�'9����)FoЌ���i�1��'�JԻ+��&�r�Fb��lPB9�'���!���95��)�Ԉ�=d�D��
�'Ќݣg�	H
5kTiA6]e�Qj�'Ȃ����!�&E�S�
JhH$I�'�h�����-i��a�+� `�	�':�)����Yx�{3cޚ��(��'� �Aw���"|5�"���	��'�����#U>Hz������B0�	�'{�U۔���=�*��tc]'O��	��� �hrU)�?8kft�%�
��؉"O�x"�A�w��9�G�@f&�`�"OH����H��*C S?�)f"OHUc�eǴ	��	�����*ě�"OrUJ�17�������'.@@�f"O젶 ȿ}�t�qm�M:��K6"O�͡"�� O��ܠ��	�?��C�'�1LNڬu��>�hAFa� �d
�'j��7`�D���sE��I1蹣���bC���G�u��54 bЉܲy��m���ݣp0H����q���F>�Ȉ����$+`m��P���W���v��$"ł,?6"~n�+n~jR�&[*:��$G��#�FC�ɣ0�A��(˺pY�P`�߬JИ0`�����;�ŀ�ݲ4�?�C��	������L�����ތr�����R�j�[4��X[��� �G�m��, �-��e 8�'ξ	�pT���J#� ��D2VH�qcu��y�t�Y&�# ��HkTQ�`��,�V
@�z����
�FC�H^w�l��m��%�!e���0��'�~�c$	YP�p��:$�S#nW�E��	a�c��p�#bY07�v�{IŖ�y'`�!&�n����*(�D���k�y�^=\(�-Y���7�|�;��¢.�����BX�s�x�#NV8'� 0���\+�5�ˇ=��'m�%�vDSh��Y�3���$�k
�9��(H!(C>!c�	Ӷ�\%f4�,[dk��Z�� )�$Z�L��u"6C3F�
̉����L�y�/E�x?N�V��H�X���ƴ��'��Ѩ�g��j�d�p��G![���8�i��jr���6OU�
x�J@�T���Ce��*:cVC�<g�
L� g�Lf��ҵ!���SfJ�6yޱ���ϬX�eY�	��d�X�'�8��¼k�CG�:rҥ�e�܆s*�Z��
}�<ib�إY�t�f�ʷJ<^�bS�]#��y��L�m��X�D��3Y�̧X�l���K�O5�'�I�n�@g*|��˚-V� �1�_�d��v����6ܒ�/�h��	B4�źb(2<8�D��<�����@�V�֢�2May�� ;&x��� -�-V=T9�7���(Oz�Q���%p汩��C�P1L�����d��C�+�E�p�� �Y�xϴ�XW��%H��C�ɒB[�x ^&��)j�@E&lF6-9���1��E��뜡 NP��RFS�`C��&�����Ӫ�7zúY�Sn�4Y�>�c.D�@S4�K�Bʀ�+�f��<������C��sl��Ro�u�sZ�,��ӡdD��R��\�I�I!��1*�d��t댃2����d�1��b��-@�z�1��	L��fE�~mB���	��d�:l�`�iQXL��f4,O���A��J�"�
�M|�V��剛o����1�O�O�:�z�z�B��v-�@���UjܑO8%y���u�)ka��XH<QFc�%�X�k�\)o
(�A�M.e61p�M�bw޹�f ��"�<��cЃ&�R�sƗ��;Nɠ�:�)�'2���RO�7f��%�ȓ|��E9Gъ�̋08|�'��Q��c�Ƚtʨ AC}�"jC�CN<��;�Ԙ��L� \���z��y8����kѯD�n��!`E5Z9���6��;�T��Չ���Bx�%c�j	n(����(^�} ��'��d#����VZ�bWdF�l68!򤓢]��p]:��b���'9�@�A鑯_Y����J�q����fд��Y!�lM�@�!��M���W!�T��M��'ƅi����d I�~n	uj�&+rpx�&�KN���waFP���ph��/چkݸ��ƪAvF>ę�"ORi�ri��Zֺ��EW1h2��چ*�,���M.ۅаk5��Z?Ѣ�W�L>1����)l�H31/U��8���hX��QQ$ـSz�*Y%�J�{��]�-6�(��S/HV�iI�?T���"�"��y��Q�R������=K� #v���hO�a`�&��};��C/�5Ą	R��_FkH9s@�"��ˑ�PK�i�ë3D���n��7�� �+҈́T�u�hC!���BMXK P��C�6Q>�ڔ`�-f<�B�b��?��]hG�&D�:6�R�S�����V:��Sg) aG"� ���Oځy�Ø�w��O7�O8�ʑa@(2րT������l�B�'S�y��C�A�B��r����B���φ<04�Ě*��yk�m�DI��u��?��SB��C����Q��ONxR$ɽ+|
���(F<>瓶V8��c�����;c����HC�I�+U�X�c�'x�l�#`P~�V�'�<��g�������f�S:\,�#�%A��Ѷg��h^C�	&��i�\�\A�eZi�$C�	�4��`Z"��&��@ެU���'�F�+��uy�g�z��	IF��@���f�Ȃ��'��#=%>� @���eF�	�p�CeŐl���"O��N<̈a�D��|� ��6"O����DXB����K���u��"O��KÊO�_;��(��ǌ[��"OD��_75�Lq  ),�Ȕ�4"O���H��u��,�Ҕ �D��ȓ��`L�H
�4��eII=��ȓy�f��\�c�d9b��җ+�&L��eEPh±�� q�б9�
�(vR$�ȓU6m33�ض+�jQI�g�=.�l��c��I�ڻd|�p�A?j�t��?���vӚ͘�A�)T�(�\��ȓA�4�	���$S�Ji��X�lڢ=�ȓU��k���r��	7�J�ȓM v8S傎�Z��]�m��Ć��܉4o@M2��JS4!���ȓ	X �"$�BM��Q4@�=�ȓ��@�v�6qA�#��J# ���d0Z���>"�D�� R�BU���ȓO:������;l9cwN?q�Zt��Ǥ���K��"�p����Z�nA:C�I*�&e@��#�j��"���^B�	�&�f8��*�@_~�$h�-�:B�	�O;�����u8�Sc�����B�	�b7�t�F Q;�,Y�S��~�B��4*�9�ŒL 6� �MF-6�B��)�j�3��8D��cՂMKdB�I:b�R�D��y��TR��P�m�VB䉸y�t��䧆-l����C3QB��Yx�]��	,4X(�C�'�C�	�=�n$Rp��'_qP�' ��C䉼��:�e�\-Q�DX�%��C�!}�����O)T7 �y�a�/!vC�Ic�Х��N.��da O�zxC䉁;�ޭP�c<��p'(6I&C�I�'����kמF��@ 3�ŔM ZB�I�t�\�ZrK�/ ^�����֩T.!� �8͐�숫P�P�HRn
��!�d��-fl��� �w����`ȾL�!�DјC�ڐ��GJ������]M!��SFEy�ㄊQ�$Q��O[!��W�G��*�Ovfv��rx!��NQ��ȱOB<c� ��b��y�!��.�첗���yh�-p��g!�dA�#`~�m�#(R�`�b�@#fU!�$5~}�$BS͂�1ol�J¨��]M!�d_�5<����Ϫ [�YGd�!��Pd��J�+3V�D�'�	k!�dZ�&'0a�W�<P�(�� �M1	�!�dA\�@3K�D_���C/YF!�$���؋�,��o ��0��ʇ)"!�d��A�B�a0��g�lCA�5�!��
�D��)�WGS;6��)[�gף �!�dĝ/C��ƥ_�Sߌ���FD�K�!��$0��͚פD+�xlYC"U��!�$Y�F<�ɓ"+�4�.�#+΋z�!� %�jB��<&�� b��̕r!��Vr@��eI7f	�JD��!�E� �82���w�$Ai��L�?!�$K
|�d4�Ǎ2@CXq)T�a�!�H4. �A�J��D��@&] !��U�<;�I֬w3��BCG�-,!�d=>v�S�하(`�W�м^!��-ou����$�C�9s�o�N!�� Ѱ M��DmqH�"j��C�"O��;g)F,)1pSpʔ2���$"O(����¡2�@��P�d��9PG"O�u�S��� ꕃ��\�PL���"O� TK��q�\�S$Y�@�(Lp�"O��1�Z�Y��Qbe�]�
�
�"O�t;�.ޔA�td�G��,���8�"O� K���Fj"� @#�d5y%"O�I���~p�(����pUґy"O��3�2Gl��'L5�(�!"O:�¶g���FeD�EGdT�"O�k�ߎe$ԣ�c[ H���"O�k���2&%��L�3 �J�A"O4��D�F7^�@�3�B����;$"O�}(� �IF͒�N�~���&"O��*�FK+y|B�1��.i�,��"O�{Q�1(�1`��#���%"O�(�� ��)���ߥ1�(��$"Oʴ2Ղ`޲X�)��4v$�`"O���.Y(o���F��Y��S"O�m��W��@��'��	ݮ�
C"O�T�Ԋ\A�v�YG�L�
�r�"OJ`3t�H.C�H\�fͦ
Ĥ��"O�y��x�nB�W�9�Δ� "O��R���7��L�'"��䒐��"O��n�!r��	.�;,�?�y2 ��?$�Q�gL#=���0oF��y��j����ԓ�,l������y� ,��@�"r^���A%�yŁ�j�F�2��ʐl�~0�@-Q��y��C92X
�	�K�!dL�y!D�4�yRi��@��ä��)�4�S�[5�yb-y:� �d
�1.�BK�yB�\�E$�+�&��	k� +��yrB�&_��e���	�x�^�!c���y2 -k���oR����jr���y�(�=ZH���/�x+��1��y"�Y�'�(���Nή��eP�$̦�y"&
�l���2f�Ό{�����@A��y�5'��-|�=�w��)�yR��\�b)����w�Nسւ��y�Y $��� a�YT�Jg��y¯��2l���ҩ[ir 
7Nƹ�y��X�UP���'KK���8����y��_J}���ݫ9j��NS��yr�1I)v���A��3�`�БhѸ�yR�E;l4^yS7�]� �lap�C���y���EÄL�T��0#^���R/ܓ�yrhœ�0��e��v)�lW/�y��P�%EJ��&U9�,m�@׎�y.H*=ʶ٨e�E%)������F?�yB��;Q����"%Zթ3%�>�y�
$��SJk��P�a���ybAɪ!���! CK�j�����#��y����*g4P	�n�kW�(�0'��y��,l�0�K�aR.Z�� ���Ԋ�y��+=$���7]r��w����yr�^3�CU,�5RJ� �����y���_��L��HP��|��
�1�y�mS�gԮ���G�:H:gIH�y�K��l�>�cG?��Iy��\��yB�Y�(�$d"�aY�,� ��'���y��?8�!�D��"��e�c��y����0�(�!�+"צai����y
� �=�FN�.�x��2��/k�2���"OT,I��]B"t�M
:��D�c"OBE��hއKM��R��׈�"-�3"O�X�,�xv �i�>a���f"O|� !�4w��9�@o��;W��Q"O��۰�0%�6��vE�l��"O���Ɠx�2�X " f\�T"Oܘp���,6�vU&`M�%���"O���6�ͦp��P&���*�Ƅ@�"O�Ղ�d�(7��#�J\�p�҅�"O�di^%M���)j��]>��""O: ��@J,�n�"b�V�p+"���"O�,if^�@lBA��/�_�!�"O��a���9��U
�1x�$��"Oء���V$R�8�/L-F���iq"O�t�!�D84� T��N� ��̻�"O���F�fC��k$m�>��-��"O��HT��
m#���L�c��IE"O�Iq���-H�2p@7J�h�,
�"O�p�c�ǅqW1i]�kU*�*�"O ��;����#j��"Iz�#�"O�D�@g��p�b�\$��0"O�$BTxQ�mQ���e�V���"O����F[1Xc�='H�V��dx"O�U����9<M��O�rqٱ"Of	҅x�@����/}lEJ#"Od�
��R*E��ܘ�䁙D�t���"O���Z�0!8��Ŋ|g>�j�"OF=�/z栣�c�71�x��"O�m�4!)s�Э�7 ������"O*�#��$zy�#P���ȉ�"OJؚ�*Ι�9@�\�w�$�a�"O����� C�Ӥ����"O��)3��61��鑂˘(�&�A�"On ��kK-Aq2�K�b1(��-��"O� T��#�`Yvn�[�fX	�"O@]˴�ǡe/���-O�H|M��"OpD�"t�J�N�/
� "O�Ĳu�	d#���GN[(d�L��"O*l�ɝ��yqFl9NA�(jF"O(y9%�2&1@���F��Гr"O
D�F��{+��S�`�{9t� "O�%�R�	��@
�/%�p�@"O6��_�E� D��)[�$�s"O(�Ǫ,���BeH��W�4$c"Oʸ��F:Yɂ]��H�s\Zl2�"O��Z�MH��;S��1C�l�[p"OF�ȉ �DbaO�f����"O4��6��7m����-�%4h|�g"O�T�b��.N�l��.�-PH��"Ox��D�C�S�� �u��N	j�B�"O� .F!Cg>�-�$B�|�C"O`���H=���K"�T��:հ�"Oҩ2'��>x� y'HH~6��p"O�Z�!qyN��ɫdm:���"O�%�C�
^����� M@:��c"OV�Jd� ,Z ,m4)��D1�t�"OR0�f��+g �)����SK���"O�x�tL�8B�9����4Q1�E�%"O.�AjC(�����F��j$��C�"O� �d��1��x���%T|�"O>5��)���)!CV>y�ѫ@"O�蒄�FP���QL�Ԃ�?o�!��qe��J/Y-"ؤ�����A�!�� 2�`e�!	�r�(�g<[(N�P�"O*8�4�V ������C �g"O�t�VL�:,{y!QN�/b�X�pp"O܁#4KO4]{��mA��LQT"O@�#��'"�`)�%]kҺH&"O�P#"S�=#�A��$B'ܶ
!�d�7X�҉)3���3\��H��թ!򤚤pn�0I��
�Vb!���
�!�D�� <Qb�Բ��(�V6J�!�T�t^�S�i�;$	� #!�E 6��@��c� kv�L�$�F�!�_�['V����Y�9�ڌ�%�OX�!򄇿q~��x�� (��H�"�$�!�dӓ� ��$o�0����`�;*!�Ѿ*�$l�q�[�*@1���\!�dC
$(9��B�T�"Tq�e���!�$X'[��Uj6NM�2%�-�`C��$�!��x�PI��a��]0]�bA�!�D�%�C�"�A����s@�G�!�dC,P�Hh��ه�0�� ��!�C�m٪Zn��A�HI���8~!�D��tD��)ʰ�����G�Jb!�ď��x�䆙�|���
�cM!�d�N2��t��T|�a��!Ի)2!�D�?Ũ�K��Sov�3 �F?!�D�& �����:	Z��!��PyC�1k��U��J��`:��^;�0=)U"O�l.�+�O\���eKf�l>�R��2�ڱ��@l}�a�*~�Z��Į4x`�
#�M��ا���H�@��1c��Gظ�[���(��<��O4͛�e���Z4��+Z�tЉ�{��U-Y;�O�OvpBV�պ�\�r�谑�L�,����w�S�'/&�GX��B4�D럶!�68��8��ɀ����
WU0��իK�W�*y���-�ޭxE%�h�S�O"�t�QO�*U`�FI�8l�3�+�IMra��+K
q(a�DmY���9pS���'��������!+-�A$D[�X��8���\<���6^�J��?�J�����~�K�.X\��i�	T?I��2���h��]iC���*�@��#�˻w[>�a4d�6}��}��)Hp��`��IxO4�t�:6���{b�G��0|�`H����\��!�/	ޥҤ]M̓/ܡڴ"=�~JG�¡]��eIE��6tf2�K�CY1�N��6��`��n�2�ا��8z�	���x`A�P�G��,`��O�|�T�#�)�'RI�X���P�)J�G_([��!�$L��O�?Ya��Z�,���2�%�1'���GJՕ�?�J>�Wj5���"c$ #AS�4
7��kZ�I	a��µ-�⟒���x��ՆbE�HX��+8�y�җ>���������OF�� 霠_�(�,��1�U�~bn�/y��O�>�ᰄ��f�f���cN�v�T�� �L�J�`���)��h�̐�����>k�<�F/	Ta ��?�
,��P:4C� o�����D�����a��D��뵊�O��$ژP���i�*�>a�t�Ыd)�U�y�p�Z!W�P@Jޖ:� ��?9r�>�j�!�skb�(�
D�<!�d��3d(�P�e �m�$��I�<)Ue��\|�t��?8R}�3/�K�<I��!��d��~m q�hI�<ѠdLd�B���X��Y� �G�<Q��M�'���D�������@�<9��ۗd�^�`6
�E����BB�|�<�� I'!���/�C|}���@�<ѐ쟲V�m�a�ڎ%Q u�!�It�<�q��bY�`p�ُ(���6�r�<A�Ëc�� A�c�+5jh�3O�n�<�0�N-W��N��( ��E@�<��� �$h���(nF��ؗ�t�<� �a��/X�cd��1�z�3"OؕAcɛ�D&�r�m�{E:ɻ2"O�LY�h�*5�����j�:,��8�"OLT%H�3:ۚ��W�P0](�4"O��V��v́3W(�J,�:!"O~`���0�:�5��3#,Q�a"O�J���E��s�L��F�JA"OZ���MJ7��	�@&¢X�pu�t"O�D��u[R�
�k���A%"O���e��̈�>Wx���"ON}"p�Ԃ'�Ĵ[�/��JP0-b�"ON��5��q.�UaĆ "��E�t"O@q�g���+�[�#��t[B"O�\R����H���A7fw��3�"O����(w�
$P׎
�6a�d�*OИK�`
8�|�+We�)�"���'�N�s�[�1��m�fÛUVr!��'{x�ə�kgR�aAҾa� M�'֕z�o���DZ�$^��,�'D,���4,�0H�L$>\s�'^�1���R�&���̶�8�K�'Rj�(�I�s�F�2T��w��1�'8�y�i����F�</� J�'��(vM�O�F��
7I~���'�uS������1�Ђ=�d�I�'~@mQ�k_�Y?^q0v��<	�t��',�uޕ�.��/�{��̨�'��̱w�ܻq�ZUy"�ܣ]ט���'R��� 
V�w����R�P��k�'���2�L/�铄���%����'�̀r%0�ra�l��R��
�'ט��1;nP��ʌ\g�}C�'#��Iw�ԍQ�(y��W ^@�p
�'Ep�������� 00�܆Y� ��	�'K��H7,?�^0��g#�Y#
�'�]8�M�}8���ݙ�rPH�'�P�i��I�2"��҆.eH��''Ra�&���2;�@O�2ر�'
T���A�5����W(K10���h�'s��PGz��pV�,�T-�
�'�(�H
�"��E�$����
�'�n�ac���ה2CIT�d
�'$v�F!��?��Uo������'��ѭ~�PE0d�� �̡��'s�y��eC+���x�E1C�����'=�$H�
�?o�}��� >��̙�'��<���|��Y3#�Z�.���'n]��$�*~�޴(S=|�(� �'��(����R�"�ť�uƼXp
�'^8����N�sZ�J劝|V����'���
GJ�"X�'ݵh��H��'����נ	%x���`�v��=��'1@��r%D)S�L���!]v�V%k�'��Ĩ��G�(�d%���)fh�ٳ�'!Z��`G�l������I1_0�P�'Ad�pӡ�MP>MyeII"�U 
�'�!���G��h�ħG�I��"O�; k����]���'��#�yR�T�G�ȅ9��@��"�� ��y2��:S'v�R�!q�r�3�	�+�y�V���QzW�8e`����� �y"�}���p�R)?0�ҥղ�ybɒ	{߶a�7�ʲ'`�a�;�y�-�r|T��p�U$���t"��y
� �1R���� ,�w�&~����"O���惫y��ȳ�(�3K��kR"O�쓇B�>\�nL�C풙J=(jE"O"t����0���<)7n�Xd"O��$�]6E�����_B<M�"OPYBKP�W�����QA�U�1"O����Z� �4�a� 2���"OV,���xBtt�֌���P;V"O��˶R�.����X)v����"Ot�sAZ�i�L��'؎�ɢ&"ON��e���>vB�b�D�Q�"O^Tbp+��qWۈq� �b"O�8��
�Un��I�|1�*a"O�X!��F���3�	l(yb�"ONL��O�ycPH��'�:.!���&"O,���n��k�`Z�LJ� ��s"O|�⃑@[\�كJ� 5��"O�����
pp%#i�#�ܐy�"Oęȡ͆,4T��B�g�o�nEr7"Oh��D�1ʒE;�%GŰ��"Oii���K�L��%ɱĸ��"Oz��E��^��e��!�5��s�<At�5i�P5"�ʁ�0��I�<id�Nz_�⊛�gsBdi'%�D�<�E"FG_:�)[4\pc�b�T�<��A�Qb�T��/��j�^��dFI�<�a �.�<� �+�#1�-;���@�<1vd��TG�G�
c�u+�.D�<2�öhET���V���!)�e�<Q�*Z�* Z'Ԓ�`����_[�<Ydk�`�j�[�cÏy.^M�HOV�<�H��D��tXq��s�|�Sd�P�<����\XZ��U�N*^��J���J�<�M�²��q��Q��p�'HR�<�nΘj��pE�5�L"��YK�<�b���B�Ҕ�$�ɉ5yΘQCϓE�<���>x��ƈ�@���a7!�U�<Y����N�"0�Ӫ� UᖅN�<�僈�Ɖz$�I<[��}+��BM�<��m��S7TP�1G��`��ͪV�YL�<Yd��2V�e�$��,
�,�%��A�<����p���JP�p<���i��<����=O��1��(�B��ChB}�<��dD�WK�A�ahK�1��+��K|�<�G�Y�6@Y"�T��v��FJR�<IQ�Ox��iTMO�D�G,�Q�<�яT�'�:��	�5��q� V�<����/G�� #�*ø([HQ�W�i�<Qbn�l����uN�2Db��waL�<i�[�=�L!s,O�u?R��)OF�<�6i�(��, '��8���Ռ�Y�<Y�j$LQ|��%(N�_�ܥ��'U�<i���"�$����ì�a@/�M�<iD����xr�ƈ"�\�U�IM<���h��[�ϋ#��ŹK@�{�)��B�f��7/C"�h�7+�\�f��ȓ&|��x���+|��xC�	
y���ȓ7����4�Q#���xB�Ň^��E��}'V��S���.&�	�p�<l�N)��*;�q��%�e�Ȥ 5b\/�A�ȓR/�`1H�%��0�ԢS>~��ȓ
� h�
�'����j3tx�xl_(<�GA\�(��E�U���g*�8�M�k�<ɑH�"� ��%�C/x�b4� k�<� ���R�1�6(p�k�_��y�"Ov����ϧ,j8|��6ߊ�"O�X0q�۷~ ��0j@ruBIx�"O����r��H:�N_:Ѭ���"O�ݠЩ %S|ŊwoÚ؉��'�!��N�CY���GR�� B��Rw!��*N��P`�)�;C��#�	e!�$���V��&��g<,`��B/X�!�䐧k���*��$# ��V`�9�!�䞩>~x%��i��*	b�үߜ�!�DA7"�p�*������X�[�!�d�@�85���;o��hS֟s�!�$�C�
���ډ%i�-c����!� ���X	B��(�"U�!�C"D+@�F�.T��@�B��<7�!�ă�S���Rqc̟/�4��V��	�!�D�X�ȩw���,�Pؘ�)	�3�!���XΦ��VFH���\Y/[)�!��"�+�� �ͨ�!�;
t���'���c��Xv��⟟4wa��'�꭫� F�JB����ȇ�~F��
�'�ti$ ��G�Rx(#N���'���s���X	�
-؈yS�'�*�'Hڿ%���U-C��p��'5���A�
�-��ue�<�V�h�'{��eH�$��p�.49
�'kެ3�l�F�h� EP�q0��S	�'����B�`-��Y��ڐb�����'#��h1�Oj\���e�SL�5A
�'B�ԙ2���9t�(�U_~qhq�
�'\���GO�.i~����ÅM����'s2��v+��~���폙I���'ڦ�*SF�p46�R�j 2OΝK�'�f��h@ H��u`��%e��'��	Y���1�@Y�gC�>"p��
�'��Y���(JԹ1�[N�R!�	�'��u��.��`��� J�� "
�'��d�E�-a�xa� /�%Hl�0:�'�NH����+=謌u�U	9���C�'xU� ��x�e�T�3�&��'�����S�ڄ/�"Sn��y��
BU���ƛ���iH"K��y�)�+;�:�I�oD�#pT��'���y�ꐈj"���-[�7�
�W��y��*&�Ф*N�'��â��yRi�'5�z k�.C#$���s.�yR#�E�����b���[��y��+nx5�s)
p�}����yrD�\3��!�64Sb���Y.�y�&FJ�ܵ�� 6SFH��n>�y"�61�t�����ڈ�7K���yb��L�]�e�2u��� �"���y2֔_=����ųCR�xi�IX?�y�)$P���A��k�.`�U�F��y"�͏1��S�m
^�(����yR
�S��t��'O�b1������y��ȨR `  ��y"D�(K���C�+3�fLh����y$� mT�1���2o��E��y�&-K `  ��<ZYѶ�
(p
�'O�m2҄� ��"B�|�F�q	�'�t@x�FKs�u�T��?oV|!�	�'�R� �]�5� �ӎK�eJ�	�'���;�C�+@>\��M��V�T1�'d�\Y�E��}�Z���8H�*��'�)*�ٓY.��g+Q�@�((��'��tេ"�%У�ֿC�U��'Z�p�� �����c3oB�Ub�!�'�\�����4�8IS�S##q@��'HP0��A9qE�������s�'��+��w+�)C�a���l#�'�:����(~�䣄h�����T���i�M��;^�]�v@ɻZ���ip�ԇ*w�<,�LD'��}��.e:Y�E�	M�%�F�@�c���ȓJYT�5&�I��	K�A�A�|نȓVnt��Z��-*3�ȟ|s���ȓ\$\lK �L{6h��g1�Є�$�0!��I.�bT�'�Q�9`���U���|f0{��<
�n,��-s0��f��R~\�h�W�c!9�ȓ9Մ��g�,�f�)����d�ȓ+>AG��&o���ê
�ub a��'h(�Y��9�J�+��G d=���ev	��2#���#r��~�^�ȓ&@L�⣧�
��-�v咣n��z?��T/&(�Qy"�4�Rć�VK`Dsp� @x�� /N���g<D��+���xp���#��r�*Ѓ8D���Qb�5o�f�FF$j�0
!�9D�xq1!�0�VX:�d�x��%�Ac6D���" .�ܵY�f��:��?D��B��p����T IKtR�b$(D��#�"�"��C�0C�Pz�� D�dhR�֗K�<Q��L�>D�L���>5,p���':�$$<D��8i��,Iz%8��ݓ&�deH�i;OPeq���=JDZ�0�n�d��T�b�P�+�!��R�>�^��� U�/�")!�m>2��)�'S�0,AR�jd�0�%!��n���L<Yի>�S�
 0�����-&��bK6U���'P�~�AV�`��pΑ���s��K<�M�+O��O�3�	8NJ�RmW;>5fqb��#L܅�	�<� �i�5e֗}����c�W�� �$"O��!�
1�0�ԐQ��}a@"O�mK�m6�	�H�5f�[�"OH"���Q9��W�@IL�Q�k,�S�OC�d*E^ИR�qi��&H�y�%�#(=@���%�??M������~r�x��	u���i,l��F#�t �kT�"� �' �x�q%���ҹ�"��>�&�޴�Px"!T�f�����N8�U�w�F��y�Oو�f��׫�g (`������'?�z�f�E�D�;���_��	@����hON6->�ӺC�Q8�I�P*ђI �̒⨆[�'5�y�*ڽPL(��
[>S��!MZ2��'�ayb�in}wM�>x��h� OH�"f`�	�'��h����z %�.��x��'� �@��I�:y�`�o;�]�
�'ּ��ȍA?$�e
��W\�}�'��ɀ�@�5��42���6>x܍Y�'�X:#,�&hm"���͞�jA.����<<OP��`ϫY!P�6O^�4+^9"U�'��L�$�5��7��aZ�O�'[fC�I6h��L 3� y��A��T�e��' Ȳr.�W�݀��b��A`�'i������ �丈"�D�]�NDp�'�`��¤:�ޔqc�C�%-\�"�}"�i��l�<I��0��1�ܰY�*��!b�u�<�5��l{@+�4V�=e�G����'�&�kD�I%:�R�T���w"��'ϊ�(eʘ5*��x$&Rk"3J>A@~�b��>���7@�S���R;nP��+!LO����5�!g[|��@�-���T�.b$�GxR��H��D�����K3����'B"�\r���8~�$J��5���ISh�/L����kӊ����}����1�˝YG�x�EՅVў���I6I���  ��aFpHђ�+2evB�ɉ~��I�V]��)§IֈB�N��S?Q	�)���8���	���cDC�Pi�(Dz��~�&�Y�����	�f���	T��|�<	4��;:�m���0O�\ٖO�@�ў"~��2@�%K�*G�J��1IJ����d�<�'&�yB&�)1F]�RJJ_�%�4�*�hO��=�'��%��)�.:�eH�l�tO�T
�'��|cԯЀ2��7�"��Y�?��O<7M3��?I�.�\�yR�%��US ��A %D�8�Ѕ��;�VE3���MʼL��?D�X3ǝ5?((S�cMZ���>D�\+gI|)9�C�\�6!Q��=D���sD�
3�����P}�V�25�?D��4% } �L{B��8�*��A)=D�`��LP+j�Vy�P.��qb�dc:�II����ƍ��݁f�ڹ�����8D�P����p����PW�>.깱�i�lh<��������V��"	�
�����k�<�G�0>�w�]!:E:��B�h�<�'S� �v�3���|~�O�g��6�S��+�`���̴7X�aY��S�_Qz��ȓ^�L��#P7*~�-9tG�=Y�%�?���_8��Ө�#��tpe�G�]V }{�5$�� ׳e�T�QGɭi_�Y��l���yi� �TD�V�^Q�H:�Z?ְ<��d�P��@˸T���s�D��!��F8P�Z`oR!:�p9pUN" b!�D�!u���cCZ�O�6h�3��Ta|��m�5/�� ��P
���S�,��q��`��\@J�v���!k}���J~֧u� ��r,X)�ԙÖ�W"j�`�#�'�����#qTJ�,���X-�J���,O��It����&�5iv���H��7?��)4,~���'��D�|Rp�O6A!�M��4A�Ԍ���W����/�.6��'qa~B�Y�G?V��C�4�������c�'�~�D�dn����� %F�=�P$�M�%�Px¾i{����+W!#�� �-�13�{r�D,�I�	��d����%T���c������$9?��'�Js�!H�$OH�yQ���Xj�O��Ӕ 8h"L�`F�aJժ��>��O�b��?��+'� aҥ�
� sDL"��<1ȃ�nØ�y����<+��RGy��)ʧD�������F�&��d�ݯVꪁ�ȓKdv�a�EZ�W4dQ��}CRl�4����b?�'�q�R�D�P;mq�#$ppX�'�%�.G�nᚐ귧H��t�@!H��x��H=xƽ�5d@�iŤl��'���HOv�I�q��"|z���44�f� �-G��^�᭄f�<�M��j`��I
h�JiSC�_�<y� If~̥� �)4�}W�[�<�Gm��'3H��S6xJ�;�&Z{�<I�'F�7�!���sb^�rE�I\�<1懓�[Vu��������~�<�!m�E\|�P"�+!��i�E<�hO?�I9U�Ld���%��D���0+ˮc�`��	��XP�AP�U����D\/g��ɺ��	S~��IjҸI��Ds���bp�Z�@jj��D"�I��#�]�G���1K׿~�����(�ɩ��A8��D�T=�h!%MԚvB䉸��:T�	\�~�t!ߋcF���hO>yq��Ҟ}��r1���ʔ!&D����o=]�!"@�-~��]`�(D�8Y�o��w:���������$D�� N�+�z���&I,q�4�&4�4 u����re�[�n}j��KN��p=q�j=: ���% �<����$b�Lx��Fx"�R8)Ƹ{��-�9����M��'��8#f��!"p�§�¨6,���'\mڤO�O�>�XfI��D�����$Y֜�B�,D��Z�ƙ���ٛR���h珹jm��IQ~�d*}J?듧yB+�}�P[�d�k��d"��?�0?�'R��pA�:i�:��F��$)�e��I�'�.�D��'���� o^�XxBw��-��O4�$?�d!����N��䬇(hH�p�I�@}�)ҧ*�|#��1=BѠ����--�Gzr�~�DÄ���`ԈS�PU�h�� �l�<�GْU�\	rA�(֌ZdF�_?I����?w���Rb�f �6)�\��B�Iʦ�Z��ӆ�\C��Z5���q�(7D�t�aB47�N���� F� ��2D��B��JA6����O��.#�LbV.D����*8��bӥy��h�B�3[�px��E"`�jI(b���*��C�0���(�Ή��
�h�$�C�	>�0x�e֑A˾��D
�Y,<B�ɏ@�a�W�V%-���PMW?%��C��;4�h��fdIjנ��!�5	H��3�c�8�n֝�!�dP#�0(�@��4����6N =D�!��|�lyc�̧J� Dg�Y�!�d�>U:��၉�t>ba�v��UP!���Qn�e�
/8H��� ʞ1!�ҩm�H�Cá�%�r�v�4[�!�O8F����d'u��i�?}!�� �� �&�$?���	V@�(Az��5"O-��]O`U�f�ǾY�Z,3@"OLs��$E��i�.Z����b�"OL��Q�8�!�*�9K�����"O<�+#̛�h�K4� ��;�"O��ɥ�!7?J૑CX�l `�"O��%�)kVRe�F�� mV�Zt"O�T������IZI� T��"OHL��d@>	.$�X��95
l5{@"O�� ��â/�rUJ�G��Y��y��"O踑�
�{f9�EYr���j�"O��.xa4�a��F|��z`"O��B�!UL��us��M{"�P�"O���4# m���RSY�����"Ox��c�S2�P8�V�@)�|��"O�1����5.g����U�[&�)�"Oxb��55p�k$NE�=����"O���Ex��t�t,T=�F��"Oj�3���0h��h:F
�9 /��r"O�,:tXWY�ƊQ'�1!�"O&D�g��~��A��)�t�0�"O�,�q�W'c`&�{$/�_vډ�U"O4��&�pr=���C�]��9	�"OP�x7 �;#~ܩc�Ҵ���!"O򠃧�Ӊ~�کx�
�|�訪r"OB�ArgO��d��PhP%N4
��B"Os����7 ��ֲq5�AQ#"O��r�-�{�N,Qv���|(bE�@"O�q���:���xE�n�'"Oĥ�&�5M� �II���"O�M��.�#^�u�%I�<�֤��"O^�pd�HVҵ�AH[$�XJE"O2H��(E+
�µ	�ޖS�t1H�"O"��e1/U�-��f&�v��f"O���R �L+�Q������ ms�"O:�7O�<�n�@D#]�q�u�s"O�5���$J�{S��I�N��d"Ot���P�#�j���OV�L"J��"Old��ʺX`dBu�X76b�"O��8qG���h`+� ��6"ODت%fO�e�R(Q�!Q�b�`�"O��)�m�3VJM R�I ��*�"ObTr�+E�W"��h��[o��*�"O�<ᓎ�Z*敓��FF��-H�"O�Ly�d[�g��YC� ����81"O�M��H�`2��:�"=E�I�<��+��?��`ENȸaz��N�<�'"�02��9�C���8�dI��gI�<A��2�#ǪN�@d@y�b`�G�<�@-�4�R��� �0��~�<i�؎7= �􊁐2"U�D�
`�<Q���� �,9�bƖkc@xUE�`�<a�"Y�Fk����b�3a<E����U�<!�̗�h��@Iʸ4�p�F,�S�<ɴ��qX�8C�,R.,� 4��t�<��F���f��d�ʂ3� }H �K�<��Z��<X�%.E�����E�<A��׸%:8�����6��WISM�<1�@��nU�3��� ��֏_r�<�W���/�PD�a�66g�����p�<)�)��>�I0�G�/�x9�Zm�<�EH�3TN�ع���,P��Qa��_M�<!f��q��<�D㍡_��Ey��K�<�g�-����w�V�@�����[|�<� ���g)�~�✻�+�+l8
�Xu"OhQI��K e�>�2�H�@�IH�"Or���+�(Tt���h���(�"O*CG�յSW��#3N�T�v�c�"O��� �&)T6�ja�[$M��"Ot����O0,�����^}��{C"O\�[5���&*dj6.궘"O��cVen���H�����"O:hҥ�4���vG��(�"O�m(d��*�(s�/O��S�"O}�e����FEQ��H "O"�P��S &cD\�2ݟf~u�"O��ن�H�L^J13�.��GN ��"O�q�^�suB�����+M<�eC"Oz�P��X�rF���AN~�(�	�'3T$h��@�DsJ��!�5�@��'��ʓ=j(88!e#�,;�����'ƀ(cqI	p����"�;1na
�'yP�	��
4n�9�f�ū%D��j�'�>��`T`�u��h'L�@�s�'O�}�Gg�,8}�X�F@٥͸��)��<!S��5�@	���/}�1��m�	y���O�6�JC�q�(]k5+ͨԘ]`�'�t2g��<=�e���
�x��'Ct�hӊ�N����@mj��'�l��l^�l��ĈG`Ϸ2|�A�'����"V���mM�&	N���'�L#�Nip���ˆ�v$���'�l�˶"�	��AGN�!���'L�Ypf�M�\�X����� b�'��1:������ �P�y��a�'����'!ۙ#�N����F��l��'�*�pu�E!E`U�����	�'�h@���M�y%��
K��*�'�򴆎�? ���,��
�'�jH"`+�+j5P��˔s:V���'��H�օ5�� Wn�p����'�+3Ö�=�:fɎ�f!>m��'x�-��BV��Õ�/��r�'H`��q�[-n���3�]�/UZu;	�'Z2���I���[��.��1{�'���Kr�A��ȼ0hD�)^�
�'Ud$���A�K�v�y�o����'x�LjE\K�1?��H�ã�j�<��מZ)��bÂW8$QI'���<ɀd�h����M¿�X9�g�V�<�P��N�����P-�|����O�<�Po�8d~%��]�[����DFL�<�vdX-W2eIW��.L����F�<�͞y �
�	,�FAS�K{�<ע���콙�Gѫa��Sb�w�<YW��8]��o�'{_^�DN�<�u���xF@�`�Z�e�4�"rD�<a�e�J	�=��
���8������'k��g�Z䁧�ݒ{� �ȓ&K��'��/7h̹�ԐS�؇ȓ]�*x!�!о3cH6m�4R~|��lc��3f�Fm�ҩ��V?Oځ�ȓ ��0cA�rp2��`�d��ԇ�Z�@��#�xJd
 �ʦ1�ȓn�&�R�
�>>�6uBA��Z�8���*��3/�)����s,4x����O:�j$GˠU��AgΕ�'����~I���e϶|C�i����_?���S�? ���. �{F�'K�e�"O@�k�,l�������DB<�!�"OĈ���/L��5�4�
=Jf�+�"O0�{����v��LyFϘ<���"O���6��,��bf��yi2h�"OF*Յ_�{{�+W��DG��1"O�}��2?&Н��-U����)Q"O����G�?�H��N�!K��;�"O�#��}�Bq�M�y�"OR=�0�R�V��H�K�!u�hHd"O <Bvn&�}sc��~
r���"Ot�yf�Q,IWh�[��>�ް	��	n�O��e��	=�}�%�rb� ��'���ap�Q�k61q�*f�v]��'�8u+��\�����M0i�\)��'���"���7f��)�RMPT~zp��'-t��uIe A)C[�N�줠�'^���p��(T�4nnH��'��4)1���*-�@{�#
?@}��x�'Z��B���x��ta@'�2(|��'����޾$JYs�a�3#�f�2�'��p���xJ%W�Q?�"��'� ��2J@�J��!�/�m1�'�HC�/�
X����_���H�'; ��Ă>: z���a��7�^��
�'�ȵgM�eKJ�qĆ
0����'��E,��+uԌ���@�2N�J	�'��!	&�]�bd���e�� '�t�Y�'X���� �4,�J !K�%�
�'�+W�W�8p�D,wеi�'gld�-�v��E���5��d �'�(��s�ĢA���)Y+E�+�'����fTA�����T
*��L)���%�',Y0�P��l&����;f�VX��)݄ )c#��+l���b9�-�ȓ;�~њ��19B����7O:0��V�,�1V�(G=�I"��2y^����0���0\}��"(�2u��Ն�,Ħ}��闬*ò�b�F�,z�P���[�+$�?i0t�1#ҩW����B��q"N@ f]xy�Uk(&X���D�V� eh�t*�2t�Џ?�DЄȓ=P�A`�Y�x�� [�k�T4�ȓk��Y'�v�lM�ІL	����qK�L�Tɐ��65�BAN�	���ȓ���@-DnVi{m��[M�|�ȓ��%9�΄+s���K R;>��ȓv�\��� &#H���R�ϸa�ȓu��bB�M$�
��'�2̄�"��U�C�2$(��逑7���K������0~z���@�%u��A�ȓjkJM��a
� )��s��V!��~��Z�+Օb�Đ�c+[�WC���nL�5��
$�F�Z��`��U�����F��"Jf��B0&D�>�t��L`L�A��LH��v��	��O�*�  �K� �V@�s��I`H}�ȓ0�:Xa̟�@��Y;�	N��nH�ȓj½�.�� �d��Q�E�ޭ�ȓA��I��^)>���ӧ�(3c��ȓ���7-�x����D>@>���ȓeUtl��
Q�+)��Sm�Iϊ݄ȓ&��9$@_?���Y c�62�@�ȓ;��L�P�7�ʸ�I5G����S�? �������^���.F"+�|$�$"OP4����>MG8��h��8��pQq"O2|�'��J��5�Ԉ��
(� "O�(C�fݔ6>�L+aA�&���Q@*O,����N݀Hcg�jq���'���c�O	y�lA�2L�_��e�'Ռ���c��D1���*PD�C�'L`\��	�&����6z��Y�',��R3i�$�T{��E��'��AVaL-/8��#�����'�H��C{<������#@����'Â��UGZ�ZE����p�0a�'�t�FAȑ8pd�ɴ�w�v��
�'e�ȣ��@}'l��Clw�*5��'�9�SC�U�TA�%�>�H��'t%����6�L�)@�=-��[�'�:�s��!l)��*��V8!Z��Q
�'���V�P=J|�1{�LT��\�
�'al�C �!L��P#��6_�>�2�'O�n�#
�5*7��H��w"O��Җ �|\ȫ�@��8�x�kU"OM�&E>ia�	��o�Fi@c"O*�y�.��5F�2�)W���z"O���RL�Y�����O-ܢl;5"Opl�P�[�t�Kƅ�4U]ja&"Ol��H�b�ȹ�"��:�Fd:�"O�i���ۇQ4�Xe�P�Ck�˦"O.��T
S��Y�1e�$4������Iz�H�i\\8�0��ڋLF0��|P`�+D/Je:�D#� n�!�D�;��Eo+P���ClМs�!��(av�E�c'@dy�Y��K5�!���5Z:����̦9\�hKT%id!��ϓc�P���Ϙ�Jc<��=zV!�d�	+4� '��p�h�GJA�-,!�$Ա�*J!��� �XkF�N!!�䛫&��U@�G��x}��t ˎdG!�H�zd��m%�2isf�8:!�Ď7�Ar�ELh���{���;{;!�_#�,PP��W�fQ�� "!!�dGa_�,��صO�8�'	��V�!�ČL��Y���"R���^B�;�'���B�;2�Y�D�8vQV��'��81i�;HB��@q��&}1�;�'�X�{��ĳ^�8*���X�����'��1x�@J�;,R���c�%�Ҵ"�'u�<���4낰{�A܎J�ч�UD�0SeN:1�����q**q�ȓs��q� ��`2�m9`TI�ȓFG��Dl�BW�hR×�k1�d�ȓ
"��p1��<늙j�.�$�1���
y��g�:J��+ꕷ����ȓuw�|B�1Tv,!��ĲL�V��m�����@�*P"T��C�)����:���`�&�@�|�W�Y8i0v��ȓP�ĸ�ҍ�*c�Je:QP.��ȓ=���s����P��A�Rp�	��u#2,�aK��6IP���ܷarZl��5'TcF��m�P�%@�d��trI��M%P�n���aK�Ot�=��Z���WiЪU���	 �&,�\��o8�H`��� �O�
z���ȓ@ǚ9�7ʚ�=}H�% �_$�5���l:(L��|R׀X	efN��ȓCn��c��s�NL� �{�2���S�? �uH�"�%W�=��IQ.4�P[b"O@�3�Ꮧx��D���&r���B��'��I�,ﴑ�D�'lG���$�P���B�ɐdH���$�~o�!B�-/4�>A���?��`��>Oז�R!�ޗf�!��N"uS���&B)P�NUJ�
�����,�S�O5lm{�E"\7b٨���Lj�t��'	2�S�E�Y�N ��A+E�&�O��H�H�dXg�R�/�q9���P;`d�����~��ԏg�m��k��C22�y	�� `y�L�Y�S�A���Oq����.^�ȹ�E!�Y1 lS5�'r�!���K/�x�Ǒ,K"	#cE�r<�I��HO�>�JP�#
�XՈ�b~yC��$D�|A��W�">娂KҫN���K�J%�D�d��t�]�c�D ��G�
��)�k �Of�M��5��МO�MEgٲDS�y�ȓU�ֱ�0���X��]0��A���F~��5�y��T�5�ȜB#Ҩ�fA��
�t��~"����T�D�x�'c[����'��#=E��FZ���cg1d\� "��yRo�)-y0�S��'LY`5q�-����N�a|"E Tp��#"H{rH����6��?��1O���N��.T�ə�o�7ߎ�sU"OR�J3�I�	�5����*�dC�������h0"�A>�.@a�nD�
�� "O"���A�&��V���p�f��X�8�����)���]#|�֊CTC( ��'@���=^�-�Ŋ J��O<I��'����$�{��̛�Zu��5���G���;3t�!9}�j�sc�\R!��:�,X��''��$��nY,YG���	��	/Ԡ"�/�\���f͇�Z1!�&B��U�
A�G��Q�"Ȫ!���g��H���:�F���ܭJ�|A��3�y�╙)���qW�Ӥ1�f���X���p>q�e����P R��,N�@��1��@���j�B���vAv �oڏ$�l��6Vg����A�7-^�����ł	xd�Q+`�O%r% |�O�J�t��t���a��+F(����D��`m����H*�𥆛�jV4uHзyh���#)��Y��~r��;n�l	z�"�&cR!aĬ(�y�+"R a�=E�h@������d{��hԅ�?�!�y�����IN�31��AV�ɾz����(?���Wx�$��� %�xx�]*4HA�A�̸O1a~B�\%�
$��"�	D����pjG�+�@(R�ێ�y"ɚ+�.�R�ER�Pƀ��'���O MK�$�(�Z�be��)<��KɫKu�|2�"O���
uu��@�pG�`!��OԤ��H%�)ڧ*U���d���S��3��4&��D�ȓK�����78���[U���T� ��ȓbϪ��4��*D����I_��rІȓ<��7��h䘥�%W�f$�d��'?X��f��1�2f��]���'
� U�@1�����7�`���'�0E οjSb�KOKD48P�'zU���mX��SkOBQp���'�n����a"H%�5�!9R���O~	aj,鸧H� R]i'b�a�o�+o�B���%�l�<��!W ���3�O��E�Ɯ!�"�m~r��r�!c
n8���π�LT��ÒcŌ(�����&�O���/ơ(�t�	#f5Z�v傥�����E�`��B�I7n�9c���x@�坶i�"=	@��5��	�K��Z�����B1kԽ[��}�*���Ѓ"O� >� 6hٞR( �RF��{�z���i� =�#
�$S�4@7�o?E��4-���A>�D�a�a�����'M��QP�,(��ɲ��Xu��D�O���҂�(�:Uȕ`&����D�*<$����M�)���i�	-}�|�/ �/��Iʋ�|]���S�I��2ѡ[�+8� ��L�a� ��9��u�؟Rz"xB�����(O^�� 0<�<�գPy&�>h����dF�M�s臃���"O�8�Tj]�aH����	�( j-"4�J��uKF$�m��A�R�V�"~�I�yy��#2'}�I6#��r�B�I�N>`�cȪF�DA���]{����o3��*�)Upʝ�7n�?�=��`Ϊm��A���	 6mk���D8���m]�?��
��t� �bݯ NH���L��0�BH��J`؟<��ȗ]gd�!(��Ȗ�#rc8ʓ"5�)�s�I�Xmv�"q���'Gܤyd/E&&�R���A^�ȓY��tr�Ghzʼ��)�h*�qmZO��ԃ�MN��>�C �O?7�G-8t�q��lJ,�u�OD@�!��F���9�q@I�ke�,��E�0�n�ɌI�I㇁,):��d�I�94d)W"^�t����Ć�<�
���(=� 1�c��aFm����Wd��hr)D6(u8 F�0� �b��: &��	�JR!G�jQ���>�Y�4B7�52V�>M{2�ʎ	� `�靚*�n���>D�����Q<p*�I��̗OᘐC��>�@��:f��"}���[����T�"�1����w�<�}�)ل�}�p�S�I�<�a��\��%ҕ��b��`(QF�@�<�@A�k��Y"H��(���x�fXf�<acj�j�� �%B�~q2�0�b�J�<qW�B�Y���ڃ�n5��c6'j�<��)vRDPҐ�J�=��|� ��e�<1u,.&1lqi�C�4����7�\�<�f>%����+\�#�%���`�<����&6�����NuMV�BSb�`�<q��2gS.��B#��%��e$�v�<��K��h�a)`�#t� ESg(�d�<	��B3�\Ģ��f�R��T.�^�<���?z�0���T`��#�[�<A���g��!���ZY� s�
�U�<����+s/n)�d �,�* FV�<1 �5]��K��Y1�\�� �O�<�F�YrV�C2���rWV��1��_�<'F�9N�`)"B/��<���#�_�<�����3>�7Ō�J���T�<aRgc$i�ץ�(-jh2s�V�<��g�?��&V]����N�Q�<��c�.:���p��	�D;\��E/GL�<�׋G.{���cD�K$.�YF�MM�<��`M{�������7[ ��CO�M�<�K�q���x1J�`�T�)A�v�<富1
LKW�M!i��[���m�<i@l���"���)���Bf�<��f��f�@ܸ�%�T���*��]�<���E�
� #�d�A"��^�<1�Nzb A�ht�p�,�_�<"Ί��V 2�'5@��5��Y�<��-\k�UR2iY�O)tD"���V�<���0"�R��7�P6�����N�<!0��@ʞu����5<�Zp�U�@�<I�b��r*����6��l��D�<Y!l� 3�xp��(���3'&�d�<q�����~7�9%�����I��yB��~��-�+�'-��S��"�y��h�t�A`EL	_fi�2 LKjL܈���s�\���L�(Qx1� �b�3m0D����ܮG��9b�R�m��x�L=D��  $�.�9�L�p��R����c"O��ҍ��&.���C��}� �@���Q@���S�:�<�*�$�>(��mX��Q�6�4B�ɘ ¥RA��3d�ZXY�$�x�C�Ɍ-¾��a�\v�4LaЪ��jC�	�|ThU� �;~�ꍃ���}��B��+FZds�-A�n��90�IE�B䉾�ΰ��J�=}�����P��B�	�[K<<1���&A�- �.��.�˓d���|��ÊY�s��ǂ�Q�DQk�<����/.t�f�<b��ХO�L�<т ;���E, �����D�<��G�= gΙ�$K5%�\A8�A�<����U�<R�C��rW0�Æ�p�<a�S�8\�[�1Q4$I��Z�<	��Y4#�P͊:�М���^[�<��_�zՆ9��o���[�{�<	��Ƹ$�yk��Ȏ��U��p�<�*SE�,ak�w�n��S�F�<"�6W^\32�>k�X��W��u�<q4�g�%�$��:8{`��i�<QЫ�	R�l�a�G��\�fE\a�<Qq@�l�كD[�=! 7�\T�<I�ѯX�fh�4韊j�)PǄy�<1f.��.�d}�Ҏ��<IKT+�q�<��/��*��4�$�.�)6G�o�<9"��8%�s� �!� ���Pf�<��Ҝtp
��Aϋ'-��x�`�<!Ѭ��Md-��?x�,�5EFt�<Y�O�O��1%�!�����D[�<��{��0B����\#j�B�<�1�}���x�MUuo�L���r�<�U�A
l|XR�ʃd�<���E{�<Q�bޮ	�x��ᅘ�U'�Ai�ƞw�<qR��.]�vUI�Ҁ'w��B�k{�<)W��~L��o��N���Q!�Mv�<@�I5!��Q֋՘&��͙��Be�<���x���鑣 o�dya�)�k�<��cJ3D�pI{o���8��Hg�<ɂh�Vt���}s�12H�b�<y�D�'-��*S�];�X�	�^�<Q2)̀y���h"�
9J���#�HF�<yƄ�%��96��J����ƮZh�<9� �6
�"sS�1$N�ңaLf�<Å�yk�  $��:�lܳ�o�c�<��A�.�쌛s�P"W�@�:b�VZ�<��[�Q�İ��vx�Pc�	�<��إϮq�3�W�bQYU��r�<�񁐤T�n,2��^6�*}1d��m�<1�%8U���unU2��sƞM�<A��2���1��OVĹ6VJ�<��l�/6PZ��6iז!��d�%��E�<i�Ïe���si�$e'x)C�A�<	 �0�{ '�t�P�w��x�<�&Y�N����@�:m,��@��C���WAFv��jsoE�
���Y�,ᐯC�3�0�σ��.���1"�L�#�'���X��"	&����Sab�<M��0벣@�PZ���"�1�c�{�85�7"V-n��M�ȓQњu�1D]�3p.��.,\۸����l+�M�+����Δ&����xT���*�$><��OK�L�*I�ȓ�fE���*j�ɀ�� ��1��S�? �}�eM�|�B��Flp�е"O|p��#ܠ�ވs���!�X�h�"O��F��7���CP����d�Y�"O��"�,ހ�&�LnUx"O����1O�q�FEV0#~���@"O�pъ΀u(>�h��NV&�+0"O�mi�K<b�,�WJ�PA���"O��1"E�-�JT��iˆBg\|��"O���CS�to*(��g�@m���P"O���A��L�M�l&\��)t"O�Lc�.	�~��k��&D�*Q�"O8��kE�>�H=C�k��#�4`C"O�Q�Ԉ����]��a
��,!�"O�I��r	�E�Q.s�ڍa�"O^0��j�3�`͙�#8f��|�
�'O6��ԣ��L'�0���B?f�Bc�'V�]2S)�8#��y��a�eh4�B�'�8�% �y�LĒ���#�./D���� B� ������/�@�r`E)D�(Ht��u�Hz!��/�vP%D���Ԇ�򜩱�T��"@�% D�3%G+=0�a)V+<CF�Z��!D���5��@~aQrG�4jV���=D��4�ݐ.����E��L�2��7D����9�A���>*t��	5D�X���K��P�����6�e0��3D�Y�Fغ\�>�y��a���o"D� �w��<mvu��i	����j�<D�����"b��]9�*�iEz�rB�6D���&ɔl�Xah�`D7�6)���7D���0�JIQ!ρ���B�?D�t��b��j9�a�jʽ5��q��=D��D� �$1L����/6�|��<D� J��^$
:��W�LX�p�)>D��GR5A�b���e&�b假=D�����J�Mތ j٠��Q��yRر�Ƶ���ޮr��r�Ǆ�y���/�rE�#c�9h�X����yr(Ϙ�DX2�Ɏ:�n 0g�Z	�y��I��\*�`���.9��,R��Py�X!Kv�|
��}��@&QG�<`F˲Ҧ\"ƠM�%�h�B�|�<��O�
/�	�G�=rs�����}�<q�e��f��i�2`��"�����G�<�NO�2])�,4��uS�-i�<�u
W�G����X�QJS�<��9+XmP�D��d?4ȊkAV�<IG զ���ǉӕ �&I��GW�<�2�"��]�F�H�(D�x���M�<!�,G�%�̻aϝ�~ؚ@p��VI�<Q��C<�����T�B���o�<9q�ڑ!��i�AÄk�p�c3-h�<y&��0�Yl%Z:�İ�Vd�<)2e]O��M�,˦I�n���]�<a�E	6kܸ�DD��^9���#v�<��)B6b�ԧY�N�L�����w�<yc$���%��$űX焐Xv;D������J.B(!bJ��Dذ��d�-D�lKAS�/�������x���:'�(D�d��,�ygl���I�f�jD"D�Z��7
	��r,h�,ik��'D�l��%�l��Ū�)�7L��V�&D��'C�L��B'�
���g+D��2��$j � g���ְ�&D�� `�xvB�L� �B�ED�^[�l�e"O�۔�>�\�ے�9EJ�y�"O��9���l�����c�@��b�"O�e� �J���C!��3tBt���"O�s�7|� �O�0Z��"O��!q��:S��� Ov<���V"O�Rr���;5T��O�D�	�"O����[�Ti�c-�-'��"O8�6��"���I��V�R���q�"O:�㯋�����&�+���f"O���M.����
Q#2�ä"O�I��CsP��IP�P:Zs%��"O&�"������9e2�9�"O���5jЈg�$+O�IjRt˶"O����	J�V)� �\�kd��"O����F޷-l�Qx���m�$�`"OT!C䋌$��1tMϿ'�����"O� �'*�� ��:Q�ͨ�"O ���ݲQ�����,�Zaxdc�"O@A�����D4���ӺP�ڰ"O�)�"�Ź|V��۟wSV0 E"OU�"/�	y\t��e�џgh�0Q"O�-�#Ե��K�ͦ1[.,q�"Ob<�sAJB�Ԕb���9B}Z9�"O��ʷ/�]W ���YY�}Ip"O���O��!��b�f
=�f�1"O�dR&�ƐN�|<��8X���S"OT5�aiS?�d���غo�>��C"O�\hd���7k�}k�'V�X:s"OfM�c��G�f�C�	� �6�1"O��� �.�C� �.K�2��%"O��X\����cą�~"*���+�y"�E ~��u�v̐'s,ҭ���܎�y�D׉<k�@3�̾���%H�5�y��2R2*�S�:A�ᛄ�ؖ�y҉ĸm����8Z��j��<�yRi2ʕ�u,�1-X�S���y�N܂vn�Ҵ�W�>>d�EQ)�yr猢8��(��#8�4���y�/Ǫp����	ɫ8� ��g
�y���D�l9���,Ⱥ��rm���y�(��T��O�.���1��y��:��`V3r��j��B6�yb���n b�a^#��J�����y҄�q��۴FW)�%Mш�y�A/R�W�]3M���!�!�y"ύz v}c��ͼ^�]�%���y�o4���`�"�xkB�U�L��y��h�9�c�B{Fh��C/�y�H��g��ѤւVꄘ%���y2�2��
rbS�Bof��%��y�NՌ�x��c�-j��A���yR��n�.����j�Vt�OG��yWmu��r�D��=w�� �c*�y" 3<����8�j��`)އ�yR�!{Q�|(En�XN�k�E��yo10�z�H�.�x�p-U��y�Һ\��=��o�~���rg���ybʞ#sp���>w�Jd;A(���y2 �,bjP��m�+Y}��[�d���yB�N.�8��G�G>̕���H�y�#��D0�sD�b�$P0@	�y�@JȊTKE�P���r��&�y���+��Y�A�����Y���y
� ����ip��1��'bCHq��"O0�QP�	5�|P"��hmP}SS"O�H+ ������)
�t�~ �`"O�9X�l�H�9�`�K�dz� "O�0��̓p��x2�Bқ]b���"Or)�q���W����#�wf
��v"O>|�G�<���c@A�'6� ��G"O<t��K�Q�`�Iv D�����"O�%����B�OօY�Z���"O���Z"F��פ��89�E�G"O�q�խ��n�Pj�L�lH���"Oޠ/48���m]�o��i�S�۰W�!�D�4�|�t�D�	��*�!�=8�KN+&'(t�bυl��a�'� D���6�Ƹ�2�9\�ʠX�'�����܀Fw���¤ܣVִ�9�'�|�IC�P s�� 2iZ�~f� �'����Sbn&;�G�pb���'��g��?������ǲo9Bc�'��	#��?�e1D�d����'Ɉň��"8pFA�3l�>Q����'*� �īFo��b��@��A��'��}�WL@<L�48!'�@�@���'�("WK�y물��R�8+����'2�)Fb�:q&�%�w"S�D<�=��'nH�DM��\��E-�<�J}*�'30@&C���>�TkT�6���
�'a��
f�t�Q��-�%`
�'��iqgHk&�)z�	ł#�B�C	�'��<�R'����կ�(��'$���`�I�!�gO�~R�S�'������#R���&���sUp��
�'VL�a����P�a����lnԙ	�'��iS���.
�@1(u�/	�bHh	�'�d%i��p�1��ߕ <��'$��8Ea\	�kmK�nd������T�͹e ^2AިX���J+�˗ h�i��=����� U�]�x�Ɗf-����H	P��>%?G���6��(��,:��J��4�$�WXv�b?%����ЊU#ƇUܠ�;��>�F�Z����H��)8��	h_�C��΄IΨ Բi�e:��Ӂv���+@?l�0�{T*��|S�`�DJq>���ʕ�w�^Hb�l��+�F\�!��,���?%>	�G�K�aDͻ$��I�+?���wH��b?5C��D��BW�N"	x���e�>���V:���H�H�`�%��&Yڌ���5�x��i� �����2�:gH�uiT��Ph�&o:�� ��G>��pd��Y�~��!�í�	BC�$��i�Ҕ0��ID#b��3�
��K�����sf���t�>���_�@����?��&'�b�T=�3FҷRK��z����U∙�{��&y�1eŸ1�H��6)y��չGK���U���N Fp&��'�{��O?ɯ;`��*#��(1AP�Z��U��t��>�ɮ�0|"u�,k�n����Nk��h��U[�t9X�c�J|ڄ&�W�x��Ո����D�e W�I�>�a��@�)�'��a�5���F�UC�(x�@5�O�88��:�)�'m��3D�:jJPCt�8c�"m�t�jX�?E�4�;P��iЖa��Z�z��vj��ܽ�?���O�S�V�.VX ��l��e���}rB�#jA�O�O@��E�F	"d[5�PZ��`	K<��J�!����O�2� QC(1+��E���4H��O@�QQ/'��?��<iRH��F�l�dICu樤�3C�禭Z�h-�.m���\sd��Ą0�!��J��4Qb�R,�A1�a�ȓop�	��G;z���ᓃ h���pN�q��2_��m1���`���L���P�'���zD�1h.���S�? �|�&�܂j�\[R�ۚO��A�"O�8�dN��M�c *��h�T(�"OR��A�H�(�J�b`��jВ08�"O�5;%�J�Ww܅+�,�5�.=��"OFP��H1,-(ujƀ%���c"O"����)]_2�+ #��x���"O�����Y������Q%�pmi"O�"������o+���"O��Z(��j ��mƎ��;�"O�eH��8^�T0��ݐ2��|:�"Oxp��o�$��-ۄ̑�B���"O�җb�U�4CK�6N)^��G"OԴ���ǶA$��%���w����"O��*N�FP���ɮtb;�"O�њ�� <�$�!�@P��y��"O�Hp!h�(��s��=)?�Q��"O�b��˺n��x�DMߏR3�K"O�u $Y�!�^�{��O=`*�p9�"OT�K��vì])T΂�u�r"OrA��K�Uռ���N�t�V"O��
����2��]�E�W�*�H	+W*O��;h�;������/'"$

�'ǀ8�WB�6�����-��*�L(x	�'` "g�l7�=�4��7'Ղ���'�D��a� =��ܡ��K�6�S�'�H�QH� �1�Q��D\!�	�'��{��$;����ˑ.@�:	#
�'�4��.ٗjj4sB-�2�f�2�'}��A���rK:�ӑ��+�p�'#�ib�ӌ"jDpf��"q,!j	�'�	� '��u��
U l��'�hY�3hٍdmFUQt�U;��ɱ�'R�*C��Y�А��02�`�c�'%��) ���|�0��
&~�
�'F���طie��pI4)S>�:�'�$��*��qp�@Gf�����(�'��{��i��x6f�yY6\�D�-D���G���uc�=������-D���s��#H�E�cИoݠ���(D�@���3C�ʃ�ϊQGV���9D��;��,"���g�ͤP��C��;D����$��IF�<����U%�ʒ.%D���$���:��޺,:�@�'*"D�x���'$ ]���f�d���!D�A��D�*���
$!nJQ���1D���H� �j�ʃBMڔ���.D��a�ʒ����"E�#%�u*p�?D��C*�	6��,��HE�Q���;vO=D�\���"3>������3G��`�:D��iF� �~�T���a�8R�:D�����9@l .K[$�IEn8D�H�m2R��-	!�|�@�6D�X��N�_m�E!��4?i�|X�""D�@(ǅ�}P���T�	`�Y1�$D�<��ꜰ�����D�m�DdP�'D��!p.Հ?�������!@�&h��9D�\�dR�Kav1PѡL�%�ւ6D�$"��.�����Nۏ'y�}�m3D��E�ݨ��S6˚�,S��`�!2D�x�s S�J���k �����%D�`r����|�Uj&�� �v�$D���*I�?�  �uK߮/�^�!"D�p*3�6:Y�/?g�.�k$ D� ��F� { vd�\�5����:D�� @C���d�|��ʻs�\qP�"O0 !�
�DHfTZ&�.� 8�e"O���s��,C%GT�V�ν��"O��SK��O����R�߲?�ԁg"O ���'վڒd3�R%"�����"O�	�V�����rJݢ�"O���I�eR2�� 0״�I�"O$M�3�ˢ(��*�rT�S�C-�!�3<�q �.T g��A��+Y�!�dҨygX�!,S/9/@9%�2x�!�d�B�~���Ӻ,�[�#��f�!��+gC�X�$H^���8�V!�DO�O`8��bAy�� 0�
!�DH[4�U#㖗NrL�8Tc�>�!�$A<E:T��#O Yl���a��X�!��+{��d� _F\xBG�WV!�d�
m9ر��0e�x��a[�R!�$ƞ2�6�/�|�GäIyLC�I�m��0��'~B �Q�%`C�	����� �?*�b|(G\�4\
C�	��x�Y��a�0�&뜽&ԔB�Ɋ@7T!7gV/Nb�"+�O%@C�3g%v����]��)!À۶~uBC�I�Rb����F ���R�D=
��C�ɛ-Z���D`Pn�H���*.�C䉆lV�M�HN�Km�	&�B��C�	�c� d�v��0K����N��C�9m�t )V�?J0���L��%:PC�I(gb���KDp��"��X�C�	zK��;�.�OX�@�t�U�&B䉫y~�t��˄
@Bz �� ��qw�C�	�.�����)WB��P�	�R��C�	�%�0ѪB�RX�*`�����g�|C�	 8U.�A�l�8¼�v�E�)�pC�ɽIFr$�ӡ�oJ��C���B䉌W���񩋱$Ȕ�z���*n� B��,\�8$��일B:��B�r� B�I�}�H�������䋒��C�I9��h�܀T|Y*w� �܇ȓ����1��H��u����dl|�ȓI��$�̒)IQ�Ԑ�]64G(��OV�=��3	\�u�hi/yK��j�z��B�I%f�::`B;l�Q�l�B�9{k&���zL��0���
M�&B��[g8ܺ`�@8-cv0���-W�HC�	HK �xg��t�@ɨ��S�B�6C�*:\�ңe^�C�)�$%��9�C�I�1���H�$A�uݮ	���ִG6B�	�q��"�Gc���	��1B�	�Z�FmzB��t9�"/6C�	�}��`�Y�o����[d�B�	:D.a"�*��Im~�"� ���C�	6v-���]�"���\Rk�B�\�Ρ�G_t��������B�I}� �TH�ʂt÷�۳6`B�I�+�f<z��RJŌ}"W�ڹ>��C�Ʌ_db�A$����0�A�2j�C䉚Ϯ`RM޿|1
(j� <��B䉰T�����,�S8�(��� .źB�ɲ�B�%�%)��=J��Į_��C�I�|_���I;/ �J���{`C��N�YB�\,4y���**3�C�	��3�� n]vݒEX�3�vC䉞�,�S�ʑ)5������ԫ�nC�)� 腱7O�!b�)QR��%�
�5"O>M�u���-�4	i0��L��-��"OL�СC΀Y�K�k0vX�"F"O�xdB@5�Z��'�і��b�"O�U�0�ܰ�D���}#g"O�#�(�ڔ)�����Hk<��e"O6��� )�����"W�(��g"O�P�b��)=V!	�R�Y(�"O��b4-Z�Ixhv�F0W�l3v"O |�n �[Z��r�>`؆�"OP�ȖC�&���@"�0�fݑ"O�Y���Řw���&�ϜF���Cf*O
��ė�_�0M��&�]�� �'�ް�J�rV�:0�C 
$�8:�'N�A���-�`�O�6�ʈ��'�Z@� �֠	�ѡWeU+n(��'����d�+a%�Q8G�۠v�Yr�'��j1��05�6�g�E-�ZeC�'����Rj �9����{���'Y�a���C�����<�9��'��i�p 
��8���(��B7̝��'��Cp�   ���)��:�8k�'l>�����	� \����>7�\�
�'�}Z��6���9�˅�	+
�'�|�eO�`�	zS)�C��(��'M�Y;�F�k�a����N��z�'�����%S�A9�ݣ!�Q	L����'�,`3F��Y�J@�# �G�l�q�'�� s!Z�<�����V��1��'�U��cE=gt��Q�`��'�n�F�uƔ�bA�"p�!��'�J�x�Eѱm��ِ�]����'��i��F�\P.��DDK(~��Ց�'	ĩȦ�$���ƅ�(����
�'��9�M>^��Y�㡖$YȌb�',JP�PF��J�e�P���b<q
�':��D��(&���6.:|تr
�'O�K��@J.|L�%B̟n_>�+
�'*e��JW BF��b胦e�M�ʓA��ȸ
S�?p�����+hJD8�ȓ5qq��&��?�������b~���R�
 R+ 7:#�H�՘g�x��/�(4��	�1pz�˒����݆ȓ,��@�3c�/1��jq	ڑd�ʌ���`��/F������4N�|��ȓU���%�I.*���#n�Lrم�a�HY
5�P*`�0d��������^��GGCP�@����F��T��=�LV���t.T�R�E�ȓp&"a{��`�¡���V3�z���i��5*S��(�Ε����Z�5��6H�L1�"�ך9y'��C:py����) �Β�/�����dRE��ȓ`�H�p�jg����G��b�*�ȓG�@�`��jTew��:_����ȓ.����U�K%jӪE	b⛳�̇ȓ?���7/@�9G�qz��߇��ȓ{�6%br-M�_�٠���Sp���G�4�S���]���`���,�NĄȓ
���
c�1�Ɛp���r����=B��Q���9=�tp֢W�,�j��ȓR�j�KD���D��܈=`ʰ�ȓ� 9� J�8,P�#(M��|�ȓo:�L1�F��RB�80�����S�? ��a� V�]��?w���*��'=B͙3Wpo���n�{��h���I��e�0��?챘���?��$��?i��?�U��!:(2B����$?i�6�	q:0p��'���([B,J�]�IYT�72��DyԔ8�H�*AN@i�n�X��;�4ha�ᘻ*YD���
!9����폞=rV!����5Y��'sR!2��?Q��O�RN�4W���si�8B;�*�OJ���O���?�� �@Nx�@Uh�����?!���D�|�'<B�B�.O��3��~�";Ѩ��h���@f�,���m*Dj�"�MK��?	���G�D��M�Cm�<���:�#�29����#Jό?�b�'/T�:P*� �lX� k� �rSdq��b���h�4�ņy��Q�CN@*\Y���6�����t�h��d�M8�,)�c)��~	؆Ɇd�̄ӂ9��|@@M��r��!�P(c�x�E�#}BJ!�?��i�t�b�����kO)#����M�D����A��O<���P�,M��/dȼdA���$�j�'@n��O�M���4�ē!���"�O�:k�@�S�#%��%��Ma�����O�����C�c�%�O����Ox��x��P!HH:�D}���y�v�	�h %��<��IԬl<��i���F�X)�`��|�䇥bp�aI�O�X���n��8h���a���J�n��`������Tk6?�R�)]a�@�7œ#I$��c�
 -Y�7-٦]��H���)�<�ݴ ����	I�TA��$Ӥ|�R��F{��$��$� �C�'tN<��	���8�M�i��'?�%�c�O,�ɚj�rEK��+Iql�qԭ�2�<�ɕ	��-�x�:��?����?�A��,��O��W�Xڤ�g�X!���.�6-�`����O)^[XAӤ@�(ɶ��Q��Ki0�V�ɧ]�]R�LIF���T���!�t��@Y"G�J����-b���1!J�Jf^�sĮ�V�(aM<��(ѳd=f��ט�"
TB@*s�U�����JI<���?��}2�5� �a��P�L�Q�����'��"=�L|Zs�_)���q��E���!��5��' �7�ڦ��'�X9�f�x���v�D����V Q����F�(r���%D��D�I!p/fp��럼�	 u��6�
�Xq�4 � [~��S%�)H�2�V&pl�bӍ�#;�L��,�\D����?o� K�=I��ڢ(�!!Z8j�IQ>g�YA,ڷ�����D8z����<��D�����4e�D@	5,��0�_(Mh�\Ȕ#�A��d�OiBw�'�iݡ�|��!ԚW�ʬ�	�0::�t`CAo�'ў�8Mk��K3A\�}G�����<!J���,�M�)O
�p������џ��O����3�i�2m�4��6��Q*5?&�~�J�*�O����4h߈p� �1&������O���[&�K��|�'&����(c�F��g�B�#�b\$��K�IN� (RE8�#�,M&�`f�P4@�ޜA�"T�1"
ݰR�-)�`q�U�R�p$)B �¡���>�I�M�U������� ��0�骝��	�'�"�'~ў���>8%��m��D�DsG��9W,��D{�O6�7-�Y'�,�%�GGR��@���M]�ґg���?y�����O~�j��  ���Sb��R\r+W��F)����@�Q����֯���ćV�&odOh��'�R�#�I)�	��&�rG�nր�&���qO��D#,O��bg_}���ȘB�i�	3�HO��D�Ħ��4��S���U�\x�R*"�q�A����d���O>��#_��\i���O��D�O��d����X07�Z��slM#p��Q�8?X��p�	�rq�G��#ƭ�(���iӚ,���aT�'��/�`�9�+�&y�ZiA�\6���Q���4����M�f_�Q`�+Ї2��;�|Pʛw>,����-!"&�!���^�b����
�=�,O���7��u����?�]c&2���8H?FP��`�[^@a"6$����,�(=3Y9F`ִ=�v���#���	��Mۡ�i�ɧ���O��	4`�6d�`[�9�E�%iV�A��,[0nf����?i���?a��R�D�O���#V�$���?%d��ynφ#'�9`-���(zAS���i!%߂4�ڤ�"�Id,T�`ӎ:&ͪ��M�H�&!ef��)� m�����m�8��ȟ`��ӑ�߆f�A�M<��C͖Q�^u�KT�<�(%!�E����I��M[V�x��'#��͝;�,50eKΜSA�YY�E6 ����O�O��C�e�E":�l�sC���hÛF�dӊ�Or���O��^ l  �)�];eȦ�jr��V̓d�*]1�T8\����'���
�Rɟ����:���?Y���c��
�EξҘɠG�Ө`J�#a=�O�O2���� �,���C���-�"C}�I�MS�i���3�̝��4�?��4<~\�G�>O'�q�t��yF ��'$���I���'`R#�#y'ޜ�g�iP����M���P�V�������]��|��Ӭ��_���:���3�V��ïY�,�ti@J%���RW�����\ᶂM�vր�`��D,~L�2��YB$���&��OLll=�~�L� REt4�S�I��ӗ�ƚ�~b�'����?��'.��33��1;����e��k�r43��� ��|z���z�7Ȑ���T@9���8�i��'b�'��'(�I�mQ( 0  �Ru��cƭ҆���"O���`G��_��M($lӀ5��H�"O U�"�.�� ����! ���5"O��
qB�bԌ�z�C�7ɠ"O�qP&�%^�j�ذ儼�\��"Oh���3Yު�� �N�趤�y�A�
A�}�D*��(���&����y�@H_�ִBeP�!�N���C@:�yƕN�̙{�o^�f֌�����y��C^rQ�&�&H�ӢB�y� =
�X����B*o��a�/թ�y2���L��@�҈iwb�x*M��yB��?�쵱aJ��ftb(�(ܹ�y2&C	�:��r䚩U҆l#�Z��ybj��t%c�GK�e86��A����y�'��/U&a�"D-3��ۀ��/�yb�R�w$Q�v�׽(� IR�K��y��Ŋ����߁ti`g㚄�yb�K�d����DS��u�!���y2� ��R��7���W��a1�@��yBe^������Q^����Q�yB��!]���
7��E����ʌ'�y�{�PiY��ݯE�t�H7���y�I�@�<���!��C��-y�O[�y2��0t��ƙC�E���4�y� кR�(�h��'r	�|��#���y��)�`Y�@�=o���[�X��y�H��V$9@���=cg�|��$�y�E�20$ȥhI�*4P��tl�-�y��G�d��N�!���7����O��dݪv�"���4�?y���M�UEc8�9b�n����	��0XEBMU�@���'*B�_Z���fI׾*��ݪ�DK(b<�ـ��Z1s���d���>�*����/�|9a��$�?F���U�
��Y�Y6���xCR�
����R�<�4P �oG�7F���C
]h��O���s�'u�.1�dl��uE���m�M�A��%Ӣ ��d�O��"|:ٴ� ��A�\�^x+A��B% 8��'�剂�HOh���ǦE˗�L�yK��Pg��s�D�� )��@�ɭ�M�3cŇs_�6�'���'m�T�N���ivDL��cJk�<�HS���X��cg�O��EOOq�yӃ۶�HPG��ѺSC�����Ih�� "�h�L�^� 0Pg�.\z�i�S��;�g&˼a�mA,r��h��J�(���?�2����O�B�j��̱C�Px�e
h�xK�O��7�'7T6����N�s�U�v�(�p�Q7�8X���O��-lO�hX��uE�!J2fK�L+v�i��OhU�咟L�I��M�ñi��'�.��>��ްo�"=[u�%:Eq����,�� �����Q՟T��蟬�I">E󎊡q�,{��ېc�U�`�۔,��D�ƨMԾ	�`Չ3�Ɉ�ӟ����S'����3��>����/y⽳�h�-��P��+��V�\(+����9�I�3��P)����8�l	�4��)Rt{S�i��g�-!:��CJ�<���MSHw�l�8�)-�%�%�q?Y���3�t$@���k.�5���,@�ɵ�M��i�'0 �r�O��	�HSr�4�D�.^��r�ñ$~`�p ϐ�HP��ğ���͟�Y\w�"�'�rB�$z�1�[)iN�����]�����+l����匔3<��u�֮�\�'��lp��T���]9�I�\ ���_enH1��!_MA*G�_��bFF
��S6�?�ē$
�oZM����I�B�h�p�'e~U���er�'1"�'��O��L>�jm�@�ӕX��<���[���ɷ�HOBc?%�6c��(8d���+�`���'}2�tӾ�n�|y�b��\7�O��r���E��v�~����לE��(F�?1҄خ�?����?�S6my�FH��7���pnH�~� � ��\ GE���8Q�Q
X��Dy2�֓���DGB�/�\Q�R�_�ot���`��>8>DU$��tO:�2�J�84fQ�pDԮ��'7bQ
��s@��K,�dC]�2���#Q�%Q������(6��$�h:B��t�O0f�0��D���@�A�^��b��{��i>9�ܴy(L`�u��k-0�96�G.b��%J��V��4�m����	r��Fح8��'w����DC�@H��S�A$R��(a����)���Cv��3.�l�Ö;A��ź�%W�_"� c!g��%�ՄL��SM���6y�y�C�kw~I!Dd�%q�I����2���JvA�j]-gb(֨%6�	�V�D����YKd�~J��DkC8g����M%y�����$[*��	͟��r���h�h!JBJ��2��q��K:%�Q�\�ɩ�Ms��i��'�Ό�eXX�bo������Uf� ��L�	D�	^X�0�� 	  �H���@�>I��d!�x�D�ݼy�d��%�A�L$8�x�I)�Msf�i��'�������D 6  �~���?D�LJ������6�*P�=D��{q�Ydv�4견;�Fu$�=D��/)N�����$E1/)=��"ON#���7g��q�R 8�r�D"O�p�: ��
�B���c�"O��V�Tt�h��&�ثF� �������8[B&ö�i�2�O��
N0��oZ(��u�3G_���p�sϖ�!�������? ��;	�,�P!�D3?� ���aS4�p
�)���0,l�)a� E��y��H�:>�'~:ܺU�\�U�0J��&5#� ȕE�T^Ɖ�S%�"V>�K���qGR��t��g*��#�:����R�'qT�n�H�Ǉ6n�
1tᕠp3V����D�O��O��$�O��Y�&mQD8hH�y��C�9?�h3ғ�?�p�i
7M�O~�m�eÌ����s�a�;�@\��oܧ*8���'�r�'���v�gr�'j2�'Kk, �L�b�����P�2=�4ʉk��$��	��.\���^(X'J��V�MZ�4�O΄7m�,]��� S��Cfix�2D0y���*aCSl�u�G,A�I�Ek�?0���՟��p�H���be�`�mh�-G�p�Jrf�� ��7�[{y��V�?�}�	ß�m�,<f�i*��J0�T�c�~1�5�*�O��K��'y��!-K#vm���,PD �'g2s�0�nZK�	�?u��G}d�%1�\��g/՚zA����B@���T�AT�@�d�OJ���O`����?���?��^�;d��0��k��Ek��G�X��(* F�	>��h�u,Z/"+���DD��Ń��2$JsM�n|�2\~,���)C*Q�<�� J\�'�Hq�˕ͦU�%B;[NZE�M���?�i�66M�O*ʓ�?a�}�Y(r��!W��j�tH���Z���'(a{`�Tޜ�����t:Y� E�	 ��O�<������'�� * �x�M�I���c��[|�� ��{�"�P�^��?9��Y���3��?��[0�\�VL�G��4�lS�'X⤂q�R�y���f�$d�XA`�7#r���j�'C��&�٬Sq�� 3��<��P*!��e�p)t�A�a�q�9;�F��QNXiCt�+��0�'T�I�pkB�c#��9ZL^`�#L]�W���IٟP�IT�S�'t�(|Q��8	��u�c��+�|�Fy6��?���K�f*������>-�]۷�"�(��гi��� LRbȑܴ�?1���	�`i6�"`�L�'�J-�����H�}�����������o�D�R�2!x��
��� �$/y��;+NBd��ϐ�$x����X��ēq;*���k���Xh
��l$��#���h���"�i��� �t�!Kۍj�T��0F���#b�x!�?	Q�i2�����|j3␕h,%;1��b썰��Z��?!˓P1p����8t�t�ء,�5=z0	��i>�kٴz��&�x2]�b%"&�֞~��Y�`�
&E��mZ�0�I🌐�d�da�������̟��/�����6S�	ل����Z�i�6��H��W\��(���_s�t�OC������?yg�D����'V%[��D�@ 
��n��B��C�bY,x]�� ��D�2��!�O��M�qHkލhU��)\$���Ϫ-�A�s�Ȉdܛ��<�7����>���O�7M��{GB$H�&B�r N���~C6���hO�> hS�s��}��gR���ҵ#��d���M3�i��'��T�O��I�+e� � ΍�u���V�B�0��IJ؟ ��    �`4x@'�-w����d�YR8m���?��j �rD,�#sn�B̇x�2���ݓ��D�O�n	�M[N>����u7�!�����+.��@�,в.s����O�e3>��D�O,��O�$���?�ش;O����J��E���gn߳(�zy�pb�I�b8"g���W����K��;N�����"#�!�����@,+ਂ4.q+S%���1#	@/6��pACR?�)��$I�{N
I(��۶�0d�5�X(�����C����I1�M�Q �~�'�"P��3V����D��c�7'fȨ��?�hO?��*Q�N�j��Y�Z0�CR ײ8_�]��4W=�&�|�H��S��TU��`c�-U��c�Y0̒��Y^�����0�	�P�ɛ+J��	ן��I�?�!��&ۧz�7l�z����%�|ĚVcݖp��Ȃ�%B�*ʓ8�rP�e�C��Er�Ɖ:h���� g�}�D��2.t��-?$c��,ݷ~��[��x�KY:�?��4*����4�P-Z�^9�ҀC-��4��e8��O���/��|rģőhB��Y� 7����"�z?`�	_���-���A��ma1�E���~�lӢ�l�py���^g�6��O���~
B�/i�H h�IسA-��%.Q� �`����'���'�1����YϠ�A�O��x �y���ܠ �V�	z���--|�>�!�j��(O�$	�E��;��!��6K�>5 #��bT�-����d�0ٝXÔ�$"V$k�S�D�$k�rbf��'>Mo��u��q�E�0}*�
/�<�o���u7��On��QD_Fi���ty�A�)��	y����-q�.�n�ݦ�� ���%�#�V���	�2E���a磇�M���?i(�8�F �O��DnӖ]@���q�b)#U�\�Ӧ )�j�
�0ƪ�*h ����G`�|�i�	E��-�OA�t��X�d<���V�ágj��ĺi�Z�!���O����j�5���Bd��,W����-w����Ţb�n��H\�<�p�	��Y�A��O��o����O�>7피d��̰�Qh�x�A;`�$�O���"�S���A�6�_;	4��8$N�!����	��Mk�i��'������e��rwD�V�G9~~I�c��`��u؞dѲ   ��M3�������c���	0ʑ�]��Qu�
��~�'��Q���)�I2�Ո� �o��P!$)�,g-Q�4��43��&�|�ٚXc��C!cX�����@��;���Q>L�	͟P�Ǯج���I��,�	�|{]wlR�i� �OA�\C8�[���tf����kș[��P���8B`|�b��׿|�"���`��G�:��'�ep惛��I�d� ����!�/8gp��0l�=8/
Y��}��� S��yx�N�d�&�	�x��1�eM�u������1� �.i���ğ�O<���?�O*Af��GY���Ԍ��Ȧ�	��HO���8���{�C4K�� �4�� p0��ָi�X6�3�����<����,�� ��i��M��0�O�!^m��q���?����?a��/�� ���?Q��^%^��q�E	)���A�q<��y�B8(��!�U &Ēdx4�A3B��#QI�i�'԰-�!��Bt�B�lT� hmA%���1��$F�9Ee
q�V�K��%*
�y�Gե�?�u�*+��l2 O�*�y� ��ޡ2 �x"�'��A������3kK"8s�� |+pCQ�n����$+ғ6B��6�.\����"I�7���^���k�2ʓ KT�ſi�2�'���0�A��ER�H���ӧY9��Y`pkQ'�?	��?L�0�����^;f�*����$*�b���\�h�9��D�z��zS� }ӌ]Ey2H��R|օ���H�~ 3�" E�F���FԠ �z8`t �"���`�m�(�^�{.	�ri�O��b��'��6�X_��Ԧ���/^8'��!�Ɇ/�b���E��?Q�ʟnc�h;s`	�H�!ѣ�)1ٔ�ɡ�<}B�i>ur޴��i5��y�+�26�(� ���pĆ��N���Iɟ$�8�>� �N   ��'̘�;��U3ʈ�u��}��9C�'Ud�`Cl�+o<����@�d�|��'Z<b�A�!	��0d �s��]2�'!^�a�(̤>є�F,<ز�"�'�����F�1�N���g��$�0�j�'�JDr�Ȃ;���snb�k�'H]� �)Vd�S��h�� �'�Zxz!��(�LQ��&�"^R~���'�̱3��_�d[����_�di�'Q޸���b�Z�s�*��a�d��'>�*��S��(%�玷Qƽ��'?��	����a�` �Y,�D)�'�P�fT(I�ļxe%]P��q�
�'�F9��Ğ�[&,%K5��:��	�'ӌi�V,RZ:}&�MM�'*�`�&c�����ub�f� ���� j���"
0R��� JB35-|��t"O|T��cW=f����V2���%"O�IBPl��p``��V��/(�4�"O�Å¤0�9��O�c���S"O���gK�f�r�!w�SJ�l��"O� v@]xw氋�KO�xKA۰"O�LI5��/4욣�_>h+�u)�"OHA�"� ^���7e�/*`�@"O y��K�&���CÉ(�x�D"O�hs�*�8��F�T�P�R!��"O2a����?&�0	S��,IԲ5�`"O~\@VBȳa��H�G�ţ(]0	V"OR��D!G>J����ۡAQ��F"O�@p���E�, ���H�bqB�"Oz8��W.$�C0l�1W�V�ʒ�͇�M����Mk%�ilYZңq����OL���O������BeT�*�"��a ];^tpN."��(t�2ƭ|�'Hk��q�Gß�/�\��B�}����N>}���XZ�aQ��Ԛy}N��S,^����-�6a8tG�ɼ�u�1\� D�",�$s����"�<^�2o�<�f��͟�>�$�ON6\�y���s�\�3`�5+E>g��e%� ������'oq�4tB�CG�-������
.�6����O�D�æ�)ٴ�?鐿i���O)��^?%���+(D5�V䈨g����c�SCP�H!�^��?A���?��$ �N�O0��O��b��M�W�W){||��5�4MKj�q��هH��5����-g�6�nZ����<12�_�=Y�T8���gq�������I�I�e�KȲ=�P���G�,$��b�)E������>Q���BԂ��B rV|#5F8!�a�I�MKf�x��'$B�$Tu�>���h�{B��	P⛞#Q���`<?J|��	&@u�`�iE��T��wO��'?h6M@ܦ��'d �"P�g� ��{��Iv;����fHQL��b^џ��ɡj:���	ʟ��I�8�T���qq�Q���^"�����hx��(�?iH`�q�'g���o]�D�^|�%㊟s���R4�Y:x�i����q.��v��"?���C��+ݴޛ��i��	Y#�_�j���c�|��ʳk�<!�����O��醕2���PW�yK��B`Aۚ�Px��I�Q�6 P�(�`D{�� ���t�ka���tz��e�(�?����=�V7�F$qv0�Y*'˒�u�?
yn�I���j�'i�h\��aK9qx6�;�׳�P0�,�����,N�x�yl1JY�a�dM��ēK�` ���ҁO!>����R�f����"U����T���n�|��S�F�U��p��G�m���xK���?���0m�O�O���YQ���_�:����P4;n��x�{R�'�ay����Bve3S/���y�`P:	��Dzb�'D�7��Ħ�'�`S��D3pY|QA%��_�a_"^��v�'���'H�X��,�d��'C��'�k,�"9��U�(2@�u�C'7b��3 ��O$: ���I��4:��b�T�O{��s�ω��?�b���!I�\{�o��&��\*�lD�Pj����P�v�iiJ1 �F`�����.�S�r(NE��w��lP�  q*���׭R�j`q��֦Ui-Oh��t��u7����?Zc�rT���>pRv�!��6D�.T g,"$��K��B)�ν{��?�.E�v ��h�	�Mc�i�ɧ���O��	!j� ��7�H$4*|j7KN�N�$EZp����?����?1�����d�O|�D��[+�]��P;����B�?/(d�s`"��wh��KW�xD�m�х�#0Gz� d��vL��eb ��Ŋ�6,��Ya��8u&�!��_Xݲ�H�$-|E��� ��I�N<��Z�]��y7����5��a�28����	�M���x"�'R��dN�9f�D��i4R�D�t`�G9铧�O^O�u�QA�;|ɰs���yԎ��2Şv�$�M/�M�L>����?����8�  �`8��l�Aa�ۧ_>��냏�iI�%�r�%�Z��}��K؂H[��J��T�KZP<��
� @�0�v	�8J��gj�����&�O$�lډ�M���ud�P�Y���l��thɵ�~"�'��O1���n�489@(T�F���pҍ��_����I�MK��I�~4�����:&R(b"љG�
uP+O0TRϏ�gg���O�'�H����M���ѯ~}z���V����c*�5?�򆘿~~F��g-��B���N]5;��s��a�����q~��X5|�Q�t}¦��(I���z�B4"$
K���P� V�0��v>��иgy�1��%],]�� �F�>��	���IU��'��O�ȱ
3f�,/��c�f2r<�M����bx��2&G�@>�t��@U�<�"�)Gj4#�Q�����MK�i��'���7x�A�@E4h���r�A_�d��`��؟p�	�f�V�c-�ß��I�@�ɥ`��'$�f��S�[�g0���·8b�C�.&��EC��Q�>�8�*ן��	ס(�JPh'W����\��T��O_'w�Z�u	�� zGI���=[G�(P��Q��?�z7�ڗf���#�w��y��7g(�3�6ej���H�|y�HϜ�?��;��'@�%g��oZ�Q4�٣v���"�����A� �|B�I�tP�`�`��D�0��\@*D��~}�Hw�2�O�)��Z�4ԠS��_�htziSa���������'�*aC��?a���?������OZ��V�=�p@p�F�$&�Q
��Ð��2��6Hiv�KQ�Y=T�>���fW14/��w剸If�	J`jߝ^a�����KP$�$dG08��]��g�+lnh�E�-z!��ʐ�ӕfd`�I<��!�¦5�4�W19��n�"Ǵ�"�`E3��/;��OH�D5�韂H�L>>!�YI� U?/&}���Oԣ?A�}��/A��jp"J���(z�k-��	=�M��i��'�"�'���1_Lj�  �%>7�_���������/�v(3u��%����O���7�R��Q/	j��9��.R:w�qO���B��q
ٴ���|�^w��$`�JK�*^��b�ZB�&��s��O���K"L�{WK�O��D�O��DYպ����M�݃M�䒒��-�|:G�&��qg���/�h,ˢK	�c�2�	�O�0�Q����7�B�1�K�M!�`�s�@$[�6��@͙������CO=oNTR��K�Ԡ��*	pTp"�px��ɭ%�0�����l�P���Yb����������M3R�x��' �Q�� �@�rѢ	��&��[�%���9���O�6.)�H9"	>^�P� k+v�0)�4$S���|"�O���|��iB��� ����#��0g��R�m�4cK��h�nx�p%o�h�i>���ey��W�,��CA��>Rxf����9 ��ŋ�}��'���'0��@��'>�'~�����["Px�v*�(n����s��J�x��F
�@)�U	�4(���@��(O�t�U,J�H� �����4Z���8�HWT[N�k"k��S6q;6	��#���X&�Z&ܦyH���n�ɵM"����]�<E��@�~��`f��Z@|�׎�t�������Q�S�ă\nVjuiEvn���D!]�i<�?Y��䟆vǠ*�ΰ32���hC%n����@�4�䓧?)���X�Z�� @�?r	Aa�Y�]�Q�X�<��$�����`�?�Of0� �7$�
ai�F�?�Z�Z�$��HO��|�PEi"�Ύ�v����~��h�f�l�^�Iٟ��	O≛�hp  �"`�\��ɟ��Id�S���O y�`���72n�)��9 Kآ?���d�n��!���ǣ�H87k	9|��ئ!Aش�䓂?I���ē]�t=� @�?��Av�J8��@�Ms�@Cd��6<�ĠWM�<Dx%+�7�z-�eGy}�Ey���4�|�I&)A�Ψ��JA�D���N1��91��>v�h���,�X���3 #�'.����UY��f.�	f�@U�&a�"2�P@V,$�D����ӟD�?�O�Oh]; ��hۑȆ�h�-�b�>!��4�r�lZ�M�ڴR����&텗!�ĩ1a�I8���O����O��O�c�x�0�   �f��v��� w>�3��R�RC�I����ۧ�ͣWX�iC���P�JC�	�~v x3`̚�&̱���T�tC�ɖMw���4��N�YAM24`nC�Ɋ ��M�WC��d	DqAAC�M�B�ɊB�>�PD�
�Z���oɈ.�B�	/D��H�E�L�f��y�t&ȩ{�XC�'rW�<�B��6�ș�ѪJ�]�B�)� ��� �_�D�R�3t���"_��@"O
���'#v	��c�<K�Z7"OH�!ro�8}I$���cW�K<m��"O<y�	Y�q��-���ՀE-4�b"Ob@c ͡mpT�A��׭� ��"Or��p`��aQ��`�6>�����"O�0�"o]�~������Z�7����"O������4
}X�gd��sR�"O4�����<)�mY�M;>�$�6"OFL��kJ +pᡅ��7`�����"O=(F̞8S��	���}��mQb"O��s��&o,4$�u��:ZF\�"O`Ȼ�+�#FUV�U!2���"O@��ł��><�Y;�V:�=shq�ȓ*l��,ۄ$�D4dN8&�����b*�%��)L�k�DKt(��;��1��7;lh���Z�w7��*"�0���ȓ{�b��%81n���
+�t���R��H[v��\ȸp�1�&�l�ȓB8a��K��pdȊ�l���y�ȓ$lY�Q�o@~�B¦Q��Q�ȓv��mB��q �
���aL&=�ȓ$�V܃3Y�[�qb��ΒR����	��(�+@	F���dX:0"6�ȓ���M]�8�P�Vn�Vh@H�ȓg\�򍉁R"c��]HH��C�ΐ;��:e?�ʴA?o����9WeH�	�b�x�ICK/B⎠�ȓQ���#$E3� �#��-V�b�ȓe&�q@w ���5���)@� ��`�.�!I�'atm*��0�V�� z�D��#��?w�H�)Kj��ȓ.&�X6,�at(��T	�2Lp�ȓ`4|��$��d;$��Q�C���х�?w:�:���o�����&j-"1�ȓEf�Mh���k�>��"� �K�(��`Fу���
��\8��٨&GrA���A��喥�P���m['KqRdE|�'T����y���?�nZ7a�2��w,�02�j�8���G#Nt����|<����?q��a��=���'��u��	�EM��Zu�^!
���؆g��I6`����+/�coV�'�­��AΥ~���K;@@����4V���pc�X@i��ٍ[ZT��ƭ�&��1�|��}����<�K?���-�
�Y��˒�L��1 �nU�?������67^����(�j}�`�e�QZ��=�IiybF7��?���i��:�&�����K��0�,Y��M�C"��j�r��aBߦ=�	ϟ�	�?���Q��m�Q��mQ��βQD�ɸ��
s�����-�:�;S (��̓�q�.٨����Ū|^w��u�7ၪ2� �w	�;+i�qP�O�]H�o�0|ޜ�``	�M��m�� [�u���M������X�B@�=~�yk��L,UFh�'����:e��)�V��-�S�R�҄�m��.�Y�瓞"���'p��'����,V
r��ڣ�֕J����'M$�k�O��$�٦%��4���u�M�~E�բ��,��,b6kLـ�D�O��d�"c�-�O���Ov���y��l �A�X�)��#�,��U����ƄL�-����H�"��1Y�O��2O%B��}{�n�t��uSC#��p�Q"u�пL�(���J�,>L1L|�r�$Ԩ2Q�4����<�½3�.I�vlB��ڴ�?�G P8�?野-�Y�(�	�Y2A�Ԉoz��)�B�J�v�2a���4G{��	��	��ᒦ���B�@Ձ�+�J���򦙫�4��MҸ�����DW-j$� Ϻș4׹cl�x �H�u3@�d�O����OV���?���?���&�@�+G�͖ �D �̙I_�Y#BI��F��(qJMy�H� ���-�
�Fy�M4t��|�Q�BT�a� ^ȴ�
�LS�VG��␤]�"���k�1�4�i�U�:'Opa��i�5�'��-G!ks��4%��@)���O�&�H��ϟD�?�SF������Ԛ,A@兏@#6�'X�#=1��dG�cdp��&E�S���􉸭M3b�in�I`�Q�ڴ�?����M;�&�5�����X�eh��CƔ�Szb�ܿ0R�'�&E���͢EV9'(��&�S��)ϚB�� `���+D0�"7n`� X��$�C�x��
�6�8S�i�p��8�˾L�8u�W�Kz�ȑD��G \X���\�H�1OZP�w�'�6�Iw�� HM�e)΂c��{����7�v�A���ן�8�ɏr�Ӻ���i�?g^�}���ۛD� ʢ� �qOp�=ͧ-��+��֭3+�l��ҏ�\��p2!\��k���8�M���?y-�"Q@��O�7��8��WCU���a��F�be�';J1V�~|�Mk$B;`W*,��Жe�(m��Q>]�;~��y�fG��8�<��|�'kT�5& *�(���^��2�ː�Uu��P���Y�瓠t���Ԥ�o�ڐ9��
�>&6�'$�� �M�Wn3�$��R�:�*��v�@�	��4"�: ���?���hO�U�H���	5;�6�s�o�!l���<1��*���Ka��O���<�Vщwh��H8���|�(�������<���   �ܝw��(���O��=E��h��xk��M���9�@���~B�'�~7�ئ5%�����?1�'��0��N��*�^A��I�@��ԣ�'�aBO՟P   �-\M�'	��'�.6!��'��@�!-\�d�/v�"xz � E��5"0��&��bfν1@����׸2W<�����!�" ʡ+1�A��5FhX�� �N��jp� $�b���Ji�,�G�Y�1N'� I0o�OT�+7)	-VB,SD���
�H�X�N��p���'�`�	֟D�?�Oe`%�&
44���Wǅ%��MbSf4��HO��H��&|ܡ[��UKJxs��O�im��M�I>���?�K<铋�* .  ���<<���z���p&=0ak�z�\ct�Kr���TA  KR �>B1�ܴ~KX�	�(O���s��<;��ęZ����$�+_�� ��O��$1<O�8�90P�HD��%D.���8	���=��{o�F�g�z�OB�)fݑ��	8s��в�E�h7�!pP���?Y����	�?Q��?���g?�.�Ot7ӭ;��*�D�G	ȴc_-iV�m��g�7C�9���+X<�w��?�j��WE�O\T�PL=|��Qa��W&���X.A�N���f�X&��/?�S�'S���Іr��g}��`�aX�@��|�"�I
2��'�6z�(MR1�x"�'x�֝R}���і-]۞Yp�ڇ�Px�i���#@�94\E�ď��5�]�s*�զ�b�4���|�'��dQ�Z�0��㪈�D�,A��F�<�6��Bc�.���$�O��d�O�i���O�D�O4�x�e���Z`Gb�*kb���	 �(����C <,��q m��T���@y�Q��d�,k�xir?H@���Q-�!��=�d,��ex��4��)���3�(?y����U�ʧ�ē�RA�IC�� 
�0�g�46��A`g��{���B%�Ы���?�������I��Et����T�L�٢��1� D�	�FN�i����U����JMp�I�MG�i�'y"�'^�'Y�i�� ��'�,8�g�޷p����Dm	5t%\iJ��fݙ�WM8N��ٵ��[�Dp�m �1��<�/�#w1zx��$DmÂ�Ye���6�U��T�t!�&I��N a�ޟ��)+�-�X���'6 ��`��&�5�I{Ӫ��f��)7)�`�ќT���8��J�(�?E��(,��-X��5��	��^Uz�O(˓P��>��ڴoY���i�t:p,K������/]��'��ӄ/yӄ���O��'mHuY���?1�4A��t@S�B�Q�{1�w��!��p+����7ʵa���$m0	/��'��I�:���``��9?�ً�f�Ox6m�-'=���P���L�� �v�F�\cH�!����Ȏ3ls�Q��G�)�g�Ol�mڞ�M������&F3<�:4蒮Ϙc��4�tf�!�~��'J�IN��򩜩<��L�G��T�ݪ%�)�Q��[�4Qi�F�|�r}r��� �uc �=#���M�=`�,2����	�a)�̛� ��t�����ɧ�u��'M�F�Σ_5���S���Md��R!��)�J���ű=f>)�����'>؈�A���p`ݨ]7�'r]�#@��}{J$�V덿t�u�P<
p$��W�ĥX� �K�F����)�$	@�Ū S �p�̓s���z��R&H�Q3�P�8ih��'�n0����?���x��'�RY� ��
8!����
�zv��*j#�l�����X�Yق�O2.�.�����@2�e�u�xӸ�mZy�	�?%�Siy���=p��Yq0��aִ��
�&��"b�+�b�'�R�'N��s@�'6R�'Ķ|j�b��5�K�i�D�ԁcB: �m��K8&����m�8���=�(O����E��VM戾��A0��E�&����h��tTT�͟35�*яQ�	�tH2��Ѷ	�mE%U��Q�F�5�>ԙ"�3ޝR�,:���O6�;��<�iݝ�'d��u��瘪}h�Yѡ�S�a�~���IP�'!��Y����Q�:8���A� qj�'��6�K��ї'� $K�mӨ���O�|���@ ЪWL,W�
u.����N���'DB&��J��S�~M9"�Qr�L�W &~�3�BY�hd�!#QKh��,C5&1�|��ǠԟxX�:�-^�_߶��f@]�zEj@�1`�4[J���D[�&��sB�w���֒x򧄖�?��i&��6M#*a�ƋC��LR����8Ԉ��`�S�����z_ĸxJ�
%�.哣o
铊hO��@٦��ش�M{�������8 �hT�w�m��O��$6�D+���V��   �a;�C,25"� �R/K�P��'�t8q �1r��E���<�k�'��Ѻ4B�?C*��׮ה!ަe��'@(��GS�@H  -w���'/P���nX<s��y��I��+̲ ��'�� @�l�,Z-�A�,�%r �I��'��+����\��ƃʿx�<��'�R���3��36(�?=~����'A���śS�V�����;��M�'6f�Aj�m������\�<��
�'��$rt��Y���z��UY/�
�'5�y�t)Gd8���,��J��1
�'�$U���@�W0�!X�G1O-h���''����JR�a��?���'�x��1�ܘ8HU����1'�J�'/Δ�W
�> �� �&!6���'O���3Ȕ�-��\Y�p�a1�'�L����i���!�ԪqG����'�q�i�J��Y��)��khv�K�'_6q�D`��@����Z�a�&	��'��5g�Kl׼�լA�X�:k�'�0�JC��5?][��^�T�ntS�'�X�� 1�d�`]}� 8�'��I��a��M��!����B�����'Lݲ��5\H@���x�	�'��q#�*�	.SLQ	�ʚ�̔��'���I&ϋ�+�R�Z2��#�����y�!�)@����ǳ'�f��B�y�L?]Y�}q��9W5�u �B��y��p*5����*b�]��D*�y򮀇7�Ա�v��[H�PD�W/�y��,]�̳I�#*����僶�yb���$��oIU3nE��-	)�yDG7h�p�bALI�����7�ت�yB��%<��ِb�Dj4x{���y�*��E>X�J�ˎ�vo���% W��y��� ��ecU�v�3�.��y��S'l�Ա�R��o`%Z����y�*E9^�JL����5x6$pjĬJ��y��!�,Y��^؜(�f@F��y�HY�[����E�?� �
KZ�y
� pE���5UH�)IE��:��દ"O`up���M�	ʒ(Č8�t�X�"OZPB$��.��0���L�9���)�"O��	���, �y��#&���@"O��Q�^�,�nE��NQ�~��A�"O�HSU��/L�Pt�4gܶ5��=h�"O��2��u��Y�4��p[�"O�ń�o�N9!��� g��\Z2"O��FL	�}��%�5�rϔ���"O���À١^ټ����U�Rq"O�Xpe��\�! A��X�6��"Os���%X�vQH���zo��s�"O�H�q.�䪅F�cA����"O�m�!A�%97KQ:+4f�B����yrȒ�$m��o�ʆ��VC��"�!��bS��;��	��~�iUc_�g,!�� �q��f@IIX���AF�2?!�DW�7�h����'WʄY��L�b�!�$��Yͦ=�r-IV�ع���65�!��O�%{��W���-7����b�!�䌢Q㲭� �W�, ��fHG�~ !��(AhM�u�.T���� � lM!�D2\[��
D�!�W&Ǡ%�!��&�@	���V20IP�*+!�$��s� )��%��M t���!�䊲����!�S�y.A��X��'}2�A��@ >����dk��~O�0	�'�;Ձ�:L�^�
���'R>] t��=�dh��/{��!��'ݐ����n!v�,�<قi��'~�P�r�0)�h�e쏞 �@��'֌{wkW�ĥ�̇q���'/��N��PؽB��-X��
�'9
� �h�ݦ���JB+fg�0��'xF(�aۥ&��M{r�ǩ^"�ի�����[�Z��Q�R:d��:��b�!�D��rWH���:��
@:3�!�Ѵ!�xu3�E�'0\�!#F��5�!��� �rx�`
�)<<�ppF�R��!�$���A�0�0-P��b�OU!��ĴgR��(� J�d.l��W���!�D�&����ܣ�P�2c�A�!��V�l����"�]��(�V$�.o�!�D�;�)�W#<�F�d��!�X�(8H8[3o�y���,м{!�$V*��c�$�!a��fl�=6\!�C�y�$��aV�RE��#���*!�$�-SI��F�'���ɐ`H�U�!�d�/'\h|���V�e��L�����,�!���[����l�!��5ߜt�!�$��(�8���"� f�T]�˓�.l!�^/���$�cq|MӰ��!�$?2�~�˗�mC��$�ف!�!�/|f���i��HFx����ӽ,!���q���P�W�\+�`zT�MN�!��ΐ3_А�rGN=��e��I��=E��']�ٹ�#��7� a蓬��,z�'��2O�y�E2��A�|���
�'�rЈ HG�T���!ɜ�
%��1
�'{><��-� ����z��\�	�'�8R!ǘ�/X��I���A���a	�',��:��

5�qC���u���'y����S#V��Wa�%wf����'����j@�\\{F�_�l������� 聑�O�C���*��"��L!"OD��"?h�j�Yj��~�`�˂"O��	��I�#KJ�6��QQ�)�D"O��Vd̅MWA�W�=^P '�'#�I4!�&T(.M��H{�m��?��B�ɛI�\���%���x@Fl;]*B�	`tX���F8+���I��J#�C�I3Fg�2G������`-[�%<�C�	$XH`�Y���z��\r�l�OB䉯������Se�"����Vf|B�	�k�ް�0� :(�`Ã��!�\B�*_V�ݲ���5u���#��W3.B䉉.O,�w�C),_2��T'�-Q��C䉥�XQV�EҰ"&�ЮoT&B�I�p� )Q����tV �`0B�ɺ^D�)8�a��a���AFcO/��B��/xSb�[(]?�j�����)ÞB�I� _(1�Eϲ^��`�H�"[d�B�I�r�d�Z�-E����R�]p�B�	�G����Q�â_S�y�n�9PxvB�I=K�3{Zps"e^7�ġhF"O
)��A�3]�� ��)U�#n�)�V"O$1B��&9���V��?��ɩ�"O��( m�3銘�cI�/<~�M:F"O�T�� XP���'�8i�0i"OTmJV+Q�]0@+�F��\P�P�"Ov""�P&H�mi�E�>8>�@�4�'���� u܆��RNֻt_~DQQd�n^!�Dt�f�"*NA�y�HȤl\Q��G{*��DXp��'�0�c�b@�Wh>A�"O�X��&p����b�*Z����"O�<zS�Hp�ERb��){�0��"O���p�H�F��tfS:��U$"O4�2'�I�V��(QeA �D��R"O��#Ro��V��$�Y�L��yR�N�
렅��GF�BMV��Heb���S��?!�ՈD�����"��9Z�xҐ@l�<�R!Xb6 	���>	���K���@�<�/�.Y���X�� �J$<�����~�<���p���K^
c�P�� �]F�<Q��؁̈���Åˬ\�q)�v�<��M�s)�%ʡ�7��Q��Ny�<YA �09ֲqJ`&�+���2se�t�<)��XB�T��@#H�j����n�<�4�-��P �IM
��4DZh�<��P�j���#���t|�B�c�<y0J�!Xk"��S�ʚ�HztH�_�<���L$\����Ôi(��o R�<��N�"J��, ���`:�Eb�<��NΪ=�J-�!��]6�l��]�<��HA�t~m�G�H��BօY�<��M�ӂ�1P���pbp$�@��Q�<���+P2|���@�ja:�
J�<Y��5$��HI\��B���E�<�w�Y�l0*@�٭`P�A����Z�<qU�ذD^��i\0Iiꈛ�C	W�<Y���N���35�,0�=�/V�<�-݇B��X@��#�&�BDJ�<��K�ni�{��Y=SO��Q
m�<q!+W-d�85���;n5:��Q�<)�?�����eD��!�h�<a�D�<4K����Hzp=zqi�~�<���<��� ��=N�����K|�<A�.�<S1��H����u�q�o�<� ű��Ű���g/T�Y��J1"O���a�6c��Ԯ�/X �ȃ"O����(OZ� ��C 
˱"O2�apɓ�2�p1X.��l���pf"OB1!�6���b��ߕ�@}��"O�cE�A7���`��ѳL����"O�ѣ@@'GK���,��V~H�
�"Oƹs�<e�@0p�ߠg�uz%"O����j�p�R��N�n�Z�+ "O�̘��3lk�	��ǣ1ml=0u"O�}K���	�.8�F�yW҉p�"O���P�A0��8��ȏ���Q�"O���1��IL��+��4��$:�"O�m������%3�'Q���S�"Ofd9w%�4h�\bq�_�c����y菙m}l�#C@.4�����5�y��J7?��\P��<)M�ðJ�y2�P(,�@ȓJS�-�tʆ-��y�M�&��F�B�8�ԣW�P�y�b̀,+��a�;6�(b�@L'�yri����|����<_*�DÐ�	�y�%�c����\�P����`�L��y�-	�$c��)E�l�CP떴�y��J�y?�t�4�M�?}t�kXq��B�	a޲=���صb���K��R`�B�'�U�4d@���ЀNX�

���q1��4hS<%y�i'[D���'��وFR�s�F�����K(���'k���pB����)� �O\2��ȓxve��%� h>�����;m�~�ȓc�F�(�M����҅
�ird�ȓ7�HH2O�2h�2ς;%L !�ȓ9!rI�RB�?3n����	��z5@̆ȓ�j�C ��_  %S¨
.p�����o���Q��FRR��t@*L9Շ�/��	��P�q�^�$K�'�TQ�ȓk|��2��y�'Ŗ&-�jنȓ,�h����|(c��E�p�r5��E�Tx�d�jHj,`s/��rI>��gU���W��fWH̓R�׺L�(a���p!1�̏GU�eCP��W��\��~��H  �I�4m�d�X�T� ,�ȓ}���`b��&	IB8a� �.?���ȓ_�ޤZǍ��U�t�Ȯ2�X�ȓN,e:U��f��@���ݫ����ȓ0H�-jE�\/L��D3w%E+v�v��ȓr����Q]N�M"f"R(���ȓ~pĸ�2iё/@�Y҈�'d.��ȓ9�ix4�	N��Yh&Aܹ��ȓ1O(��ǿ�6]UL����p��u�fI�<��4�Ꮇ:1�4�ȓ�X������W�V��j�!5�<�ȓd���q�ٱZ�ܣ��G�f�ޅ��r+.�8�� mRH�S�̌<,��l�ȓ�qa���\�ˀ2@�.���}��&��/��]ǗO��P�ȓIIY��Kl=e�4�G�����ȓ9VLYa�,�	&�vi��M�8���?�T<ID���[J��Y�7/����ȓE�\(%�U�\��S`@G����l�p	����K�X���"��{D���. t 7X%	����ም��(�ȓ'l�$��˟d~"�A������>:uZ厔 sF�y�W/�$���S�? �����.;�	��T%�pٔ"O���`D� R@T�D,Z��>�� "OH���*���h��Uʗ>2e�혂"O��YEN��&�aҰɍ�:Fb�p"O��i�%u��4��BD� ��2�"O��:�cK"0F #DoR @��(�"Ox��%)՘)�쑒0.�q�֠�"Otҷ&S2n���Ox*�y0"ON��k�6Z|��1�#� a 0``�"O���̛V6�m3��G��t�2"O��䎔�+���ghˋ'0&Q�"O�5Ώ�[�D=c%��&oN�Q $"O��{6O�,0|�I��� � �a��"Oجjd�M�9!^=�%D�#8d�Kr"OB*�)�A��%P�i��"O�)y6�V�4��!��&?=6��"O(��i|t�����B� n!��"O�4q����L� E2��Q���"Ob9��BC�J1�ܱ���:1Nt="�"Op� `=ig�M?���u"O)�U���}j�p�Ϙ�l��1�"O��HBu���G�
o���I�"ORU���V�=F8�1r���]��h"O�+�4g߸qk��ҨW�R\��"O�AB��"kt�aؗ1��T��"O��S�13+��)VbA�f�V�1v"O���%EY��銃g
�o�(h�"O\����N��Y�h�I�^ػ�"O&( &Iė>��)�1M�z[
%��"O��m\�úՑ�Eǧ\�t�C"OfT�bh	�(2�K��a��C"Oh��k![H�D����!I�F�ɵ"O�a��U�"�F��V��)NNP��"Oi�0��$T�vp9��:~��"O@�"� 	m�e1M� (�p�8Q"O�pHE��P�j��6k��2���"�"O���bfӖ`1 A%O�{�	�Q"O���""��|u��EE�P
VYB�"O���.iڽ�u!�
mRl���"O�e�F[LR�Y�a�-[4V�KW"O�|��Ѣ7�8����j:��"OFm�e��;�Y��n����"O�R���f$`�M��,��m�u"OjȈRj�(�J��
� ?�� X"O$R!��:0�@I�5��}���d"O�=(@(�ö�؂�L3D���P�"O
��A �p0�AD�Tl�Q"O�ġ���gӄ��4o��� "O\�C�͉yo��3�\.ef#"O���Ҥd�(`Sr	�m*v���"O`�V�ި:��c�ܶ$*n�+�"O.ru���F<L�3��5^"����"O����G	�~5�mf��,e�"Ovy
X3z�XAd��<%5|@p"O@�f ^�G�<h�@eQ�:�I��"O�q�DhD?qV��P�Μ�9��u"O�t��]ZL1�w�U����"O>�0A���oD�R�ϖ5�85�"O�!9C��?�(��R/8Ѐ�8�"O^d�D�Վy�Bt!��NQY�܀"Oj�R7��# �(��e�B�gC�8"�"O:��Q�ډQIwk�>zQ	S"O���4.U.2J�����ɘ�P�"O�Q2�����;�k�*W �A�"O� ��*"CڦX�����#E0ȡ�"OlT�Q�Œ9� �Q
rN~��F"O,��`CH2r�lpR`��f�2�"OFX3B�Կ1��ɦ�����[7"On!PT�Z{^-H��,pVR,S2"O�`p3霪\�D�I0�Q7_5��"O�D��)SS�����/-40JF"O,�R���3����B�Q�H��ᛓ"O�t!&�ϳ�a`��r��Ys�"OV�Z��@�,�q��aE�p^ @�4"O�	��޹�NԠw+��-�Y
�"O�8���7�@���H_$BQ�"O���e
 �-%o㤡jr�(�!�هk޹��"Z&cx��q�u�!�D��
 ��M�:~��bv�߄l"!�$���@�2!S5~ݾ3��0�!�V��`���m�%k5k	=>!��7k��܂@*��-��uIG�V*!�و!�!iBf��`�Eʞ�!�$Y15H1bR�R�9�i5CQ�!�$F�@J�p�6�ĕa������+r�!��3��T�7@�7ik�|Z�猹3�!���Uq�0nK*HN��X6I�C�!�d,mP2�aH+ y�A� A�!���{xJ�����2�i��*\/!�	p�� ���g�~���썻^t!�$^+	g�!�4G�dj�T��]�*]!�B�]|9�Pk��C�ՎH7!�d;�D�SDK/SV��HS�89!���4'{8J��^:,��#�!��_�Bɞ����Y7FPU�fb�+	!�䈬5�⵩uEԇqP��
�����!���.f���f��TJ�y�bM�|�!�D��>�^-�D�&3IVԀ�N٣b�!�z�8��%B�!�$�@���zV!�*�xY��GZ�_���B.\|E!�dKr���#�k�*MsH�D�9V-!�C>��h�͖�OeP`�Te�*!�d�1�zy��g��v����֛y!���44��
Hr2�)3C7of!�$ކ K�5[�CA�zt����"W5#`!��P"�Ì*hƬ��q�M�fD!�ĕ<Z{��G��[�T�dM�XI!�D)��0"��/�0�
4j�� !�$�)od^�i� ��mȅ�ʕ!�T :�B�iÊ���<��ۣ0!�D�!lC�ܛg�G�T͐��6�!�d%����S'ߛ� I	���H!�d�L7�`��m� � P{c�!S!�$��}d�a�фۥz�����D(�!���#!���/,n����#?|!�ӫ^�xMq�\�@V|m�F�3v{!�ă�)d"�%!�UMT+s�Ė#E!�$ژ[1�X"�Z\H%�q�M�?!��1�P�S�Q�=0��QuڥL!�ě�����k�d ����,�p!��Ôo$��0��".� !�P[�"OP�:'#I�6s�lY����  �L��"O`�j���������F�9,�"O&L�7eΥ)�%�P��=�JY��"O����\�>���mZ�.r�i*p"O��p�k.<$)��B�~S֨�v"O�pjD�ص8�J��1��h��\�4"O�=����hj|�8A�/���`"O� �ȉ�I�J����
�L.�X�&"O�`ĪA�%&�y�6G�M��*6"Oz���Ӎ8�*`��U�9�"OZhQ�'I�����䎘5��u��"O�C��?TR�Y��]W�ˤ"O��a	<
���!�4=8A"O�+����f��M�a`�1 �E��"O�Ĉ����AP��S@FWA i��"O��T��Px���N"O)��y�"O:���+P����X����"O@=��J#j��-��O�~Dkg"Oj�Q�`ãDm ̳q�5�Ι��"O������^|*582d�d����"On�rA.��Kø����ߟ.���S�"O �0eNF�.��hP��sw:�3"OF@+2L���A�Ƀ4@R ""Oօ�#�U1]�� CbI�F�d\�"O�	�	�&�^T����u�i�"OP�Ar�P��ⴘ�CK�&q>m�"Ox)�e#�Rȸ@�R�[�~���"O̤�P�2V�a�T�E�Jl�ۄ"ON	:/�6 J�����
�O��c"OJ x���7)�&����|��ɋ&"Oj�(�,+Y����*����XG"O�@sb�ۨJZ�{R�=&�,QE"OHQg*8LH1�g���ق�"OL	�'�L�>�����"Wܚ��"O�#'��v�p�DG�'/����"ON�+2Y��9UϠ	(|��"Oh�i�A�5���)���$n�ű"O�%�Q��1���`U2)+��@"O��ڥ�%W�̣�,E�zo�h�!"OD�j�N�f�(}a�KI%�2�Q�"O���'��rߺ��KۋN���z1"O�l�(A/=zĀ��O+���S�"O�9�6N�H�\-BQ�Z0}����"O(�"���/T�����96�j��"O𡅫�^ʤ��-�1� � �"O�����Âu>P�Tl���XZ"Oh�����
)� Ѣl�# ��ٺ0"O�SG�B;\x�ӑ��Q����r"O�����	������|d�b"OH��]�@W�ISH'o�4j�"O�E"���L�i�F'�d�]�"O�<Ӳ�I?�Z��ǧ�52�c"O d���
^�Q�2F�
eٶb�"OR��*_�;�������/F%޷�"Ov����̠E����U�M�Cl�cr"On��'o�
�򡒷�[I����"O�AbI1X^Pc��@�����6B!���=�ڼif��`el2k� �!�Ěaݾ��tf�0Jܸ[���A�!��Æe�XB��pDD�X�ƙ�!򄅎E|p�)�'
�U�|�[��7a|!��QP�x��ϕX�8)��3t!򄌮wI,�`�
G�*���wU!�O���ТE�l= �!W�� |!�$ޘ0�̡rTI�}�E`� w�!�D4����G!�HAE�R*!�!�d[��f4��O�l
N1s�-��!򤁟zFZf-6o&�m��mA�{�!�D�{��r��E;2zұ��B@�V�!��޻m�
]sH����M�H�=}Z!���s�fx�h���y�&ʉ�!�� ���w�I.:��1rEn\�,]BIcV"Oh� �CA�����V3"x@ ��"O�|�e@�5T5{��$ma��"O��  A��V�"9��%��$UzE��"O�P������0�EF/5�MPv"O�Pj�B�!��Tqc�@/�h�a"O�H��ǆ2oV��UkE�w i��"O����#�gs�[���2�� �G"O�I����� ��KӃw͢ـ�"O�Ё
�Z�2�i���h��)�yRI�D���B�hJ�q��0f�.�y���hstm$�J�ezN4"��F=�y��.��B'Q�[���Jɶ�yR �%Pl D�@O#Z��$;En]'�yB*��~�� �o�c�E���y2����\@���[dp� ���y�P�8��!��
M�T����y�/��Z��Sܮ|z|�!�H���y"�;t`z!�p燴z�)q��-�y2*\6�V���ND�a"���y�K�k}�Z��̶?�nY2�N 9�y��ґAM��Bg��==�p��Ӥ�y�@��~�|i�nG�2d�		#�K��y2�l�	Z4�N$�
�b��y"��6��\ʓ@�&Lt�@{B 2�y�*�SټIJ�#Zp�����y˞0�@}���T �JE��L]��yr^�_�Ҕ §|��Q��N��y��C��d�s ��� ��y�(-z��(C�c>�jefk9�y"����b��q� �xEB�I	�|Z��ŭ��sɊ2B�I�F��a�� �0@&�yw�
?!�B��.0"9��(K�d��p��%�0B�	�J�u��	t�!�!�H�&�^B䉼U�ܬ@�,�,,8�	`��۸r�@B�I�B�*,A�
|�:=����2%�C�Ic~.xAg�? nMxg��)�C䉐tS�5��O)<;�-b��	;`��C�	& � �r�d�<S�p#�(�0&C�	=D����L�xTR���8|�C�I<9��Ը��n��)�����B�Ƀx�<���%Az�]C	�� B�I9E0�����U�|M	�'O�E��C�	">��*�F�0��Z�bM�U`B�	;��Y0�KU�h�4�M�;Gu4B�'1�ppC��6����"E��C�I?#2q�G�q��0ѡk��85�C�	�<�H�S-6��`q�Iں;\C�I.it�\�
��4隐�ׯV�b
0C�	�:�
�B�@)��dI�HS�nu�B�I�?B�5Xw*�͆p�dE�� C䉩�Ҽ��I��f�X��tぉ*�C��eJU[&*\�3:����� C�	�d�YzՄ�LT��z7%ކd �B�I ��)KG��1Fb������x�B䉧Cp���d	��^I�hdዟ#�<C䉖	��G��� =b�3@�N4:kC��%J
������Ql(Ҫͣ[�B�1x��ӥa\@)Б�̍_?tC䉽K�&}�CI��8�0�d�;V�B�I�:,�Sd��A�_k]�B�	:_(|5)'���Ns8���D����B�I58	fE�b�@��j�%+Z!�� fd��L��kV$�2ů��}�Tઑ"OR5��� 	�������.�*���"O�C!�U%L�b��[�L���"OZ�p�f��P~��c�C�e���"O�h0�'l����Շ"֌�A�"Ov��A҂w���$��>�ʙ�p"OH�U�\���� �{v�L��"O<�@C�ɲGy2��C<$i:���"O&Xx�-8F����J({I���"O�](�ˢ  ��.��/@5��'�p$��ʀy/�Q�6$$o��0	�'lf���g_��X�F�s.��p�'�f���Um�l�u�R�t�V���'����G��&��Zl��b��X�yB���¥Y�j�8NX������y&��<����%�"ȢHR�=�ybbK�9
��f	�*}��`1g���yb�@�0�p��'l����1c)�y�FY�F���j��^B�	�4`���y2X�Gr���mB/G��)GO��yr�ыB%�g	AC��p	I�=�yR�?d�������.$��ޜ�y�ȱu��@�!�� �t��%A��y��*�"�`MҗG� i+��y���oHxb�Pd�x����y���GWf@�e���2�K�*�%�yb j~�|�Ӌ�>/�� ���y2��F#�@s'=zȱ��+�yR�=�@�
��93���!����y�k�)cK:�k��0=j���fƐ�y�E�rF&t��H�2f�@ ��T��y�!BG�a4��x�y�qn�-�y"A2~��p�4|Svu��l	��yr*ȵ8��0Ud�y{Ƽ�V���y�/�4E����&ő>io�kCmQ�yR&�!ƒE�����5 	)#戎�y���%��� m�
.����.���y��[�F�*|:$o��w�Fx�u���y�%٨ht�@��f'`]�1�љ�y�k��dc2����ՙX:�\R1� �yBB��T,�˗/K$�2Y��^��y�2mZ��w�V�|(3���y�,�1׺�20�Z("<)�".O
�y2��3h�|Z�	�=E&�q���yBf�0��ؐ���L��Ue�'�y��V�f��l��=t�%�T(ɩ�ybC�2N���w��z������y�
6�r��J׷3�=AT���y�NLz����9}�ڬ�F��y�l�&���
a(�?BC����V��y2!E%q�@�Ɉ6:|X�B�R�ybޅ(� @���axD)���yr��0w��,`@�k�sfe�.�y�`�8��x��ۍ^yc���y2�� 4}"j"��\3~�!c�H�y2��vJ������BB,�x�	�'z�)���S�!`P�c "a��]y�'���;����8�>q��oa���'��h(B.��Hԑ��DC�V����'���#MFJ� �n�N����'� KA�D������ȹw�$�	�'.�ʔ#ߏ`JX@QDQ%n;(P��'�H@� i��:q� �h7���	�'Xܨ���/� @ڀ�D8h:�	��� La���^506���/�I.��"O��B��mh���D>E$c"OR��U  mQ
y�f��KZ���&"O4�� ��s���W7_I�Q"OV���'i�ܻ�-�a<��� "O�\8h��+�:X�抸k/���"O�l	�,�5��ٶ��!A�*QQ"O��c�߄e��S��W��QZ�"O�I�Vh�F4]0�y����"O�50��Q�px ${�#�+��ڲ"O8a �)̂W%��Y�o��^���d"O<S��$>�ı���zU�U"O��Q�"K����TN�U��p�"O��@�	جg���������ӕ"O�B�oמ,� �Ke�H
�<��%"OFPS�^�\��-ɕ�ښ|q��g"O���r����v֌� 5Wi�"OdD�Vǚ:Y�E1'"T--���"O:��P,Q�0�8CD����R���"O��b��v1
��.¦&ꉀv"O�yJ΢.���qOOI��͸"O�	��� �Z�heX����l0���6"O*��M�=�v�8!K��~*���q"O�����0��I���=�r�a�"OX��Y(�#�]8t��7W!�d!<{l]eKE�
�q�ϻl;!�U�ʨ��59�\ipʌ�,�!��E�|�ڑRqa�+���H6���CS!�DLoOܰ`�E48���H:W;!��yH��	�%	"3�d�A�ط5 !���q�b(��i(��1b�n!���P�ĉ�A�J����Фlg!�$Z�*/�tcցG=>�D qU��,!�� 3��Sq-��h�(Pì- !�D��7�dd�D%�?oV �E�R�`E!�d3<O@Ip0ß�<l*<!�J��h[!�N�x�p��k�"'-�j����*F!�d�75�t)���w��`xUF)x!�$H,^+l�t�[(Q���hD[�!��gY`ኖg��|�.`�"�(A�!�dنBV^!�g-�>���A�L�t�!�DH�z���z�# �)Ҁ±�!s�!��=uP��ZW�,r ��n�g�!�dW�s\u�����DZ`�{F��1!G!�F+�ڤ#P藨|2I��J�hB!��t?�p��`A/J���D�P(yR!�$WY���d ~B(Fk�>A!��Th� @�$�!2<)��i�:=!�D%'L(Tq6�����1.��L�!�ċ@�2���!@�>�`�5�'�!���Ťyo�6\֬Q�v]5�!�d bZre��-� �.��#j�3`|!�ՙQ�Tm��@E�_��x���Ӷz?!�D?(D���e�Ծ_�,0QY	6!�$�>Z�U�0M[&��/�!��S3�� �A҂'�&qK����!�!�Đ
~�s @י&�4���-q!�G/7� ���� ������6r!�$�ϰ�c�/�!o�ਠ�W:�!��?s�jx�F� �p1�Zn!�ċw�(�!'�<j�D�@��!��ڍz*0	����80���]"!�Ę)�Ji�g��c�.	���
{!�B'�t@�EAܿ6��@�&aX�Ss!�� R�@��,m�Ć(&���"O�S�GK; Ub�����.�
��"OX��6)G�
hu(���H��4�G"O�T����Bu��r�AY��T"OQ���<W�t5���i��G"O��×D1rڊ⇬�.��qR�"Ov�Z��ٞ�0��1.,V�v���"O1a�_C9�+c�O�NYr,�"O�]��$����,M�D�&!�y���Bi�A�FX!A0m�F���y"��.�1��G %w�����J��y��0v'$*E��x�;F�E��y`P�zkt5s�NS��l@u��>�y��}E 8���H*UzL³h@��ybk���%��fo��*�(%�yr%N�p�x$����d��S2d،�yRb�R�0[�VA AL�:�y�� V�l�eɐB�Zĺa�S��yRΚ�4F �5
I� ��y�M�Vc��#�צT(�0��,�y�=/:�d���TT��E��y"�t��8�Ί�(�h k�(/�y�˅A$��d�Z�$�`�SBn	�y�ʂ�8�Ru����l�4B��y��<wp|j�+�SL0g��y��G���Y��摜w�$��eO�yb-E}��@жjZ��Mk�(S��y"��#~�&g��j)ھ�y2��;nE�O	�O^h)	����yb�{Ԓ�8�]SP�
%��y�l�+j�c&��b�@��?�yҭ��gf�UR���\��ď��yr`ӛas�0�%O�D}�Atl�y�BH�`�X5s�CO'C ~������yr�Ѱ ��XKƪڤ-�~�����y��Qp�<Т5۔O��y3R��y�i�1��&��7K�n�1�΂�yҊ��_�Z� q$*L�� � _�y�
��eJ}�D�	5�4q���yrmY=&�@��|QL-�N��y⣑�I�aA֤�+p�&�F�y"�ϓ>=X�R n]�lv��J���y�_��|	�W���_d�&/�,�y�N�=F�(@�D��W�z�����5�y�I�v&�-��MصL��lz��֕�y�l�ԡ�D)CȊ؊Tʓ��yZ�6���U�ԗ8�&���ω��yR �s��J�C�4�<�:�F� �yr&��0bX��Y�3�*���M��yB�A�6���x�䎀'm�
p�?�yR @5O�v����L�1�ҁJ  N��y��3Zi�%
�������穛�y"f��(�l�cMЍ`��[��	��y�)�=�E�fl�#4��3��_<�yBe�1 ���蕁��l�����y2�;�x�Ta�"*6������y�i?)L4��N�ÈU!�"�y�C��\�3QDԕzb�a�Q
޸�yB�K��M��Bw��D���E�y�Ē�~�	!�$Ń]ޜDR�n]��y��!T��w̙"�9qw�P�y,��Z|�P��� �J̙�cʭ�y��ߢ\�FЈ��0	)� �����y�jՔ V�hy��v�\ՓTG�!�y
� ~�-H�a!�Y�LK B�xxi�"O�A{`K����ED�Tp����"O�а��ǭ7�h!`�/lQ���6"O��
�Um���7O9V9�M:�"O�a�aeǽ:&��#E.#j�"O�� bB�D��=���5"O45�m��@�Rm�%�dv�m� "O��� XH�tP�-_�_S
QyC"O@er ��2$bz���.ы4(h�"O��!�K%�(!.�6F2��hD"O���ud^�6[���mA�Q%%Y�"O��ʁ�Z����P�I�5l !�"O��	5e�(���&#y�Ei"O��8T)Y8��ݻn��p�"O*�¡���u�&����M�Xk�"O,袦�B>q�U+!^�w+��:�"O~�����?M| ٲ�ʌ��:"O�!����(D��(=n��C�"O6��pNV i#��'�d�8�"O�$�7i͊:��a���	�TU��3�"ON8Ig`��BV��A+P�4U�"OR���ȝv7����o=k�R�"O�`��� �l|#q/tG�D�#"OА���[=��i��^0l2�y�W"O�%�G`H�Q�mʆh6�&�ӥ"OZ���@_UyQG�#[��b"Oj�3A�ɫ����s�O�wV�Y��"OZ�Z��K�ɒG��4Jڶi�D"O��Pd��;3"h=��Éu_4�[�*Ox)Ӳ�˖sv�%�V+FN��'������LVU�$��qk�5�	�'d.�8�KS�Pf|1���-i `���'p>��#B�	R�P1e(�q"H��'{T���I�2��4�:i��A�2�)��A�$Xnn%�'ߤ5�8,��4�y��ƠW',d8��:��q�e҄�y�]�K�00R��_�z+�u�4EJ��y2N��Z�x`��wu`�xT����y�mN�6ܵ!qL�i�@MK$ƕ��y�LS��n�Xfh�*m}(��S���yB!�&).�B�$ܚx����0��'0ў�O� ��C�w!�|���[86�.I�'�<iy�K�-M�"�r6#�([���'s>�c�h���D�B�1e�5��'.v�14��g�ř�Nێ
��$A�'�$��L��B�����kʿ9Dm�'P�a�4M��cИ�I@�*�s	�'�dАM�D*�I�v��V�j��	�'��= e�� o�1�c��T���i�'s|
�j�0��1�EaU�#R�`	�'h~�Bp�A�8Y��L������'�\�ńs���i]!����Y�<A��ήѺA� �;g�m�Q�Q�<�e)#�[�e  nvTU��P�<��쀲06@��'�VʄH�-�K�<�3�Z#l���{#ʛ�z�&����J�<����%�
�y���0:��+�bYJ�<�`�L:3T�����)�:�!�'�0�y�I��P���Qʍ��Д�G�N��y���<"�2d�gʔ��9qv�8�yB�5�����_�5�P��Z1�y� G�1�RgDN�A�"����\��y�E#'�q�����A,�@�e��y"!��~���:C��5��PUΆ$�y
� ޕ�!��"#�e�u�E���f"Ol���KV�PN%��B�dV�"Oޱ�">R@03LP�\x`""O|�d"��;�%k�H��-��P�"O�ذ�S�r~\][���nk"���"O@<��e�.GK�ܡr�O���"O$���T_�v����=� 	{�"OJ�(�*�.o\�M�0F�ƀۢ"O�1ibgِm6�5:�mH/B��t�D"O𘒳�Ƃ=~V��k�,k�"Y٦"OpѠc�LH;d�����qw�� �"O�X����t�T�qW	ܗ^k��5�'-���>"��`
���(��ʖ.d�C��.tQX��v/A�i�ʄ�FG
?g�C�	0)g������Wn� �B3^�VB�I�{gb�#&̝0�^X:si�k9tC�I'gƽR�*ߣ4}�-K�	<wv
B�83�֍�G+ƃ
^x=�����X6.C�I;�� ��уg1���a�I�s�B�	"fQ0h�s�P�;��a ጟ[�B�ɯI� l[����25h�����t��U�E��#6O�,����bG&s!��C|�@����I#=�J +�oP6S�!�$ț<̈ɀ�ܗV|Z\pp�ܷs;!���"9� `�kT?��`
g%8!�dZ���.K��8��lA�p4!�P�}S*)xQ�T�P�w��&!��F��<X��˛Y]<����ϲ2!�D�T#:��A��oAm���!��\k)� %�ȇ.��%y���	8!�۰2����!O�#�J�`�a:yJ!�$_�x@*�;42�����O&4J!�$��&��q���33!�s��P a"O8�W��>zئI��u��l"O�c��ܲ&d��'`H�iVV��f"O<�4��3)e��/՛IM�}+w"OXA����2j'�u�Vn�aB��iU"O��JUm&tflL�b�ԌF^,1�"O�M��B*L�z�N�A��"O����P��[��ty��)�V<!�Dʉ?�����֛r=h��bjE!�dH+�©��@D�0;�qٟ?+!��S����(W�M.�YHe�]n!�,3���d'�E�D�H&��h!����y�,
�?�����*NT!�D�@���Za�Mv�L�I�^!�DP��P5�$&�-M�yf.�
�!�$�w��qZE�Z�!�H5���Ī2-!�$9��iP`�\�V��%��F	!�$R�!I�xPe(R�,�"�dC�6 !���Y'�	�5k_>z� 䁓C�7p�!�Ē� ���*K�Ll���F�o!�d���h�G�Q�sN� Q�Ϝ�U�!�2�r�16�Ɍ7�2��um!��F�8�@��&*M��f%3k!��)4�\!���n�|	��9dN!���,T�봤XOqᚳ�ْW<!�Dۜvˬl�g��0I"��	�71!��9QV�����#�"�!ȏ0]E!�� �������;�<�b��7P!��ɔv���'�2`��å��\!�d��%򞔠�� 2&�Q��Ǒv<!��4�<k��mƠ�Ғ�ȧ{&!�d^ }��!Ô�B�5�ҝ���0#!�� ��s ��W��h����W{ޅ�"O��A3��0�^����Edy�ݸT"O�C�̌V405�ȥ��{&"O����e�[���E��K���S�"O���uOM�w�Y*#��]��DS�"Ohѱ$2��Ђ$���&��h'"O�PQ��f�0B&�=`��6"Ota)���j���� ą�H�rv"O�ڢɍ8	E|�E�Jqh�f"O:����H�k�b)	e;��c"O�H��j�H����"�/$�"e�"Ot��--O�qR�
fI���ϝ�y"��p�xl��_rX!�v����yb$Q),&�4�J�U�@�&���y"h�9h��IY�,]�S�
�{�����y� #<2lH���uP`�$	�ye�:q2�����$b��`	$�F��yR��'*��Q O?U�1�_��y2�Բ	�>�EC  VDءx�;�y�H�!3�x\��Z�m�(Jí��yjM9wC�5�BW�r�y�R��>�yr��%@��X� OS�����r�A��y���:wn��s�k�"z�.髲�U��yRg�<@��Ip'�xz0	[G�Y��ybD�L��G�,	�ժ�ǵ�y�H=�.р�i�w�6��eL��y��X�8���Ɩt�pq:�Y��y2��vt�@ )I49E&Ȓ�C��yR�
U#<��!h�8�D0����yr��>ax�&�L� ����1�y�f�5T{�sJ��D}�<���+�y��ߙV�a��+�$����gǥ�y�MO4,H�b�I�!�z���*��yr��rI�r!�q�����Q��y���옰�Hq��]����y��$;j@��IK�\*<��b��y���[����4�X%nq����.�y� ֊(�X �0"�#2��C���y�&[ ��9p�Ԕ
��X�LY�ȓ%�r�I%M���fkՓ.0q����PdlCC�e;-��Q�T�ȓt������'3�Xp`�*�&lx��	���P��(fId�d�V��d��ȓ2,�z�'F�VмH�&F՟.��H��e�6�C�C�_ h��.�?�8M�ȓ4�����Ѻg �p�]�z2����>1�v��.5��IwG�VE�@�ȓZ��ٕc+?���!���I��Ʉ�9�Y�WkS
 �qb�Ű?i�a�ȓ8	��Pa ��Cڴ#� �$։�ȓ0�v���L ��}�r�X�'�ZH��m�F�����<P(]�Ģ��t�ȓ)�p�"���6q�6�	'��lpf��ȓ�^���Qvv�k0��^�Ѕ�<�HaS�!�IL����ˎ�3�6X��\�H��զ�X���AXpՇ�dLu����1FZԊT��r��̇�Q;��jA��M�6e�7���"�2���{y�l�d�B��d���7N��ȓi��}�FF�s��(ڡ�ȏ%"
�ȓR�v�`j@ʠ�v�	X'䱅ȓS�<�"���	pxA�$�́)̴��tL��h\�lR^Ĩ�g��_eJ���uԁq� Jt��
�Mxp|��S�? B��f�;fl��MNA�fH0�"O�U��@�*@�zj�B |B�"O1�ƀ_�S�� � G���"O`=ђ �/S�H��#��F�s"O����۰C�,xP�#�*��Q�"Oܭ��ϐ�j�`����ыزA�7"O�qj%ӑ +*Qb�O20�v%:s"O,u*C��*Pmf��BN�j��dI�"O ��� E7x�UC��S#G�q�t"O��yCjZK�f@9{@�x�"OHU�0Ń�:]t�����$:<�x(�"O�-wF�?z�L�����+�4H�"O�`�ӡYnT:��k<pCp"O�t�c`S�YJc'x��=	"O�� ��;*���+6:��Pv"O$Ѫ/�v�u '��`<���"O�@��� !񲰹��?d)�IY�"O�0z���vo>�8GE$O𑺰"O*<����5R���c�3"�|I%"O��XV퉤3��a�锑7\�1"O0�x1'����B8H%�	J�"O8�&<�^�#��S�6��a[�"OLiȶ�$ L�a��-�؈�f"OP ���R&��(��##��	�"OV}Yt'�@0C#ۙ�B�w"O���SM����1w�F��%�Y7�yQ�v���)�?I�A�D
�y��֨~�N! O�	1��%XF	��yR�0~�<c��ŇQ�l�pj	.�y�F XCR�ʗ�I|�50�F��y�[�Q���I2�X�:����& ��yBF��f� '��9��,�C� �y򂏀n���cH�*.�j��1�y�BS<��1�&��)�d�ReӅ�yb�V���QL�6��D�!�,�yr���y�e�BD��D �y� ��|0��ҡV%�IS��(�y"I������� ��Ezp9�ᅲ�y2�X�_i�@$o��JQ
Y3�y".� 5�.�ժ�Z��U0�$��y҂�1,A A�QGD����;�y��	�j/>��b��S\fE��*I��y"�]
34P�P� �+N�Yc��^2�yB(ܿh�x�5��0K���a�V��y�l�q�.q���.d�\;�I��y��
����0䭠Pة�y"�\@���y���	�xP·&�y�F� >�$h&�y��`�ʛ�yQ�0��b*ė.� ��ƕ�y��+A�@��N���Ȟ7�y�V0%�4��Nx�h!3#/
��y�k�DT4y��Fޱh�r��B�N��yD֙sZ6����o�ZT���-�y��I�h%�0-��jpv9�qɔ(�y�k�9-����*�d��p@����yR��;0�e#1L	V�̬PlF��y2J��6�����fX9L��ThA�9�y��]�0�gD�;C�4��-F�y�!�N���z��Ov&Yf,Q�ybN� ���"��0tt���
�1�y�$E/Z$>�"���lX�+7l�(�y�H�����R��&j����fE���yr�aK�Ph׸^<95c�y��G5g�p��ߌ^�l��$���y
� ��06��)�!F�$�"OT����S23���3h��`'\y��"O��CT�� u��@��i��D�r�"O�Iې,Dw%�}�vJ�|lp�`"O��:�D�#4^�M��?v�f`�q"O^�ȃ��>G���f"N�7ռ%It"O8�A�:v���P����PИ"O`�:Q��KG&��FY#o�X���"O�{0���_����E�[�.��"O�!��θ|���T���6�B"O:�:�&� c�6��@� �Q��':���S@4||����A��e��8�'?vab�E2}�pi0��o|�Q�'iu�o�2�)өa&h��'�0�J�!̄��pH5��O�$c�'��'��x�	3%��p�J�'�δ˂K
yo6��E`Rz�h�H�'�V 	�靘d������Жt�"���'.̉��/��f����AK�C��m��'a�b��>�"΄4�У�'�ԹE%��M� �HT��A�@ �'�2�'&&JvZ�p��Փ8���8�'p�5�O�,N���W��zJP�'p�X��_�ȉ�FƋ�y!`��'��5	 ;[�4r!&�9v����'P��� ��3��q�ڨc��� �'IRX�0K;�H}�p����؋�'�(��uյ3$��e �� ����'�^`Hg�3_0�+�,v�6;�'W��6�ۦ����,X�kN�Dx	�'��ص��$1z�qTEF�>�%s	�'<C��\�$��M�3�́gy��	�'� D��,n��<Cd��:1.= �'�����-�}c��9�Js;� ��'�$,Dđ����:nQc鈫�y�/j�@:�$-�\��,�yrE ��Bp!瞑ya������y��$;{�x3�!وjZ깊C�y§ݎI"�K!%��kp�e%X�y�C�?T��J��ĭ*�qׁ�/�yrD�l�&! �B�RE�3W!�y���D~u����5P5�P�α�y�._3$R�́��^�;S� pA�Y&�y���g��鑪##���[�c�
�y�唝Mz ����P2j�CZ��yӏ!��d
v��֚Q
�Mә�y"n\-T#��cL��ȴ\ȴ���y҆ۧr�tQC�P�3�ۆ�Ц�y�������ei�*���y��Xx�]���H'0�(9�p�ص�y�Θ ?t𬉵��b>�SЬǹ�y��0�*�F�R8�jq�����y£݀#R
])�[#-�%��	B��y"-��%�,����Je����yR��t��dp�E������Ƈ0�y�:>��)�������C �'�yf�9H�R��@�*ݜ��w���y�m�s�:�р-Evꄚ���#�y�NֆKh&���E;i���;��E��yb,ƹw�B��6l[ �,��y�+'N�cd��S���Tk��yBK8m�����5rb�I1�P�y��7�~r5GZ7�pY�3@��y�-�?t(�#�眓��ܣ����y
� � )6��`x�;��� �>�0f"O
�x�Iº!R DL
�,�Ku"OF(IQ�2~��I	��̦bҞL�u"ON�H��5e�PJ�O�G�JUse"O�5jG�˧5�(t�Gi��v
�"Or&�5S����@#ә:�\�"O�y���+Lp�#)
1P&���"O>X� ]>)n4(G
�h�Q�Q"OX�ׄ�yT�9s�EZ�ao�!"O|���ʞ�	�z �c�	f\Щ؀"O�pw�,S�r�1UL](O�T3�"O*����?y4��2�B�k�Ƞ"OI��DTO�d��t �>
����"Oh�3�杜�ZE��\�Pi�!�"Ox�C�E�}����Ƣ���C"O��R�d��e̸���5W�XthW"O����%��2���Ж���Ϊ�P�"Oؠb��T�*`�4�4��x�Ib"O �p�� ~O ���T2j6% �"OPh;,;/��������&�f��"O�ls��Yfd�	CD
�G�T�j�"O�-c��3&6�:Č�����s"O�<�6�[<`�2l�41�b�*"O� �f8W_V���I�&d�&Iڳ"O��rG,��cAJ�AFC�,	�"O�M��G `�X��!2���"Or���5�5:�B|/��:�"O��yf�˅!)� 	 �T3�Py�n�B%���@��D�����E�2�y���>~w,�wfhR�ܫ�+ ��y�#��00�2bK��gL�a	�B��y��,4 �9���dJ�qF����yBM�{�jL��HVt-��ƍ�y�ƒj$��s��<;'NA���/�y2��%^@t0��/���2q���Ɋ�y�Dza0D�D�ټ{�,y{2����yB�U
<�hL�g��*R֘2ポ��y2��3���#+��@���"���yR�м9: �	7�̺�������yB�2[�Pi� ���4�1��!�yr���oۄ �'��ؚ���G�y�Eē<��0�/]�AɮH�5!޵�yB�M�g���/ڹ=vde��L���O`#~:!Z�;��af�A\A�q!@�8� %��K��G�\���Lf#�ȓ�/D�� &盒��\b�(�Yk�X�\�!�D�6�6@R�j������0b�!򤗶}�"=)V�D�o|��
ԅ�H[!�$�-5��\:�-�'vD�aP���gz!��
��q !bPh����S�_�!�D9. *�h�a�TI�T��Aj!�ũ�
-��.��WE��ҡ֖3!� &6�^=,y�.��Ą��:H���'Y���n	-t�~;�
�T��'َi+�(�Tt�3�D�!!ː�	�'���#�^i�XB���o� $��'��{��0���J�F�g��,��'�*��C�]�i�8�a"O9Sf`8K�'-P�� '�/plh��\�EO�|�	�'�F�P`N3+��ط��:/T|��'��؂ 
E��p�ㆬ@t�؝��'��$��� �<uP��ㄟ-a�x"�'����'$�!v������].:���'�*�������i��nG�B�@���� lD�P�N�!245��'i{&��'"Of+�O��Ȅ!ׅEl��i�"O��
gm
M	Z��a�C�&�xd�Q"O����N� ��]��`߱~���3�"O�� ĩ@"s_��gm�a�Z�"OP�4oīO�|���mq�"O^4�q	�2H��ahA�E��٠e"O�|3׬ρv檈��/�%.���E"O^D�CW%�Z	W�B@�
}6"O�8�E�z�a/�?���ѣ"O����M/'o@� #��-���W"O2��f���Y��=G�ղ<���"O��D��0|�R�� ES"F����c"O ��@@M��:Ac�Scr<a"O�ũ!oH:^�Fd@eґ]]�� �"O�I�"a��]�V�&�M/nVzU)!"O�1�uT�V�i�u-L [D�I!a"O�̙Db_)��gl�!/�E"O��ZUl�4O��C�k��E,޸�6"O�jU�̒X�H�
1Ę![�0`�"O��:��_Ne����(�W��`�"O@���o��x�B��5�
�}_��[�"O&M��I<<�6���5OLIY�"OJ�q���2���T� MB�@�"O���D���L��X��±=�\J2"O9K1IN�B����`�T�N�"O�,��nޅ-��!Sâ�n�8�"O"0� �/�Fd �'F�|n蒀"O0\��K�~'`#a�F���l��"OYKU�T"n����߇&��1��"OR,���#q���b�-`�إ:�"O��bV��lpB2��M1!"Or�B�W'O\i�A܇*�~���"O
�'u�J}�i��J�~t!c"OJ��'��G��jE֗w��y��i�����p�¤ua!�j>3W"O�4������]�-"WBl�sq"O4q���Lr�Pǭ��.B*db�"O��y�O�N-�J��E���&"Ob��G��7�(��։�3 3�8��"O����JP3_��[�
�,q$����"O��QCf�'��51@��&�E"O5	a��e}�}+w�&A���"O큁g�~Z�5k��4���ˡ"OzH7�+T�l�rfD�:��R4"Ol}x&iĊ(�:Y6��RqFz�"O�]�g�=B|���A�4>>�I'"O�x*e�$���J��O4��*�"OF!�W�u�1q�,�9hDt�"O4�sSTj@uC��4c�N��4"O��rw��?1\����<Y�7"O:5���.q}�J��%�ҽRv"OA2Ui�#���9�Ɵn�Ġ�"O�4���B�!>��B`6%��Ds5"O�$��C�#|��u�@E�9a�h�"O�1f��S
B@�b�h�e�i����$%5,0�0��?��1PǬ��E!���B�c���i鈵��;�!���`5� Hš�a{`�ր>�!�S��D��g��g�D���B�^!�'q�ȈZ ԪK��������k�!�dԐ?����W'i�d��Db\% !�Dǩ3��Af�O} ʣ[7)!�d�&&K�U��$��%\t�s� ߯e�!�� ��8���d�0�Ҵ[b��"O�]������A�׹{;��"O��7	"BRd$�@$V�I4"O���o9Z HZѨ��'�\`)T"OҐУ�r����tbĜ:��X"O���e�	T���b4Z1S�x;&"O������n)*����v�x��"O��{7�U��ȭb�aR�p�Z`"O��D���T���ы)�܁��"Ot�t�^��<�D �Q�r�@�"O�T��ʅ8_�z����*�r}{0"O@�j�,E8�\���;��ف�"On��D��V��a�HL�e��8�"O�ݙׄs�JUxw�58�\�P�"O�D�� ;w7�A�6hA�Z�:�r"O��ec;4�v���ܚ�R=x�"O�=٢�K�~j�B4:����7"O8����)��M��kI�pv�`P"Oȕ�b��*i���)���vBT��"O\��1��o��'�U�"ObU(S���$�T�������$*!���=8-���S�}�z%x��0 
!�dB�^b���/f�~��`�4Q!���&1̈I��X)6 ���(-VC!�DH�b%��fT!�Rm�gF�,9!�䕦]j�w@�>	��=�1��R!���8҅�F2��ΕdӼ��0"On<:��Q�~f�ҕ�d����"O��9��9��Bp��_��U��"O��B��ųN��"��U�~^�u�U"O�q��ć]X�4!Sn�[Vd|p#"Oz���t��5{2-��9:R� "O<��ƚ�w�x��잘r8�|R2"OD�n�}�䥰�lچv(�Y�T"Ot�D�5PxS��u�J"O(� fa�B�z5�.�"�9i�"O4|�,M�P��`@g�4
�0*"OtTUl /Jm� �QE
�x1fls"OT�:u���uh��Ѥ���r�"OX�9��U�l=0� ��� Vd����"OZ�f�Ԃ
��U�g���ja�p�"O�ITF��#�Fm*�F@����# "O��9f�����s�£}���"O�h�*$6pQ JG�hV��f"O�!��i��[G�H�L؁"O��B"�Ԝ8����i4i�p�S�<A��6�:�BS&=�2]����R�<����8v-��%7h�m�d�Z�<Yab[Y���¦�J���D$�Vn�<�b`��0Fa�L��̂D�d�<Q�%XU�sUON%'��۔��T�<�E��'H�@�j&���u(F���N�~�<	�K�;vn|E����"	��q�R�<Q�����,*�"
 u�m�O�<i�/��9�"�#�+T�F+f\�
]�<�T�d�� ���p�h�k�Z�<aV��0H��t�&)�3L���cDW�<��a@9fR"��ui���z�<�t��L�,,P���"0�=���1T�t�QH�;l���E��0c���J:D� �	� :T^��E� >�g�8D�$�EH�`�"�J�.�-�V��!+D��:gi	6�<i 4��� XjJ+D��Z�mB�j�1�M�o����*O� l�y���K�]���W�7���p"O�����$�p-ȄN�:���B%"O�\2UFS�tuC��F��Ґ�"Ot��B��>�X��+.����2"O�Y�Ќ�	j�tR d�
9a�x@�"O��?AU����d@n0Bhò"O�%q4�CX�`�0��\�IO�)K`"O4�P�ԅ 0�����B�DG ���"O�8��g�L9��J7o���"O�!����+�p�맭 VRP٫p"O�@�!�Bxr�ub�3P`Nla3"OLK��܈1�b!�6bɞ?�@U
�"O�ѡ���)P�=s@?5�΍z1"O�i��E�6M됡��E��S��"O�˳ ��q& JG��C�0�"O�ёȋ�8Nl�3�T�
~xA"O� �W���l�1��R'>�� ³"O�z4E <k��t
U���Mj�C�"O��I��Q�jش�#LP�`)��"O�+�,G�.��)�gj�N�:��p"O`$��B��<�c�ߟӲ{p�'�1O蝹R����(��ù�J��"O�0:�>
�T���ǜ����8�S�iȒN�`���²2[�X�v�Þ 1!��;h��˟�K;��q�J 6+ў���I�Oۺ���G�&��.(B�I4i��K����:�
X��Ӏ=�nB�	47.�zH	�ik��27BQ
S�rB�I4z�1�Þ#��l8���H�B䉶nx���B׫c���U@	.4��B�	���\с]��ց��	�%Z��C�I�Y��	�6���F̐*�H��yE1 	��V�"G�z��1�Ѡ�yb/C348�}rO�?M������y�jFg?Y�`W�4k�(@� ��y��Č��=�CF9}�}r�"H �yB�U(L\8����7����/���yr.�� ����cjI%#R��be�̹�y�gL�rLn��dMɘj���\_bC��;}��h��|�6�P"�,B�:B��&Ǿ}S���L�PA�f�)BTB�>s=,��3ȑ�1�$0C/6ZB�	�1:�A�@�pl�]��W*7�6B�I�bRx�˥�\�J]�d2�B����C䉪$e���P�њV��,S$eŧufC��^�P �4:kҼb�e��A��C�	 �ԋ�c
�=p��0��_
XF�C䉒��2��׽ܜ�(RH_�x��C�(kPt¥韲1<`P*�	oC䉌<��A"�p��nФ^�C�	7�&I��D�z�Nx�S�P ()�C�eW
dpqF�		���MK8N4JC��%5tH��i��%�l��'"ҁ'�tB��*p�!�0ybx�)���_$C䉈&�FTC��Ì}�*���L$-�B��	-���a��|�dJ��ȴB�7bd�p�E�Ì
ό���!;�C��(M̵PV���y|��@g�dC�	�e����s�ߝZ p����zxC�	H�j��.)�йZ��	�N�0C�IQ�} ㊅�*�L�0̒�/�rB�	�Y
��ᦂ�#�A��g�?u�FB�X��LKC%�X��a����B�	8k{ґ(� ٭++�Xk����Y�*B�)� �պ�@29Bpk�f^��A�"O�\ K� �0�7$ ��4�"O��C��W�>�.|%H���T��"O��7�ڔo�*<q��&>D�4���Q�a����7Cƺ1 �������	>24Ju��LG��r���1/���-��E����餻�H���Y����'�J��eP��*$"�d�^]���I?>V �,ʓ�hO���"�R�	U�k�X���Hޙ,����cœ@�?Y���B�j�D�0�2xE�)D�Rd�K�W�4x�_={<u�g@ @ݬ�0�{�T���A��L�5ŀ7~��F�0D�H��*J:@��\�G��1k�zg��O��[�)߰>�'m����ɷfk�0��E o��l����!\] ��Mޅm�čr eV��P�V��Z$���'��U#�⌬J@,���aZ���}�8D�t�zf�2�.	�����|7�x��ɜ�o�Z�ǌ�h�!�DΛ6�&��`�h�:Bl�2~�Is� x
q�� ڡ"�V(c��<ip�e�"lRAdM8-� �b���_�<!A�7Y�Ak�ҏa	2�R��>V�|���5$� �0֠��o*�+��D[�]xf ���M�N\)r�º��y��#L�FH"aB�������� s��i� �؜^��0�bb�'��*G��F؟�!��"'<�
#OS@�.����!�d��dM �+�bPn#$:�*c/�A��dJ��Pb����Y��V�Ҙ��yV�+��($�z0�T����(1�׀�=qop�z�M��LQ�Pi�KR�'*v���)i�;6���%h���#�"*�q�!)��r/"�T��n	"n��	*A�H�G ��U>
� �F�"S���1�� ���R��4d���W�B�LPC)O�)�&�.�5��
��fA`�HG ًҎU�� ���2F8UŜ��pm��_����4 ��`�ǆ	�s����0#�IS��= 4��eO$Ц Qi���ރBV���OFɩp�S�{�B����w��PZ�';��R ˽7ٚ� ��o�i�6�,P
��#[H�H�m���l:�O����Y�y�OGjF�\kюK�y=���ψ��x�/Gh�Tѳģ�"]L�+��L�q�`սN7� �eA��D"����і
�X��T��<.ࡰ�O*@�`�m��B��Dυ/y^�8R��9j�`8��ꈃ�����D y{z�Zf2.����ڹK�B���'�Oʥ��9g]t��B����:�����W�D1��ņ�� �CW��x�ND �s��h�V\<@��$��!r�Tv���yҤ�N�N�H�M��j�Q#���D��,E�#����&��5S�4�������P�>���w��ȠKӛT��z�aS0rp�'���0gF>����6"�,�4�(u,I�&sbh��h.~ɹR��W΂�QR��:�ў����VS28 cF	tP��u�&O�������u<X��@BN/9H�׋X�&��"C�Ē9;F��\�>���R��-0�L�D4�S�'%<����1{F�Txd�ǤWF�u�'������M���`FE���k��ɟ	�D��Z>�k��S�i�A�a����o#���<G	/dŲEy��)$�ᩃA�?t����L�"`��jb��:��O~*a�8��ϻp| �r�b�3��!��J�d{L`��p~��d��2Us�ku
¬e�lZ�*žOGB<��O�S�4�
v�ɤa�^��4DD3�?1�r�����	�Y�r��$͖>�0<�M�����m�����?�lb���6<
\�ZB,6'z����'t�Hd���hO1����-�m���L�8�<Q��>!�i�3u�)@�����x]�h"欃���IOzt��i�����Z��QB�2]0�V�d+<O�����5��5kVl����#�`�b�i�2e�jQY0!AB-�O��.ʃ
�b�'��x��9F�&4�j:z�C
O>y��+H�@ Py��IB�B���1,��$ T�6?�*��a�<bZ4�ҫ�������ɿ6�<��b�,:2���A�J|d��D-9:�:� ��Izh�C�jS7fG �ХL���Й!Hˎ^�veCFDP����.�S�'.jl�B���.��Y�E�. .��<Q��&���fV�v����Ҋ��j����&�+2���Ɲ�G}Z�Fx��'���c��03�,�z�g�=8�dQX�;��CLB+Fx�ыCk���(��I�2�<|Bb�z�$)�E���+(���\�t�S�f_"g?IJW.��]��oڎr���SԌG�H�̍�+c8�,y�K��<�J��R �:�dh3�;�Ot���ݒ4��cR�AY��$��x\0tc��$C�)� �i�J�P�9�׌��!!��ۦ"OYR�LT+l]�6%�� ��f�<�bDP8���� A]P��[wĔF�Q�7D��"g�S3a�@LH���	���ء�6D�hd�JH�|�q�@�+��Q��7D�h�`P��r�i�l�$v*����3D��04�	�|v�1#��J;�H���uӤ9��)���$ r��l#R�T,FX	��a2D��iƤ��`b�� Ri��A��P3��/D�@cf��;J�n���$7R$�<b�h8D�p�Pi�?8��;��(�x�A`7D�lqA'�$`��`\'��,y�'D����#�q�<4k���l�rXj&'9D�8h�B�(�j����̹78 	��9D��!�E�1exTXCd��$D����3D�d`�A�;�4c�HF+:`�$�"D����P )I� :C�
�N�~��"� D��#���'�����.�F�lu!B?D����%@�p����l��U�:D��� G�fi�PP��d�3¨:D������P�9b$N
H�f�ڳ�9D�tA@�A1�Y��H:�nh�"D�|C��	�j����@-F!�L|S@>D�pѠ�_�5�s��L����w?D�����ƶD�D���B�&Ԟx��.D����
<4�4����G5 P�#s6D���A��J_�"$��:F"�|X!�䀒E6}���F�+����L��M?,Q�A�JqO?�ʷ+�X	�^.��%H�i!�D��-+t� ��,:���Bǔ�Ya}B�Ωu��D��v���Z�旅P�4���7��awn].�HO�����O
��u��=>���N�>@��"O���i^3�t�p�m�<�E8�"OԕS�c�T�X�;��`���"O��ʃ��3%�ne��*�hL�"O�`6 ����q٦ꙸ �-�B"O��+d��:�Y�ǉ�z����s"O@]0䪋�V�zX*��f|�xRQ"Oxp2k��M�4y&�߃.5���"O�\P��U'=�N�j��b&Ĝɖ"OH9r	S�]
\ a����v!H"O����!+Vh�'�D=`_@��1"O�HhT��`T�7$�"%���1V"Or���I� �sWb�(~�Vi�"O \�G Z7F��aZ'��4��"OSsB�r��k�7A~����"O<��B��C|��,N5���"O�*rc�d}���,4��
�"O���GY+$t�1���!60�I�"O���I�[�`���(A)ҡ�%"O0�xR	[�!�Ա~F̊""O�E���0D=��J �ATl�$��"OŰf�3`="�\I��T"ON=$A��{��D�.6�1�"O>0*�J}y�/ȯQ��H�U"O�E������"N�3TH��Q"OZKf��?b��aPW���zb�G�D�<�LQ�h)"�I5�N�L�,Ae�Z|�<ɴ�!�T��"ǒ�i<f �GDG�<���$Cɸ�W�/6(�x�D}�<Ig��0vt쳗�MD0����\a�<1��3A�~�#⡎L¡��^u�<yC'�T7��j��){�w�<9�"E�	��L�SF�E��R�MJZ�<� D�ۆ@O6@�����0~�����"O��eFV4�8,�c�*U��5y�"O2�:�`9pa�qK�:h}�3"O^-	��_Y��ШF�I(Z�p��"O�y�,�j�|��R�MlE�9�B"O�tH�[61�~���S	P!
Ly"O�d�#ł;�JT !a���lL�B"O\e��`���f�� J���1@�"Of�)�M4! 0�6�ێiq�0��"O��Y戓tо�;��Nd�i"A*O�LhwG�u�rH E��Z�*	��'�6�ٳj��8ܠ��L�&�$\�
�'Ll�i��� S
2�8P��.�IQ
�'9���E`�5+�~8Ѣ A�� k�'��\{�ҪI~���-V�H�#�'��8J�E�!��M�J��1ڤ��'��B�+҈QoR0�q� 75|��(�'d�ԣĕ^�P�2�H7)H|��'u:�)$�8 ٸ�aE�D�)�\l��'RBhKQ!G�@U���,�B���'�1JV��h&��{D�^
i���'\H�r�؈?1�ѦjR�f�
`I�'`�q�f^��t��ֈ��7��#�'_��2#��w��ܪ�-]���X�'h�$8%d�	��P v����60��'�|�Ʌ@� T8���T�L�dDݫ�'�`è�,0�觡�<c���'���"�I�1�ld@���#/t0[�'48���J�4v���8���:1Gb���'�>�8B�J&o���1�Y!0�`s	�'�����#ʳ)UBi9��_
]��Uc�'VaQ6���),��@'S�_�`
�'��8wB�R�d��T�L�i
�'=�)�f��Ơ*@ J�@���
�'m̅+4�� d���+��B3�-`
�'B�]ptj}st��f ��;�Ё�'k�4�V�;TL��Z�m��0�&1J�'-��Id��.��p[ (�PF�9z�'��t2�I�8u�]��Y�~��X��'(��S!�ԔJw
�
Gr(�${�'.�����p���b�a^�+�'�Sg���{��3j"0�'�
I9q�1�"��B�� ��'t8:��ӼBB0�jq@��p6��'$�H9���%��Ѱo�0F��z�'.�;�dY"l+��[(>���'�d�0D�aдA�c��?�μ0�'�"��	7�F)U����Gz]nC�I�B��[�IX0.� {��\�B�I2��a���O/?�)p-��C�	M(N�����Vƍ!��;o��C䉆��)�cP�C,��`'`�=w�B�	9{��=X��Ȗ$��Sk �`a\B�	0��yv�������^B��p&F� E,J=d��!�W�]*J(�B�	�nX]C�8>�����2��B�I5�qc'����9�-�z��'��u��̏/k	f	�J,�4�'� ܈�ş�H�Q(�j�;2#�A
�'(�y��'W.z.��X#�����<�	�'v,�"%��pjj�	�h� �`���'�T���`M�nO�i1�=!�D���'�j���H�f3H�� " � �L��'B�M�@f�b�0a�D�
��� �{D��5sK���%.ŗ�Պ�"O���$`��N^��8Cm��>��
�"O��@�jA/<�"A�L�1K�$|��"O�(Ʌʼ*��LC�N2 ԈF"O���OX�+��pRTjŬz>NpC�"Oꀉ��]�%!"U�DX�`��"O��a�'�4^�b!*`���h1�"Om0���E���a������8�"O8咠bK��:aB5
ļS�d��U"OH�zÇC�r� �S*٥�x�xb"O��R�M�b$������E�&�{�"O|XbЦW:��P �[#S����u"O��bQ�:A�Ó�T�(]
�p"Oԥȳnŋ���� ��hQA0@"Oܑ+�ɪB��|H�o�:�� ��"O�,�	��J�&(2Q(�-��qQ�"OL4�%�[�>��y+��B]����w"O���B-����C	l�}"O��b \ FlXU�&S� +rq��"OxÒ��:��1j�K�04����"O6��EC�y�0HѠ����hš�y2&�����w@�!~��������y�LM�f������aD%�y�J�!z��c����M� �B
�y�AW9���K�ʋ:�̩�p,M��y2-�)m>ZQ�DS�,�N�Z�M1�y҄�(Y���a��˯-�x��+�2�y��I P�d-��fN0HИ���X*�y!��r1 ��'N�� �Z��yB���v
�	;$)�(_
"-��G�;�y"J�|���ybi� �������y�%�z������W]�8j��]��y��РyD4�(SȡJ��y󌐱�y�I5��q�%+�2�p�òe�$�y��	f���
�D�9����[��yr-`�Z�8��[��^���o�;�y�K��y,�S#�cT��&iS�y� ;/�������,����\��y2[k�y#i�>��Hԥݨ�y�x�B[ Mni���C>E����'�$4�L�(.D����43���S�'�,�I�j�+V�����/���'��&o���|px����ީ��'MB	ҭ#pO�`��N�ԍ[�'��[2@�+SN��`�A�bG����'4h���X*r�$!P��Π6Ҽ���'C&ԯ,	�f�z��P0y�P�8D��P !߀cl�|�����Q$�-D�P��L�*>*��s-�� 1 ���*OJ,˗�8\@���E�2" ��"O���ee��"�8a�@8�p��!"O�K�'��t ���J�T�3�"OT�R�M<I������:)PU(B"O΀� �		j���S��X�:�"O�u� ��9+R01 hB�*�)��"O���F �"���?x`D��"O�@0�E�<�r�*�b�3j�t� "O�-rRB\����aa�:~�~e��"OZ87��>n,��!�1 ׀�("Ov�5�i��Tq�ͤ~�^i�5"O2���ڋ[�����Q|�l�J�"O�%�ǔ�k����'ƿs�B�ɷ"O޹�hK"8=���'�b��-H�"O���/5c���I���:0��D"O� pU&*�4�Xp����'#��yɂ"Ov)@g.��{�t9��HŊa�"O
�ȓ�I��ZDCp����4�	s"O�!��S� =>�C��$��"OօI�d�v<��8���;k��|�0"Ox�#f��;K"�M�%�1��i�V"Oz�����9��(p�)Χ
ü�K�"O
	в�\��ݹ�g�2&��0�"O"A�I�rth|Ҷ�	)�*U2�"Oz��a��z�f�`�_�r�
���"O��╯�-�~��d뒺(�V��c"Or�[1*�*6~��p+5Q��r�"O0�t`�?� ����~=��"O� a�6 �Ll���6-�� �"O���E���T�PZS#�5�V�0�"O��#�a<]�t84$K�M�`+�"O섊@�6�$#c��5�r��"O��Fk��2��s�� ���"Or�ѭ+L�����aV$A���v"O���m�D	И�|(���^%�!�䍌d��uYg�M�X\��@o^8
�!��ժc� `��̊�v��!h��O�!�D;5���Ϗh��!k �%O�!��$5 �]���[,�h���J�!�d݇>��̺&���W���ԼD�!�D7A�.�1�.@�X���ǬP"1k!��'�!*�K�>5bhL{�.�'�!�D3@]�1�����,:��!PF��S	!�N�,HLDZCH�=<���uF�g�!���B>l��@  P"�xӂ�"�!�$V)�����J<J�pɉ#K�g�!�D�@����PO��+`d�
A�!�U%8�TA���#`�PdS���'^!��.�MPR�TǊ����M#b!�d��R��F (K�FL��N�� Z!�d>��a���.
~�s�� �Y�!�F�6ʬyr�._<o�¬
'KL��!�$��1�@�E�N���U�ˆE�!�D)�zՠ�� �H:�ı�IъO�!�Ć!p�2�+F��^$ܑ0(�2e!��H�9���jU�3|	�M�4_!����D�F5�$�a*&OH!��.vI�H��D�;Pa���΃VO!��R����",NH���H��9!�$O���"Ce���sEsC|B䉍V�\-)�R��j�����PB�ɶ��q+���? ���%�9NnHB�I��r�a�e�?,�Ȇ!18B�	�;�P����@�J�>��B�0Q�^B��z����@��>��K���laXC��NŰW�o��D��;W\�:�'��[v���"�,%*ꂺ)A�5Z�' �`�&�X�#�>����A�.�&IK�'�u�`�/
^EC�+��&v&Y"�'~��\��{�F��2)�
�'���!�� �&9C�.P�H	#	�'��5z��%
��H� Fت�'��:���Z`�CW@�h�'0�U�'�U-i}���U��-`���J�1�hM�c/�@����'LA��6�����Y����UR} 2Ա�'TPy("-4�)�iD�3�	��^� �z�������v ��8����f"h���)�$D&xP̤���~�$ �O�>Qrrn�%J�ΉQW��Bp����B�'�TX�����E5+��諤�.:aؓ-�d�^P�?�?�� B��6o�>3�X�� W�Z��؂���-Len㟒������<=����%�%�!���>1�k������O�j ���@�W�ꄐ�.�2k�*%;�'`��D��S�5��$��Q�r���5O��p��uS�/������s!�G���i�)��G���Z�k�|��_Jx��K�O֕1D�Ϻe�Љ���r�A=})��$;b�s�~�SD�ӑM����_C���D�!OU��Ʉn����� '}��h�l��ek�,���C�([�s�e�G�ƈ^��l��(~�S�OG<��S��1������,t�!r�9�8㟢R�͔Q�z��D�&+�fP�@P�E!�O
Bç0_�|7N�<o�N�y#�-o�d�=��ַ�?��i:�6��Q+ɼhc͈��	?��y��8�����\�[l!��뗴$��A!5�ê�~r+�\��O�>��	��/�\�5�qu~�g��P��lr���i["kl��qg�ȫ��U���" ��!�?Q 5�T���L*M��ay�	��sX��W��9 -D⟒��b���q���)��ۼO� ��$�>�C`7����O��p���	�P�
� 6�ɲ �|�k�'L:�BE�%��~*&��2 �~�cc�Hi)��:b��&�$}ru&F�}I��
�'M�a��C�V��1�*�v�"Th�'��[�LŎmY�X�ec3�L	@�'�X�r�3��-k�f��y���'��A�"H׹L��t��k�4[fPj�'�4*��-K��prT�H�Lt���'L�Xb��@��d�-|T�颦/9D�Z�+A�r���@��IV�a��2D����X�R��,X�-�yBV1H �0D���¢K�	UA�8j�4�R�*D�,�S ���M*c�E�dD{��#D�����E�>f�#���.��s��+D� Rg��x��|��eNp@t)�(D��Z*@�^����(��v*J�ZC�&D�0�oW�5.��rɜ�p��`�u�%D���AI�=0���Q1B��rȀ,i n(D����k�"��5��Gv0R����%D��X`��@����WFʰoKH�s�-D� ��,�9C^y���9�k�&D����ϓ4�r���]��!�d*D���D0	�9@���6S���A�&D�(��jQh1�Gf��逹	B�8D��냷T$�j_�1��8d�\&8�!�d�t��(JW$��7� �I����!�dBU�\)��J�Bܔ�֧EH	!򄎽
!��0���dˤP�E�F:	!��
� 1`�_�Y�1�1�ʌg�!�ě�y��}갆ΘQ���1�ԇI%!�D1M�i	�+Ǚ.�H��@�"*!�$�#��
��6.��Xc��7!���9I����>s��� �
�k�!���=�8Q�$j]2�c�GܬJ�!���d�(� �uS
�!��\/%�!򤁈 ���ბ��:����!�$�%4F�H[��T#!�|�V���	�!�D�H��I�1JՓqgx5��JI&=�!���#��H�@$Y ͓���!��$.��yKs��|Tt!Ec¹3�!�U?8�ZAsDC��u7p���B[�:R!�ę�0X��uf�^)$l+�˺h8!���Z�T��m�>2�D���	Q!�d��y	�@�5�#�U�$3!�$Sc��%k𡁬t���HR΂�{!��Q�-&� s��C�}Ҫݘ5��C�!�dV�D >�ㆢ Ӽ��\r!�dԏ_�� �1o"��+�2pT!�� DP	G�6Hl��W	P�p$i�"O���`H�%�|����B��	�"O촪��2%�5�&æ ��=�"O$���n���� (�<p:�"O"�#���o����AeفH�*�R0"ODYR�$�%Ip9��+�0�s�"OD��$�:K��On�"��#"O��-E�2�I&��-3��Ѻ���yR�=OeD�X���=,y�u�R6�yҢ�R�A3d�#iX@��ֺ�yRG�8�f�åjZ����Ԧ�y�V%M�*`���S
S��W���y(�8b�H�@j4LL�br)K��y���/�&���!��Cڤ�������y�$=�<��+ ��	`��!򤓺P�&�ðCL�k6\��n[�P�!��R?3�.(�DHQ�0���gK�n8!�Rq��O����Q���1	4!��U;,�D��C#&{J���w�ל32!��]�5x�������T�V,�Q@��\�!�$Y���T�Ur
�)�O�5�!��:��p���2n>� �C""�!�N�8*�pxU���n����� �!���m@�%�3_&ĩ���Z�!�d�7|1���͉{������R�F�!�D�����դ��{н���e>!��d�U��+�U����P
�P/!���GT�(5�8�J5�2#�4!�$W���,��{����(�n!���W���XD�8�d]H�E/c�!�R>g���v��'`�X��/?�!���	���:�& *�}R�N(x4!��]��9!�m�8�,�W��	1!򄉸hg��
��L�i�@DC��!���^����[�0(	����P!���[����*�;\��Q��J!�DL�OZH2��/N�A�c(�4M�!���x-�<�ÑW5H�Krl�5f�!�䅆��0����:q�d25�O�!򤄄SO�y�Ƥ�#������1�!�d�DLT����y��%�ϊ'�!�$�1��!`0�S7d������'H�!�}��n�6@�P���F��P�����'�����LC�i�@��S�F���'d����G� H���)��^�<�6�
�'aZ��#$@D�\F Y�%�60{�'�f���� �5�$	���۩M����'�<|Q/Y'+����$P<v�x=�'�(���Ζ���{e�W�s� ��'���iO�}� �R%���9�P��'̙a.�W_��K�����J�'�B}�󨌀,y�AЍ�VQY�'�~�J_$N�{ËU$~)`фʓbD�hq��iZl�@b�H�|���^���#�e�9�@m��ҁD���ȓsOn,�F+ۋ �Z�{���x m�ȓ1V!Y0�VX�֐;���1-%��ȓ�tH�ҡW_�TCA�Q� p歄ȓ">(X�4f'XG��e��#S�p��B��Ev�ͶU���D��v�P�ȓ"Vl�f�ǘs�p�
c�Q ����5���Yb,S���&mܫS�Ĵ��
��a�$��B2�!`d�@� ������,��QMF�� ��!]�|)��S�? R�ʅK����A�D/��Ӧ"O@�"���&6�؁���!,}�D"Oʍ�'��1s�N�PD�t��H2"Of�BP(R7vh07!��.���"O4	�/L�`NZ�E*1�P@"O�)`)�B�.�@$V�j۸%:R"O
���ZCt�Q�i�'�x�r"O*aSҨB�7 `e��-۷�:� ��d#�S�OLP����R0DV ����̔X>r�'�z�h�O ��8�bQ�<^c��*�'����Jђ�h�+`�F�Z�'Wz��Af�#A�����Ȓ[����'�Jѻ�H�)l�iia�[����'�r�i�@K2.�����K*���	�'z��8���#�3� O�ܰ		�'�n��&P�,���$���p�f,h�'��8a�e�rS�j����'�Ѡ�JT?���KG��<`��9�'Nhi#,��l	�)9�F�06���' P�r�!��������{;|�C�'wHl � E.E�(�Să�N�A�'�f�Tj�*(=�`Z2i ""�t`��'��Uc5L�΅R�#k���*��yD[y��*�3ޒ�;�K�yr Y%a��xA��tQ4c��
��y�F�"��h����>�~U���y�ۉ�Lِ��"����+͐�y�hϋ1���c�����(�����yb�p� LC i��~��� �Q�y2 ��N84�[�o@,<A��O(�y��N)&aF
aI'g��	�&BQ��y��ȭO0
���K�nj�L9����ybň�
�� �̒�5|�5(���yg�3
.� ��B�+���pB��:�y��M%�Z �tiX?2=�002���ybL�!���Q�ʼv�N��"���ybM�5/�x�bj�$v���P��y�
W�6��`�0V�u��H#BE��y��ÑtQD|q Fmu���ro�6�y���R%ʐ#Ɉf9(��4B��y�gE�l�6:"Ȋ[�θ9��ӓ�y�HO�����$*�[f*ٰ�Q�y¢�:��`փ9nh`��$�y���j%Q�B�0 Ҟ���K���y�K��$����1��1}�V��/�*�y2�@�7�0�y��O4_���3����y��;_�<a7�$vX�t(���y���S	�踂�H/: z��S��y"e�2 ����eԑ
ݖL$!�y�/�,4�,xZ& �{|h�kdŔ�y�B��F~�U�&䁪%~��E��y"�>N� X�K0P.*�!
� �y�k��(P��� �Ǝ9>�B����yNL�'f��1�f�*� a�p��Pyr�E-K�����T�}�D!�#)X`�<�aS�@s�8��ʴ&�P�J�d_�<�b���o����KV�p�X�"�mT�<ac�&��\R����T9d�VM�<9��)%�$P!�ֈ�0�H�*P�<�*��U�Թ�f4�L��"�`�<����R �b�İF{>9��g^�<ug�D� 3��+R�
 j`�	]�<��B!�Y�g�eh$�!$��N�<��h(K4�����&?�ċ�K�<� ĵ{�L<�li��꜕G���"O�u)��2�4�wJ�+c$�Ċ"OJ=�T,̶7� ����]�)rH[�*O�Y`�AZ4RKą��ŠV�8)�'�I��jJ�J�1��R��b�'6mK��X�<�Th�n�;����alN��FEf�(�� ^�@d��/H�YȖe%3~|q�'�2;����X��к��?@�,$�������ȓp*�4�0"+2c��1"��(���E�]���#�lyq@�jE��b"O�i���R�#��X�Y=-�"O�@�2�� j�l`j�S�"�� �"O4��"&��@�S�S0��2�"OZ���c\;,
�A8
Ӥx	n���"O�l�T��r�)���\%y_2���"O"�P헇>�`�3�h�FM)K"O&��E�Y� �W��1-[��%"O���$ �[�Y�'��bJ0�"O���	�)Th�2�&(&��Р5"OXőM��qC I��R�P���"O�4�3��. d.Idk�����"OL쀢Ê*��!$%�6���(�"OH4!�    ��       �"  l-  �7  .B  N  �Y  �d  �o  �z  ́  Z�  ѓ  Λ  ��  ��  ظ  �  c�  ��  �  p�  ��  ��  2�  r�  ��  ��  : {
 �  G �# �) s0 �7 �= �D mK �Q �X �b �j �q Sz Ԃ Љ � W� ��  `� u�	����Zv�C�'ln\�0Jz+��D�/a�2T����	#Ĵ1%�9�?Y�� ��y��%+���Ɨ�Tvv�[U疟bhd�W�N.
��&�
�ct\�`��խ;XBX��'T2����yj"����� )< �7�@@t80{���4j�8,�F��9�y�B�%�,ɸ4�� �T���D�D,P����22o�L��@�L���2)���	>�n�Ǟ)A`�XٴE� �����?���?���+���-�1to�p�j�@>�iR��?�6)ҘHUX|�-O
�dϛu�$�9OD��T2m������i�-��
���d�O��O����O^1k��i3��z��_>g�)B���C�Q�!��;�a"v�]:8������qxP�	{6��fc�,!D�H�s��*�a9�W�͓��'E�h�C�QRa�1O�,ʳ��O�����A�j ���'��'���'2��'��P>A�;<Z�`S��+x����ğ�]��\�ə�M{c�iA�7M�����ɩ�M#��U���&+�=�DP��٥>K��	�������S�R #=��_�O���b�&g����3� N�������	4.�]r���iC�<�Q�?�?��i�~7m��Χ�2Yw	<�3ԍ�.2�y��GшP�,xۂ�i&�E�E�Q�	���/�o��l���9J�!
ަ��ߴ��I~�
%hf*�9	�.ܪ�`�3`�Ћ��7`�P��p�b�̩m��M�PH�0a��txp!�_k2	�DԼ7�Xt�piʖ<���0u̎�
�(��D� ��l�v�oƛ�obӎ�nZ%KШ�W/��c�z4�P٩X&>eh�"_�_vJid%B_ py��)�M���*U��qH�+U�0p�{׈��?Q�Rj$*&bP!Q[��x�}#6mX�aR� ���'~6�����iD�_�"T�%$�o�f�DU	�2��Q��h�Zk	��*��'��	ȟ ���h�����5�RpVcV�M�8LT������:,冈��ꕈR�sÓS�(Ƃ@ێ�۴s1<E����K������G�`��0g$�0<٦.PCy�B�<AAA<;�f��b#\3`H2y��E]����	埨'�|�	�X�'��;z�<;�l�UHEa'̅7DR�'���l��	��'�������O�䈳΍�}"�`Q�M�yπ��4�'��	���5-xӜ�D=��ӼahS�ݸX��U�'���Ī�ϟP��g��Iyr+'cؐhq�4>bb�0��T��B���L˩T�<�J\"��c�>�y����ӃfN�R��S]�S�J����I�q���N.�"��65����M#��|R��S�_F��EGB�z����g��A�؟��	(�'O1��-J�F\3=��y���?��3T��؟��ߴvě��'4.6�n>���-@2)d� �)�u���Ђ�ئ1�I]y� ZX���'t��'�	 $Dz�9����H"�S��Y�V�� ˆ�M{G�O�%�A �R�����qO�U�#�Ơo<J��BH�5�$����!��3�� /D��s):[�1�  *�O�<i�Sg��U�c�Y(2~��Se��M;u^���C��O���$&�����x�
���L`� Cf��}�'�ax��+d�"܋%+hBIŤ��?q�'��&�i�\�O�)��b�J��arIG?���E�`��;��X.�����my2W>%�'E�8�P���
!.:�!�b�^���f�'�,��_�M˂GFi8�p0'��_J�����(U��%yHP�h�q��5t��PSd�V�f���%GL�fjQ�Lp�&�)
up�Z�_@i�ƀ2/���릉z���<q�Ob)�w&Ta%� RBn -�!��'k�y"�䖑M�R�je'�j�\�
EX4�d�����5;�4��醈Z���n�L�Eb�P���5.�f�) m�=�f|�IEy��'!�?���:5��H���G�b�,�s ��6��eA��Q�9�pԓ0%�}�����B�>�Zph�A�O�!J�h�F��-�WIG�T�@��A�2� =y��թH���`���f��'G7��O��ڲ�3����v*@�x�R�<Q����'�>��L�"u�Θ��)J,N��A�6�Ih����dm�t%�4I����`�.Tؐ�!V�y�'�m!!�}�j���<��'���.�����EOq���G&_)��i)��?�����L4E	��ЏdΛF����!��#Ӥ]S�HDd_�&Ϫ�K�,(?mJK�D��G*(� �P�O��Ac�дͅj��	�U֍� $ۙ}� �:Pl���	�2���$���mzK|Ҏ���&BvE���ٴo
��r������?K>Ɏ��i��Ĩ��J�D���wp1����O�Un�MSO>aT�v�QJd��V�ժ�F�`�V�'���'�2 u�3L���'_�';󮑖X�ر��,S���sUHOjV���TE�]�qV a�4�uS>e�3�uղ�H�� ��M�w䍨<F �0D�Ֆ4�� r畋p]���ʂE�Z5�O@*�`���y��
f�h��7�
5d�zp�4�<֛�p�'�~p:����?9��?�� 	.0���ꚒR!td�'�L/���?9ӓXf<�;'C�EθR2��I⟨�ٴ{����'OD7��Ol�I��J˧��=����:�L	AC+"6h�u){���' ��'��)��,Z�\���!؀;�u��	dނU�w…p±ɴaQ�;���qu�'B&L`��3=X�Gޣ�T�����-n�d�y3��k8��n��[s�㦈�j^y��|�蚐������0A��d�=D�|�p��?����'i>�b�[�7 �8IPh�0 !A�� 2|O�b���Sf'5B&Y��+�	G�<�b�"������ISyB"BPN�7M/�g��
KL�t���y
\+`#ş�'5"�'u�X	��#����3��`�ҡӇo*� d�����m��A�P�nM@u�'���!Go;�
�'�7w�x��Q�b]T�3ц�<�U�	4�9)&�Y� JHh@�|r�Y��?)w�i�P�f�x�Tm	�f���SuCI�]���$����I-s���w����,��A1}�6��8��!��|���ieы6M���H 0��t���r �pӒʓ'<�"��i]���ym+(�bY�3Aϊu�ȽB6$$X���'v�d(�6d,���wɁ0����3���U�x�pu�ϭ/f���I�w���z-� � (� ����W�%��yȶ���ڠ@����5CM����	�
#��В%IK~r���?)�i�#}��O���3O���1�6������DH>r�r��D U�rA��0�ўL�I�M�w�iG�'8�q�P�T�6�P�ۏL�Z� d�'j�P�蓠lXퟬ�	p��zyb��;��}a@�_�(�>x2�k3O����S<\6Q����=dކ��t\>��3�1KcD݊[h�ݹ�'VQ�ш�$*5����`R7"ٌ+_�ĖO6����� �y��ŰN�&}#�\�b�8R`i\�T�v`�<��Ƒ���a�L>�*�6��4���U \h���T������OR�D�O@��Г&���.F���	��(ݒ��'��@g�֝n����a�4��	�ʧ4D������!AK�.�.@�&�{u��H�I���?����?�Ѹ��$�O���+^�|�����J��D�F$*�RVu�j��ac1��{T
}a2(��O�ޢ<�Vk�XP��!��(���x��*����6E�)��-[bitښ�1��"X<��<����:w��Th�V�$�XL�T����(����?qt�Q�Z��{���y�&�I�JI^�<!v�2�E ��[��dq�#�W�	�M�J>�7��>��S؟@D�X4"��Zd��ˍ��I�*Ͷ��ϟ��'
�x�1j�)DBhI��3w�b�%h؜S(H�M޴	y�s+��l쑟�kfW�Y�x�I�m�a��jtK�{ت�Pnכ7]R�!g�([� �˄�3�100�9�I�2�����O
�W��)����P��h��#2�7�Op���ꇜ9���{Rꇧ&h��1B��*��|�s�'��� ���D�`�W�yKR 2���$O3��)m�Z�Sc���'�x}�A�C+IAn��hO��B0ڲ�'%�L+O������+	߲�Y�$5IQ�H�A���<w�#珜*��AY�G:?���):l9#1j��m���D� �6��0^�� �R�'pC$��c�;;�1� W.���'s�1��L_�--�'�����d����`�N�[�"}�G"����?����?!���=	��&G�0�l��4�éў|����Mӑ�i��'	��Æ�E�?b�CТU0��!y����<�1F� ��I�4��Ky��	�:�p�0v
H𷅖j�a�R,^"˘Hp�ȟE7�ɡ�_>�3�I6!��ѵ�ޙTX 3��K�L<�a*B��g�r8��;0�j|��f�$O$�O�(8����y'��bٞUӵ$06�P�AQ�؄ ֛FG�<ٴ"L�����w�L>)f�9Wi |��0y)"�Зj�)��O\�E��[�l1�``�Ƅ	=�ؼK��� �?���F����|� �O�i�$�yrr��*�K���4�A�ЈRs�n����'�"�'{�)�����v5dG<i3C̞-b�0�5ʞ�X+0�ru暯�}��'␨��ʝ�TK
e�#�S�=��u��&i�΁�Ղ�?7��5�P�T�X��L�c-JA�p�|r,��c�,ɹ1�!6�"0�*WN�{���?����'>ҏ��.�����\'V���T0|O�c��3���5=*@2�����b�,�d��i��Oy��}i��'�?���^�Y���yV$ġ(qJ$p�a��?��-И(��?y�O�\q��K�*
l�rǂ2c.���*M�_�RY'��O�*�`jޑ�"?�eL܊w���U�Le�bpie��5I�!���R+L]�e┮R@���	�m?r���O��h���b�GW2jv4:"��'p��'�|��I����R(L�`
��Ѥ��L������܉įti��8sĎ�dC2LB�+�OX�U�]�0�i�"�'��S)�f�I���H��5O�x�+H:�h�����VZ���Ң�ʏ1�>\��(O�x��	=��ϻ��u3dDҕ,�є!U~,��Y�Y�/ǌ�!P�$%Z�PH�QC��<��O�R� ���J�œ'��4&n����O
.�?�ŗ|���^�v�heVv�`�s�Bb�!�DE�[ۼ-!R���{�� �&	�y�ўX�	��HO���V�X
=y�xՎX�^�P��A�ڦ1������جp_���	韼��ż�π/e
�ۇ� �7��X���-bܜl[Ň�"NH�@c��A�eCja�|BI>y�@Ѝx��Y��J�(�q���ƫT-�I��!d$���{E, �|�H>y1
�XmΥ���@�w�J8����t�J �	n�g���4�l�|j|pA�] L-N<�ȓL# ��G��*�d�1��y�t�'�T#=�'���<]�!M��'Ǿ(;J�-/����������?9���?�1���D�O��?*5��K��;FH�(8�l�F�� S�M��(b�a�H �n�̡� b�⧥�6$=)
��Y�RPJ�(�-T]��ې�߻7?tE��/�@�l�V��l�&�9���}�ݙ��6��8���O��m��HO�"<q���1�Z��I��<I���VX�<�kʖ
��	p�(9����A	I�ɴ�MK����$��V�6���O����+)v�E{�@A�t���G�����O�\i��O����O�I��vl�E�q��$��2/�d�F�a��p�f�B�!O4�Zs�8mD�됭�%yr�lZ5Ui���j�>�u6;Dи���ԷP�b�'��˓#s��`B��|�ĄA��;�Q��Οx�	Q�S�Ou�|g��{�.8���| ��/V���L�R�|`F_�e  J�N	Gb�6ͷ<y�@5r˛6�'�2U>���d�ܟXz�!z�R�����AK"��`m�؟��	�g�cW"�":��(�DP M�5�'П��^-Z�1��?o�l��f;7��'�������Attq�62P���+�O���`N����&o��<��9X�Ă���(��D-!V��'��>�ϓ[3Z̒��8 �5iS'΅M`�ȓ$���#�lJ�#��u��� B'^F{��'v#=�̗PZ\ K�L�v~�)2���V�'���'��Pp�B��+�R�'w��'����&��!���G�I��}�5h��uְ0�PmRS�@8IY�a���X������\�	�Wl�< `��!T�t0��ME��iƤF��#`��@;�ݙ6��cz�''�vT;��@�3wȣmZ��yŤĄQMp<�Dρ���޴�?� �	��?���,O4�i��P4:�����z���cxKN�˓�0?�q��DSр�>)� ŪpH���̓�Msw�i�Fg�pʧ��)��LP�G��KAƴ�Qh\�;���lJ�qX�XƤ�O����O��D����?9�ӪZtJ�3H��	�+F�y2Ä��^E�gI��P&�8|ay2���5�8�4BD3^ h�+Em�P�p��F�;tH����X'f����d�
w�j��˒�3`��W�W�y�����'��g�(�d�<����'՞�ڣ��e�`C�g<�ұ�V������v~Hy�7@�z�@	�E��5HRʒO�To3�Mc/O�R�
���	ߟ�{���`�4d?U���`���	),�m�	˟�ϧ'�� ��:r	�ag��}a�XPf��0���ã�1�B��Ί}���T���(�xeeK�X9���d��(QJ��E�_������h��m�����oP*#<���䟤(M>�@�? ���2/�&Z=VX�/�C�<��G��Z���Z��\�`Ջ��Y��lR����@�!�4Z�-f��d�L�&����3�M����?q(��1H���Oh��eO� �HP�	Q|E�m�aJ�O6��H�"��7�̪^�KL��- ��Cԟ��'7�H�f!<����)٪*����'?�50ߴt�f�[U��6>�x�)W�~�'jlƠ��LH�A���S���t=�'�\���8ɧ���F'F�yk�=J��B����"O�0��|�
Q���	�)K�M��	��h��$	t �k6�ѓ��TSe�Շi����O���J����*�h�Ov���O��$���<;��`釃��\#�A@,��P�P��h��GL�����
2��c>U&�x�'���k�0��t@"�i��`���hŔ��R�G"�c>A&��gP�T�*)��ᄒe�tp�#
�O��&�~��	�X��d��APX��w�9yg��	�o��*�΁*�'��}�t��F|� ��ҽ�>�1,O�Fz�O!bP�p#��ό��c���$���+F����P����t�Iܟ��	�u��'�'x��0嚽n�!1m��ENE;@�X9[<�֏T;4Th���L2Xs��Z���ЧI���t��(��1uFm*>�kw)� ~�
��A�h� p5g�', �[4�ȉUu���bO�t�<�ܶ�?b�iBўlExObG���Dc�ı�����hO�����|�@ � S��r�O-j$\��OX!oZ��8�OsBl���'���'�P�j��y6�*Td�\���
u�'���E<DI2�'��N�N]�J�c�7k��\tK��D����*2��H�A�������%�*�&��@#�oP��5�3$�:|��Cw�YѬq�. �`O�"5�A鉺	2�T��� ٴ�?I��(Q�=��N�!8�6��(T����O�⟢|B��6�tL;W��Ass 	Px�<�ɯ�M����`��'��$S���	6M�fU�t �`��(�d�O��'8C�T{�ecn��A��!|`��ڏ&R�E���?��$�.�veaCA҈jC�)�����)��Ȅ3��@cF����B������]J*����E(J�&`;"
8ڧ|B�����,�Zu��#�7P���'_�R�Fx�F�=�'��cMø	��q��kFs~��%F4�y�DԘ�<	�5	E EZ� J#��O��D��*��l���;:p�u�HV�	����ɥM=<����Gǟ��֟�I��u� ٛ%� �� �49F9"���^=��eL�d^8�T�����$S3J�襒q�w5@����%���F�R�-��;sQD!���� N��c$�~��!�o�Ԡb��'t��	:�Z���O��=1�a�Ȯ��s���5-E�DD��y�����M) �Q� ܢ]`[;��D�W����'/�I�����D�T�Qn�+�Ԅ*2�92��.�VE����p��ǟ��\w@r�'<�I/ 0�;v�[��Xi�0�I�i8�PKC힠sHt��sK�~؞�j7)��G�ŢP��(��8��Ѩn�6���58ꘁ	��	![*\5 ���*�!��H�͟l�	v�'��B�k�~z-�3-��`����&7D�ܚ���c>\sN#t���q�3��ܦ��Ity���%C����?��%G9Oʔu�GcڰJ��H��C�?q��7�|9#���?��O�J�3��;u���ae	Ne>�@BGKA/�")�&���f�!�#��u��pS�i�'�"A��a�.' �9B֥��\��� �D�]���q���+��@ե� d��{6nTE�'�@Ux��*)��<���L�Zd��a��L*�^@�@o�T��ڲ�N(6���y?��h��3�O�P�	9K���G��z��m	ba�@+�d�<�#�ٛ��'��T>}j��矄�7cͪS��m�G+� kQ�t���ޟ,�ɂSۚ���#ΜYm5��eI&a����˝_>~p�O�6�ѵF^�U�"�ݎ�qd����b٠*	�h2�l\�o�B��Ŭ=:��r�~r�f��N� � $��g�>���
l~2(���?��i�X"}�O;�#���T���Y(N���g/3D�Pk�摾&4$�L��q+�9S&N4�8�>uIRE�.�&$K���4��͠P@צ��Iܟ��I:Y���TKܟ,�I����	μ���"� YdaA,@�69���B̓c��IO@(��Պ�N8L��!ϸ	��b��f�#LO8�×�3[�쑈$ɁT��cv�!�$�
T���č#"�hy��2:��� �D�P?!��p�g'�!Yh���I�'4�I"�HO�	+�f�ۀH��`0�\�g�F�)����#�|���O4�d�O����?a����C	�8) 	_�I� xHB�� 6�T-밭�5���'��J�) �8�N
8h!`^�5|hd$��@�Ib�.�$t�j��M����׾q�R�h�f��\��CO>Q�f��4�M��R�C�(Q�K޳��5�	x<��"J�4����Ѐ܇ ��!{2��i����<��0wT=���4*D��Nc�ɾ�M+N>Q�ٕ|��S��SP@Q?s�t*��ν~���Ƌ�d�I&B'���韰�'$�[�$�M���Ս��6�% bE�>s ���T�]��x�AN���@/�	�u3u��p�����'G<�t��Ȟ�{�l) �T�v�N���#��9���R�J�I.8�P���O(�1�"N�|oJ�c5����$�Ї��
pJ]�a� i�!��,�47nJ��F{�Oڨ��U�,��\��'�*f�)�w�Y�[;�X�p�sC\�M���?+��5˥��O:yY���p�(A�7"T7���8���O�����GO���SI�30��I����OF�s�	�T8#>���bȈI���唟\+f�&����2͍�Y :��,�'kT�I�P�����2F�@�'xaQ��?a ��t�)�\��ɖ��'x8����	v�'.2�'��8Ѓkڨ�|���S�M��-��}}r�yӠ�nZC��&�tu�b �<U*����6l6�1Y�4�?Y���?�ᆚ3&�6݊��?���?A�we&�+6m�=v&p�/@�7�J���j���IP�?j��J�3 �8����y���P��m;��T$�h���'�@|(V��+w{�iqΕ-O"�5��,�j��S�k�����i��C%�ޖ
��d���?�Z�k��O �|���	ϟ���P�z�T�N@,5u|�hfaG�%��5�	�',���5C�168 �)�)E�i�H�{Ѳi�2�8��|"�����-R�����A[���a��E�1�*��C �O>��O����<�O.B�80���j�-i�^9�e�~���i���m�:\�D.ث~2�8�ǓS�^�&�@�X`/	�+d��;��V�NxpS)������`4OT�:�c�qN�8��H3$��Ұ̈́�@���'�ў�Gx K6r(+�`I>K�yb'*؊�yb�RY�j�q��ج}FM��a�������by��_�Xԓ��qS���O��Ur�΀2,��y�'������I䟐�Wb�+L�\E��¤T���B�-<d�`r�ݟ|~����{l�m��	|�,X�p��,$�ej0M�(Vp�U�F$x`3u�^�o��j%�9O,̓@�'�"��t�C���Qq�g����8��=�O��1�����{�Fׅl� ���'�:���!��3��BN����H�(q!�P��˓)ayʟ�ʧ�?��u��1��O������$�?Y�i8"��R�LN�y���q�������S�V��Ԙ�)Ժ�x�u�0N��I<BOι��	�,p�6����Z�,�Q>��%I�/$}8�Иƈ�'g>?�@f��D�Ip�O��� \e����5�X+@g�R���"Oܭ"�g�n���A�M&x讄���	 �h��ab��~aеò��/G�$�A�yӾ�! �<	������4m�B���-մ
��J�@����H� ���:�Ph��9�w#3�3扫y$�@([9��sC��4�!� �:�V1"�F�/������4�3扰V/�PG��=nL�<�g�܋v�<Do����>c�b�O��3�d�8U��
4���8dl�hŸC�ɓ0��y(��׺gtlrvI�kb� ������om�p�t��A�T�S�\�V*@ q�Ǧ�c� \O�0q��"\|��c�N�Wh�Y��6��( 3[�ssS���p<�`������x�
��VV��
6(J�#����ȕt���&b�0T�P��L."s�1�
Lnh�:+A�����'#�6��i�'��p� �.e�T�ɕ.w2&�0�0D�t�r�3G��Jf(�U�TqK��-���N}�S�8��W��M�2m�`��]�p�Y��)g?� ��|�'��(*>�fM��t�6����Ch8�2�/O �ቐ��#KG�B�"�[�#�f�����FY<��?����r���I�r������!򤂹[�Q#�	6+�>��WE����F�Oh��C��v�x�z�W�j���|�ϋ3�6�Ͳ/�Q?�۔ �-<�$�&�<!�H�x3m.?a�)A<M0B-��䒅A����`,�'~1��ڃ,ā+�MqV���m�}�'�Zq�R�z�v��A�ȭcxaE��U�W����Ǜ)���aU�]&���N7'vB�hӸ�G��5�(J�<�A�
��'��u�<Y㫕�8�.���M
�Rܼ��Jx�'��}�H�	@��I�'�%�Bs�D<�M���(���;j���g�'���I�.�.���YP�9Jc��y"��"�0=YD��t� ��9~��rG�d̓]��}��	=v���	fe�Ԥ1q���'�,Q�.�O�b>c���3K����A�mY�^<�B�	/D��s �ɐCPA Mͷ�z�!	�<���)�'-�(1��[�#��0��$P�)�p|:�L21���%�N�(�&=���I2V;1k3ʀ)y��L��;V�@�G�/yN�Q�b�Np�H���L������?�4N����B�F(�q qBw�HMC�O�0,X����B!��n��I�M��O���#�ĸ[�Z%�K�'p��c{ݭy���	�64��a�'QԌ�`I�_��t�S��J�ܥ��O0��5��^�HfH�.�"Y�&O��K��ʓ�0?q�'�X:�0X�� K�|��%�Y�	o�����<���V'��ɒ4F�Y�Ա�BETyR�;C��'s�T>M���\�`�IkmUb���	r��3P��#_����I!"V��X$0冸�V�ڝ[��O�1�zHZE�5]v�5`n�8�~R!2O��r�!�6�Z��q,�8Q��C�]+]:��i�Ҙ�'?Ft\T/6	R��K�M��ΓC����Iן���'����R7� ��+��W�Ltz&��-�!�T���p�˔P�Ιs$�ƚN]�O�D�\���$��g�\��WH>[=��PC/�?��'��L��p4s��'�R�'�"/�����?�b���␻R~ڥ�R�]�Հ<���N���'�;��SO�J�T/"�	��_�.��Q����Qj�Hi�猑j$"�����O�Rge-�"����2�S6�<9q�}z���c�p�K��b~bmǌ�?���hO�牔�^���ܲ%�|A����
��C�IĲIT:
HB�*�j��NS��*d$�O�XDz�O�"U����%��rW�l���+d���AJ� �*�#�<��ܟ��� �u��'�"1�"�A�nQ"t6B��/,��QK�8)�)B���	efy�2��.�p<�T��<IHX( 4.��� BTK��M�3q���鱮ތz��&C�,i�0�7�G��j�0E��	�HPӢ�I<g�|�P3�4u�	x�'��4{��X�BTv v!��B���'2<Oz"<��\�l��)Jvƀy��!`CGyR�f����<� `�x7�Sҟ�'f�����܆W:d�	F��~<>��ɮ,��)�	۟��	N�H�!.�d�5xU�<NR���'���H��"_��)�@,��\E|��,%��8:��O! ��(6D�z��,��G�$\9���q	�u�$&�2P�����mN�I�'�������?���d�5	�DAVd��c�L$��)P����9�O.z&�ؘ*@R�sC!�/8�Ԅò�|"�i>��,Ov8�Ԡ�]|rO�Q���
�\����	���\�Ity�W>�	�����/�<���hO7
����Oܟ�J1�
�Ȓ#V���d��	h�O��+B��#l�	#����Az�A��'�0�x1@��U�H�Ga�*1F���G(4$��)�	3m50��P���y2"��?A������t���  ���e�`�ѵ슯^�8�C"O�$�ʏ=�dd�f&������	%�ȟFD�b� �^����F��+|�{��O>ʓ>�b̀��?����?a+O�I�53ĥ9��I�-��MR L�7?��r��P�1�<hy��T?�X���?#<	T�#n�b��ł(���k�w4>���dJ,N���Qc�I&C�L���O2���E�-���'ٗ� �RI� �7��O
��,��y�iU�H�(,㚁!\f(A3�V��y�U�?���F���E(�?��i>A��IyRiq�P��F7PR�u�Yh<����)���'Sb�':�)�
D�N\���Z��0l�D8�>H`0N�	{hK����H�Pn/O�P �ʀ�:UX�4e�<���p!�Qqfiaq���i2�����A�p<����� @%N��N��IV�ץM�b���g��(E{��	�r�ZU��7M;�8��c��6�*C�Ɇ,�Љ	��I�be�l ag��h��ʓY����'���'u�6���ޟT���|�QS�R:nyaEf����$���I�	ftI��ϟ��ɘ=�칛c[F&�$)*Vv��'d�$	��)����V��m�Z�G|�h΍4n0a�s"\E������0G��� �[1En�@�׿A�0�ʦF��E�~#=!�+Cş`Jߴ����'��iW>ވ���鍽zX0*��D9���'��O?y�Ч&L����(j��p����	�M���i�R)������Q���1HqR���	�~�Ƥ��ퟤ�	��`�	Ry���H,:1ʆ��&s���8���	ax¹i)����i?QB[SM�+w����"��:�<O0b>%���4T��!%R�3���1�JZ
�MC��"$�D`�'OVM����?��'�?�'�\X��
�I��s*�4I�(�C�A˛&�'HN����'�b�dظ|����u�������Z1��fZ%�M!�a�8k(�f+�?��c^Ⱥ�'��n�OH������Dx���J�<x|�
�N�hv��E��*)�V�d�O��?!�'���	��M��R��,��'����Q��B6 �Z�c'�'}�5+���?0H�=w���ޟ��I�?����<��d��G�:\Z0��dH�6����Zt�P�I��k��L�`ϓ^S������u���5&H��jE�ޮJ: 1����M��'�<ً���?`_���'&��O՘�ч�^MPpHs䄊)G�D�b��
��4�"�'����D�&��禥�Ǉ0��J3�Q���5m�-���0�M��'�[��i���_���S�?���>~7�Y1W)
p$��D�#'��\��4*�6)��'��l`��?y���?A�'A���O��,��Gu��|��ɐ�|K��k�i!t�Ё�'?�	���4u���Y��I�X���ғ���>�NA2�M�pO�D�ȓ�:<ò�6aԔ�JaM2z�
�n����vy��M���d�YgF�h$���,9[��Tg��6M�O���<���?���͸O�:�@��_�	L�k�l]�J�$ s�}|�V�p�OZu9�䋭:qF�p*�0gw�|�%�i�ў"~n��}���+6��*b�e;��ٵi��C䉤*h3	)�56�$v�RC䉔� Ac�.]}�	�t-M��BC�	�y�LԺ�dA�Ahl�J�#�)C�zC��>�qC h�5�ZEcfoƂeuvC�ɺ9d�P6��HK��fN4	/pC䉻	�~YÂ'�#x �l��&W�jC��hY|5��^�[{���`A��MpbC䉕!�TeÀN�P	�Ѐ�[�"?9��?����?��`��:�/�#,�zsi�Wf��ӽitR�'n��'uR�'���'���'z��� Q��M���8bt�w�t���O����O���OP�D�O����Od%����kC6=R�X*����$���1��ٟT��ß��I��\����������'�]�z|H� ���Q��4�M����?���?���?9���?���?��K�g1�1eP�m��a�0*����'pR�'|��'�B�'��'�" �5�|TSw'/_r�E�3�:C7��O��d�O*�D�OZ���7�O�$�O6�Xr�Q��hӲT�l��C7�@�M��ܟ���������4�	�D�������1~PڐqR��.��pAU���M���?a��?y��?���?���?��/ �suި23CJ(J�+�HB�����'O2�'2�'���'U��'�R�N�Ai�	�t��<6�\�X� �+h0"7��O�D�Ol�d�O���O`�d�O���9r�:PHW��Q�Vp��h�4J<�mΟ<���x�I។�	ԟ��I�� ��
X�tM`N��
S@,1ܥS�4�?����?!��?���?���?��:��\���� o���æ�2kn� 
�i��I۟��'?����=c
8�+Cbʞ/T�,�C&���9��!�Z�'x���6O��z��U3r>��I��iI�)U�n�8�n��<�O������c��0eT�$�6���h3"G2����S�E� @R�_ 1[f3T��>�ў�S�<��(�a�F��EӜ9^�D����l�'r�')�7���1O4� ���ѪH�Z�����fW)�Z�if�$�{}҆h��|o��<a/�.�ig�������E�όh�a��My��G�e"�Fƥ��4��8�ăc{l扟���#�[�
V�jbk˯mx"ʓ��D�O �}�.���j"�I7P��PS)���I'�Mk��EP~��c�8��'vn>��dϙ�x�.P��ײj1���I*�M��i2� mڹA�Op�z$kV��t��Yw2n�Y��A�Jt�Bo�;����$�O���Oq@i����8_^���s��rQ�)O�mڒC��b�����e��8�E���V/�(���I�����M��i��$#�'-Qh�K��ް2����D�8�S��}�J��'=����n��ѣA�I� t���L2m�m�rc���J���\y�]��'���4m	>���}PcDͤZ��Z6�GA������M����y�GyӒn��<���	0r,R��2�H ��̅-X��+a�y� )���2n;��#��1G���u��$3=����gP�q@� 3ΐ<Z@�V>u)�'�Iqy��iޮ$���C��%�`�
�"M>Ѵ�i��<��O:m�f̓2!a�%B�WZv�҃��iֈϓ����ަA��4�?IF�# ��0�KƬ�V&�!p)��l޻)�\I�r"^�zN)�7���D��J��B�O�ɪ<�'�=�A��.el=r��_�ʽ8���0�v-P��'�d>�� �7	W�M�|����:!���^��y�O�	oڊ�M3�'M�O���4{.�	�B���;���c#�@�.�`� ���<ٶ\�O��I�7|�u1�8�4.�T��EK�r?�]"��Bh˓�?.Oj���ɡ�MӤ%�xQ.qT�p���	�sDL�w�'?ѕ�iI�O�9O��o�"3�tHBe�T���b�BP�Ծ�8�4�?��oL H�\���?���%�L�R��`~����V6v� ��f�@!��A^�JRS���#�(���.]8��$�L)��n	A(����矨��O��`��3O$�1b�a&&pkFiP�B�48�p�`�Ƽl	�?�On�)�z���_�lpr>OF�PiF5E�
�CƯ�C0���O*T���F��Q�4FF�f���N�){��2Dh��t��Tm�f%�'���:F ��`b��"�]뀬�8/�,�r0K�=	@��3���
B(����0��
3�K�m=#�����:/�p`<Oj�Ő�(�����E�=��eP���4Թ*��7&"lp@NTs�y ��Ei�@�(�4E���[�#w�,�@�z�8EA�@��S�f�b��C)� q9tʜq�JbbR�X��i����Du�A@�f�@hZ�J����@"�Irf&���!��?A��?ͧ���O��zކ�#���fA4w����'��6��y�%|�Qק�O��h��O�( ��qc[�uDlbo޲sl2��A�H�+���EC* ݎ�����"�d/��u���A/
ɶ�{���Hl\�Z&
 ��p@%�&a_�)��"R&{�v؂�ꁙK�x���fY�'����e�jS��I�M\� TaKF�P0�f*�6+��{�W!ބ�]v`�����Avҍ"C׮sz������p%i�kQ#�� 6�}08豍U��.��RCv��q0���� � �)iT?�ht���U`��cO�0��)�B��t�<9���� ��r��&�Mk���?���3�x��'��=,1��1�B��o�c���?A�M��<A/O:��-�ӟh��턻$�e���>L��V��Ɵ��	����� �$����`�Oj�1O`E2��ϛ3]xx�-����������'Q��P����'g��'�>e���E|�82��� 2�2T�'u��3%q�It���'a�'q"��'@���#�Ӈ]���R��Q��B�1����?����?���?��#J�t�kT���be#�Ř%�h*��?����?Y�����?Q��	�@`+��L$ĠL��U8-�V�S �X;]�2Y�'2�'���'{b@��p�i�0P�=#�W-�r� d�� +�B�'�b�'V�'�r�'��(CC� �rT2u�ċՌ3ЎuR�, �#���;�\�������	���	�
xN(�O��d�s�d�x�$]����I J��.f��'\�'g��'hZ����'��9�"��#��4��3"��&�8�d�OP���O>���K�&ʧ�?����
������bŅ�;[\P�$$����?���f:��w��S�SZ���fh"���/|(�m0�����l�'�4k��h�`�'�?i��F�	���q���2> I�A��^���OL���r���>���J4J�̛�&A�L���
r�O1xwD�O"�$�O:�D㟒��?���M�p���h
�0m�Xg�ļz�����=�4 ���I�O�PT*� 4�Ԋكx*��'�Ox���O��$�)8p���?i��?Q�'��I���JP�$��¼S����(�#IV�'���' 2���e`��E�~Z"��uIӔv9r�'���W��������IV�.w���ᖳ�����U�W���'u��q�|��'K��'���:b2��K0G�vgv}��C�$�hT�pM�ty��'�B�'��'�R�'a��( �PsjN|B!�Z��@�WhR^�<��џ\�	yy�&��
g�dBz�K��v��q��VN�r�'�'o�'�'t<|CF;O���C8L*co�9xy��Z�������	hy�A�4����j��V�s��@�fμgxp�� �IH�I��	5�:��<Y��:Bl6��A>b�!y��G쟰��ӟ�'�nU	�^>��Iӟ杲p����'(<uR �A�^�G��%�$�	̟�᦮�۟�%��3� ,HY�@Y�!�>H���[ה����'�I)�t�I�<�I���iy� ę@:t�6.��^������c���'��
D�*h�Oq������A٪lEHܟH�(�Q�'���[1�'�R�'@��O��	�����7R<d2�'�9g �"f�/,'���]���ID�)§�?)aV�"bi��eE<�8��j�>�?����?���s��;(O4�$�OX��d�|{�$0<�҇�K�Δ��C!��*#�~ $�X����P�I�]�	B�7�5ٴlAHWd��	џ�;��Q)���|J���?�+O�8����C ���� ��8���O�˓�?�+O���|�+Ob������$�Ju.��d�:���!�7^�J�&�d�	⟜��Dy��'��	[��5*�*�1����R�	N�'��Iן�Ily��'�f4��4�F��V�ׇ��l�䌌	[0!1c�'��c���?q,O�q��� �F�!�l�!�]C>��O��D�<��C�LES,�8�$��	qX�A؇�4$ڢNR;0�(��-�Iş��'�쐪H�h��@�%�P9�ߞi�м�Ǧ�O���<I���0(����OJ��.�䕳�4ck��&mL	��O��D�<i�!�d�'�&E���M-��� ĩ�(���SS�t�	_`���I������p��jy��Ư^ܽ�6G����xB�ُ3���'r�I��
[b Ìy����V:O��qA֠ݾ$�trD͖��?bA��?���?����/O�ӧ>��H!��rj]��5v�����VrQ�H)�)�2�QN��C'��(�!75�`(���?����?���ڡ��?��'����"�]5i�v�!LC��z�D�f̓	8���I~���?I�-���P�߭(Y��#'K:9��h����?ik�:�������9��\y����
�Pu@��\81t� ;�=i���'��P���'b������Ɵ��'�0\[��9R��(�KԺ!xk�3*OJ��O�d�<!���?1�jD��R}To��T�vUr�$~I`%�J�&����ҟ��'SDU�R���LX��J�.��]���p�@�R���	ʟ�	Hy��').V�B�w�fH��JYW:޸�U��q�����Iןh�'�D�%�-�韖9ѐ���L]�p�=#�k�7�
�$�O��d�<!��?	�@��?�ΟP�+�c�0�@d��Pf�s�'&"�'��* HCL|���y��#~XlPXdc�.K�J��0���?�/O.���O��rE�O@�'�?q�w/ʉ�$���8�(Юc������D�2���mZK���'9�a�<�g�ڑ�� kFg�O�,��A�����I��w!�����O�b�O���@!!�4fǥVO �4<YfT�	��l��埨�'H�T\����5�7(�"\��J�~Ȅ܋�!�dY;bD�S�O����c�*�,�:�z��Be
-��7M�O��d�O�bv�u�i>%�	џl	��-c�U��D�$+��)sDN^şl�	��H�ɼX���O����͓N-|9r$�ӇO���⅁5�f5�I����`yr]>	�?yTiB7$��\���X�G�!�G-��D�d>���p����������Fy�+��E<�(e���wg��8�B�$ѫ�>y+OR�ĵ<q���?A��iL�1j��ǖfɠDb+9*��"ee�<Y��?Q��?�����P,A��T�2V'֑	t��#]$�a�$N�EO`�d�<����D�O��D�OxU��1O�!�ԨA�L�����J
VX�$�`c�O�d�O>���O4�Gl�R?I��s�2a�B/��YȪa���O2@(�IΟT�'J��'8IU �y���|`���n��DCêYn�����O�D�O6ʓM��PquY?M��͟<��NLȘ�b�WQDL0t&
w�V��'`�')�.C+������'w5Fxg�b+�l#������wyb(�>6��O��$�O��G}�-6j~=��mL'F�6Ms����'�r"L�����<���4B�
h��5	��˱"���ҁD��?���Q��&�'2R�'�����>�)O�-;�`Z��r�ct$��g�U��O�4�u>O��d�<�����'�t[�jZ9�\r��*vt��A�!g��D�O���JE����O8���O�D�O�QE$ˡ d�1s��l	L�˂H�O��d�<�c�Z)���?���?�bgLX>Ց��%�T��L�?��S��m�v�iv"�'�r�'����yB��E��d��]��;t���?��pWd�͓��d�O����O��O��p�׭Xc� p�тc,�
[.D̊�nП��I���I����<���4��a�
̜���	>�t��B�<���?)���?���?��Di|A��i7j�ŏUq���c6~�|1�'���'[��'0U�h�I?f��ҁ����T�2���X��'b�'E��'�BL�,|��6M�OJ�DջG��AB#�țW�.\���Z9T�d�O����O���?aQ��|����y�@[ ��<�!Ν����B��?���?����?6�u���'��'V�$];W����h�=Ar�{�*vb�'v���`�rea>��IGy�OW@�SrK� W�>����R��9���'���',2��{����O��d�@�I�O�8c�
I�c�BH��ݙ� ���H�<�JI������?Q*O�)":��V��ni��3��ث�#֟�P�E�$�M��?���Z�'�?A���?i֊�-g-��hve�
1��mY�˙$�?�A
�?)���4�������<� ~m��� ���+�A�<���ae�w�h���O��D�?J�����O�$�O���Oh�	2��yZ�����F�Uh4����OJ�$�OF��@�������O���+6L�AH?|��� ���.&&���O����Ϧ��Iٟ��I�t���4�ɀE��Uے�I���d8�Ήy�$�O�0Z�;O���?���?9���?Yak�6�H�@C�ƨ@�vҲ�4-
Y���iir�'S��'��'����OF}zѡ� J����P�{��l�����ro���O�d�OJ��O��'S�,�#�i�D�Q�O���Jd�!��Mz�'�2�'��'��W��	�q\N��Sbt�a	H�-?H1�cm�
i�,������ٟ����x�I`�R��۴�?q�k�P��ק��3^2�b� d� 4 ��?����?�)O2��O�W~�I&?T�L%R���l�|�upr�K֟���x�'�AZ�()�i�Ox��N?�.�BWI�#~��r��� ^�D�O����O 1���O�O��\
W���3���4l�tB��ՈV �_�4�����M[+�^�$�$��'�`�en��2I;�2?<	����?A�a�Rl)���S�'pP���gB��X	AN��)O���	��<�a�4�?9���?���N�'��cL�Tͦ@��)g:�I�)�8e�� ���y��|����O���_�YS�y�b�hJ�������	����I8Y�|"N<�����<�SOC�4�ļ��l�M��d  #Pߟ�&����_�Sǟ��	՟��p&ʥ(�(���T?9��]�B��ޟP��,�T�K<����?�H>��i�u.�bH�����R(���<Je�$�<y���?A����	�W��(a��l�D (��I]ς!S�/@��?,OF���OB�κ7+"��F��t4$���"�dQU0O�˓�?����?�.O�p	%J��?
3G�1,����ǁ-��)�l�<���?1N>	��?I!!�8�?a��[!)��P�6/ɼfj8$1��Q���d�O����O��9�X�+�����`�ض��7����d 3*�b�'��'�r�',~e
�'��P�̬��S�
2D�3�]�=(�$�O��d�<���H2G��O��Ov��`��!2�� �Jԑz�>��@�|��'��f]
�y�|�Oqp톻Hi�lݒ�K�G�*�?y(O��c�ަ}�O�2�O���:���eb�<6Ub�@�*�H���	����I�:T��?�}*�n��H�����U�Tm��"��� S�)���M���?��rB�xr�'�J�pү�7R�	��Jw�����'Y���R����ܒe6tjhB��ɇ�^��ׂ�M���?��?<��'�x��'[2>O�U���ϙi�=४U�=�����'O�'F�!����'	2�'L�0C��^=@a��j�/cd����'�R��@��O����O2�O���7gRVP�T��dF���)R*�<ِ�����?����?A*Oa V��ڀ$)���-mN$$��m��8�q%�T���'�P���Hy�A�ZJ���4�Տ�p	rț#o�4�	KyR�'���'-剅rb����'��̩��ųW�(e�Ȋ�%Id0�'���'��'���'S����'u���d!]$-��g��"�
 �'Y�4���l��dy��K5v~��.� 7�R�DD*`I��r9b��O��=��;׮������Ӝ]6�RԂ�?Kx�qe)�g�b�'k�W��KV�F-��'�?��w*(�8P�
)"7� c-�DSp����'P�!���'��z[$��f���3Y�I ���U�����xIt/Y៸�	ԟT���?]���|��ǁ�K���vV4H,���!R����ϟ0��iC���b��>q�"i�'-�B�H�đ�`C�@4��O؀��-ʦ��ן��	�?�XI<!�����b�
��)���+U^��SHFHFx����O���-V| ��S�
	nv� !��ݦ�IğH�ɡX�^��K<���?�'Q�AG!a� /B�L������+E"՘'"�'����"�fԳA�:	z�
[�3b"�'�6���'��O�$<���	&�=�օ�hw��a�n��d�ʓ&��<���?I��?���@�`�`P�
�BV�90_q����$�
��$�O��D�O�O��d�O��z�A�j�@�������t*c�+=Z1Ot���O��$�O����`=��SS��m0�
6"-���=7���d�<����䓨?��r�\�r�/��u��5I���l���	�#~��:*O��D�O<�Ĩ<i�dמ��O�� �.�-n�t�K�fѨU��q��'�R�'i�OVY!��	R	��
o��h:�ҧ菟lq��'���'��F��'>��'P��!�.oh�
�o�:]ش�r�X��'b�'( �i��������7�����_0�I
b���?q+OD���)P�Y�O���Oyl�,#Va�-ٳ)>���;k�"���џ8�	:I�#<�}"���P3�)�6z�n����� ɤ���M���?!��rg�xb�'��;�@ɧ)T���aDț�l����'�Ĵ(����4Ye�H�.���� �I
&�FI��/K�Mc��?A�G�0Pi��x�O��8O�t��-ҪY?�`� "�p��AC�'��S�\��K^�,O*\���C!ILDK�쀿u.�a �!���t	M�<#w�[
47�噢��+@�P8��B��H��ПT�	�<1#�[6y��̲4���'^���uA�W��џd�	��	ly�	�J]b� *�{��ݵu���hᬆ�(�p�'���'���|"X?Q�S��?�'&�@Bhd�cI��ey����� �?����?N>A����I�����vr���Rís�H�!j�=��0#&[,d������.����!�O��8Gl�!�Vy�'[�D�J����'Y��$��7�.�h������m �מY�0̋��O�u�P�q��(� yD�űb��;֊�
;p�`��ҔM���J�D�Yр]Q����i+�8&�����L9xFȥIVĜM��+��!p�@(�V�i#Q(�)˲-W`\SdኮW&
-��_�HT��&� F��2���##�P!�&U��?��Z��?���?���ȽDpu���ǟB�P��uW���������Q���/����O��� �E{���K?���-��H�:D�xXR�L[=�"?Q!�D���I^�8�R�F����X��T�bҕ>I	�MU��P%��$�J����ND�^d��		�~�L�'_�x`�2y�� ��l��ɔʓDLE���iP��'~��I�y��צ�QD
%.t�Wl����Y�ņ�?�"���B�Hs��._�$0P��#���$���`&p_�04F�6����N C�㎩}����
T��#}:6�	����Ф�n�������\}b��?a��i�6M�O#}b�'G�L�sJI&m$�]+N�W���O0��DخH��DZ����D��.r9Q�q���R�tߞLR�fʣCĄ��hۆ.�������O����O�Y�B�Ҽ�D�O�d�O�ʚw
2HP����D1�QJֆ ��tk#��S�6�;@I-Ѷ�y�jî��g� ::5���B�=hU�DLC��I��_�I2��)��U�NT��$�N�˧h`��B2TU�ôai��b��(^+|��3�0W�0��'�P����?����w�d���2.�b�@��;;�D��'t�ȋ��7d��k�k�\�!G��O��Dz�OI�P���3��V���cY��S ���s��,8�Yڟ0�I�����u��'R>�nUr`&�
69��/�&FP��봌�M��!���	�N�c��7<O*��A�?�(m�SMŏ0�8(��cۼ l��bO޾��x	�o�"~Cax+ϗ�M�tL�>B�Zm��e�������K���	{�'�.ĉ4�ؐX�fs��9q�R�
�'��k�H�	l,H���fH���L��kݴ�?A/O �&립�I��lZ9b�^"�J��D�(��l��d��� �,(��?9�b������I�u�ɧuW��`�,,s��$nPY�.����Oؠ�G旻W0��>}��g�3vg��U���Dq|�q�K0�>��i�������˟��;���!D�B� 8D ݶ��H��?����)�/h��C����B�# � 9��~򮱟��$.E�N�>]�"��CȸI�#���d4 :Xlҟ�	k����1X2�i�,��2�ҽZ'��A%ַ֌����O��6�DSq��:�iT)>�0��|�M|Ҕ)�%0m����ߗ���:��d}�jQ�9�b���ҳR��ͻ����&HKCA�V�q�o^z�"\�qU�B���On��$?%?Q�'�NEp� XY���C ��4���A
�'���8 �( \�!��e�)����@r�O�p�Q>�hغgNZi�T�C��O����O����M�=��d�O����O�Pћw��IY�e��i��]"�`U`��׌4J%�	o�7ܷ9L���')jUq�<-վ(1�Q"��@���( ���4�&�+C�8����'��ЂlϞby�:�S�/��D!?�U�Oş��)����?����M��bѨ*���xw��	kr`X8Ď�U�<i �P�W��|�Ƒ,f��Ux�dv?) �)�/O�tR��A��|���Wc`4sA�jKԐ����O��$�O��� ����?ɛO?v�x���*UPP�
��E��`��J�b(�2��7Ħ�BJ_�,`*"?��ş.����ԣ�7vdl0A��4x��e��Ht�pk������ي�F�i�E�ס�n̓j|��l�`,~9�2.]�@!�$��LN���9����hO�"=!��
�9��xB���,lz�bv$^J���>�g��,?��@� 0�f�	��E����u��py�C,C�'�?�4`ۜ��@��r�ϒ/��xb��?Y f��?����?�֡D2>Q���K���%�s� ��(!k��W���H���BV�P�e-+�ph�c�ʁ�lP��#A�^�[5��)�$1�D�k��&g4��`�G�yQ���1&��O�5mZ����(m�&�:AJ�,UR�,P�)N3�v�'���'!�1��BDp��t#�@*���	�[�:EA0 ��U�~D�<��-D��̖'j|=�q�>����iY�Y,h��|�*���-��z�����l�ҁ{#��򟠁��ٰlS����U% ��+F &��I)�I�|W\T�!HO�"���pKXt��	�p��q��۟K�p$�gFN�.B�����O@���JT�U���A4Q+�ЬO�Y�"�'��7�\�(����e� �pg@ W��\�� G�c{����"O\��
�M�b2��،�����h�,�B6�	�o��@EP�c�h���d���'��P�K1>=)��'�B�'`R!e݉o:� Dİ��ߊkߘxi�b�FU:�RW��(6	��iA�� ��d����O���OT�Flz�JU�R]��AZ��TIf�i�H��h�1����Or5�vc�3a�}:��;���U-��<�I�+�)�Iϟ���d�O�6��5�^Kc�ӉI��(P�L=a!��ϕY?N�I�U�h��dV"FE���m�'r�x���D��H5�]���N.`�­�B̝���bp ݑq����O��d�O�Y���?�����Ds�Ļ�d�	1�\��q�n	�B�e/#N���h	&.#���D�nZ��3M� ld5�c�ة&R��C���9%����
�b=kb�> }�,�!�ɗD>�7-]J�>��Mζ[��r)y��u�ܴBt�'���'��O����>@5L����
�`C'���yB�W$5�|!Ţ�)q� �&��)��I:�M�������em�ן��I�����1����M���\�K5"��?q'+��?���?��H�A����"K�)%��:E$^�R���:`�Ôm:�{��2�.�#�9���Dy��@�[3�a���(ru��
����(y���"�KS�^�f�ap.�$
f(�剳O�h��O�����,Q� �e�P���=Mt���H���~�S�O�Bl�Ȗ�f~dh0g�;'Ƭ(q��T���L/B�4�˒
�#6�X1h5#4va�8�'�P)#v�uӦ���OH˧ސ���M� D�_���6G��1�";�ߌ"b��[Ą /v���e��<�O��OM��P"��i��Ej�L�Xj^u(�O����(�U��+������?�������D1�;1�.�3��>	%J����ݴQ���'�>ͺf�Ĺ��ə)����H�e���?�ۓ\�����ەD��x*Rm�@�=F}�d6ғNLNq+���"a0��$o�R�͊㬰�(����P�W��!��ן��	ş�y^wD�VO�&����"{y�g_� ��E�Q�埜����X(]K|�>��B�	:���f��7_���q�cA�T��)�O����� \�'>c���PHK�*�TX�d��<��z��;��$�3Dxr�'���wj�B7꒹1�X��*��%��i�<Q����OC*�DU�]*$��_i?�������<����q��d�p ;S�Jd��aʸ{,R�;�.5�?����?9��u���Oz�$d>�A�i@�J(Q'M�:¡�A>�d!� �W����&�2��<9�	nӚ���-�"`&�q�Bm��?�&���ђ��	+uDT���48�"���n�4M��u[�#K�_���b�Տo��I�����?����]?�1�H]��"������M��;b�7D�TQŤ�#j�-z�iũ���v,)}l�x��<�7��>a����oڣch ��8�Z �gϽ2�&<��������?)��0�Ⱥ�F�	�,�AB����+sAK�+b�]��IL�L��"�56�Q�\���3��^7�`̰�GEy'�ĩ5b��8�R5�k͙a P�3lP?J�F{bH�9�?)T�i��Of� b!XI���Q��ɝB�b�H����P؞D+��a��rdl-��T@��<�O.����6}+�1qI�� éޞ.N� X�|a4.
��M{��?�,�0�� e�O�7��-5�0	�f�v��D�s��P�Y���F	���K�)�0Td)��I�OЉO�Єq�1kZ0�F�X*)Uh�#�O*���޼S����Aw*Yrϕ5�������`�0P���(�H��o0�+Ă6��	F�'n��'�>�q'�B�	40y��D�s����.}��'�a{���+2�	7�e�R��/B��O��EzҲ�*� -I	�f`Y���Y�d�1��ϟ���ڟ�D�ˡ%�0���ş���˟L�Yw4�&�K����4ˉ3>�L��ئO+>�G���M�3��z���5���}��J�}A�u�����FjRqR������5'�['�Z� ��-$��I���;��t�@�T�4ycp��[̶����'��7b�{�����O���O���|�����&�P��L
"$�|��"O���B	e|���țZ}�X��O�DzRB�>�/Oa�2-đ��m��$)��5��Mʰ!�D����O����O��ĄQ��'���AAF$�d��-{q���.��z�����)�6[�<���	/���"�� 0��-���9�F�v�;�����)�I����'�j<�ڴ��<a��M+E�b�S�A,���xp�'���'�����?��6+ L��e�8F�]���>n3.B��)*����zj�Bf�+ �'
*들�D�$JPn�֟�Iڦ�"$GBuK��	B�:Xq����-�?�����?���?!���h!�
�j�b���uwFS�J���M,4��Qy�$�1��OL��%M}�!�T���B��h~����k �3�:_�"?y�O�|��K�1��LQ�l����d��M��5ER���?i������^��(�3#.4�B�����~R����3��"/F��`�]Aɀl Q��+��D�
!o�˟<��^�d�)ҷi��(c��#�&X���9*P�@n�OH�x/L�e>tY �i~ �@�@OT���� 4��h��?����1 J�C��}Q%W���&��>V��GK�"���S����f��<�Q��\�t��!��V3u}�}��U������O���Ϧ��IX�$�i�"_�Mz1K�:1i��	��;N���'n��'��0h�N�<#�`��&��l���QΦ���4��O��!�6�A+t�ic�D�s�����'��'�ay⭇o�R���JF4d2�G��y��_�́�����IC��;@��6�/ݻ/�����'NH�AM��eQ%DN
�y�'e���2
H�j��x�Q$x,�H�'�<HT��I�H���d[.v�`��'!�U��լ옡����;kZ, �'�f���!�.�������?2)4л	�'R6h�`i
�i"@�k�j�-j�m�	�'!�P��K��w*�ٓ�.��x	�'��$�S픡+��8e��=HB�dJ�'��\IB$�8�F�8%���E����'�~��$qq�Qٔ��#3��� �'�y�%�W�6�e�� �\��'G�����_"��2�杓S�,P�'9�A�w@�)D�*a�)J�H���'�Â�" �h�Ed�@�
�'g��ч��X~��P�'^��6��	�'5(�'"��c�"8E!�7H!��'\J�9���5�X��%F F�l1�'�n!�� O�pyk��Q�С�'!������K����u�Hi8�'�r�ab-é>A�D ��7>d��j�'e��Sq�Y%#j\���˅N�ֱ��'J����Ǝ� ����bD9x>a)�'�	�킜=�R�Q���$,���'P�}i��^+l4�+�9K\P� �'j��z��%�q�gс�x�	�'-\��,4�� 05��:`��'+���Ah� c�E�мO ��'�t�7
E7{*��䈀�}6({�'�4�&�ԨQ9��ঈr�P�K	�'М-#��ǽud8� !H9q��k�'ጝ ��B~U�]�5@(w�� /O���[�3�@0t"���4���P�nI�}�|p0*��8�~�"��!w�:)X"i;D��C�����,�x��1� o��hO��𩈕6�D�'�!6殠�$��D�!�$�
\��@�W9�p|H@�-<g��)�'��=�1BΈD�(9#CD%1���r�'�شqB5���ƌ�b��s-O���d�#�:��t��.����LS��}�X�FƉ$-��t��+l�� r�>D���D� ��i�`��	��H����O���=���>��o��8����녶"h�t��w�<�/Q��~ic�ޫq�J�PE�ЮQ�Ip�W�4�a}��É��\�5���4|��#�e���0=���͘;��9�⃯���0� �5aX<��!�*C(3�0D�l��l�Mk}5�ɩs��	�n1�	)p��5��Pj�Q?a����82�� ;���\���"0D��B�E��V�8h� cơ)��m���D(R*P�>�+J����©~�z��%�V&  ��0`Θ�=~!�d�=�ԕ;� �Z&a����I+�8&v��A���C��ٌO�1���܇�	� ⡠�
�s�D�|���r6�E�6�t� �� 8�!�$��(�.�3N�idD�B��\	�1O@�z�*�
�<������;uh���� ޘF���:db\�I�!�Ĉ�E�t��҉53�h��V��?=��@4-k�	�9Q>�(���+�
B��b�45��ZL�s��8T���zB&[�6��1��S�? �%�W�ݥ\�Ь"B�Ӏ3JB*$"Or�B�ʹ4'T�B�B�^=��3�"O�<3�O�}�  �֋A^`A�"O6�'��"�8M;%	C�тa��"O�=@�!�G�^�!%�31�VKe"OХ�"F��y&h���.:����"O�ܩ�)�q����o
0I���;�"O�Yr� _8c��
6��ƅ0�"O�x�!���FW`xҥ���: 	�"O�=H�MN�o�p-�𭇐N�>���"O�]����{<�s��T�Z�f�YV"O��qboK|��0`�3���"O�؋OT�2� ��Y��"O��c�LĊz�{Tx#�jJ46AR���/�TQ+aݠ750|���\�~����ȓ`	�0��HsbLY��Ҭb�4\�ȓB��	��/D:ԑc���O��9��A��]B�\RҸ��-1��E��L�D{���#Z��ٛT�E�&��,Ez%�&}����}�"�s�|U#�2��=k�bƺ{)�0��NL�<n��#A:4F��5��e�AEĊA��BC�`�R
_�QN����*��� 6+dc��X�,L��U"OF�+cB����aU�$#�@�Ǐ�91 \�qp�N0B\�B⎄��iU��(O\�9c��R�=@��4D/�m�S�'��9:�-Z�n���Q���,i�X� /J4ʧ@IZ)���M�"�����i5��rw�-Jk�M�dmZ'5$=�v��.vv�ɵh��(�$�[#����kr.mۆ���yGkԈb�$�3Cʎn�\�&Ň��Px"*D0~�[c"�]縈8��O�\L\�ڇNH�2-�m�eˊ��l�5D�-�K#�Y_㼌�O��&��[Q�h�q�+
��P���0<���P8VI�@%Pq�B���lʚ�b��1e�D��fk �.�4ժf,X�D!P43��:i�8�R���|rDB%ʓ@�U�i2���F��U#��$h3?97A�*~�R0ȅ	Q�H`UY*��*���&D�b��E�NϢ���Ül	��n�+v�l��Tl��2���;����A��_p��[/��l6���ݿ)�����T�\0���>=����R��Y|��s%/�2h8��ϻ<���	ƮN�A�I�"e̠���u{�aYr�(\qPʣa�|���ȃ͜>隬¥g%>�8��h��8��-��.	+Yv`�c!
�~���:�M��C��	��ݒuǞ��	3�A�n�'?���`�^/_{������35
���'b��g}��T���@3l������!{�.���7y,����|����#�8�2!)�N�=�!��.D:�ӯ��9�,P!���� �<˧D�`�zK�l�lf',Cw9+6���$TҔ��	�c|��
D�'<<�z��Z22�5��A�(JZ��8�,ܦ13#OP�Jd��4EۏC;2�J��20����fӤ`�8���Y1b&� g��
f����	cx����ɢD�l�9�c������AO�H�Z$�� ��f0r�1�M�𬳄�ĠYcW ���:�z��'�>D
P�� t����M�4�M���_)��냀�(vN�m{�(��nR�������5ό�X݆��d���E��y�Y�Ȗ�oFF2F��3ғ5��0��G$8�-�
F�%8@�ɏ�pd�s�1X�t�c�C�Ħ��!BWO�O=j�Z6�՞5a��3f��)�"�I�F�g0^����$M�e�֪�(���7`�y�AR]�b�j �øG��P �V>ѳ�
h̓4*J]��	\:k��c��
8���	4=����7y�&K#M]�	�э����  o�<�����&���Ɍ%Zޤ׬@��b��� wP0�=� �	�3��K��½���%@ݕ	<�tYs@��9��){)U�yA4�ѵÛ�y"�X��S$]&v�<t	5dž�?� �1:M�M2��BSF^�'mZ	]����+�F�:)���[`��`���^�!��مu5b��b��!�v0%eW�[s�QHߴS^`32�����.�Ĉp̓a��
�L	SV{�:.�\��I�i-���N�
t�Z�{r�&,�|�{��A �(�p�/��&r�;F8�z��Y/�� @�I��R�|�ǎ@���O�-��/I�f�3UK!�	�b3�|���9^���S5 �<!��Y"��p��	5j~:���K\��	�O�]��IP�e\�S�O�J$��䉶XhԨi��L�\����'�UAs�S"X��5�#�K[Y����y2��Z[���	�9�5 "�݊�,];���0�㟼25� ?3r�?�h�ㆆ5#�h�o0r�&E:�-'D��Q��8;Y|�"GlO"�8�9���G�Z����|��$�g}
� � �O�bE>U# �G#V�:�"O>�t#��઴�Cl�+�:1y��@2���pn
:?�a|��ɿ!X|88�#�\cVARwoE��p=��ךP���kQ`d�DQ'�%a7�m�c@���'�)D�,�f�$N�z��1��vĨ�s��*�ɻ`S�	��%ȵ2�?I�c`���K��U�L8�L�5�*D�Р��#~�l�rKQF�,��c�<�V�	��/}g�S����W�`�6G���iɀΝ�c/!��ޓ2�e�c�I�c�: ��,� '��5��^5>ʌ�6�'��03�bV�[4*!1l�05�4@!דKL�%���"T��	�@�Bݛ@ C�k<jI1s�Kc� C�	�%8�rB�׾\��tD� �8�l*r#�c\8ё��!��<���&X�&�bc�Ȟ(ZB�'\FY���c����Ý_��h������'��"}�'�E�u����#LE({�Y;�'�n����!B��\[��Ƒ�N)��*��2��,�O0Y�A�9�Ye���� ��&"O���/Ԧ+߮a� Ɇ]�>��"O(��HI5����o��.�"� �"O�X�Ql�?$���� ���bֵi4ў"~n*c���z�Oӻ>�!3'��2
��C䉵6� �p95���*�[�[����~rꄬowjه�I�-ZlɁly��HI��W�@���d�9��4�lJaGO�,�jr~�Ѐ��=H4C��.(p��Ԛ��a���9��"=ɇ�i,d�e"���%?�1FnϮ�jl��M�<z� �)�A/$�Ȕ�&��]$<!K�!D���d��)l��7���C#> �(��@�O?7-˨5P�nǻ6"Ȕxf ��<r�woL��l #+{�6��~�Ӊ��L�oט�AS����,�W�N2>���Mڦ�sѩ���8���	�H`�j�4�H��[�!�ļ������~���U�� b�,�S��yB���;!ֿ_�iK�o��V������L�h���ɸxE��s��Ah���܁!�"�%�dp�M��g����]#,rb�r��y(��ZX������@��t^KӜf��H1�%V7�0<�q���ۖ��0.��QQ����t���=G���-o�`t�BD�L�~�dL�c�~���F&��)�'\�RŊ��U8�j�
�Ê�;��\�'r�ɠ� ��t{����˟�]���p��Mܧ9t93��"|;�#�N�:s\�=�I� �F]�v��kN|�>y��*e-���!��B�Z-x��HQ��+d(����H�3>U��◫�W̧=P��ɗ�ʽ�ӈM[�|,���Y�Ug�`�&g�:��@��ɝFh���$õ^R�� �n_�2#'N!:BX(2�[-*�vR/h��c�]?�v�
����h�	;r�ԩb���)r���Bg)Oڙ�Ůբ�B���9C��c����ec�Fq^BI�a��;
lH	�'��5cp�8eP$��!&~��2I�L2���8I���u��9d
��;Ǭ
��OHd#A�Z=V3R(k�NT�A<� ��'�Z�� �>.����K�D�|�����9��c��R18y����cP���'pFy�3#��@�CE�	9a6���'W�$A^�R@�����)@x�+M<�#��Q���˓y��л��T�*�̡3$�M�!�d� ��"�nF�c.�완���!򄖽P6�ؒ��8^`�C��!� 8}�y�M�,f������o�!�DO/��8ڃi�~EB�S&�U�w!�DX�d�X�.�<RSC�5�&�
�"O���&ʝ	��V�@�Fl�&G~�<��F��"h�$�7g�`Ȳ �~�<	7�sc.!��1o���{��_S�<'��W�J���� .a۰�{�!�S�<���;n{t�Ҳ�2�v���$�P�<!��in��� Щ2xD��,]`�<If��1�l� fd��}�0��c�<ybBʁ  N`Xs�/c��)p�ƙt�<�Ѧ��/�����زeu��c�oq�<9�i�{�T5��gL�i��<ÂEs�<Aq�ͰlF�x��"�y����O�V�'m�a;��m�'[@�� �앜=ZT)��J��-3ل�S�? �eRp�|�����ϊ'&R൉�"O�LӴ��D��#�FI
�X�"O�E��H�(���z��:�rU�"O��J@)l�pt�"`�aT���%"O�(QAWU�����y(�H��*O,Qy�j��u�N�SRН~�q@�'�Ha0�$0.�(0 ^g�`��'b`���["b��� �
�'�r�X��!�X[W�6=���1"O��S��<{��ehd#��F1YT"OҀ�V��;���!�X6��s��̋k�$$��N�������;.t���K�|�"ɰ��րy�!�D�h @��C�4X���54�!��'l����7Ɍ�<Z��	ع�!��4a�֭�Q�X@��Ȝ*	0!�;O�55��-	5^)��GF�3!�I�4N���gnB�^��qS���!��~tE��E� AC�,L�!�d�.=	�8�b] wRH�`?�!�Țu���d��%�*�(��[!���.��I�)ʄxm�(��8H�!�N�9(��`�xcVÈ[:t�!��G�F�*x��+Mt�bT(۵b0!�Dц0�P�`L-r���􆈻<!���c�E�2� ~�i��(L!�$ ���DCt��<>�E{�䖛h�!�d�#*> ��
O4���x����L!�$ b�*�SE_0D�<ѸUb'�!���z��UZ�O�7y��蠊[�!��>��
� �*pj�����!�$�B�~�bP΅�*S�)[ЎB$(�!�$�^��t2��	rK&!9�҃~C!��,�	4�ǈz0��x��	5u!�ZN^�[A���F{p��␛!h!��ֱJ~hxQvl̈�r��d� f�!�$�,Z�|-�3�j���%+��!��4.L @U��|�
��o�!���s��%RAM��L���V�Q�!��'��͑RO��Q
4I��*�aBm��t�
2��%��p1-%+>�t)1IE�`��S7P2Q���']>��!aK�?t8���)[؜Y���䓫^����gI�#�\���ŉ5I�bGڻ6��iX O�1<�.�;գ��y���R/pu��+ڼK�Q�7��
�~���Q�\�рڝi�VIkt�J��?E���~�\$��Ȍ37M��r��8�y���-@�h�c�� �oQ�j�Bem�� 0��F���&�$=ZJ?���ĊI��=�R.[
W܄`ᣃ�5>�~"e�/k�$���[Mk�q2ɒ/<R�,��(ݖ��Ұn'a,��'��B��LJa	���D�A�È-dccc+�T�1*$�\�Y<��6�Pv��M�	6;��v&%4�cC�^�_�C�I��8�S6���#��%��HZ�m����y�+�'�R�mi�Q$7����d*���E
0c�15�V�'�v�I�jo�����n��22|�xc��� �.��hE�Hmx)'˗Ꟙ��,QV�׺�Ӻ'�����ڳUԼ���%X!wy"���� �O~�:��#+*& Ѡ�VNC�$���۪ݼP��j2MZh��Ib?��]�Ј�aزD�2pYј?�Q����K4���Ӂ#�ѹ�"�u[(�[�L�NO0:h�[� ���b���"b��i*�m; r M"*O��*��D�\��DH?��y���'���"��-ld��Չ��z���5A6�lc'���=����O�gyB��e��ᱭ�	e}� �I�-2t��Yb�:�O�4�EL/y�8Y0�b�>�`˅X�t������O�p�wI�X��O�^��<?��q���\�7	}�$:E�~"�^1,p�i��e�6C �i6�
�^jn�P��Y�F�iO>Q�O�j�d�5~=��͟�D���(5���QG.P�E�V��F�I�;�~W�6��! Ђ +�|!d�'������1r�к֦GA�~���+� ?D���O�	�d �;�����>���4�O�Xb��(��_T0��u�}
� ���c]O�����Ԑ]�$Y�ǁ���T��ɏ3��I���u��,��a6:�*4�4ߨp��R��u�i+?�:�]"+_0�Z#���mCѩ��4���$�	�}���R�* ���ٱ1w�ȃ�"ğ�OX��W�݅0�UBF���#��Eh}��Y$0�&�H�-�<��	*����O�D �a¨d[Bq����Bhb��'KH��&�sǺ��B�7:��ڵ�D>��|2s��,��x��	M�KH#?�BI!w� ��@n�8��bP�t?aM%2K���d��r�\����۟T�?1�L� �dp3Aщ|��%�r�2cI�T�:�O�I�'a�7͈��2	�z4F-s���:�FMsׄ�Op�=ͧK���;ߺa3��#n�IГJ�(o~v|F~���8<s�F����o�T_�&���a$�� ��0Q%"�9�\��O��D=CHI��G�!"JEw
�N��D6z�|Ju�Q�Kly�q�?K���C�3*]�d�C�#>�XH��;}��Ot�*a^	� ��"}n�ݩ�#$9?���0K@�,���ν
��@��?j����Ѭ<P���$e��w.�t��P9^Mz6����'p@pE��h[�P����R�S=fT�L�0䜐	�T
acM��p=9#�p�ma���,�V�fꖖ4YbG�+LOt 1qC�O���mO��я��$=nI��)�0{��8ѕx��C�!v�(
u�۰ ��p�����ԟbJ�qǚ���		�*���eG���'%*���i�A6�H3?"�X %ٟv%�JD@�FE�+��	��X2-�j)ӥLT �T�Ɓ� ��ԟў��%�����l[�0EL��L���D/hL�`ò�!O �<P�d"��ӔW�\sGI���yM]R]�}Ɯ�D�  pOS���-��M���$�HO��I�:嘲`X8Z�3[c�~���з.9@�� �φ)z����0��I�����*�Mh�l;s�"&��p�GP����'��z�(���4��]�-�4@(O�^�xX��r��*A�L�<b(1�Gb<��\ڦQ`��i��|{���!70J�oZ>�"56OZ�ЫB�%~��	Q�˦h	� 5�.A=*Z�/��Pe�˓�hO�Z�Z󴩡����%�i:0pf���1G�:
:�)*U�OЁ1��(O�n�:v���� 6 YT�×E��i'�S2�]&��h����&\79L%z�АJv4��F�(o��t��	�]��.�>���Rg�1~�`WiQ(%����Ħ�B��|ZB��X�2�
��<V|�u���O8u\��~�'{Z�a�Kn���T�E��	7��G�<���ԷH��������;���*^]�����?1dN�+,ѫ��ŕ������c�ɇEQY�V��.m�F�:���n���ɖ2�th0�ǹM�>qI!�ӂh,LiSJ�+n�����j.�Ą;��䩓�(;jh����U�L�q�L�zy�����&9�`8X�֟ў�J򄎋3��{^��F\�d��J4+�e�PQ�gE��lfԅv���֝��O��s�hXY&��Ȑ�L�Хc�W�4#ߓ�yw�I.`�������9�����O�g/��BvX�lU�ß<KW�;���G��+��9�,�|It�Ұ�́.��#u�ۡ��D�BӪr����b�ĭ.JI+O0Y&�,$適c�8B6E�s
�l@�	� E�����!`[��d�h8�bкv�lSgΌ"o��i̓�2����\�g`����N�X9�'�,�����*�:`�h׍Lx��x��� �*Y�B���f�#����"ƌ<��
�*B8��,x�b�*ŋ
� ."��gҮc��;#�V���D`#��=�\9;�#ӟs�j4Z��\2�JЙ�˜�w4"�y��G�<����O�v9�	�5{���e!�<�6Q@g�#A�]��Nl6P�w���*���y7��x0�G!^�AE� �v� X��3O��Г���?IwN�x�i�ּg�6%�I�
|q�}g�G�'}ZŨ1�I���`�
O<"_�X�ݴ<}v u�F�"�^J%���%��9`��v/�tj`�D�P
~��'���yկC#��P���29��2�'o.}�BQ��x�hd�_��8���h�D��W��^���g��/�.|l��L�0��W��9v�3v��OXm���&W��$S#�F�2$�e�"��6i��ip��_u�j�(GJK&m�ax��Y�g�����GB#���a�������{���ަiI��ӪD(pP�GޑpG�)��&V]��i�DZ22ߺ�rJx0K�n��{"��'0��#��{ҋk��,qJ�hP���#���$ߐuo����OaHƁ.tX����K�Rю��,��L��d=B�&m�@₠8T���/gӛ���6-UB(�*��%�f��Q�԰v�8��)� $�bi�i�,��I:����0,�����OP���ɶ�Rd���y�j�`6�'�m�U!U6������)&�P��޴	󺄋D'_X;R�rEdȟ��u�Y����ӂ�f♰� /}2�}~��1e�Q~�a!�ny9�a��#Q8\"��TYÂ��'�d���<wA�-KFJ	�h�U`�M��i�@'���1VmXv�A%fZ�x%��V�Z�i����� t`�� V#3�tJ��
���;�B��?1�.K�p����O�0��6�*��r'5n�09�ᖭ`T��ç�{\�U`�&;�n{*�y��ٹL7l��B�>~��<��� u���qS��3rG�C�m�qOz�au
��4���)�瞻zv��9f�>��Ǌ\����o�6\H$؂'b�x��Y#�:N|&h��L�x�f|��W>m����X�N�Y��ԭ�T�-,6�"��V'ڭ�vK�*	�Є剋�$�r�L֌z`J�b��~7�H�F��'�����д�E�x�ʯm!�R��2tz�y����;�azrg	}n�\Zt���~�� ���'�M�P^�Bm_!.x�*�6O�5�'T�4Ra��j��+�* ����G��S����OO��L�2'��L�`c��x�-�N���}�~�$>��X�B(�k׉Ycn��C�%V3��$���l[�H�&�U�%2m:0�g����~�5���3`<��8��m)��'��;�	�Ӛ��ɶB
�,�g�2�;�8D��um�,C��!xB"ӝq�Y�G�;W�̈́�w;�)�A A�b)�f�<S�\扲\���#���(�ʐ�]NZ��'�z)��L@�
ԑDƊ5 ���'\O$�����$'�֘z�bt��
ֵ���e�-Pj�%J�)V'/,`\���1��O]�ӌ �AI����������bBr�xSgJ!(����D�?��S��߇mD��x͟���'�?Tv@��eG޿8�8�5��e�"5�=BD����J�{r��Ct�YM�2��HSD�I�88�m+���QcNhc���̚%���ɖ�~rJ
9(�( *O�4%b�	�?1d�e��xk$���`%��G�+Cf�XS򧟗Һ���A�8�ay���,`e�4� o�5��4؃�(�y��J�
�V#=����P�w�X����� h$\MyFA�
��Dǁ:��2��P\��X�7���ڔ ��^MPa��L�<%P(�y��I1�̕�W
��1��ؐ[0s���wNF�0�O=d�HT%�4���^ 1Xu�%��j��9#+E�}���A��T�<X�f�Ҭqz�B�T�X� Г��'�8 �,��
3��$�*��QI<�ԫ+j�&-�� o&� z��,	5:���a�"-�b��3���У*��d�QN��=�r�˕�m���)��W�]e�8�A8\8�_��p<Qd.��씣������(�@��ҐI��O;�"=��"h|���SKE<eQ� ���6f��^Qy�dS$	6B���:<k`)�!�Z��m�%ď E��y��ɖq�B��B+�`(�L�0@p�̓c�n�I����vb�h�'�K8f�# �*s�Y�#�ੁ���]H�6�%kbY1�/�5_<��Bcǩ��Oh�8)$VŰfO�+>x�)"�>�E�WH�[s��x�Q	�hK�� 3L��uG�.���e=�\ ���B>57�2�B�\�l�s���.M �Qw�P	����!цx7�����'����CʉK�)�k X�t8
��\�82���t�p�'g�O��
b��fN1a0júB5���ʌ`��y2bҘZ�R�5�V�)$�ŧ{7���K$  d���;��@�R�-�
�8���1!�|��� ,�n
e�?��``ř�ą�	B��y�c@�
F��t;>�x���O� V6!"����(O8�v~<x���_�@�6 �Ov@XP+G��܃�^�[��ˡf�A=b�Rش;�6��w���>��살�F�^����?�E��|P�W�آ\�ӎ�]tN�Sh�8ň,�M@�~mX���	�,(�=`��X�4^�*+�= �@ʆ
�b�c��I����'�&P�V��9fljiئdN	���Y�e��<�"l_+Ew��m��֭#2��ZL���/��}����*�h޶��a˚5�f�X�lS�8��Ô�|=ԙ�K���'s�Pk�bְ�?q���,ffݩ7
�"!v-{��H�'����6��f�f\S"�Vz��БD,�3<�H@�A���(�O��H�A�1R/.�����e�ĉ1ɚ�`�9a�'�j��Z�\�����"#$^]���S/xK�`�k�7�M6fą)�t(�t��!|��#��]d��X5����C����0<aHG�$��)U��S��;���"	d�n��<��X"t�J�y�P��$��P?X6�E;��4�|}2h��x]���d%��r�Z)(�Lّk�)��I�%5""�i��Q�L�i���Dڑ�2�/=j��B�H�0YNTb۴QJ2�	0G�4�.۩
��<q���'B��Q�(K�}$l����Ki�'��]kaF
q?�� Z�9�|�oڷn�1�0J�g��Ӆ�� ������P5w#�=�t���*	r��(�0=����G��(�%F�9��H���y�x8Tj�>Q �F8 =�͈W�҃K�+�<A�~�AV���hxC��9)Ls�E٤.�z<��:D��&��f<�B���:% 〸>�1�Y.PJt�
�!9GD��Ӂ.�(�����W�.Qɉwk_��1�"O�tAÏ\'F�j�M$`�ȩ2�"O| b��p^�i
�(_�(| -8P"O��6��G�\})�G�+y^��"O�H�d/˝i��e�d Ou���"O4pk� ��J�O� >ց*"O��I��۷=�I�!��D%`1�"OF�@$�o�H��aU�73�Q8F"OX\B3.V�F}l���������*O�=���%{ђT��O��D�<�8�'M�]����#z1��N!;���	�'|�����1vxRh��$ĉ7rb�+�'E�)ؓH�?whzRK�F�D���'��UAǧׅ?�<i@�#͑Fr�K�'f��g+74^�����?x���'�"�ÁI��s!������$6c�{��� 6|�"��$���s
�,_J} "O �q�j[(}�hC�Q@*&���"O,��͙�[C�hy1�N���"O$��\y���pIT�	�5"O,�i��Ӕ3&�:�G�b��"O��y�oA4%��`�P�7
|�� "OR��kY�9����Dԧ=
I�"O>��G�	y����S�'�z�s�"O��;��$P.eY7oÉG\�P�"O-�����T9� �ļ :�t#"O`��%Ԕ5'��qL��~�lH�"O"��#_q���Ӱ�	�_��y�"OT��r��=�r�ei]!KS�01"O2�M�$���#S�ܳp`�P "O�q�b��d���dF�{9���"Onq	˝8$b1���A>����"O�ha�]�D��%;�.E /�!C�"O�<�Ak uf\`�&,��t,�Aw"O\�oݏ{^>��,i&��JC"O��ju�8F�J5�X)K�X�q�"O,��� �4bR����D7{n�Q�"O����>� �r4��9��!�"O&}2Gf�1r�8Dh��\d*��B"OP���b�"�I�%K�-��"Of@�"���lH�@GaB�r;0-Y "OY�c�O6 �-����I�\* "O`Y�!gω?jf�W陳[f��`6"O������w�~`���
:��B"ObQ��Z�S�T�!�����"O�I�gJ��,{�ogt¶"O��Q��ؑB~hĐe�T_G��d"Oh��m�,�ƌ��iH<709H!"O,	��CV� ɠ���ț�}Pj�"Odp�4 R�Bz�L��&�pCB��V"O�)�$E�g�J��W S'�c"O�(P�
�XԈ(AcP�Z
��"O6��ܰ.w�!��a }b��e"O�hj��+ ��3 F(To����"O\u��V1L�d��BV����"O><�c%	�:�a�k誉w"O(���쐧k(�	e�E)u���Â"O,A��N�"��U���K�D�Ó"O�ȨDD
�.�j1"QϐG��t�"O����V	.�l�s�1Z��p�"O���4O��rM.	�C�Q���s�"O�5S�N R���	G �1%�x��"Ojs�"т&62�e	N4�ܑ�"OL�
�	��y]�q��EO�=� 	�"Ox���e��~�@���j�<���"O΀"���T�x���@�2ĩ�"O�0����_��x��,�5E"Ov�+5��6֖Aj�RTܘI�s"O�-�V$�(\�F�x�ͲA�h��p"O0�9\�v��!�ʺ.K���Q"OT�E���K����ӘXB�c�"O�|����s����H��� �"ObEP�kO�A	֤h���F���Q�"O�T2���!z�����(�X��"O�����2f��\�p"F� ���Qv"Ot<��m��-��պ ��.j¤�`t"O�<(���9_7��!�ፕM�6�!W"O�r$A�&Y�lѲ���(�<i�"OL��B��~�*��4 �� �Hͻ�"O�$YBg�]�Z��D.F�`�n���"O� 8�k%��+x�"1������LCU"O���&�� T���q-��9xA�"Odi�&P�jjV ��̇�HU�!ڶ"O�uX����L�8��Y�v��9�"O��+Q��X�zh�WJ��I�`9�"O�y�Q���VQ!j�a��@�<Y�
�z��1��\��,�R�<y���;Y �X�#Ju*歟O�<�U�ͪ �|�s,�%�J`fDJ�<���#N�P�p�?u��B�E~�<AcO��T�*Ԓ��Y���^u�<I�'�T��$�6��5�f�.�Z�<	IH*i���k��e��Pq�<���;_�DɘB�,����f�<1UCڶ"�^͐!�I�jK7�^�<!'$G�X��1b��=��3U��V�<!�,q��	�%�O��
X���S�<��Қ{b���يq/���d&CH�<a�ဢ0OPyKt �3hD��|�<i�T�e�v����J�(�ĀR�<� EV���D�f��(]��`BQ�<)b*�!m�P����:��`h�/s�<�V��4� 0��@�*B���s��i�<�e�
C�0+�3@P((��A�<Ѷ
\�ԓ# #m�a�v!�{�<�!қ2u>��P>���Ǐ�v�<Ѡ�_X����8&E�0�@n�<���C4:����GҐ5��T(�M�h�<�rD� d ���)z��P!@i�<4$^�k�U�MM�?h�sa�p�<�5��$`�� ��e����u�Dx�<��EͯU]�	���!A�ɀ���w�<����1T��t�MG���C@�u�<��U1�f	C���!0䬰���E�<�d$V&=^��ޒYp�C��A�<�5�""\��B/^3%����Q�|�<I�n�%I�^�`���8��bNa�<y��u�j2B��Yq)�d[H�<��8`�P㔨V�3.�|�i�|�<97�^�gHPH�q��^�\��f�r�<)0��H������
?��p�n�<Y�K��Tkt9C�B
;$���Mo�<�Gf�3�l�A*��Jo@y���g�<����1%�D�sě�4͚���b�<�@�"OS@�!pJJ�6{� @Tk�[�<��,� K'�Ԓ��Oj?T�u�s�<�Q����pM�/6��Ż O�C�<�q#ɕw����#%�;{�`%��|�<Qc�?��)���^�Y���i{�<A���/�6Q����R�:s�l�<A%)_j��h��f�n���bc�e�<�QdE8_p��&�/|":9)�m_\�<�?e���Tf43�A�KX�<���W x���2r��8d��K�<�0Ɩd�(����R\bA�I��0=�FA�8?��)KD/,n���w�F�<������ �'�'i>i����}�<�SiӁB	򕢑hS+F���*�y�<�&�	�~}k���'<u6��3$�y�<	c���|k�\i�B�#zT�w��a�<	#*�h���*�BT1V�*�K�^�<�fEu���:��Q'XF�ڕ��`�<�R��'s��d��aA�8me�Ƃ�p�<��A='�ٗɟ/� ��dkH�<� �-���ģp> 0�B�E�5"O-P�$��[[�qs栙�<ȷ"Ob�qf�N�X�TX�*L�S7��w"OH��.Y>Cl�����"b ���"O��
'��{
|�c��(2�$�2B"O�z�MP&z���%�_/��@"O>ի#`�+
 �u�F�1�@��"O �b"σ
Bu�@�%�(O�*5�A"O���Cm����Q*�$Կ%�p�"O�m8��»kH���d5�,E�$"O�!D�!�+���3��=[��'D���D��	m�d �!,@�X�yQ$�'D�4u���Fk��#j�i�#D��Wn9��KC�{K��C�!D�h
�I�4���{�ɒ���I�%D�D�����(F�X{�ℇs�i�P�(D�H�&#��9fJ 4,�ao��`e<D� �3��H"4h��kJ*:�H�ZU�9D��@�
�Rk���.
�i�0�bc�8D��ywI�-|�"�9a-�"W)�H��#D�����U�!�-9wH�F�z9z�b D�T�Qf��R��}���5d���j<D��q�Q1G�	[�)G?�t�P�;D�`��b;V���5.��/!�PI�
;D� �M�J�`�K��Yx� L9D��'n�6c�$0&�ъ��R�#D�ɱ��r��GN�3q�\���)5D�|��LGI�4,[7d����fE=D�ʶ��8��a���ߛ~:��Җ�;D�(�g��	|:\Ȃ���q��ɣ�7D��R��	:cF�y[�ƹ �^4
�C5D����	���ȴF�`4\�K9D�T1����iA�ϻ�T\�bo7D��cwDH�3ƅd��Y��"21D���5��M�T�P+ޭ)���.D���FD;tF�tPpMOJ�����+D����M+A����0J�Z����0>D�|��I�25(9�$��}κ���>D��[ h���h��MA!"i��ka@>D�4�5C-� ���
���UX�o!D��Wk�>mR�}С͇�`֥�B!D�� � �Bǔ�ɔ$��,��9Sc D���� 7���P�!Ӑ/t�]Äg?D�dѰb
 
Z���M�VMz���;D��cB�ί}R!��V��V�iGK%D��Sv���,D@���mmX�1��7D���@��q���P��63�<���3D�T"ֈ �Nu�y�Qf�PQ4��d�2D� �@�վU�^P�!�B$L�98! #D��q�h�5!��P�"k�04�Q�+D�Q�_:>�|��I�{&`���+D����^3y�F���6M�y��)D�P�TJա����e�A���'�$D���ce�m��!�P�u�d���%D�����+nw�(��
,lf�w�$D���G����9��I�"��	C�$D�$��̜z��ɩ!�F�\<��2�-D�L�3�ȻU��	�6#�?�]8B�'D��q��;j �PC�*�!
xмy%�'D��JB׬��C'ߙ����f-0D� ;���fբM!N�Z�l�Ѐ/D�t �d����taK
b2b��2D��Q�Lӟ3�h�bWN�̂�B�&0D��:�d�6�^�C��� v��-D�� �$��B@..����F�bN��y�"Otu�����I+� �"H��5�E"OJ�� �όyy:����M�V`HT"O�1�5h:^��sG
����"OjȢ6e�>f/iSU/I
f���"O�����X�D^�(ӡM�PR��c"O�������1��D1H$�h�"O@���ձ_����pd��s��%"OD`�&H2^�v{� B�K�r�"�"OB����J p�宜�ap2"O�ñ%F�h�C�٢qd�j�"O @��9k(У�l�� b�h"OƠJ�N��,y�u+�06YHY"O@� �M��.4��ѧ�]4-�L��"Oj|�Uǅ
*m<�A�ˤ_���i�"O��xQAD#?���1$5�����"O�q�Q�%1�J-AD�M�e��k�"O�uA���?���AL�G,
�@0"O�ȐG�R�4�A�*Os��"O������?~�,��"B</d�!�"O(̰��H���b�a� |z3�"O�]�PȂ���H�q�ا"e4� q"Odl��+L��kr��""�6���"O���Ԃ���K�lG4>��Y*&"OP�$
_�K&k��8�F��"O��YU��1��= OFo��H�7"O^E�TH�snh{"�T��H�x`"O:�����(lh�:��-}|��W"O 1� )�Vj>��d!�v�B"O�Qa�B��:=�S��X-IP�d�""OδqLO�8x��IeӾFI�
3"O:��U�}+8`{�ă�	B�� �y�`�0Iz�������|�# ��yb��;44t��ڬ��`��@��y� 2��M�SS�U��P����1�'Br<��N�"q�P)�1`#4��'K�QRP���p���擙\M��'��0��EB�_���9g��<���'8(0$��wn����Oöy�'R�j ��VN^x��E�@ݨl��'������J�)� Bתo�j�{�'b*ȱD���IZ�
 F܄�H�(�'N�Hr2'���Z䐆�N����	�'��@�zW(�Ҳ�_��(���'�6�ۣ���\3��6��0A���'��Q a�ڢPY�%�f'�)fh��'H���+A�: bt�ᓳ)ZPr�'P�8r��Y�l�qaŭ79B ���'��[�NʚN%���-]�a�=h�'C��HR��l���ZcDH3�~���'�b[���(�>$8 �'o�Њ�'Lhk#�ndl8�Oؽ�.D�	�'�yi�g�>qw�%�0Ҽ�����'�b���-�&_wfh"�f^�9�`\h�'�tp���?	��hZ�,4�9�
�'���P�T��ep��� -g�`�	�'b09�e���H*&eÜ+'�qi�'dN�w�C ؓ �2)J��c���2��|�ڴ\>�y���Q�A��K��E��P�ȓ�-��ϙ]��k#B
9�����n���!�ƽ_�( ۗFʉC�pd��!1=0��d�2��r
W�Ȅȓ=�� �� U�wU� ѷ8m娍����
e	P?=�.4[�J��X�H��S�? �Db,X�d�0� �1;�\L�"O�y�F��1kd��2�*�`�h��"O�H÷Z�bWl@��װi�&�jW"O�`�u�S8�,Jt���FFku"O��b�f�2P���f,��k�њ�"Oұ��9++� ���U�`UTP9�"O�qp�K13~��/�V�^X�"O���P(l0�AX�I�(�x �"O�Z�h֎���͋�K�
���"O`���B�MD� K��?z���94"Odʂ6�8�"��݉R�5AU"O.�[�����y��Bתz%�9"@"OZ=:@"�?Qg���"پD<� �"O�j���3:tV��$ ����<�w"O8�ʤm��R�+ōIv��v%�1�y� ˄(i�`�@Nޗx$����#B��y�EK1s��<�C`�2O*��
�yB+];`5���*4)DZ���X�yBFC4S���ʡ������-��y�N� ����4��T��S�ֺ�y��ֲXҙj6�D�I���K��y�k��L�t�Č�#�Պ���0?�-O�KS,��B���ɰ@��&���%"O6A��[��;���?�2�J!"OPe�M��BE���CC�J����W"O�}nM^`�B� m ~����s"Oa���?U$����-�"cC~!�%"Od���=l,d�+5lI�7��!"O�	�L�^��@�*VO<��"OJ�ӶE� ��-��)Y�p �9��"O ʣ.�8>/>�3"�f�*�"O�y��Ę��@�AbBLN���`"O��g�ζ%��T��Ƃ�@���""O|��&�Ј͐����فe	��"O@d9�����H�U�	�"O��yFO��&��B���	�`2"O���JU�<#"�kGaI9]�%+4"O�ժ&m�hS�9��C�]��)9"O�`�th$J`Ɖ�|
�� "O.�37~2xZ�ַ'Y$P�'"O��b��+L�!��b�Y��"O���4(��Tg�|K���GdX���)lO@	Y#!�%.��`_;1�]8���(�S��H�Pd���ja���r�W:l��B��j�����M�2��
Eb�B�	��]�p��N;�1[ëӴ/:fB�	���@���[;�-�tD*)�DB�ɟieJur�E��~�sԊχ,� B�I�e�VT� N[1n�%eM6	�VB��u�����C�j؝@i;n��B�2[������qH��Qc��B�		G��G	^�2P�i@O( e�B�I�r�NI���D�5�ҝ���M=ETC�	j+(�i6�Cb��Z2C䉹{(Ԁ' �9L� �(F*����"?��)
�\�6DB0\�,Ŏ�:��Qn!�dV�>Y�<�
�D�L����W9e�!��Ȕ�ΐ:�c-@�̐���{?!�8!`|\� ��"hݲhZ��ۉ{;��?�S�O�^ ��7z�9fL��S꺩B
�'T�yH^����a�M�Nm.D�	�'���8dT�;��Y)��T�o	�eZ	���~/�=Vt2�`A�]S\�`�Á6�yb�T��$xak\2Qn.�څ���0<���� 8�� Y�&u3��D�x:"O��s��a���{���:9��'|����©�>��r.2(�ʁ	�i;D�p�	�3u69y0CӨՈ����x2�$,8�z����J��l�B��n�<q����Hx��K��|)I�M�<�ɉ�8�^�������o[Dy��'<�����1x�tm9�P�y\��'��2F�� l��#C�c�6�C�'��A2�kDq�ڕ�2W[DX�J	�'
�;��[)6Y	�� `��x�'�|�!�a�ynT	5͂�,��'$��\�Iur�S�^&%��@�'�tՃ`����=��
	#p�	�'�NR/Z@�a0Ӭ��)�� �'f�xe�U�~�`��"3w�d��'8��h`���a�����z|6B
�'�LMc'�_�?S��#���cj�l{�'&��0s!�b����0&��W��:	�'pb��w���;��-�W��I|<s��x2K`3pU��L�(wn��cW�I��伟lD{���,	�4`X�i�/ݖ?����*�'�y�ŝ��`��I�%��9��E��O QEzʟ�����5��
x�.j��-�yR��'��<�1�"o��h
��y����r��]Ӧc�^C6	9G>�y���9x�F`�~��U�	V�<��R�Q�nCc�5�����-�<َ��,�R�(w�ϩS�Ћ䬒="C�ɀ��m��K�	/L��a�b�0#8�B�6H}���J�nݎ4q�h�f�zB�I�V~���D��Uʰ����x�C䉿$�QC�m��)��� �`N0�<���T>��j�?O���H'�߳�dz`)2D�  �D	2����ޞ��� J�>�"�6�O��ȗHN� ��k��R6)��(�C"O�-+���Y�,�oY�~͉"O*,B`���`��D-�3K�j�8�"O���4�lAX��Il��h6"O�-�fdV�Uˮ�Ci[;"���"O�q��#-��сJΫmp��0'"O\ȡ0��0 P���Ɉ�5p���"O΄�F�\�65�ػ1χ�[z`�v"O�e^E9�d@ǢK7yHx8��!�m�<�mO(I.�i�.(��M:3��j�<�1�
�.9�� �Āq�����i�<ᅦٌ6���X% �9�=�U#�k�<٣o�g�RypblW<f�aa梒d���=�J�4i�ł��Ǭa���m_�<	�%��f-����)�hh� �@�<1$�׏J�d�&�@.rD�v�<!���54�( cA"�f=�Ju�<�'�'�n�{��B�K6lh7�F�<qrEI�������v�Qp��Vw�<�3k�7�RX8�"�vF�L1�KJ�<)��_�L�8��՟H�e��o�I�<�cl?C>�� �$6\�hDE�<&ٿk�|�Sj J�hC�{�<i礊�b�DQ
S�zP܌0��{�<��ڌiNp`!�%X�:��A w �t�<sm��3(~����*4b4�Q��t�<yc��-`�H���C!����CO�W�<��Ƙ;��D�G�zz	iT#VV�<i�KQv|z�B����H�SEQ�<� �}B�/�,&L,�R`C�af~h��"O�Ԫ1�؝0�ԁ��h�0x\��#"O
e��*i�� 
�h�[;��"O0�`��2|+�4ғB?�hp��"O��Y�$��	��i8�CA�]�̩+�*Oj(1c��^����UFA-<��Р	�'����ֺ.!ֈaDX("[�X�	�'���ꃪ��DQN4�N�H�j���'�HQʃm� �㓦/(�0	�'�r=�� I r����(D�:���5֒�y�/�'N�⬒G^1�jB�	�/�x�P ���Ęq�+<� C�ɤi'����PL��P�f���}HB�I�1���ķ+r�-��X:hB�	�E�f�H�n֡9��5�GC#y�B�&1B��X��۔�X�X 
7[�B�	�,X���.wg��X�`OyNB��0cthձ��B)m��4��NT�C�	�OFT�1�N�a� "�̲+8�C�Ɉy���R��U��H ��Ɋ��C�I�FǨ���DN=#[
�	�&%��B䉫m������6{��cu��?p�B�	9!H��	_�n��q�ˋ�M�XB�	7��R�cܜH֢IQ�!�=�LB䉕��I�C��{��e�˘T�B��
7�R� W.B'K��M:q�6B�	D��dR�cb��m�!�$s�FC�I=PiEK��G59�5s�Z�f>xC�I����HȷO��#�/�MB�	�3ӈ���Lܡ��
�mC�I�SGDP@'�ÒS�mR�	���C�ɳr0�h�a�9�X{��Xİ�ȓn��iT�ػ@F�uPP �m��	�'���)� E:��7�ͨ�p�'�\��c
g��(�F�6�6���'�v�`S�6n��X�!J�=�N��')��K�$X�.Q�t��8l�"�	�'�}���	o?.p#�Ӡ^���z
�'�~}���|~�q&c��"x
�'�=��^�$�y���37>b�b
�'|��a5h�[#$��u�B�}f�K
�'���(�)]]� �c%�_�tb,ij�'�PT�V ^rX�{��r8���
�':�)s�o�-8�X���[�dG|�	�'�=����|H��0&u�iY
�';L��BI͸.�ȃ��.P��
�'�����Td��옗oNN��A
�'qfl��ⓧ0D�uі�Cb5h�']p�p!�O/����'\�'܂���'��Sca[�\�T�Au�G�$8�$��'-�H��K�=rʔ����f(*�'��eo\2t�: j�N��L)���Jʆ�!;�zh�!�
FϦ�su"O�h�盛z�%�%��5����"O��z��Ҹ3$+Wʆ6�T"O6����F(�J	ױ(����w"O0q���N(�J�CԦ�4̪u"OZm�@�T|��'h��"O�Q�*�
h(ctaƲ�`�E"O(@�B�6ʚѹe���)�� �`"O��h�c_�d^~Y26#J�y��!�"O�<B�����	a�J$:��U��"O��	�� X!��I�/��B�"OD��W��%7'�6@^0D��A�:D�� ^���.NL�Z�FP ]�"O ِ�+ދ!�u���l��Ѱ"O�Ԡw S�@T��31���`��"On����Р��	�� ��6�i4"O�ӱĉ2L��O
���R"Ov:�N+S�H0.^F����"OV!R��r���ʅ�����`"ON�xb�Dco�
'�۬M�Q(6"O0��4�-X�2��gO�mA�ɇ�kr��ɠĞ�\��A���i\��ȓa?0�E�E2FF|����?W*Єȓ0ErE(#ΫKY \�I��d����ȓ i0��ļd�ru
6!ʩn3>�ȓ*��P�d���K"���%˦3J��ȓ{�6��U!q7R�3��)�d��8�d�b�U�8k �[嚌6���ȓKİ�%R�_�<͢b�Z
%�e��Y���@Q-y_`�����R@l!�ȓk&lP���ǘ%��5J��	�|�L��B�6-�CU�)7>�IA#�b�L�ȓ,Ɣ b�֎#0��ōN	#DPЄ�4��ԁ� ޜ��T�_�]�A�ȓ���we�y%�l#�܁Op���I��9�3�ڹ1>�d� B � ��ȓy�`�"m�/�
�(b�9T`�ȓN����"!B00ȎA@��ر64ꑅ�[�h)���&^��� Sc�,A$JL�ȓtZ�A8����f�B�h ��!\����:֜�9���@F �UyD ��x��1���=H�Ez��D0,��cH���1��G��鶍Xvl����
�̬�d,42����ír����[�Bđ�]-7�2�q`D+s6��aR�L�Ӎ�-:Ș<��L#%��Y�ȓ����c�f5p���>Z�i��*[~`k��4#f�]`���o�֐�ȓ/���I����]�8 ��[�@$\Ɇ�[�(8� �?0��\A!��+b !�ȓ ZA�T��+o�&�� ��8����O#���Cʗ�_�8�k�%?��E�ȓX��Q�dID$Mo�X�����$��~
��c��7s��1sv�P1Ҏم�v� �!�M	]'�a��B�Y^��6��<2e��!,a��)�-j}��g��r 8���A,�6G�8�ȓ`Ͳ鐶Ȋ�� �0n0�݇�

z �ffJ�r�����KY"Q��7&�xP��#�T��B퇝xa~���{�-/"錅�Q@I!rɇ����+�VHtq
���@��ԇ�U�<�Z�-��Zl �w�4S�ч�|�n����X����_�}Ұ̇�(RirN�P��ܲ��I�8�r���\���&�4����Kt�Bm!�$�M��%�Z?��1Sf/
k!�*��x�/�9d���e��<l!���1ec��x�{�dY�2O!�D,J���UMӷcD�Q�2d�!�$�|8L�ã �<H�����%�!�Dەk���G��g�,��5fS.'�!�$��!:ଲ��>)\��e%K(!�dC0C���%O :�0�sI�=�!�D��p�V]q�eܒ�P�g9�!���J_������C�d��F���!�� B��­1���PwIO<����"O��Z0�<~-,��eb[�W/���"O`�[�O��P��Թ@�*	�
"O�� G��}j٪�/˸���"O~�X�A'J�BMBA�kE��@�"O.
�ϊ�T�t���Ɛ�a@H-3�"Oȹ���K`�������d�v"O�"�+��U��M)N�V�H�"OZ�UFu�H��W,H8Κ���"O���Z�i̕㖫�7u��b�"O�,1����h�ɓl�����"Ob�i�l"J|��Z5��*~�:�q�"O��(b���B�`��h1����"O )�� n6�df��{��%"O�`JcǞT�� ���P����e"O�@�S��E]4�-�ĥ��^?A{!��*θձ�#
+;i�l4�8a!�$�j�~]�E�z{d�BR#��\!�D�N֪Y����?dH%���==!�X�,��|�GDO�|{�i�)�V!��+g���Q��ʈEi�`� �O�'!����xprŎ@�8�VP2���(|!���O���g!F�#>�8���2�!�dڽ8��H_�\�4ڒ��%�!��O�^)&��h)_d�D౉�n�!�,�.(�c0�"�IF�Q�l�!�dK���q� /�>u���>�!�N�@Sm�"��DL
:w!�Z$3��Ń�f�j�l����6m!��	�qu>`vgQ 6�M���@%c�!���:_p@-Y�L����2�F�V�!�F{�L��6̟%-w�$Ç��i!�$_	m\)�d

"��H�gd�5P!��A�Lə�G��E�ӤE!�ʫ;T�Kr�^*ybnL)Q��!�D�1��D���V�d9���+}�!�$��tx�=��A��d�Ę+`!��Y+�t��.԰z��b%���!��B#&�@pk��ɀu��3p�_&a�!��V�g�\ ��1Z��a�fIϜ|�!��8b?��8��M���D�U�!��>���a��>4�@����2�!�dP�x%�p!�Èt.D�ص�#!�Dͦc��X��m�u�T�\,�!�A5A�>�"#�T�	�� ��G�	$!�$��_6�[�KUusQ�!&��)�!��ԘL��MI�����¨R�!9��X	�'Uj�y��K�:��r ɺa� (��'�$����B���aʯXAFL�
�'BR	���בl` ���J�?:��p�'���R!cС{� T�"��5�@�	�'7�12��f�̩����65�(�	�'H �BS��1�*��W.�}�A��'%��P`��'7��y�#Hw{6��'_�U	6��^� lqA�J1$ߎ���'�z4THL���]�� �0В
�' pݘ���2�(�R���>_��� �'�I؂�K-����U�Z��Ez�'�����S��59E-,�\��'��iuI�VF��DƗ!v�,���'L�`B�H(A?
a�2h-a��@��'m!#���5sz���E�S� �	�'�H!�C� ��4kq��=Hڔ��'_r��%D��6���`L�@1�A@��� �Xr�~�SÊ Gs&��"O�!���a*��K�)رU ��"O\�1#��9L�\闂D�	��"�"O�5��,[�^ܢ\S��/C�Jm�"OV�����Ye���w#\mkS"O�����#]���$1<�1"O�BQ*A�o��iB�C�-N�3"O���	I�hw�l	Q)/�"���"O�t��d ������g�>zH�"O�`wI-Ьj3�Z�wf��A�"O�u��bĉNB�R627�~Yq�"O�tg�6�(���wy<ջ�"O>Q����-��wAU�9mP�"O���K�#4]��	�O�?e���"Ont�� O�B�З��X�,J�"O�`3ӮQ?��J9f�h#"O~����X�> RR�(X6msf"O\�k�OE5F�=(BM�!�,��t"O`Çl� 
��E�#A�.:%�<"O<�OY�{�Ȱ�� �%�hIx"O��f)ۅY��f`�t�@$D�<��O�o^�<`܇K���S"-D��	�I\Gx��*�#ǘW;���0�!�H�c���
��_	v6re�dB�`�!��֒-�j�j���@'H�	eC[��!���i&4�pe+!�HP�B��8!�]�f'4Q��@X6�������$!�ՖwO�t�!K�|�|e
�k��3�!�$IU{�]U-�N�X��[!�կP�n,[4��8y�dm�Q�̺�!�dX�Vj�D@�ڶ��H*f��n�!��*`E*аգ��c�\��4�Ӿ)�!�$@�6SDf�@Ҕ���b���!�F�{��QI�g��R�8�Y�V;�!��á*�D�9b�A������˖D�!��Uk$2V�آ^�~����'�!�$αZ䠄�� ^�)��؅�L .�!�E��1�e��^4��R5}�!�d��{�"��`F�ߔh�gL׵A�!�
�Y��,��ʻٸ!xc��	�!�䘹G�^� @E�.�²K�`�!�0`�����>��&��!�$Z�bA��xv�չ<�����C�� c@�, ׽P�aeN�NW�eo'D���&��R@�HQ�@�g1��$�9D�����m��%3�����]��e;D���S�Y�'�8����ѥ~2�Y (9D����D=f(j�o�&|t�A�F�6D��y�EU�,cg#�%s�I�S(D�(��� 2����tNx)�t�'D���B���s�!	�&ŗ<L=1P�#D��[�ʋT+
i����p�Lx�1=D�,Äŉk�xI[g.�=�����0D����WQ����	Tth �/D�H��f�d�ڀJ$�� @B��XM-D�|��)IҌ)��
״�ѻ��*D��)��Y�	����E��t�Ҭ�B�'D�p�с�H�tأ�L	6Uʘ��2D��z�S!*e�y��CF;;u�Tڐ�*D�c��7s�
�(D#C�pj��6D���&�	�f� _
Դ�4��* �!��7Cѐ�2P+��B� �&o�+z�!�� )���4�^�(���[�N�!�D1L�xق]�0s.���C"O� R��!K�`y�꧍�+� ""O>9W�Ϳw���`�l�-)��	""O��0H��N0"�"Jf�	�"O��2�G#tI `)ka��t��"O�<���fى!,j�r�Xt"O����H���\3���m��q"O��I��߼=����nI�:"O�����5r�����g8�h{"OpqkV�11�tes��4d�õ"O�l�e
�� ��l��L	V>�v"O�Hh+nH��!��a
���"O�S�J� 8�G`��jy�W"O ã�z�.�Yti�"/��h"Ok��٣{�	����}�ܰ!�"O���? �!0�I6~�t!�P"O�ցA�b�D�� ���a�"O�l ��f�L1�(3 ����"O���nN	u}��`�
�m|�A2"O���6`I6"bĀ�f��8�Y�"OZ$�A�t�|]x'��qЭ!D"OJi��_�B��r�J Flx��"O�a���&n�P�E���,Of""O��2����Y	�)c���;4��Y�@"O,1B�&� tЇ��2*`�#�"OTآ�J��¥���93i"Ox���I�>z��jaH���E�&"O0�aBεck"��5E�b p���"O𨠠l<B�νqu�Ӧq�l{�"O��سL�-aGpԳ��C�\��"O$]���	0 0�@c�@=�hܚ�"O:�HU�ݯ8�=�ĉMl8�!�"O���5��+V�a{�I��oh�Ҕ"O<*�̋�7�Z���H#bU��r�"Oh,h��G�b"�i��BO>N�"O�1���7�dT���N�����"O�p��8]1PL�`���hUiu"O�ȃ��1[j����O;x��y��"O���"�9K���@�O�H|Z�"O�� ��U�?�f�'6]j��r�"Ox��$O
�EkqhЮ1���i�"O��[@*�+0uj��Ǉ�z�H*�"O8�`�,��^�>-;��L�*d�r"O��{R��r��=����j�"O�ؠ��a�vqI6Ю`��5��"O�=�� ̳-������n.�5��"O��!5���Q8}A�d�"%����"O�\PD�Շ���Q֤_�dLLj""O�t��hT��^P"�hO�Q�Q�S"O��y$�+�xt:ӦK.`
��D*O���FQ�H]���9wL�5A�'�Xa!�&l�E1�#�?9f���'~��Z��K4��#'̈�	�'2���ԟO�M��C��L@	�'����@I��*Q�(_*y��'=8Ĳ�A&o�������?"�,���'�e;��a�y�q���!��D��'�J�� o�C��5���B���y@�'v���p�}�L�����:\P=�'�:�H5�T�9�(�R7��|ip�'Z�T��d�n)����i��	�'倥3QF��&ZJ �c��5Y�'glIj�̲D���b��6�]��'؄�x�؋8�`\2��XP$;�'��x�^�>��̻3���Y�"����� @$�t�	�^��<*�M���C%"Obq�͔:�`$�qdZ2K��L��"ODY2 䚪!���rLO<�F5��"O��u,��%P�����-�p��f"O*5�J��<��Āt�Ѝs�"O�C� �;�B��P���P��(�"Oڝ:��Y�
L����ҳ<��E�"O�8h1�7gڄ1T���:�h8�"O cD:*��Ya&R�,�&`�"O���'��b�H�䕷k�@܁�"O�RGIM*T���yrJ�;��y��"O*���fX�)�����#
�z[6աa"ON���2�.]`g�=V`Ek�"O���L,;Y\�pϝ� [��C"O\aYv�_Z�r��%��9@7"O,D�w@�3�J���ߛK�\��f"OxhI��J�]�h�jw��%?����"O}� V� ��$Ӈ1+¨��"O��"Ӫ�	zTyiщ�35���a�"OXz� �>ވ��ǩ�/���K�"O�)� ��0ʡY����/�l�U"Om�Dp�z��̼��]��"Of`�V�ْCL]�C�6��i"O�ݻ�n��93�-x ��.f*`�"O8��2�-Z健O�]cPܙf"O<�y���STpAI�,�JLP!�W"Oh��Y)��Kt	V?���_�<a&�Q54
�Z���m�b��q��Y�<a֣�N���y���2�����`�<	Q$O#b��*��k��H��g�Z�<I4�;���C�2r@X!�1χ�<��+@)p�ԍ*C��q@��4�y�<���݌r��8f���hqH�)���i�<y�A�z���ӗk�6@�(���$�f�<��;u��peEM���Mav)f�<a���3L&��a�V�Y�4ɘ���V�<����"6L�@ؤ��:0ۊ����R�<�pNV5����ʖ�v(�"��i�<A�+�r�\��`C]���M2d�Hn�<��6r�Y�KQ.p.��i�a�t�<�V��'�x��"��
����2��I�<1"ıkKRQj��5b���B�7bz@��.ZwxXY��R:lC�B�	�VҮ}0��U�#kN�+%k�ZB�	!h
&@���Հ�*qzÆJ�~�B䉭�Z��5�ت�X)����q�B��]F��m�Z[:54/���C� X���+���'d2L$�����_��C�	�Z9*l����,.h:Ph�ㅰLjC��{:�}i��L6h��Z�ý��B�I�TC�!c³(�,�ّn[�R��B��>��E�SI�fE�����(O�hB�I'HL�AU'�-��9b��I6$C��eo�!0c��&<�ԩ5+�n�B�I����{2�wf��,DG��B�	)�"E�Ԃ/� �@R�Ì5.LB�	&�XU9	F?n6���e�G�	4^B�	�B���ƣ�D��R��?j�~C��JPK� ��%��K�z��1�'�R��+}'�=3`��b���'*��6fY[�$ܡ@nq<)P
�'�r��F;o�dh�L˼?���C
�'�
�C#�Z���LB'$J�c� ���'����4d["��ˀ/?�1C��� F���ޡ(����a�ה>'����"OJwn�	U =���UAsرS "O*�WI/N6X���	TH�0"Od,��	�>i&��jQ�� \;�Q�"O<��v�9S�N5hM��e!&@(U"O��r�W��S�k�G}�8�"O$F혈f��@����jr����"OhM㣒�a]�mC�MP��x���"O��Д�ݬ0x�ဋ@<F|���P"O��yA���J�(3*U.a����"O��t�<YF�Dn�%`>�s"O�홢닖>�*y�q*ղ-Y>��G"O=	EDR�4쪘��B��t� #�"OL�W�	<`�(��
(r��j�"ONЋ�	Ǽ:a�mK@��J�j�w"O��3턪2�*A�!�J(�K�"O��q�%B-�P)[|� �9�"O2$q�Q^4@Y"�>"X�x"O����Mٱg5tq�\�uv,!G"O� ��+��!F\3�fS)y��h�c"Or�k­���vr��^��4�B�"O<4�%��h���Ss�47"ON8�C!��L#�)E*^cH��"O��3����i��0;v	�wZ��ا"O<��8U@ s��Ǎ|�|�kv"O�[�)<z���($#�D�V���"O̍2R�H?���2��p�i��"O����%6K�<��%��y��i �"O��c
(��Uc�'����"O@.M�.�b3��|�B^8�y��O"WP�ڧ��`���֦^��y� S�R2��#eܵBl�A�ŕ�y��'$�l���:#˾��Ј���y��֕6���x�%�p�*��%��y�!�8X{H<����5k����'�M��y�O�4L���.�pY�}��M[��y���G�R��Ꮝx�ഒ!�î�y�@�7PϾ%�O�i���!�H	�y�Bq\����-ܭeb����d��y򁈊~���U��S���wc�y��� )�"����&b\8�Wl��y")X�4EzC�۱F1T-��Z*�y�ŏ"w�t@����=�x,��gX%�yr�O�܀�ϗ�<�J�[�H^�y���+�2U+[���%�'D�k�'J�p�A��"**$��c�Q� 	�'v8yh`��L��ܙӊCC� ��'��X��Q�O.8��m�:?t����'Ԇ���E%qz Z�P;	��+�'���sl9=�!��f�7�"���'�9j�A�$\�H���3+���
�'���U��o���'S#��
�'�5{6&��d^\2�#R�)�����'\�BbEE�A}�t&T%=R���'פs௅Lz̘� ��mQ�h2
�'S���ԍ�f�0��E�f�U�	�'����V,�x9|��!ɉ&(F�+	�'"�IB@Y��m��̓��' vXX ��
n�ŋE���Z@��'� ZAV ��)lBj���'u>�����3t�f �#�6���i�'��,��a�>����@�ݳ:�,���' !�aB_�o츙���"`p<��'BHT�� ��,0���a��P��� �;ѭߛrf����B��C�"Of����1�FШDC'.���"O(d�S��nI�!��H�2-���"O�a*���C�(S����ѱ"O�$�FH� �>@�E��$J�B��P"O�����7�����ʍ;�`#"O@\R�|Q6 R����P�R�y���C]��K�P�Y��CJ"�yb�L��`0V+��FI
��O�y��#���6nG1����D��yrC�%guF�q��S¸�bł�y�H�wH�1#d�FB�����y�� ()�)�̓<CZ�Ԡ��y� C,_�X3a֊F�D��-ͨ�y2����lʥlL>�h�XD$�4�yb$�6� �He��9�����#�y�!%q�1��ߤo�T۴m��yrg�.hk���S�ZDYį���y���67�����	����߮�y�
]<5�L8���f�U3��yҦ��2M�q���h�N�Ҋ��y�螸#�h	�l�Z �J�+��y�n\�m12�����Z�@5�L��y��"H�-�u��D\���A >�y�'�sQZTb�-׀C��2����yRo�5pdZ�J���3i���.F��y���;=��92#��'\��"3��y�%Y�X'��`�+i�� $(U>�y��
Pn����o(`�>�Rb�'�yB(�MH���(�и'�y�JT?pJ��UJ��lnн ��y����A����Ыlp�K����y��#nL����J*u0\��-�6�y"T8�Np�W�KzO��{�F�y�mP�c�|dY:t���[6N��y�c�_���`-"ǰ5���.�yR��$���'*�� }D����L��Py�e�0�Z�'cs�l���K�<��f��%Zȁ;�%�%J��N~�<y���57�$��ԇ�3Q��GX|�<��F��X�� C��j�v��"&�S�<A���V��q�@�9]�Uv+�g�<Ѣ��57�h��@#nl���H�f�<ɴ� �t��\�oC�%la t	�d�<)�I��Ы&�K+��)XW�X^�<9�'�mJP%�G��U��p�Br�<ae"3m	
�w�E. :v �ge�e�<�SL�I1F@��?J�FPKeCSc�<Y��?-w.,�+ͺ!sd��5F�d�<���	+8��IԲ%��Z]�<�4�$��<�K�%9L�P����X�<9�G	S�����Υ|�zlB��U�<9r"��l�M���#�҄(�E�<)pÆ/��AkG�X
9p91 �@@�<�৒�ۆ��4�C��08�F�MT�<�cC8e� "%�Z�g[�y3�X�<�2i�;'�u��nG�mct�j��Q�<�t�V5s|б��������G+	O�<�r nZ]SV��6S����RI�<�G)�`Z���+�*�X@ҵ�D�<A@\�V���1#�=HK��[E�<�eC�i���c���:��u+_@�<�Wbpb��5MC�l�u"O���k!w��w��:��Tj�"O� ޼3'�J�5T��#큐b�Vq�"OUQ!��*�X�3�f2|sh
Q"OzY"s��t���7�
>���z�"O�٤oJM������p���Q�"O"=x"i�41|��#���+rȱ"O�)�  �A� 9��$��,~� �"On�������ئE�xi,x��"O(�1r�Bc�����Ȋd��T�E"O��Bd!տ5 ��Q� 6����'"Oȵ�s#+2�}��
�F̚t�d"O �B�`�"���^=,�~D)"O��F��|j����e�M��!��"OFP�S�E�5Mh�I��B�>r���e"O"0���J� ���;�+C6se��Bs"O����١/���q��P:S65: "Oޡ��*b�F�!�
< �IhE"O��@7�S	����eLW�@x�(��"O�x���M�V��J�꜕gs&���"O��Q��1�����Y�oF��"O��k�K�i^�M��M&:8�[b"O^K#��z'Hq[f퇑�B�P$"OT�y��X�p�v�)�	�98��}�"OEC[�%:��*ri�i�@�"OLH7�� 6���ǎ�6��@"Oz-`��[� .Tm�m���HPt"O2<�6�Z׾-�%lA
<�^Ƀ "Oq#W֟)���Šy�0�"O�P���ՙ	�n�*a��]�s�"Od;e-{�v�aS�*q����P"O�&a/*�J5�pJHh�M�t"O��K$e���(��'�)O�i"O�$ 1+��57��w�ל0A��� "Or�)�L�_"�}а�;]!��d"O�l`�ǆ(&�`�`�%u���Ӵ"O��S��6�lQ�@(U��~�Gx�<�CKBWnA{�䏚B��Z`�Qz�<�I�:Lb�R@�!F�)*���Z�<YV�\(e���;��	�,I�w�k�<�S�s��`��[%�d�IW)BA�<��͓�%��a{�
O�O�֍�Rn�t�<1T��r8�W�E�Lj�CQ/�p�<���ݷq$�왠/M#E��sCb�a�<I�aFm�<���B�(K��e�PDY[�<��!��/�t9���7svHC�+�U�<I�NÇ46ҹ�S�N< saLf�<���:c���c	� nzj�A�W[�<�pK��A�'�c�e�f�LY�<���AAL������8dm(�W"�\�<i@�%N�ty��1(P�A�cMW�<��#<@����*�8YtI�]�<Y�;c�J�bBƂ!K�Ys�N�<)%��$[�z���lB$<{X�����N�<���a�9H�&h$�	��V�<�I\�Q���8%�*c��)���f�<���L������H�O� )�D	n�<)��ذJ��x�c_8�F	�#Pj�<��K�YxRe�pA�6�&I����`�<1d�;o>ҭĦK�b�4Dc��XA�<�L���Q��׉�n�
&�A}�<� -�>j�Z�I�NM::�u"�KBC�<�BD  L��)�,�pT��vI�~�<!���,�����A�)VY�a�&_�<��+�?z����K�>��1�p Ss�<���;��836Lm��Į�o�<� ���b	֗@\��2�.ʻG��q"O�� iF=�}��N9FL�h3"O8kC���%:"Ђ`.	T*Bs2"O$U��.�2�4���F��3E""O��y�d�c�b�2��@�C���
$"O�L�b�˴	 4�{ƅ��T|��"Oj���n�<4&؄:�U�t`2d�!"O*��G
r�T����(#2v�ZW"O��Th���t%��-E�49�"Ox����4v�T� �\/9<�f"O����aͅ֢푇/.	��P�1"O� +��/�V��c��z���"O�V��C�����F�X>��2�"O�����H��-G�-%v���"O�U+BLYi#�`]�MrV	�S"O�LB m�w�T�ӂG��D�T�k1"O�UX��ۊd��p��tU[E"Oʌw��Kݺ!ؒ	�g�j�4"O��e*��
��l���S�d�<iS"O���<�����6^\�1S�"O��#�啸��T�q�K�H(��0"O����B����,p3��}_D�R�"O�[��݊4,�=���Y#B��Pr"O~=ɶ��3K�Fq ���:<:�"Ob�EM�:3�ؕVYv��%"O��pâB`�LY���.q�MJ"O�AE�h�\qI�Bлa�5"On�#�`�$�zvd"�$���"O���%�F�#�j%��"�"	�@<�"O���WM�sញ�F�W����+W"O �aT<(�RX*�Y�c�4͋�"O aX!Aǎ3�d8��4�r}��"Od	�#/�n�f9�ךa���h�"Ò
 s�VU�G/�Ly>uQ"O-�ЪY���3�_jDL�Q"O��Z��܀(����M�����"Oؙ��/�/p� tc"�oL���"O��XŪ��Q�(B1�ζP�f\��"OVd��ŉ*�ιp�NA8[t� �s"O�5��k��l�N��rV�܉"O|Z�C�h��vL޲K߮ C6"O��:2��grRP3��^�)oV��S"O@H��W�o�4�)���Hqr���"O�Eȥ��	2�h�5�@�pl�ĩ�"O" ���.I����֝%zD�q"O��Aϝq������F��"4"O4	���*q|�@
�ϝ�3�ք§"O@�H#�^�$ o
<h�͠�"O:h;���}@p:� 	M@m��"O��`�
B
$���$@[7B�ኄ"O�3�G�(��sH��{�pq�"O<q��� d�x�{��M�i�6���"O,�zA�rYX���
�<!����"OxY��� 3V����rJ�]1r}�"O��RΝ�*�4ۄ�*䈻"O&��cf@�CsNɈ�GX�$�ձ�"Ov�9�C�nTr�W&�l6�5s"O�r')�
�M����'� J�"O�qr#�L�[�0!;�C·h��i"ON )��W##��"��ͺrf�Z�"O2���޹|i��j�@��I�����"O6���-��e�M qOTrX�ʔ"O(��&�Cƺf�éDT����"O�ԩ��H�]��[.��bPxܢ�"O� �|���
��ã�S1�����"OX=�bCA�W{t)��΢����"O`a���t7���1��'�6��"Oʽ��nɢ��1@�Q a�1"�"OP �VKޠl��|�'� �p�)"OB��6��)8+��)�aF����"O�Y�%N�7>�rE�VF_�X���"O
��f	�4���i׆�=x�ph3 "O�!^n�NYj����Ҥ�A"O���f�5o��P�7��k�"O8���
Ú9b�I[�*"z h���"OP�0#K@�2���K��$��$"OT�5I�-��9b�G��)w�l�4"O��#,�ܵ���X�Jg���"O&� h��aX�|iL�JT�,h�"O�P(b)ÖkT`�8 �;`��ř�"ON!��%J�{q�I*`�P�<}B�(G"OXE�t��3M�D�6Nŧ!ʒ,�"O2mB�I�rt`u-	C�Հ�"O$��J�NU����\�X�l%ض"OJ�3o�K3����O7͚ѩW"O\� &�ǅp�̀���U���YP"O�	�&V��B4b$���6����E"O�|[ I�b#j�C�f�H�b��"O�Ӏ�V�W�Ŏ=q\6m�"O�a�paS�q.e�fDY�^H0��@"O~�S�U�w��G��M?�-�e"O�����7A0U#�#�;f:�Ԓ�"OL( /���0�$X F,�麢"O1{��+]�x ��I$|٠�"O$�3@�8uCX����D\U	W"O�r�h���E!����"O$8�qN[��4)ga�%l�
|[u"O.�j��� y������-3�p��"Of ۰-�l#��"%�H=d]H(S"Oj��)%\,��A�A.7C �0p"O:D
O�H*��q�V{��`�"O���` 	^�`����?��$��"Oh-�$�T*{Sh͊�ܿ;�p-�"O����F> u �+��R�7ھY�"O������4Jپ/�h���"O��S�R�ʴۄ�,�h�h�"O� ɇl��Z���fL�!j�x�#"O��F
?pɞY�#�=]���)a"O
�:ǧ�%�ȱ��I�"���"O��c���	Q��P��ja���"O�U權'\1�m� `*|QR��"O�X���ͼU�H�"�/˥	��)��"ObM#���)_��M���~��k�"Ojl[��E�����J��Lnt`�"O��Cg�D!z��8ap$�� Q�!q�"OR��F$7G4D�M�>��1��"O�K��: �p%�� g�R�a�"O�z���+Z!`q���k�0��"O��"�I�&6+��`�#V=	OPh �"O�-�t-!d�ڑ��b��@�8Ԣ"OF�x�@M"(Zp�4�(�l�"O�l9�	��&N\��O��| ��"OR���!/:��9S/ΒE)ȑ�@"O���PȘ*�����,g�x3s"O���Q�7
&�� G�=1Y�D��"Ot���(�%#�PI�(Ӿo����"OP���aΐx
�I6��1�u �"OP�CB�7�r}�e��i��� �"O� &ݹ6h�?vP�,����~gn�3�"O�u#�-�G����u��:b였�"O��� ��@bp$�P�ʔ�3"O|���*@�5@�"]j���h"O�<����G`�uZ�`M*g�~���"O�5�$	+eMνuM�+q����"Ojl"$燾��t�`�ra"O� ��r�r|:�/�6>nmh�"O��䭊�$l{"��	Jܐ��""O��A�� d�]h `Vl��yH�"O4(��%��C��d5�;K��'"O,��@��3T�ܪ����}��ei�"OPY���yKz�ACc^�Dee��"Of�9�.���e���=W�xYD"OP8�ݨ,.4�s��"V���"O�h���޻튉��B��Iq"O�����*��]�`)͞*nA�U"O�4�1eL11>���ʫv$f"O`�ɒgƣ�Qp��5u*�9"O�m	�A�$ʌ�FCIܤ 6"O|���C�d03��/*�r�"O�=h� 		�x���O�%�"O�m�o%sY�-��aH��"O��2�/H�=�w��qc����"Od��0�_1H,��@�!���P"O�Aq��E���k�kS�b�"O��0�hWIVu"�i�14�У"O�dT }� y�GR;�ȑs�"O�����L�Z㘔�q��>o3�I�C"O�l��P5|�~�Po3�t���"O�e9��C	l����T��>] �"O�%{�)]?��J�nA%J|���"O
h�s�D�jb�`8�!����$"O*t��㊑/��-�J��t(�"O8����&2�9Tn�;����"O� )��M�g2��!�L_��Ԁ"O�d�7J�!�X��ָ$�l�[�"O���V3-�X�Z�i��)"ON����%�����+?�:�r"O��z��5"�`Qj�f��Dp��"Oz8����vmZ��3%Oc�]p%"O�Pc@��B�L2%�ЭӅ��g�!���j7��kë��ڄy:�Ŝ6�!򤜝A8؉��߶g�lz��#_�!�Ļ�~�B�A�9a�xA�B;x�!��'�F9Rl��!V�8��[�&�!��iI��ÖKPp��N�>.�!򄏢XrʭpQ���34p�k�l�/�!�d��z(&�B��A3�h��k7E�!�d�/ N0E�S�=��%أ�Θ?!�DZ)6Z��"����_ݐѠ�O^�/!!�d��v���2c"3aǔ�OمI$!���)��B�+��)��E �!�d�W>�0SL��u�♒�,� $�!�A�g�Z�Dg
�$��O�]�(E�ȓ M�a�0ᄹ@o�93��!u8p����Mr�Eu��m1�D�I�I�ȓmlX�&�T��T9��P( d�ȓ'�4�めΌn��0�D�èE��ȓ7�01��( �B����֮�����C������P$F����?n��t��\]�Q �Ѥ}j���@�i�䥆�,�!�d�G{8���2P�Ȅȓfi:� ��9��904��	v��P��S�? >0`��
�O?�ѹ��l	��qW"O6�0�cߖQ�.M��ˁ� Sb��""O\h"��H<	���%J�./����"O,��B�	-�j��iŋT�:�j�"O�ă�6W2t�	V(Tw�J���"O�U���cH�gQ�h�N]q"O|5�L�?1���f�^�M�E��"O���eΉ_.���E�B�j�[�"O��ڱ��(z����*���qIq"O���WE��#�V���*#;��8�"O
���!$�Ԉp�	�;��;�"Oθ
"e�:A��X���X�(@"O��b$ǏHJh�)�F�9@Q>ti"O�dB�*ʏ8�4��#���DAA�"O�E����/#̸".L
O)�,�@"O��{�
D

xx�����5�p)"O"m���%G��p��ػ[��EH4"On�����oH u+$̰6�]�"O mC����"�\q�+�aɤ"O�i*3d
� {�|zW+=Z�j "O~�r��TnHc&��;�d*B"O=�4��!e���	_�XԜ�r"Op|�f�Ɖ70��i[�
Q"(Z6"O�ȳR	۫3���8G��9"OdA��{G ��.�|�7"O��Z ��4ϔ�р��]��9�"O�A
ѯ2ym�q�ΒS<h��"OpJ����u|��`�m��<XyKf"OH�"D��QT*�X3m��G �d�3"O��K�@�(�ȩ���m{��rP"O���E��D��u#���]�-Q�"O�I�,Prq8�W�'uf����"O�ђ��>v��E�a
>H:9x�"O��2�K�|��(�AN�@D|˖"O8���-��R��x�1�5@���"O��30K�d��X��'�2ʒ"OL��t+J%ZĘ��Ó2�^�V"O�qq&G[���iU�^���"O4Ń�d�*k���x�J�Q8��"O
!9D�'|�\yZP��3ڽ��"O���0�A�O��(��Y�F��b"O<�Ђ�A�Z�!�	.���"O�R�����I�V�D�9�� ��"O�3�+�D�ҁ�a�M/b�Ց"O\�9ģ�,�d(j� -9��L�"O����3�&q����1%��x!U"O���D�14,I��`{����"O� C��	;q7~�k����4�@�"O��y�Ր��\�3���^���;�"O��0�cP#��8��L'�Ph�&"O�����$K�A1' �.`|L��u"O�,�2`>[-�H��d�3fBj��&"O��+�� k�q��� �X���"O�}{�/��(ߴT�Tb�=;�a�"O(tY��N P.@���5[�� +W"O��h��Ņ0̠-�#*҈
V�i�"O�T�������B�����2P"O���u���|4{�gF����W"O��Q�գ���!h�\{"OXl.�8aP<.t�����4_�!�R�%�$�7䉆
�dq �#Gu�!�<��y����La;"	�,k!��� W8N���-`Ժ����Έ,Y!�D�)�B��$\��3T.��M!�� �M0����q_���OM-w��q�"O�iqh���u�ҭE-�����"O�q���4\Cr���&�^��P"O�,;�����rwE�D�<��"O��+vl�"�b�1�j�ix%�'��bxp�2!Ñ�Bf�h!�Դq|�HH:a:���a6>�xa��B�2��ȓN
$��N�����tŝ,4Y��ȓm_��zB�Y�������[�'��ɇȓ�\q��+q튘���n��Q�ȓ��j`́�*x9�1�Ы���ȓ]7� �����ܰAQ'�^�@�&��ȓ"�<T�ca� ��l�'�����xֈL!(��w��8X��ܥbʉ�ȓC�<l��Fț�nhXը�2x�T�ȓyeȨyg��� #�P`	g�نȓ [ZrI�3���m˟�
d�ȓK� "�ʟ�4t3 ���n5.��<ߓ]qJ�{q��2%)�9�2�O*��E��I�<���N�$��G醥D�X(�-�h�<I�hȑ!�@��E2n1v@Y�' a�t�@/Qr\��`C2	�d0+�[(�y��:@Tz/7�D�CF _<�yR�X�a�X�feM�yur�� �9�y���3w�ƴZ�סz$��ٵ"D1�y�*�?�Z$��wu�)�����y"b�| "ܟz��)b�JN$�y­ƣ3���e�k��U
��\:�yr��3�� �G96�L5��!�?��'f~Y��]�G������:B۰%�'�m�J1~y�Uj婆)I����'����h��3�HT��@�=�>���}�)�I�z84S@���$)�񌕵0x�x�	�^�6��F�'&!��"�K}#�#=11�'��0����:����V7et��M>����)%���u�\�Ib �>)?!�$ţ�MSw�¶h���J�V v=���)����B��qx�������A�`$�X��4)�t ���7+v�i�
�9k��\���?!!B�m���@�	�g-�uf�{�$DZ��Z� 5}���$��r!˞(8*���C��y��jWڥ"��?)�&Jq͔��O�FyҐ?Y��L���:��1� �8fa2D����iO��TA���1;��0B3�1D��3���1�F����g	Ni=q��tE�ԥ^pt���퀢EI7��>�y�%�F,!3N��~��s�I��y��οh%�E�gF�p��\������y�É�D��@m8x�S� ��y��6+;�%�Th�g�bH��9��x2��f!N�X��ֳ/�2��d�ŏ1�!�$�h����R풥,�� ��H�=�az"�DB:8���x dַq����6��!�d��|�؀9�'���l���ˀ0�qO��=%?�B5��	]+xdҗ����� QAI(D�L�G��D��s`q� ���&}��)�1D xs�W�7��8񡣄f1@B�ɬ��Hj�Ʉb<~�:� �T�JC䉫W���q@�;�D8�U�����$}��8Ӆ�&l�����5.I�D�-D� i��B��)$�\80�"�R�)}X��'T�>iy��B�2����gE��p����5D�4��σ��� ��Ę>O����E�����d�<�|&�(xv�U���wj���<ˇ䲟���)� �)�΍�9Ǡh��(�7�>hy��O���YF�脬=n�l��s�ӶyW(Q���<D��B�� ������8�i��`�<ي��S�G8�P�,�>����ѫQE�C�I%M�������$�e�N�y,~U��Oṫ�	�Z�~qQ��	�H�E9J��#
���d^T L"Sȱm�0��ڏD*!�$W$AM����]5}��bV�P�-I���F���V|@��l�3,��a�1��?��'�4)9#lѼ~U� kBG�%>?V�b�O:����hO�O
��N�?5>`+�.��
0�e���Nq�	6q�i��p��R��["�ؘ���!�DY ^x��"
�JغM8.��Ir�	V~J~�'�r����W�(�Q�gM�^�\)�'�0�BC��y+����A6[�e�'�L#=���� �\ P*YМ�p��+G��|2�x��M�@���T+���G�Z���f�����y
^�C��O՚< '�����"<Q�����mq��	�D�fI�C��w�L�狘�a��B�I�7
|İW&�(.{�!91O�*�ZC�I9R ��҆%�� È]�V�R�sabC�I�L�|}�d�B6Gm��V��!Bb���'[�pYhR?��PF��q�j�É��'��͐�d��nE ˖NX�(�|�j%���F{���J�9��4�5M���-�V뗱
��D��)��TK�C��Nh�v&�,�r@X5D�t��O��!N����%B�16F������p>�Ď�Q��,���A�v��D'n��@j�'����a�� ���p��(W�
���'��Y'����
����܄U��$��'Q0@�
��۔��$�
K�|��
�'�@͂W�49��)r�C�C����	�'�f��p��fl�l�]�4�`y��'<�A�ԏ��̀+� �>T�ͺ�' )�*�� S�%y�/Hiz��i�'�D�ip�P�yr���4I��+	�'D��X�-K;H� ��ȇ=B|�T�	�'�S���Fx�LI�ݐ3����'Q*���M4&'`!��d�u�&x{ד��'`.�Y#�iӶ�� ��y��Pj�'����b�� ~z��ơ��t��
�O6�i=ў�>�J��Y��
WY����'D�8����$s��V�Z:Koz� �
9���^��yR%M%s�&�� J%0,rū��ū�hO"DE�E]�k�|��L�	q����~�ў"~�2����.L%x�B��D��4H�t��hO�>��FD��9Z���*��[#�piQF>D�jȈ }L,h`����9��^�F��"<E�ThuӖ 00We��2��7�B���"O�����S����e��f�|�S\��Gz��	�g��1���̓T?���F���v4^#>1��I*S����OE���F�|�ش�hO�>i�J̸&�RQ�@�e�Xx��HE���xO�(�'��"~7H��bҔ+�M����4?����<��)lO Yʰ�՘(�.�����2�z� �Ū>�J<)�Y?]$� �z���#m�1���cÄVG���ȓ5��!$��>f]n�� �
q�B�Ii}W�&��g}B%��^P;$�7�f581S��0>�J>QTG�>'�P���[�`�x��J̦q%�؇�I�%�0�Th��9���5mB;9X��?�	�,|�S����fT�C��^����d��.�9S��^������ay�>/O�A�"�_/h�)�Ď�f�`$B�"ONP!���[*J!��-'2�|A��ɢ/�:��� .����ۦ����.q"�ie"O���c��|>fX"BI�Lx�Z���?\O$(
�@�~�^�8A��P�t� �	�HO�;\�&\��B-)�
I)���6,8��O����%QR|�Ӄ-�!�/��ԛv�)��}:�ˑ`���j`n��.�a�B8D�̸wE��CD�P	���=�ēE����铒kݔ�Bt�G�M�KGmIu{�B�	�0T�صē"?�u{#��9U�HL��6Ȍh���͈Z�T��b�5���ቍG�
#<��jQ�b�l Y�U']::TSr�B�<I��� WhD�QB 8nˤa#�Q�<4��-��0��E3.����S�<�n�`����0YCz�0�k�M�<I�@��0�H=x�䉷t����sl@�<����$f�X�i�+��'��vD�<q�
��@�*e	CؚC����gZ|�<�#�eP��K7>�=�+�n�<a!�v�`D0�z$r=�3�j�<�pCT�9�i���ܩSk� ��e�<�$˂lZ@ի�Ìq.t��.�b�<i5D�7۶��)m2$�����x�<���HQf�{��Ɍs<:U��s�<�#�ۘ"b�9��3*u���M�r�<��T���]��F�j��+tK�n�<i�ݘK�����o�"~�:��s�<i��L�n�Q�K�qA<Ъ�a�l�<y!`6V�t ��$L�D�>����d�<��k�^�(J+�02p�
7�{�<��N� @�n��D�I��y���t�<��/I�iYj�q��D��`'R͌C�I%e,F @b�r�s�A���q"OlQ0�ߛ�
-[�6@���1�"O�(�a^�8��q���.$�B	Q�"OFQ�Fiĳ+Z,���4��Qf"Oڝ�uI�>j�A������(�%"O.a�@ͣM��!��Ō �n��"O�A���[�jm��_���2W"OvP3q`D(��ae(@1L��P��"O�u��e�Ŝ��$ÆS�p�z�"ON`{�ǭy�&�8G&��Di:1y�"O�!�v�Ҫk{|ᰄ%�P���A"O�qkW�zB,����@^�<��"OLUزFթS���`�U;wE�K�"O����Ɨ>;O4�ct�=/���4"O|�@1�̌2�X-q���R�E�2"OV��C�0O;����@�d�P�"OD�"d���X���jvL ;�,�"O^ŰC���Xr�,�1
V���"O,�1����x%@4���^�u"O*�B�šg�삣��*l�>0��"O�Zu�-T`��J� �>x�"Oh�`�K�3�� ��	�=&t�郀"Oph`�ٽ	p`F���SU u*"O�Xc���F1`��KL��jS"O,L�'�C�(�l�(5D�3&JT,��"O^A�4���,1;�H(=�B�1�"O���C�Ph��M�<|�:9a"O\�H�+��t˶MظiQT���"O�RwĎ@����=3M�yh"O��9u��Oc�h�'�#Cjt�R"O���A��v����FB;b����"O���Ɖ�
�1�%�q����"O<ř�	^YCP�&�>>�
!;�"O� �IB�-V<��y�	�,.qp��c"O�̑	��hf�I{���;d(�Q�"O��@��2k��ȹ�g�?W�Cw"O,���y6`Đf��uB�`�*O�9�B�?��Ƞ��Vhj�%��'3xT�6�΅@�@�����7\�*�;�'*f�(��d��T)׎��T��'!���f��Ov8y�%��Ly9�'�ڥ����{�ja��']Cgph�'o���î��yu�u`@9m����'��@�Dܧ��M2%�]+_7��I�'���.+&LЋ���Tp��'E�)��'�c��љ���!J����$,OR� O�p�\�e�����Õ"O����gP�_h�c��F]h6i�d"O�-�<4�8%��Ð9^�s"O���A瘎J��a��CX APd9����"�(x�d�V�WC��p��F��y������D,;#��s��	!`
 �T*�1�!���<��c��.{� q�AC	b`�I����'8H餟��?��@�^%E�ȱ�h�>O���p�*�OP�ɕ��G�{�v!�vB��'�`�O���Ċ�u��T���?�΄�g�_�S�!�$C������,��d��j�&�!�$	�#:j�v��3W��H��i�,O`�X�%�)�ڤn�Xl�/O-���ZP�<ٲ�0���R�
i���1�N�-�ݔ'j��e�3�	�nW����/�&fu`Ҳ��+*�C��z� t ����r��"� ���O\��hO�O�X4��NK�C`��3�D�4b��k�'��-����\��e9bb��.��Hx�'5�ɠlF�I:p�Q#��.��mJ�'\����H����Շ}t:���'������+0,J�� ʋ-4��I�lG{����)XC�����A~�`E�(ix!��4WO����9���A�/Q��hO�q�臭W�v��	,
p�ȓ`�Tp� �|2f��`d�R�T��=�	�r3��Ԧ��~L�f��&�6�'}ў"|�,�|��w�W� �6%]�<C�1PW�T<���W�<��DU�D�8H5n	Y��Em��x�bc�.H#�%/��w��&��2���8�S��=v��D!E�>���?`}��4�'��"=9"E�3z��(�/�!/D���f�'�xr�X%-�m;u� �~����f���>qO�`Zu�Ұ#Yl��q�ܷN�:Ј�,D�p�S*�		l�x�\�+�\h�'ғ�hO�����T�ؠU �U�QF��k�fB�	�
Ԙj���,e��Bb�S�EJz��hO�>�B�
{�
Tg�V<rU�6D��� ��&\��rqgS:3q��k�?D��S�W�Z?&��5��$����0o=��ȟ� �@�o�$؄�N�N
:��0"OJ���E�E�ƈ
�E@'A���"O(����ǁH���s�­7ɢ��"O̭����)Y}����  �v�R�"OL��3NI�k�&�;��@"�:��'H�C�J!w/I)0�V�R�@�1!�I,���
'�E06��Tj! Z�0�������B��p�j>YJR��B�\< ��C�	se���EA^UL�k$G�Ko���hO�>Ic���} ����� �{L�����&D�("K��Y�ʅpfB�Q���𣲟|'����h�� �;cȆ���M��cW�&�H4�5"OfXQ(���K�B= �~\���0|O�3e�"p6�Ƞ�E%x�`��"O�]��O")��=� �2�1GE_OH<����|<0� �l�>q h4�B����؍�D+�B>��ْÎXJl�����4��T�ȓ5�tɑ�D�L���"A#V%x�0[#�'�L�Fy��I�B��x�%\&}y@���Ä g�fC䉜.Ȁ)��	f�pj �(��B䉡0�`��&��w�v-7�_?�B����K1G�%6^"%Y�A@�B�I����Pe�ʖX��˲`~�B��)t�d�:�ܝ	�괳%$�8B䉠i���:-r�ps�G�!
�d6�S�O�&]�'�Z!h������e~	��O 2�̑�K&�7GE�b���9D�T�qŒ4�@�)7KZ�Lix�#D��Y��[8g~X2����o+�=��E#D��!7G�D�p|3�L
G(��2�}��Cቋ=��$ۣ���j��5 ��B�&���d<��
=��YA�U����FWzBC�I/d�Lp���+X�zʙ?�C�Ib��3�  �B�T���J$`�B䉩MF���ч��� �
�>�$�h�	V�TӖK@;��0���S=���Q�,4�ع2+�u%�l8Zu�ź�/�W�<Q�*~�Zq�g�ѩ���B�AFU�<A�oI�u�@H� ��_���Q��W�<i4�ݣ"�֌��jyJ�EiW�U��2�S�'&���
��۵:�<i�Ԁs�)�ȓq�ڰYG䚎e�`�Q�?݌����?yw�9!�HRr��)yUJ��A�K��(͓�����*Ao��鳢*�f	�ȓi�p98GDG)z�@t�M�-̎�ȓ����cLK�]�*$ D�� Eɂ5��[R$���
�{Z�}��C�gL��ȓ��y�ЍOs n�4��J{"��EMh��U*j�ji�lR�0	���'��}��d�^��vmR?^�8�F���>	H�(0g����e�^�ɳ3?D��h�/0�������s���ѡ2ʓ�hO��o�:ö��@Ϣ��0�Ģ}�&�G{��9O�ar���՜X�3ro�l���iuў"~n�z*�Q8)�T5�����!!B�I9�銲g�-w�`��voT�W���9�±"4�I	���]��p�)Ga}R�>1�̞fU�A۴�RJ�B$zvcW�<!���/�Jta��E�)m��r7iن]B�	�CB���'X��SKÑ|�b��'�ax�D�F��91t�4g�Ppk�D�~��O>!X�	[>ba�g�cm�Ri�OtB�I��ĈƳ1vUc!�_�b�
6mn�����&+T.a>�4@��ͫK8��X�"V�y��^'!���I��p�>)������B���j�f���.lH�������O?���8 ` b@��S͎�.:�C�"O��RS$X�#<���&\�TNU:�"O�Ғ/^�(ւ����b	$�0a"O:�x�P@�]xኖ-��=H3��d���i�O#bY���[����n�;q�a}��>��[�b(��դ�IL���c
n�<IFыi�b䃷��:�~]�s'Js�<�C�x�9�T�I@[�� �I�o�<q�c�`���*WnI�<B�e�RMR�<� 
!�#E�*
$�2AD��U<�$�jX���q��O�T�#�"�|�<����;4����_�v����w�Bm��y�Î�)aZ!��[]X����Va	�q�-A�A�!�d�'�=�p�O�Z5"��ۙ~ia~X����cZ�tS�Q�"`>�@��
,D�0��N1p�d�j�?bL�֩(�	<Q����EJ�fi�l�7yujl��ե�y2KՓ.�����j�x=�񏂵�6=i�'��';�>����7=^I�Ձús�y�4h	5-!��;�XP�G� O@�Q��X��d'�S�O|�I�2�]M�����H�/����	�'�ڨ�K����B1�H�¸��'x���f79�m[A��#�h�C�'#~�D
L ���[p�8ʼb
�'��}b�G/�
Z׮��z�2���'۔<�5�+{m��97I�;�X\��''��!�X0�^ ��o��D����'-�a��τ?a:�v L0e�B���'�L���( In�a�`M�Z���!�'��Id!Y�|����Xʞx�'���♱s*�C���U0�P�'I�uk�$S4Z�2�i�-K;�P�'���Jӫf�1rse�+F���'��A��Q,^8`���,�d"O����!E2��Q� $�@�W"O����ʖ&�bx�7�V"l��؀"O� x'KZ�~��9��
��YU"O��EF&f2	��ǒ�L�2AR@"O�����%=� �b��x���"O�\FAB:�ȼxD�Z>y�v"O �(�bˡ)ꘑ!�݃5�-�0"O��ٷ&�f%8�M�\�a�"Odhz af� 4� �R�zLv�R�"O�YB j��������jMX"O�x"Z�`T��bC<`�v��"O6�A5鎓�B���� 0Т�v"O��8dM�P�"���(�?%�����"O �e/ɘy�(�z��&{�9 "O� S���+9(�8p��-�!�"O$H�$��K�̵86�D�W�h(�"O���3%޿3g��0��]�̡u"OZ��w��5H%�0�
"�0�9u"O�h�C N"5��"/*�t+F"O [��02�4وE����b"�"O�):�&�@���NH?���J�"O�IY�뚫&�2�I���]uv9�@]b�����Bs������t�&�؄��%B���c���$c!�ʲXђ\y�#��H���ɨ�!�$���)0Տܥ[����>�!�$Iv���Sd:T�lP5�ҬLw!�ґiT��L�P�Hũ�`�7BP!���kr!8F�ϻ+�Hl�6`C^X!�X�B�ֵ�o���p�'!W'|[!�䒤��Lr�A	w�hAqa��	,!�D]�er|ࠦ�=Ej�Ԁ�X!!�dGrQTX��Ԍ��=	T.��O!�dM
X�(ؐ�gG5=������ӼP�!�S[�Tp�ׅ$Q$ր��LUR>!�d�I�R��!%Ċ%vm�q!�=(!��P�µ�Į��V��� ���/�!�ęZB&%��H�@+���-N$\\!��k��`���� ���'��3	I!�$[�hJ<�Ѣ�ț!Va�AnX.H�!�� f��d�ߣ>!����B�#L��i�"O���*�)G�x�g�B�M�F���"O�u�b�]�s�����Z��X"Ot`�2-/,#�=����7�&L� "O��s�J3����rN
3�L���"OB`��C¬r�l\�U;J���"O8��1H	I�����|�l��"O��t̀�/�ک;Q�_ ~r �"O���`'�X��%��o|:N�
�"On��d&�U�0Hy��
�]��"Ob�ұ�3DJ��&K�f�,�@"OF(���I$��k�ȅN�a�"O<3w̉*���:��)3ڥ��"O�WS�y� #�m��9�H� �Yzy��'Z�e�e�\ �8�ᢗ0	���d�#B�Ls#%*�`$����!�$�KzX�d����n)�ρ$a�ў���S�]BL�sn֣<�vչ5��!-�C䉺jrj�B�o�H����BڤHW>��&�S�O5�is�$��#4r�xv��M��)�"O��a`��.�B���P,(�<	CV������'^�����LM�D𩷫U7�����5?��c��z�g햅~n���W�<q����BH$�Y#�V8>Ѧ�R��e�u8�{�)�g}�k_Zv�t�r�!`������yҢ�"D>�$!���f���K%�ΐ-�=z���a�����Wa�	p�N9H���A�i �azB�%n����D RF?Ee�k|�G��l;������Z�<��0ԴI�l^�%���P�K[�$���(F��g�~E��:Q��5�L����S�NV�<��;=��C�-��H-����׍-:��c*}��-���I-5��#��VE��hg��h,B�#q������N���hљ4&)*��$t�t�'���ٖ)��dJ���E7 ��|	ӓ$Pj����ڂow8�	����Y�g:9�E��0J�8B䉂3����q�I:p��`󕏁�R��b�h��oA*P��4�S�G��u U��!_��Aq��-E�B�IЌ���/)N��S��NhQ�����F�|�'��I�Ǚ>-|=�E$_Ab~���'&���O~�P��=�3H�d�!��պBR�q@׹k�dP��h�t�!��T�#���&C��Tr`iɦ��7u!�6�H�c��Z
S���7nH� �!�$FB�1�Jφen���̑g�!�� ,!'L�E��	ZL5�)O)�!�đi �x�� Vc��Б�0�!�­_�H����;W"�̞4-!���C�����Z�O5A���=$!�$Wy������<c .�#�$X��!�E��u�f�K9W%��#�C�!��H!
Y:�ch�|�ӡ@!򄅗;&~)�I%�L��3�Ǜb�!��G�?��Y��̖�O�t$�Ə%�!�d�"h��%�r.�
[�<�jd��.�!��y��XZ�,��M�U��|A!�d7r�Ҹ*@��=F�B��S�X8!�$4Z9"`��=�Q���$:!�ϿX��(��ŶU����N(!��P�Z��PJG��,:�%��x.���cA�ŭka��N8�@�+�N�Y��C� �� �W�]���;�"O�؅`N9f(T��Gk�y�8��Џ\�K���\�J�"9
�D���f
Ze���oF�R��ͪ���� Y�W�ђBTJ����ǧ8��HK��}�54ET�Hzt�Sk
�|�wi1ʓd�j��� �a*@A��~�6����\,ݣ	�3�V� x�I�ꄿ_%(q��X�2���W+��ZЫ�B6�p>�Q+��!a�� �Y �еɇϋ����2f�<I�&߿-�d�jB��%4�S�H�re���<�(�b*�a��7�Tr^�}��
O�X�B�O�����!G�2�`��޶[)$��tj�{pD`sMW�zL�]��BB
M����ס���iŅ����L�5�F93d�K��vuɢ�'�Z�QD*Y  [����kT��� � �j�냖&����l��>x=��	«S�&X9B�(\��ɸ�O�*�Fy��ޅ>(�h��ލ.fduo�(��d_�3H䘠*�Tt��G�|bqリ~!P���C��Ղ1	�'j�0��b\��ST)�/�$]��N3�O�L��ȉ�a�`��W6 �c�*M&���!6��O�I��A�#��|�Q(�b�P۱D�W:�B:� 9� �Du0 ���Z�2/�����'PVIZB���9���.ñ2+��;��O�W65ɣaȋ3�80S���vD��Q��S�>��@�²7,���OO�6���_.\�Ⓢ'<x�BՌ�23�Q����BU�=�p bc�/R�� 3��&p@�V�g����B�5�EȂ%l�A��N�g#j5pC
�)[���6ړ@���T���V�bUh�b��9n}�L��HB5�V�S'")�c�Q�H���,�^��(G�N���C�Rq��	իd���!d�ؘR�a���w؟d��+9�J��U�O��̜����Bf��S�Ĩ\�����ύ��zy!�AV*8�B���iN��M{ס��!��O�v��5J��kڬ�`�ix��p���(M�� Y!05��fXF8�����X�\���hS#Ho��I���N#�I���+�>!���D:���?ACE�]>��ۄ�0tF�T9Юm�'��Da5`%� ɨ���9W
���OJ$�T%��e��f^t�|)5�d��JF�`W�F�Z����HOb�%� �U��Yc��^/w�� �u�'0�c�j]�@���"GoJX��*�s�>ɸ���@����`�I;E-��;c�ʠz��a�V5�y�G�l4�d��5�V�YC'XrN�Pч�1D��3�-\�ģ���1O��&L�c�lhy��4^��z��'\��B,�m��Dag.Y�$� �� N��ddAk�s��RR/�Rd��'_�� ��(�6$E(�@���$6�6�)�KN�a!�9/�v@�G|,QKH�f��0�@!ض[�C�I1ub*lb��Ps8u�ы�0����B&D��y'���V�KN�te>@2��0�S��vu��N�$�2e�2Eƀ�Z܅ȓV>t����|�Q6���{� �I�w��y�ϕ""�V��ۅ��i_�GF1On #�&Z��pB�dC�rJT�Z"�'�p!1#��)͎�	�$
|(��
�7&����,؞b��T�	��t�뉍0/phr���$z2-��B�1�N�>�b��e��c�GS"��'cND��.��za횕&ي��ȓ%��h����~�AуSL ���'��PP��
��d�O�>M*�+L�w��,�0I̜�181�'D���*�/Y���L��C��TS�g8��C��\[��'��ӖO�h]b}�L7�|I��f�"k@-D�t/�����C�^�y�׏�y�"��xa�	�y� =�v�݃}p5:ʐI��H��	�J!��(�8��AC�%x�C��!~��Y�jё8�č��1���*&��h<�O|�
���2!���T��<
p@x�'{��\d���dv�4Y�F��&�F�9$HX�x���Q11D�ܛ&��BP������$U�8C�9�	*R��	C��C�?9�G��nK�`A7/e�;C4D��8W,��X�8}:cI�K��Sd�U�u�:0�5�3}�h�j�����
!\AKE!��MVo�#t4!��/lrD�S��E�.\���K#j�زfF=�x�rt�'����"g��	��u*F
Y�O�Fx�	�o�����ҩZl�I:�R�9`7Q�ր��`�/�:B��"r���G�%b��!�ra�<��`�`H�f	�c�%i1,���b�P��eLLj�C�I��\`����<����6`؞*5���h�.�'4�#}�'��1ξlm�:2�8��MH{�<I#&]�4S|\�P�ُj ��H2bSϟpX�G
�a}�)E>2pd�
��P�yB��~��ΰD	�Q�W��y�CY�MaBI��a_:>biQ`NI�ynՒ(����B��5c)�ċw���MS���sӸ1S�Έ���`�֭Q�69`t"O�E#�$V;�D�	��T�idW�������B��1O��J�O��W�L|�������Be�'N���5Xl��B�!R,L��a�
U�pɚU���- C�)� � ��!e�+�)S����T�	%�M+�O�f��	3��	e�̘����6)k��;
nay�g�)!%eBƔ>ѷ��Z�J�Y�%�76��	9g�OѦ�شSc�A�G͌�tF��)��9�U���Ij��ydc�2����$}�Ɖ(`�1��Wɦ�F/g�(�CՕ{V�y@�o��(, ����ػ�4%��p�AB� <u�?i�*%�F����*�@���5{Z�Zb-	j��,Y�B��E�|J�2OQQs��)7
��UjXb���x��ܙg��`��>C��=��A�"S/zTY�®�Xhv-����,�<��,�t!��F�O�}�MR(rPU�J���4v&�aq戔)��Q��_�5����DL
0M�|9 O�L�v�yU'�	>�Xx�̄(-�h5X�$�5�ń���?��LV���`�`1}���ȧAHr �S#T�}�NtYMX%!n��(:�Э�r䛳OE��DHH"z~����	�v���%�ƳS���b��\���'��!��Y����O��p�V�)0Hb�f�1a\������l�c0�B'pe�;f�-�1��+�'ה� `�9v�YQ�!!�~�� #ľp��Јs�'l`��s��$�x]jǂ�v �D�9��d���V�t.����KC���O�&�c�G5�I6=9��Q�ˬ?|L��������� hYh��S��E��C'n��)�@ ��^"���>\����3�PxbN�k����D��s������ɀ�6���������� ���[�L�L�td g~��!�R�y���
��D��U2��`��Cbnl!^�"@(�
�?t�h�U��x2�� ���i�ŀ8T��	׆ʂ�y��L1|�8T9f��cvo����(��><O��;S�S'U��� 뇴z׆<�7"O�0r���!RQ (Y��B�ö��"Ol��v㍎j�F݊�F�W����"O�����Y�<`TG��L] �"Op���̧p�I#!�F>��ma�"Ot��Q)	.7���#؄E�J�;$"O�g�Y�"6�8r�U9 ��h�U"O<�Rn��
������C���(V"Ot)�G�,��&OA�Ɋѐ�"OT�v�ů)Ev�k�o�=�Z)��"O�<�`��BCD�1�[(+S�y��"O�e	����tK��4�RW"O�}�w�;R��2uoӅ3�����"ORI��ʯ�^�p���n�z�@�"Ox��ɑ�]p�]#�,�lǴ3"O�:���V���$+D �H��"O�e;Wb
 �f�q�꒽�����9R� '�)Ń@�֐����B��֯�*{�!��B�2(�!��\g���dM�-B!�ė�'mt�O�%_��z���-�!�<BKl ��GZ*L�����8�!�d�l�Ha���P&rK�M��=T!�$G9Z3����
Q+_&D���� '!�$�0j�	c%�^8t���Ā�!�DC�?�P�PԈ�c�P���  �z�!���=����% �8�8���#�!���;�Ԡ"^��8���֧]�!�đ[�t��E�� etdZ0hΣs!�D�/AF�ܘQ�G��QY&�3:a!���D$dbs�5EwdA� ��^!��O�E�6rqi/ j8l�C��?�!�QuPVa���Ǌlkr,:�)8+�!��T��+@%G�+k�u�w��k�!��Iez��d�]]�e8gHߩ%q!�,qL�@G�Ѱpfֱ9��҃m}!�K8.�� ]�	[4r�<P!�)T5ڄ*AS�(+~5bs�D8*!�D�h_fKs!��J��d�J����exT�H%B����awM�����6!��M� 0H���X��ȓm�,�/?_��aDBǋ�n8���� ����?����*؆zɅ�S�? b��U�	m��pXR��H�UQ�"O�81�U� )���,�n��"O��k���3<��lM+x��c"OДY�,K7z?҉#��ѽ@0�;�"O�бf��f�6d��
��Tp9"�"O�
#iT;B��-ё.\)I ���"OŀFΔ<aTl��'�8��"O���
���H�&j�-,Umz�"O�e���#& z'iN�;^�!2F"O�\��&
#5�0A!
�5��@ F"O���⩋�#�}h"΃=Y�H @ "O���5�C8Sۜ)HW�ގCRhr"Ox@E�![�>�@s�k�T]��"O��H�Lg���A`���	���*$"O��H�톪Z�Tp�!ǝ%�ٺ"O�ECp��Z�j���?=�L��r"O6I��T�|N��ϝ)\�,�5"Oڭ�W�K�f�)��.2U4L���"O�\Cw��)l�������*,��#"O�+Q���_JT���B�*���"O X�@)͎)���3\1�"Ob�4�I�L�� `A��<H@Eؗ"O��h�A5�E97�1f���t"O ��F����, k�GU��4Pg"O��!���v�h"�	�Q 8 ��"O�E�RAW�<(�a�dU,E��"O����Oư���G��w<1�P"O$�� �ˬU h�"��(M��4�#��(A���	��Y����d�(�� ����U&�Y�A�*D�`���5QF@��Y�@�������I��M+䄊��>��A޲�l�:Dȃ����s*�M��
���~����O�١� ��I���5ܸh�"O��b��k�2�R�5�����Ē�0���GEK������U�&=�,�ELU3=2qa@"O4h#a�J'j�t��
���}Z#�)�h�N�p��'�g~�&�6�:�l�(Q"�	0T����y2BИ,T����UՠP�c�R*'
��Q!�'|���Ʉ�ЁA/Y�)(~	C�M$Gb��D���qufS��~�E�]�N��a&V�M�	�b���y∐%*@�Qd@�]�T�+���'�H�b��<�QF�4a�r��s��S�xuty����~�<	&���.K5b�?n�ָ��K^a �c��|�+^M���D�{��\� ���hkc��?Z!��_^����� j�5o!������|A0��,@/$H!�Ǫo�����ݒua|�c3IS�x?!��T	c9�R�ʘ�0{&)X��M8S<!��a2x�
	�HM�ѣ���*2!�D>R����:���E�7.db2�"D�T �͗L��,�vn^�TH|!�&D� i�I��q:�������� D���B������b��ƫ3Z���C�#D�X"R	�V{\�����	���3R� D��x�j˄g�����Ձ�r�0��!D�L뗄Ž*9rd�bc݉eS(�zq�<D��qWhͻ^C�`K#n��*�1�DM>D�8��ޟZ�ZA����(Y��b0�>D���H��HP·��=N�p���&D��F��":"H��CL�ra�P�#D�p!�B��I"(:��B^�E�i D�[EkW�K�j�9R�Ȉr��2so!D�t��G�5�� +�`$w+.��rJ=D��k5�C�
^h
��ĽG���b"=6#ޫ  ��2����Q>�1��T�(;�hI�Fϩ���A�2D�� ����HG'Ӥ�a��j�1z`�˙^�~`�q�ڟd�� ^"���E��;k�p,�;=Ľ��C�0#gj�ȓyT 3'�Em*� �$hZ)�7E�3!p
�c�F��
2r@���|:"�0���zg�2@$�����fVi��iU�!a�A(	 1 e�:t�5�V�-vO�	�'T�xc���Gߡo�8І�I+)`<�e��%�pP��%��w����Z|��*O�,����P^6�@�k��M����J I�j!�;/#�$թE�B����Ĉ�\!�M��F��$�Ιx��A�#��t��dM>A��'�ϑ4<@Y��M��TaN�z�� a�5�w�Zf�-0��PP�̳aF�����ɑ_�t�����0%v�@���4� �@�'���y�n"!�rѸ�$W�pz	͟q��=:bm�Df��&%�Q��� �-�41Y穜��3�'>?q�S;<2H
��>t�4�-���@U��:�ȝJ0��W&B�h�ʽX�m�y[8� �i@�tm.Ě�>>\|��*Y�(Y�H�-^2���CCĄĵ���4�����_�82DT���������Frv���ofޡ�'�Uh|,�o��DL���ԉ ���W�1&~1#�fQ3Pa֬1Gɬ%�(3��ױ l{��Fz��rbh�2!	j-s�P0Ufܤ�OȆ6-�m4HH�p�M-^�i��DN<�axb�6`*X��Z� ~V����'w=���F+�]����M~t�.D 5�)اC'�m�qݑNyz�Z�O�ў�q�"a���Qp�|��#?1bG�+�Jِ�jم)"�Q,���KeÏ�e敨�&�& 6��vO='I (2�c�&i��|*"cNN؟t	`��6ZT��J��ҞKM��r����q����詄�߮%�>h1�7[U��Z���ޟ�J�/c�e �&�sV,�E�� Hp4iCo>�XS���$���#t �ᷤ��:�j	s���>,1�I!R�>ƀ�]jt��}��A5��So���`'�R��	 ;�҅�¥AL��M���;ge�<��x��nf7F��'��\GR�{��U/aq�� �F	u*(��ɋ�yr�vZ�����8��v���y��	n�&�$搊GV�&"�ybA+fF�*5Oźs�dؠ�!L��y���=����)�v搥�����y�$ϳoqh9���23hx��"��y�N'D�`,r��
�����cǄ�yd��R;N�ˢ�[F��уʵ�yBb��O���QLZ�%�P��PJE8�y"FR-KfJ!z��2%M����m���ybH>M����,��nNN����ybm�-@��I�cMW�K����g.��yR���G|d���/�1:Hu�!��y�N�.V14��/Ī#��5�1%�y"&�4@�Vep'm��(x�m�*�yҮ�?/Z�[�m��������y2��5���qA����2�����yBb�b�DUٲ`Վ�h�k"˜��'L�i�3ƄH�O����m��V�㶊���.i�
�'&9�Bۧ<��ÅǄj����a�Ҳ3.�y&�����Y�L����?:Zei��'?L�x#�1D�����9�� ���Ӊ_[@�Ϯ-�R��#Ύ#�<��$��r�M�a�߈gJ�R� ՂWR�z�G����`�<	D�4i���	QC:(�bvL�<��턂s�v�8�AH���'�eܓq���s2'o""~���ƘK���ґ/ �U�̜����\�<Y�)H?0�c)C'{4�Y�+��p��҄��z����(��/L��h�e%�-cDAS��'a'`C�	��41����C3�t�����:���Id�)�Oą��-�ZU�P��/o��8���'?\y�b��8;Ȩ�͓Mh����͂P[�� ��Y=�؅ȓ�T�!���<X�R�aʊR��\�=���(GC�����:�Isr� ̀�A����"��#�t�ȓ^Hq�[> ��p�τ9�d���A�5e��Of�F��O.� ���	
ȥZR♑R<�U��"O����
i��X���N�؃��'�����@�NX�;�h̨W	�hRL�q�2���f D���U+єF��c2U u�>`��f?D�����_l荋�3��12;D���M�r�0|Aǁ���Ƚ6L<D�� ��1��C/4�T�����"OY����ut1)V	γC�h0Z0�$N�B�l8R�sr��!F�	(4�1�7�^���rv������]��%S��0�8pFb��;+�}���> �@!1A�& ?L9�#`�>n8��G~�DJ�
�:�1��\����	�IG�~6���_%���$�]5�d0�!}�ݛ[��u��K q��	��3���6[U��e�Ȗ��)�',�`�UV�0(�I��D���O�i �ӟ����4 ��z��5�S�}�t��mׯ#>`�a���%�9}�AçJv�I�$���W: RE���|l^2 ��v͈# $P�RTᇆ��������E�<�a�<l��³aD���	��e0%IG+e$��G(m�T�	��R�� ��-l"����Ϸ�4Xk`�
�"*`]领���?Y�� Z���B6}Zw'$�IF)��mn��.� " ʙ��K�
Ec���p{
������ N6���1�K],��xCC^�m���[K���Eȉ��)ҧ	6,����f R���	 4�6�'�J�h�+@�dqaF$s�j�p���JܧO��B��Y���0&��̡�L���5��� ��SM|�>��`�N.���(g ��a�'N 8�����ԩZ8VNI�|bV�q�L�����Q@�(g� j`0ez����|��QEL���BGCo0](5ϝ�D����Mڃ_%-aTFR�V���`Dʐ԰!�u�O8���N��Ҹ'�!
k�}x�8�l��L�ÓX	�����~��lcĥ��u��1��=��S��Dr� h�ҡ
,P�|CቸI� =rq��"&*�����P���'MP�	$�Ų�x��!D)�,r�d%�69�X���x�Ҝ�� �#	BXB�ɩ-B�P��́�I�+7�P�3�"��2�i��)x`ɜb��R��D�g�+=��$z"M�%f~tK���ݦB�I�F1��9��$�|�A"eP�ul�O��J ��<�"W���Y��X�
���l�<	UEaaL �Y�G�Љ���i�<�A�C��y˝�c��:�a�S�<qN?Fʘ��	U� 8�MJ)�y���#6� Xʕ:h��O�6�y��ob+�;?���B9 B��ȓ(kHd����_�P�� �=���h�
l�N5��X��Z����4]Z��#�'�h!����`�1��wu�љ�D�=6 x �+(�2��ȓy+�h-il����ӓK6�p��:D� ���u�ԑSLn@�M(��8D�X` �-�xy4.� �xF�6D��PK.hz,�i$Չ%���n5D�L�)�15t����̮?r6���	3D����
Ȫ|��jN�H��Q�3
/D���]آ5�ƃ !8HE�!!D���(�x����b�9�tz��:D��"�)��8���v�*q��`$�$D���g�ڶ�*����sͦУ�� D��+V+�	P�}GJG�%qn`J�I>D��t
��~c}�$�/t,�J#D�<	'J �B\�AȒ&U�-���@"%>D�����IǨ呃'L����v�<D��aS��*���g�)\�ģ�<D�`�0-M���`e�8GRB�8��/D��3'��*Zrq�G��}�8H@�+D�;��"I�	y҉@�OZ~��7/)D�l���/PW P�щ�S|I�d+=#��z�Ń��4ũ!��H��	�hH����$څx�Xe�6j
�@�>��\)�M� �\+,�DI� h�����sӼ�hQ���<$@P$h��v�q��i,H4;��Ä��D��"B��ol	Xp�֥G�|��T�܍�D�f�v�Xr�=O�ل�S�Q�d(7�Q�Q~���u�Q1P �rB�'��� %���kl��?a�(7bĽd����A�<�t�r"D�C�N	�L�O��>i�¨%�`��5�HL�"�XDy2�<G�Ը�=E���M	�陇΃ F���6��.�?ф�)§��ś�T�Z�r��3s�=9Ԧ�+NP�5�I��HO�I��W�jq�� �4V�̐�DǮ~�O*�Dzʟ�� X ��
1�8Ա��
�|1`=r�|��J,|0b9b�O�4�`��L+x�و�J?fֺ`Y,O��v�[�S�OSX�拜/_UD��rC��c*ʅ��`����E���#d	D�h$E"r�נ�^;�=J�`Ta��(�x��sӌ��*�A��	@�F�8�e�#Q�v⟒����7���;�ի.Z�䤰���O���%p��O�>����H�5��rF۾(Q�y��b	��M���סR��'�pE�$g.^b*y@)Թe� U�uĂ�Ms��5��G~R��Ŧ�3�i>mӕԘ6��p j{�>��ɒv�W� ]��S>A�����%y���+gaR�P�b��#wAQ�S�'S���a�� >�a��'��x�O~2��i>�bI��Q��U9o� ��b^�g��}��E��|�i���اh��I�3�BIZ(�$Γe7�`�"؄>, ��}����[5ޔ����2T���eB�/����'�	/�哂?ʱ�tU�!eN%\Rz�yDkK��-b#�'S�P�5��G�� ��ϐ�6�vQ�)O����p'�~��a�j��u��T�g"O�څ�Ҁ@�@�fL�.��8�0"O��c�#[&`�;�
��)3��"O(��&�Z��L	�SJ"���"ObY;�ۄl�6d	W��4m��v"O�HC�h� >%"�XQ-�?M��@��"O��2�@t�<��'�N�m����"O<��7,�#F�,�" ���Z�(�"O:%�g�C�'����1^�K�"O�M2Q��(4�R�ې��D� ��"Oȱ
�jF�5T��%ҫG�H�1�"O�}�B!A ��(�D#� d�ň"O�b@�N0OC�k��d��[�"O��jL&{x&%��l�_��"q"O���!�옲�"q�"�r�"O��Ku,��?�8첶��}Dp��"Or�e�OsTQ;Ũ	�$딕yV"Ol�ad�[�ːhɲ� �S� ��"O�Y�g����C� ��la"O�r��>or�J�FV�Uؖ�0"OH�xqA�(MR�;6f�(�D-c�"O�3���
P�k��ޤ+آE�C"O�����4N��E�@�O ��3"O�!K8-q�#�� ��`"O�Q2VH��f�3��µ(����"O�H;Ui�N�h62{�1��"O�<Ph�O��d`��"r=D�`"O.Tz `�:A����\>9/���"O��HP�)������ZD����"O��3��[�U�ٳ��9Z&���"O�\iG̵?�b�C�K[5/*I�"O��(��w����Lhr�q"O(���%��oPz}�r�)ob�8'"O�p�v
A5>; ���*ثrM�!�5"O��5��& "��22�;6���"O�
��؝P�B�26	�d4bܲ�"O��i���Ȩ�񑡋�x�\%Hd"O�,�� :o���V�����"O�Y�B��{/l��I9K7�4�"Oư�!��!��!ύ'\,}p"O �i!�
n�2�
6-ޙ;w&aP�"O��3��:k7�m�Ì���m�"O�9c4Fלm�0� �ʈ;��"�"OJ`���۲\!z0Y�
P^���R"O��c�@՚Bw��"��U1ݦb�"Oy����2Z8��0F��,$Ӡ�2�"O�t��`
. ��\�%�'t��䲆"O@�p�[<ɭ]��&� �81�c"OΥ�o�4��%)�/�=*�$��"O� 8�`�
^�ؑ{��h� ��"OΌ{!RaC����
�&�@0�'G��NL�.1�t��032�!�
�'nQ)7�!C��1a�/�,@��Q
�'��� ��V����ѣ>Q.�[�'����'�
�08���Ԉ:Β���'~dP��D%Q3
u[Bg�0�P=X�'{���@Z%6t��9���-�f��
�']"����'�4���)-R�k�'p2�Ҡ�Ñ%�^��&J���"�j�'�^�h���2��#m�y�Du��'�0�à-���lы�3x�`}��':�}�B��/fj���ݡ��ɨ�'���y�J�+n��2e�L�c־!�'��S��_8/p�\X�F�.]m��Z�'4��Z3Z3 D�Iဍ�A;=s�'NT�ǃ��vdx�Π0���
�'WJt�V���K�6D_0e	u	_O�<&�P�Y�:��R���4��p�<�D�D%��d -P���KE�:T�D
�U`Tj��2�� E(0D��{fEu��H�ƭ˃Un�%;�b-D�`��'�\����� �z5�4�)D�$��)��p4����4:A`'D����bҊWlq��B�,A|{W�&D����N޼{��1@WI+!�p��W�&D���c�֠b4ܻ"�X�(hZ�I�'5B\Z5�Yow&��n��L�X�'x>eEb]�DD��9��� 1��'p�9B�T�TC��(l�z�'G�<3��26�f�����9C����' 1K��-4\�iN�i<� �'Ҝi�vA�<j�:TxQ$�I�.@�'6����1/��yrĈ��=$H�
�'D0��7�+w%� bw��Jx(�{�'�.@�#ns��ڦA��q�'�$�ʅ�@�`��գОC��'�h �
�*�x|�p(�96e��'8&4q�¶c����ׄ�1&�y�'�t��t%��g�v  �K�._;8��'��p�K�|sh�+akA�#��H:�'��@�$��#J*(�+͘���H
�'�4C��*51
���I#����	�', h�P��n5�� P� }E2�0�'~�R�ܤ���'bЧ{�-[�'��,�!�((��2��ކv]����'T��� 
���KV��&q/���
�'q���KH 5�r;e�F��	�'���5�}|ЈrD�w�p 	�'o�h	�*#f1ya�4;J��'��0Q��>R!Q��4�z���'!�W�!H,��ֆ�#� ��J:D��C�"�6X'�8�&S�,c��9��8D��@!��Q�[�f��@��Y��1D���OR�
]����,T����ѥ1D��Kc<o�hȧ�$����eC+�IU�����'\����O(6���!*D�4ф�94iIz` ]*�SEa-D�L �M M)����FұDU�G(D�LjN��^���!�N��a2D�@*�(�&e�^��o�w�
T�	0D����� �̠Y�	.`+��Z׉ D�(+��~w�ͪ�aY���1�j=D��!'�L�VgHQ薩���a<D�� �� f�5��8w�M������"OeJ`ș�gL���w��	g����"O>�J��Y�&c lc�ę#x�TR�"O:l�hө#^R�0�N��QuH��"O�q*��T�;� q$&DY�A��"Oh@�p(M*���'m%y�vq"OZ@���VC�@"N�Y�J�"OD�T�R� [���P�S��th�"O���EȘ�.�JpI�&H7:���"O6$�wFWnD���ꖊq�$8�a"O��f���hZ�C��bFu��"O���Iŀ*�q�B��,��Ykr"O��k� ��I��`��0
숧"O��FM̿,4�2����4FJ�ȅ"O����8c�����Lްq;� C�"Ox�94F�2�&�Uꑉ��}!�"O6��˹�YC��Q�_���C"OxXJa��.�0�q5�^B�l�"Ovd�7L8JF=�d��O�� �"O�= f��Uf��#�ɫe.P��"O��[�"V|Ct��0	d��"OX���ㇺQ��逥�4#J��"O�X�R�2I���p*-H�7"O���#�]�d�^�R���Kv�6"O��j��Ԗ���!^� >�H�"O��0RFG�~��Q�c$���"O��
`��zD��5B�� v��7"Oӳ�ՙ(�R��Vǀ�&f"��c"O�yk���;�Z8�G�j�l���"O@�p��_=YO�*`��6 �"O�=���Ύt}�冃�:�2��"O�dq�E�;�B�H�4nX�"O�`���qSh�:H�>��Q��"OX�����f``:I�6�\$��"O���P���x� .�!t�-��"O2E:DU�^<�ҏ�|��P7"O�yPG�P��tJ��_i��D��"O(��P"��v��3�Z�7�Q�"O��ƄY7G�N����:-1���"O:u2U�ŒM7ܕ��S/�1� "OzP8#��(Ku.��a/�"��|)�"O�M��Y��+uk���0�"O� bVo !{�x���y���+�"O�h�� �:���CpNG�*qyE"O0����B�|3aM���Xz�"O�M��l�?Dg*-�&+�*��T)t"Od�J���y�l��
D{�F,A"O>�x��ڽ 0� A�H�=�r(y�"O���D����A�w��(ԚJ�"O�u#O$|��(�v&7�]�"O�e�ġ���B 6`@:7�z
`"O����$u)Z��F�F���q!"O��3��>��1�	w�z���"O(|i�&�/jv7��ur�� "O�
�!W8A�64��g��j���"O���3	�
�xJED�
@\M[!"OV �d -b���C��K1~���"O�bC-_l�l��"�jl��"O�mI�L(Y���٤A�!v�țF"O�Q���5|ɴ�W��>���"Ox� 7�?�J����O�5�(��A"OJ�|��{`�"{��0�"O�Yb���`q2D� ���̽2q"O��x2�D��2D��2pK���d"O� �\���݆{S� �RA�S0b��"O`��le�LJ�dܮq�]�R"OB�bV,�/��.��)&`��"OZ$�1�J"��ّd��Rǰ%1�"O�1ۡo��n(ީ�v��%C���["Ot�(	N�H�r��G�f�<99R"Oh�K� 1F���͆=a���["O�D�歓�l�p ���7�dYa"O�;�C�u��$��Y+G��R�"O��R)�9D�4�É:&����G"O�d#n'���ơ��u($�"O��'��?�t�A#�,gf��""O���E.��^e8�s7#�nK@�[�"OI�%��a�h��tcZv�0[�"O`�KF��"�qBpC��6���Y�"O����׻:p��%��/f��"O���/��7�T�1׌M�ylH(�"O>mb���}S�+
|{�"O��r �N�8�p+�~��(F"O��1���xkX��2a��Z�6	�Dd��~�����4����O>�iȔ2'/5�F8UIu�^%���=c�@50ش7��uc�iؤ+�x�h��?Q��*~9�nʯ$��P��u1�A�,}tL�����z@�e��iZ�X���F�b�jǕ�D�c��ZE� \�"h�G�Q��񱠅C��?Q0�i�*ʓ,r�F���߁ I�/�(%�'h��Z$�Ӎ��?i
ϓ|Q�%l��S���$�xA��Q����=��i/�6- ������IiӪ|�2I轨TX�-�����O��)F�Q����E���ծY:Jtz!�@�"FM�ǍZ)]�Xi�eC�/';�4a$��J��E��H��c_
@�?!��	�Fc�!�Z C�≂eA�.UkҔ�'�t84EW�ӱibVQ���]H�d�{e1O�e �i^*�l1f��R�ҵ"��i�>͋��QW��Kg�D�O��$>�$�#(�˕�f���:�ZSB���
ǓJIdD�?�d�@�hˊ�C�&A�y�Mq@ʒL�6�8��Ӧ]�byB��	�6mb�������"fG�Z�ⓔV��3��'�b�t7�����D�p����&&k|,)�����9�-Pz�`a�! J������ċ��L�xs�\H��c� ���25���ۚh0�$�,V{�,p�� }�)�U�&��?���d����1��޹���p��&y�l��뙝vL��?������O��9;W�P����#Gt����RI?���7Y�x�p!L������,SrMx�j�&�m��@)ٴ�\�x��i��]�X�SԺ�p�d��i�HW/M��x�f�X~��OD�`���lU�劃��6;��u��N�8�D��4�O�~����):h��K���g,���}�J��22����Ҵx���(@�X�~���;jޠ1)�e�0�P3��D�G�L@�E��'�a��Q��L9�)�~��h��;2`Y8� �hp<�hf �L��'����剳l>2��*=l$�z��u٪�������ߴ��� #`d:���	]�k�8$�2 �#h��iD���M����4����'�II�`,�H�����',�x��1g
���i��G��r�Zs����O��dE���� ���5�XNP^%£�F�.@�xrOݳm�ʅ��#X"
����1�L='>�)�wv�騂.�/x䅻P*�8
(lCb��O�n�
���;�>��w�E-��)SPA�7��@CC�:���'R��'��A�D.W3D0��Q�%eAvя{�bq��m�{�I�?����-1��!}�V��)�n�Ɓ�g���2q����M�ϓ�M;���]��,[K30�����ڰ#1�\H��:`0X�* ��)	�p�:��G�d��r�"υ&�lZ�MS�{ˮ��g�&-��`���!~��1�g
�Jt��Yw8�Y��.]`
c��ǡЉ&u�x[!aA.:�mۅz�>:��'�&6Mv�̟��D≻6'(�@�&V�S ���.:�̹;�'�`5���K�66љ��G�E����
�æQ%��ܴ�K>i��ߩ��h   ��     �  �  g   �+  s7  mB  *M  �U  �a  �l  Bs  �y  �  F�  ��  ̒  �  P�  ��  ѫ  �  T�  ��  ��  �  \�  �  ��  E�  ��  E�  ��  � � 3  P# �) I+  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*hE}2�S�h���3��˦Ђl�g�K�'[�B�I7����$B��%������I�#��B䉯>�~Pؖ/�mg�9� �<I�B�IA��rFMB���
P�� P,�B�I�E�pC���>"�����LPB䉫]̠�Q��/�a����	{]>B�ɂI��5��@ғ�x���F��B�I�z8�, 2`��Hr��/)\�B��$<a�a�f�B4�L���C��^��C�I��� E�d�pcd��<�C�ɥ\�<l����w52 �d��)��C�	jY�)"��
R��qG�E�0�B�%��1p�K�{�� � ~1Td�ȓ.�X0�s�]�Qk���˛����IZ�'�r�;��	3 r��#G!	�2���'s��3�$S��\u�Ay�N���O�=E��!Z֚���`��2`��EG��y�h�#b<A"���{��	�f�$�y���FEi2D/?��P��Ƅ�y��ܫ���rV��c�p��,���yb�.:�|��CA�,F�]:�b�>�yr��0��p�K5$�����ʊ�y�噐|:��#֖ôs��İ>O��
@+(@�z���BM�;�J.D����V�H�0��$	���p�*D�d(g�BbB$��S.ʤ�*D��v#;g����:��Q�L��hO?�D*al�[�Η!2��uҖD\U1O��=�|�֣�s%�(���&i�CM�O?�'��A��͒�A���q�D�T�>0���=O䴓�FY!lb>����G.X��|�"O& Y��'~�ډzQ�R~ґ��>!�; ������B��N���F�~x�,.O��S�? ��V(�X���IϜo�9`�"OP�[gN�	��䢕�0*���a��I9(�R0:��ԟ��!Ԩ�E����fl��ft�j%"Ob��dB^�I�x�
ˆWZ>����'��<����d�x�P��1�V%ҵE��_H�ن��<��#H�st)�C��ZɆ�n�:�`�ޮ"R
�@� V�h�O.�=���C��!�{c��g�����f_M�<y���"���2�E_�,���I�<�E�M�y.faӪ��Fp"�4/�P�<	��
R�� Z�	4����EJ�<��N҈O�֠����IkY8#�D؞�=��a4��A���̕;#f���K�<5*48A�th�N�6P��P�n���hO� �=��J��`��b�8E�i�� ?�����na��"�F�_1�"���s���2E7?^��痩T-�ܫ$"D�@g�T�d7�1$%�"{u��96��<�/T�z�h(�����yJ�@g�q�<�&L�����d
�g�HpC��j�<Isd
 j��1q�ډpzi[��hX��Fy"�Yj�:����֨�Lؚ�yb�p@w�u:>q1�K�4o2H�����dt��է���D�Nڰ��6m������6�!�/=z� z��0����P�P�|82˓�yR�	xyR+��k�v<IG��V��3���0?q�'��];��T�����S%i��8E/J?�g�'h�8���@;{(2�� &iXP	�'\������Z�/K�
�@j�}r�'�T��,L-(�b ��yv�̑�����<X� x�^#IP�9%āo��(�
�'QT�c��4[����g:�؁��hO���%jԸ+��a|\�aڄ"O�*1I۟u�$����+\D @��>y������j5:R���=�4�Q�ay"��Q9�M� �na��A�N�5h(XC�H���ў"~�	!wu2�j��ǙV�t�jG����OF}&���R�-a����$�(�B<]`C䉲H1r���OG*?F\����ڴ/3N��W~��'s29��,ڂti��R����x�^���j��*�� QW��GT� �C^�<-�OP����w\�=������I��؇+�DFy�;���Q ��N��,��(<��Q�w�!D��9��RK?P�8��9�^�У��O`"=�§��k �(�x�'ϙA��e(M��L��!D�dSf �X'�i�L�~⌼���>D� ���̤8"�t�w�H> �|$���<|O��&��{%��*#�\Aj�#o~3@;D�@�a#n~,��B���i1r� V�>����S�<Z��"TᒢO�(��k^�߬�\�鉆z�\;������u`���Z6���$ʇVH�x�BL�E�U!Ђ�t:a~��'U66M +��e�$ꕄ-A%�0"�${/!�,2{<=�&느95�%�� �< Lax�g%ғ:*���ǳYyl���ݾ{+��ȓi�l`��!�Ӣ��Vg�0�����d�tack�6Rߢyp��[;Q!�i�ȓ3���(�'\�z��S�+�5����ȓu���{r+$�Jt��[�x�|��ȓ4p]S�fUVN��$�V94�l8��Y�*P	�%@ڤ���a@�2NՆȓ?��t�(H��e�筃9x-H���lsg��u0�(��À<,L(�ȓ�6\S��N�P]H3���Qim��S�? ^ac��*8Q���,?RAX��	c�����(����@�,Y�d,����S�~�j��\��hR�]�d��`�,@j���P">��p<����(%a |;���#rJ�]��m]�<��S"fp���]�e�L����;t:1��u�� b@��A6RQK�A��2M�u�'	�#=E�dO���| �C�4|JKc,˲���0�O�#�[���|�ą_8]l\�Q�#|O�����>��`"DO�`��"O�I��%�( n���+�$@p�#sV�p�Q+;ʓ��'��4JR	
�Y�]���,sn��
����$Ai8�����ʎ!���cP/� �1On�=�|��[J�z�۲h�4�b!Hs��By�~I<!DH׻dn��P'_�	�j�	4���d>�O`M�Aaԇn��A&�-5T�	3VM}�`H>��)�,O�	9��t�ْQ�вŠ�y�f�x5�'����=i4cӮ
��)q������~|�\���L�
E(Ƚ0�|�g)��f��� U�'�[�jq�U��_�P��,�vq����䓛�<��<T�tLZ�z��tzl[�'�qOZ�|�E� -iA��1�םK��xh2�PH<��KӬ8�>H@�¹qx��m�W�'�ў�'
Br𱕉=&������
	䊠����i�Ƌ�(1��:��M	@(�x�=iK��G��N	�b��o�9J�p0Q��yb�ǌn'H]#�Q�;_&�C�_��?�pB@L�����	�Q�ą'�>�����KE���#3D�p���՗|�Z a*!ndy�H7��x����N�����Z(0�>�D��,�y��&�S�O:��䢚�tl̉���>&�,	cŪ+D�X �ˡGC\�;�J���:�.}"�'8�\��LO:~�豸wf\�gQ8�
���d�0y�J��A�̣~���)�E[*FKqO���ĉ� f�c����t� �%M�;Fa{���,�U)�ӇK��K�$�",!�DV�X]sp��0KC�����t*�'������)��@W��̓!-��#E!�$��� {a�	�H,5�勒 !�ĕ�]�Ԡ"'L4M۞hے�  41!�d��<�E�3�Z�s�2�Q'S�j!�d	�Jk�My'&�c�Ʉ��!��\�o)��Ƥ���f�@����!�ā�5H����O�$��p��4'�!�d�!����Ӡ-nx��PbL)�!��3���u�\�OR�u)4�$�!�J;P`��hN D4,h����)�!�5TeB��-�Ac%�D��"O�����ͼF 4Dh���.81w"O
MQ���&u8vH2�C%8+�d�V"O����Cax�p8��Y7	 "O��(�l�h���H�$ݯz9Z�J"O�H�G#H<y�[�D����"O4��uB��B�"u""R�2! B"O0���-�-K��Ё�@֬�N�*U"O��%k�q��@�ĺ��xJ�"OD�h�B�OX���`��IXX4C"O��р+!>@°��%�D��"O.���%L4�U��,���f"O�4��b��/�z�kp��L���Q�"O��k�#W${|�؁����+�`5�4"Oڱ;��g)	�eD;o���摡�y"�N���C�mɄ���յ�y��~rᖈ�]x8� �C��y�ޣY=�������&���ͅ�y
� ��*�!��<�ʍ���ߊn[$z�"O����m�$��8Z։_�c��A#"OX}��@
�^@���)�t�}JG"O � �-�a:Eu�	�D��u��"OH���M
|w �:��Hn��h��'"�'z��'��'��'}��'r���m�,�{Ԅ��mv��!�'��'R�'��'�b�'t��'��@+-�<_���R�+T4v\�DA��'~B�'8b�'bR�'�"�'br�'�&aX��N��0�����0x�'��'�R�'���'�b�'�r�'��� !��S&�Еf��*2�����'�'��'!"�'���'[��'����ղ��t��I-{;&x��'��'��'�'5��'v��'{�(���o ����<�@����']B�'�B�'ZB�'��'n��'��pH�d�0�+p�B*)j��5�'t�'���'���'r�'&R�'�v���C?%ʊ%�'A�Q���`�'��'r�'B�'�����6-�O8m����<	 v� �&N�P3(8�$g�O����O0�d�O(�$�O��d�O���O�L�� Y9�Ƙ���0�{B��O��$�O��$�O"�d�O����O6���O�d��&�Z@1�� j�l�An�O��O��d�Oh���Ov�d�Ox�$�O-��䉂{�5�C�g�p�v��O`��O"���O���O���ZΦ��Iџ�k��ѧ!& *qm�VX)�E(���O��S�g~��h� .@9p��k�CN_[�H��c���/�M#���yB/p�"����WҬ}ipb��<N�*J��	�"$4ٕ*?y'�A7WW|��%��m̻U~���QY���R,ʨ˘'XB\��E�����u��БcU�n��1�[/�,6�>'81O��?�����{%�bzP��� ��bML�GP�F�a��B}��Ԡ�5(i��9�'�ኄ�ۍZ8�RG��<^� ���'B�]�X#I�R���i>�I32|����&��2��p��)�e&�I\yҙ|"dl�$�I�3q��.6�r��� �?�ʀJ����I}��u�X�nZ�<!�O"��� %bV� 8�H���ඝ��p萆�T� Ѩ8擘���0��䟤;�o�}x|����&4�d��Izy�_���)��<���y�0���/����Ҋ��<	��i�����O��lp��|��� 2��2'Jח��@�B��<6�i&F7�O0f�I�.>���s�>�`�	Q'@�5)S�rL��f��>����^���D]��$?� b&�G�h���E�^i�q�4E9?I��i	zY��y��	V�vX�X`�H�1R!R$�_����'��6-M⦩��ħ����+�Z�����[Z�����D¥��5W�'��$x��0(�^��`�HM���g~ҫڋF�@T����e�l�Ȇ�K��Z���'��'�n6m��@���p�����G��+����¬J$$��$Aߦ��?��<Y��i� 7��O�܃s�4x�\rBȖ�[��q��=aCI�W;O�}�%�7�z����W����O��4�V�~�y�%  ,3p9p/�u�T����n���Cy�Z�"~��H�-��i�-l��d�֮�U�u֛�����㦭��zyB"*:�pz��ݜ:	<�����/1�D�>I��i�|6�O�)1#���9k���O�A��\�N���wt��c�╠[
>]�Ԯ�Qw��=�'����O�T����p](d:��κP�Zy20O��O<�n��jhb���O@��p��:]���R�Qz~��>�D�i�6�a�t'>���5Go^�㣥"����C[�qs���p��0G:?���4.*��A�4��6�Nl�Ӣ�4��8��)5z]���/���g�$�AH���mD��`gNɣKL�i��'�B�g���$��O\nZm`l���>x~�
A��b��<@�4a��Ã�ey@P�']�OB�R��9v�n/��4J`i*f�UXS�)�g�w�H!\$ċ&,WVO�yC'Ia��1]�v�
���g�<b�<Q�6��)�Q�5&�UZ@��0��H��KދT�����M��B�K("��8����(Z�(KRM� _Ԛ� #�Ѹs�
�:킷.�x,[
:nB=[�(�I�V��O�
K�����ֶo�Zaz�/K>B��@�P�>�f���G��|jTBcEX.�4�
���FP�X+�$@(.j�u ��U�*�< ED��T:��G��9ǜ�k �6��fB_%�P	p&E�~�v�'���'E�T  ���OH�@+֯��a0�����X��K�YQ��x���'$"���O��#��� �ꨣ��Y�"�L�s�*���	ܟ<����D�'t������Lꄥ�$���q�(`�%>*E:S�D �nAԸ%>��	͟��ɰ�4�b��^�0�AH� �ڴ�?���(�?	�"S��͟�$�0n�$.����f�ʮ2ŀ1�C��>���ݮi��c>?Y���?��?�� u^m�hT�*pm����4 {*�:�J�5��d�O����O|�O����O0ͱ��X�' h�[U���V��4k�f*9Xph�����������I�0�	�h���Im��R-�
o�|EQF�\��q��4�?I��?iJ>A���?�5�ڲ1���o�<"N68�u.�nQr= �"�TYj��?Y���?����?ٵ���?i���?Q���Gf�A1�b������V"=���'8�'{��'Π��H��ē-d!�˕�P�ƭZ��88/��lϟ�����8��|����럜�	㟈��#�rP�;��41P�#fy�:H<a���?��M&~���<�π Zeys ��a�2�����$�$|[��in�I!VI<��4,������ ����	#�1��!!���rR�=q�&�'c�.��O�����i��L��U���"�Ļ��is�x�@�'��'�r�O��IџX���O�֝��g�0"Z�#|^	*�4�V諍��I�O��J�.a~ $��Oxu&�����Οh�	�`&�8�'>��'���O���� @�"�FEpG��� ���Ǉo/��O��d�O��ӃG�V���Qr�P�s��x��Un��d� �Iy��'���'ɧ5F���v	N����3bd��ޒ���ҟA���O��$�O��İ<��NZZm�m�QX�9r蓴2��,�-OL�d�O���3�D�O�����n��#��=*��#�� b��M��O���?q���?�+O8|	��?��b��nA6��r� Ő bn�\���O��d<���O��ߊ]FL�	7SH� ���=����L҃s����?���?�/O���|��+��x�G��wD�̃w�>�0����iu�|�'t�ό�N�qO�a�k��R�C�>`�$��ֳi��'c�ɽp*�OgR�'c�W3h �vn� 	�ĥ�G\�u�nO���O�)�g&�O�O�Ӡ"����ku��ɺF��2d��6�<��⊶�?����?�����.Ok�?R�r�J!��!�"���V�'�k�6##�O��l0w,0R1z��Ŏ�h��1���i�60i��'�R�'�2�O��	��T���c��A+sJ^�1���3��TA�v�Kڴ!�|T
���S�O�®�[�81�	&t���Xw�W6X�6��O0�D�O&�Z����O�D�O����� c�b�O����ᖝx��b�@��.�e�I�����x��(%&�T�I�]�e�l�����M���3a�����x�O&r�'��I%&KI
��z!�U�����ڴ����O
��?�-���b��ިQe2��q��� jE�#z�'��'&"Z�|�IS��)+��Q�@N�&�L��d�Ҧ���{yr�'��Y���ɾa{�e�'h[��ʅ>�4����,TL�m�˟d��V��?�*O8�zF�ivl�Uj��}P����N�6LB��I<����D�Oa��m�|������X8O�ॳU$��vn�馲i��O����<I��DX�ɅD}t�vۭE�2PI���(|7-�O�˓�?��a!����Or���k�\r���o5Z����Y�4��M<�����H#Y9�֝�A��\B��ݕBL��s�'�/R���?�D�Ð�?i��?!��R*O����%R��/	 �A�#X>m�6�'K�W/׈�0�y��b�4���Wlؒ��l���B
�M3�L���?����?���(O��4��t�0��z��(�eT�Z���4-��b� �c�S�O� ��W�S��%���6���Z����'���'z���aQ���I�V�㑩��1!*u�G
�{�D��yRN={��@���Ox��<jb*�Q6���ig>���C9��l��h�rC�=���|����?�/O(�A���%���8���'���ŬRŦ���\r�h�IVyb�'4��'X�	�}^����|�䀑�LK����A�k�;�ē�?���?i*O ��O��`�HN�0��VD�4$ �y��І~����+��O>��<�d�� 7�Ɇ7� I3�#<͜��0mŁ:��Iɟ��IğЕ'$��'� �I��'#`��²Ov@,���U
a(��0d��>���?����d����&>m� c�Uʴ��%�J�NѶ��k��M����?�*O����O\@H�g�OX�O�\�W"C�n�4A�D+Ų��4�?A������� �'>!���?ט�,)؍�cꙡ_, �95	�,m&6�<i��?�S	���?i,� ���k,���(�vf\�v�l��H��op��R���T���M{W?q�I�?�p�O�a�e,L�J,� �FT�]rTD��i�B�'� ��D�']��'�?��'��i��x�q@�=��`�ǢM�9K�<(�4a�ƽ��?��?�����?}�'���ܤ
g��!(��8��cE�M���+2��<E�4�'�j�Ѐ
�a)Aq�˺?�*|h�h~����O�dY�}@��'��⟈�I<l� ��6�έ!$y�B��y�&�{ߴ�?����?��L�b���m�t�'����hFb�� 5���ّ�$4��v�'b�z�V�ȱ��F�@3�lѯ)�Iv��ȂH��m���$�;D�2ݻᛟ�Iٟ<��ty���& Q�rm��x� ���*D��F�'��Iܟ��'���'pR(�ְe�@����M"4��u���'b�'���'��P�\9W�\���d�R�	X쩡v��|�����\�7-�<a�����O����O��>O�L�&���J�rԩw�,;?> x���9�����Ix�'_�MЅ)�~�������`���
$j�I�|�Ra�i��P�H��ʟ@�	�^�l�Id�d��O7p�e朰[� ��%!A(*��F�'�b[�d��������Op����XFH˾���Y�L���T,�~}r�'�R�'��@ϟ��`�f���P?� ��I�P�=��aB��1�'�|��2�y����O��$�6=קu��G$
�h#�e!D2����k�?�M���?� �t~"Y��}2���Q4`�")�?��J�,�ۦ������M3��?����U���'��c$���,c��ǭL�,B�l��Mx�6O����<	���'N�� ��'�ʯ�p�0)\9Byj�i��'bґI5�6��O����O���O�Q�e�d�!'lN(Qu���W�W=)���'��	�B0��)����?��e�h�"5(_"g����EK�Q��"�i���ǌ9Bn7M�Oh���Ov�D�m���O��Ұ�M�cJRp��j��T熁��i��
:�yZ���	ȟ\�	�t��; _�UX�G�[q&�:f��o�p����\;�M����?����?�R?��'��+ "A����j���%y���'���'h��'e��'�RJ��1�7�s20�S3� �D�:5��͖�#br%l���8�	����	�D�'�R������_3�P�E�.�x��dA��*o,��?���?q���?ag�K5?�v�'e�W(���l�&D�9"!�1;k6�O���O�˓�?#��|J��~ L�>
娶�M�	��C���M���?a���?�a��F���'$��'��T�C�i�xZa�O��D���D�z�6�O�ʓ�?��|j����4���Jy�8
�n�6M̄ D���M���?uo�z��v�'q��'6���O�rH�27�`� ���U���c�ڇ=<��?YV�Ԑ�?q����4���O�F��!Z;� `�BZ��شT�(t�Q�i&��'���O��t�'���'\~Q2H�<�B�{gd�:9l<�{�b���
a��O����<�'��'�?I�j�	?�R���CV�>�:8v�D�f��'rR�'S#U#}�`���O��D�OJ����|�C�, ��@l� W�]�Q�iu��'��ʋ�yʟL�$�O���;�`eS�ʜ(z/�"�Ǹq�0o���!AD	�M���?����?�AX?��H���6cA��6�1@�׶4J�n�՟�@��y�Ԗ'���'�B�'�Rc̍Z�J]Y�OP*0���B��PvEÅ�t�����O����O��O��Iٟ4Q`@Q4h��h����%V�ĚP��:R���ןd�	��	�|�OE� �tӠA#�i�0m}bȅ��")��	P������	Ο8�I��T��`y��'Z�ʙO��EZoS�!Rh����#��7M�OH�D�O���O��$�,>��}o� �ɾM�T�
F�$Dڡ��`�S�̐0ܴ�?a���?�)O���� 9��I&}"�����P�I�u�n���L�M����?q(O�!:���N��ޟ����eZM�����v�`�{���<�ֵ;J<����?Af�0�?!K>�Oi�L�%&���3� K"0Q�-K�4��$�vU��m�����O�IX~"&�3��0���:}�\�yUd<�M����?q��ڰ�?�O>�~ ���cvb��bG��j���TM�����!bO��M���?q�����x��'�t�Z&��? U���D�\b��|�`|a�5Ot�O��?!�	1~��U	� L�up��� �Ԑ#'.�A޴�?���?9�D�&Nˉ'�b�'����}?&`c��V>אpiФ�� ����|f	8@��&���O��D�Y#*���<U��LL`��mm�ş@��d ����?�����3�͗�$�4�� �Ŧ���H��|}��S��y�W���������^y���[����k��|�%��/s��e�e/.�	럜�'�2�'�r���[f��{��V� 	���*���ʜ']�Iß��	џp�'�d9 �h>��iޟM�d����
>BH����>����?�J>���?��O���?�4oS�:U+P���>�(�$߳K*�	��h�I�X�'�2śU�#�	D�U#>����L�n�R�se�� ���l�ߟ�%����ߟ�
~��O� 	���q,)�5	��zu�ᚦ�i>��'��{���cL|������
y���&k�%ys���"F\�7P�'��' ��x�'�ɧ�)לgo��2�CD�1�Q��W(��\�D9�#��M�R?�I�?�a�O8�!�ܶ] �ղ'!
>z,��;u�i���'H���d���T�V��J��Y��,���>��iD�X�7�O���O����c�Iʟ�P��x\`h�*��_�@�pej��M�Dd^���������f� 䒤	�#I��R�B�M�\��Ob���O|����|����|��Q?��Q)Oo� �
����,q����)&���@Z!�ħ�?Y��?ITjI
|Fٓ��)/��`�`)��ћ��'��i[eJ2�$�O���6���Z���*`n�3�HW\a �@"U����E�Q�Iϟ4�����'.Tr��7����)�'�8�U�qrvO���OĒO���O�J�ÎUd�S��\3f|��Eb�=�>�D�<���?������,)���'X@R���[���` ��o�kP�h�	��$�l�I�B��ٟ�`1F$��`	:BPۀ\�����O��$�OPʓC��p��ɀ^�"����+'��ű$B%�7M<ړ�?�u+ߎ�?�J��x�� @�6�eeSQ� �+��o�����O�ʓu(�	t����'��\c��Zq���@5&|��� ��O.�$��B���O�>!�#-���Щ�Я��.>��ᓥ�>��}Q~A)��?�.O<��<�;Y"t	`Z�\�"�C0�39t�mğD�	6z�����(<�)��S��I���
��e�Z�}U�6-۵v po��\��՟������?a�.U 6�� �B�Qr8(CS"�vs��D�6�O>E��,�X�2�ʠ\'�ݙr�_�Y�0e�ݴ�?���?i�D�P��'v��'����-�.u�S'��a�$�;Q�*
ñO
X$���O8���O��㥃�
1�ڒ`I����;7�M¦�������H<)���?M>�1[�z��A�$��L��$��t�q�'p�i0�y"�'i��'��'ir� H���	ɜ_�����oՒ��@j�gH)�?���?q��?�J>y���?9�H�� �>,��Cѿ
��Rb\6���<Y��?���?��d
0q� ��I�⓽M��軇瀧z��c%�iV��'�R�|��'���ISzh۴8(d�Q��;���1ž<J��'Y2�'qR_��@�̆��'Yl���'a����Éc℉��i=��'>�O�4�5�)��uuȸ�b�>�xl���dF���'n��'B��a��Sޟ��	�?�ӏ���x����O*�������ē�?���$mI"��p�S��k�!.���p)����`���#�M�-O(���&�ۦQ#�����2��'��I��	-8�1�����W0>P!ڴ�?��A�d�Ex����� -,ѩtO��i���M��
�&[��V�'���'"��2��O���p��:1F�pF��	|��%�ަ�--�S�O��M]2A���С���j8����G[�6-�OV���Ob�R4hV[�i>��	l?A�a��]�8	ssR���a�I���Igy�)#4d���<Y�D�,p�ꡉ�K�I�y�bX4Ɗ8�!�)��	��K��@AV�J��"eH��dN���I��fӸiF�I2����zbH@d�T�w`�(<5 j�I 9T\�pd�>
[*qC��@UB���5/�s�N.tF��S)	�8"����"QL4���z@�"�%���fi�������6���B�Jٜ��)�j�Z�Z1Q��3�X�x���B�b���'�.��A�X��T��^�ly�� a�'��F]�'M��'��ɒ�>
�{3"R�HMI�n�4����_���`���:l�A[��'H��R3@�}��� �z���R�*���A�/tQ�?Z����n:��'X�	�~��y��T#:$6�1�o�
b����I��`��Z�D�I�	ބBg�C���Mˣ��(�1��A��V,Xe��<(O���Cc�Ѧ��I���O��1G�'�RI��&;0p������'|�)��l8�])�RA���O�SG�DƆ*Q���EN�:.���N���_���K�mD&�(�M�;0�8�?�����/�,U�F��\�u1i"}r���?ip�i�l7��O6�?y�6�� !���$�	wR�z�+�Iן`��	 N=�m	c�R�:e�$	C���G������g�'��aK�.��邱��-~���k��"�'mr��/��=	 �'��'�Bkh݉ �A�?4?=x&����woC>�iJ0�\T���Q� :M����|&�R�)�d�44�A	?:@3�^;V�r8HUkΨ aAB�4����Ç��I�to4��w{|��s̜*�ڈz��U��u���'��	�:�
�4���=��Nr��/�uZGC��d�X�ȓ4n�(@�	�(��� �7U<�Γ�?�&�i>i�	Lyb�ԣN��灺o�JZ�_�K�@4Y��O`��'���'�]ܟ����|�#� 	&�p2V���|�+�#�_���$�<PE��i���'��<iq��7xؔC�!�>�yJ�j����dKM+'/ �a��Cd�Z-��	�Zj�4�V�,�&�R��
=ZT@���O
��$ړ��'��%���E#$�l�@�N0S
�'�jU;gȆ@��1�R�=
�bU�y�Ce�����<I�ȋ+��'�҄�7C\���q]ऒPdR42�'��`x�'H"7���r��V?ORa0���vl����E�#	T����'�
`��ߐ!>�'䘥�ڽK���qG�  r���i�.e�	ȟX�I����t�ùHG�h�_�v;���%�Hy��'��O>I�v���*+��:�����k;��H�4��� 1e�<^6MU&Sx2����ӥZT�hlz>��	R��iW�X&�FU�����-
�\�Qf1-~B�'m�l3�B�	ڑ��a�a�*�T>��O��i�c��,6H��n] "��3J��+r��78��怒'�mF��I_��~�@F/�0~�&�E��-��=`�����OP�}���W#�l��DX�f����T#�-N��)��po����N��x���P)EB1��I��HO���VM8h�h��-�?6��� tG̦��������<���$�����I�x�i�)ZQ�!s�4�/�ax"X+co�&u d���?�ta��-Y��L>A�	���!Bf�P�h�XUN'P�@�τ�6��/��@��L>	�bF<6�rp�d�]���� ���?9�Op)Y���?I��?٧N��$Tl=KÀ�N��@��H���x��\�|�4�;����8�V��w������N���ɷ<i��]�����d�����.RD ��jF-�?����?��Y
�n�O�$n>QxGep�|3u%�?d ����!�3��|�D.C(y"��'|j�E@���Iq�� ҕ�L�˒�(�I�C+�*y(a�"�����^�T�E���ޝ%�1O�I-k�����@=S�p�e$ԍ2�����?����2��(`heQL��VM:5+A�	P>��d>�ĝFIܹ��M�86D�"���G�1O�mZ̟��'zY�S��~
�����J %G�RD�v�U�0;\�+���?QD��?a�����/��rR��сI� ��	]D�? "0���3D�B���T	��̀3�'�֥r�aFekdl���$c`�T��7�Ex��_�s.�D�@�r8�X���O�lڬ�����d �Ǥ��P�����1J&1O���+<O��L	�6�Xո�B�uf\@: O&�l2R>@T�W��q����Rl.��byr�)$h��?1,�>T�!�O6!��
	"��<�֫�K�I(���Op��'X�T��7/�BMƥ�,J����O������
�-N�pժ`Ŕ!#��'�.)ӖG��t Vx
.f@jeB���0hfD�O��qH�g�%g�&��d�U�HM�xZN�P@���O�m�H� �I��B�(��3,�&�6*�
���C��+�YR��H��)�b&E-���m�':T��G
��,��fۘ~�2�� �`�N�d�O��D��@s<��E/�O���O��DG���"H�,%%b� +��ܺ��i!H�Dx�k��}�� *e�Z1��',�����y��y�RjE8DX�!�%@ X޼��$�증�a#�q��'�DY�$�M�Q���S2(�/ ���h��'��'���������d�O�$�`�� Ѽ��.۪p�B�z�G*4��F��F���g��]�D�:?����. !�d�<G�݂?����J�~�8�cZ�Z�七���?A���?)��=�.�ON��y>]���!UFhh��׻' ��K��,P��STEȜx�uR�����<�����yd,�S� ����|��b��hAXܻ��E�ab�Y3)�cB�Y���$KD�DFxR�Ȗ@���ڦ��/�`2gǯJ,!��r�6�#�d�Oh��3���V~T�f���.B$�G��`?lB�I�R%�9c�� %>�S����Mc����4�?�,O��dcŦA�I����3��E�X$�26n��]���Ɵp�I1.
P��֟�ͧf����sL�X�ɰ5�G�����%)����\�-���Ӏ��n5�a�G,ʓ> �jP�Tpڳ��]5:q�EA� ��۵BܖYU� ��+i��g��2az�<	3�����Ty҇אT�k�i�?mw`ay3�O�y��'�B���2�3��ɟS���PgM?)��C�ɲ�M[�д	~ � ��hPPA��r�	Hy��Y.6�Op�d�|�J-�?���w���dEN���'�ڧ�?y��9�|ط�G�.�#�BM��y*���'3Z�X�`hR�3�����#��a2T�O�y��郑+�Vl�ARp�>�3b�,7���#��(a$~���h1}fB��?�!�i:�6M�OV�?591
��+Al��2��3���k�o0��џl�牊A�|�l�0ƶ�p��J@(��\c�'_>�#�h
\����UI\�`~�ʧ�Ck?����?�f��=;��%8��?����?���֡ñ�Pu�f�ʛf�[���#[ޡ�d��ye���C��c>�O�‭S,N��!hP	0X��\7��A{���۟,y�玾(qq��'�� �@/�VI.i�O��fj���'<�I���4���d(�ɭytH��&ܶ1��P�u�B>s�B�Ɏ15�Չ��	<+�\;�Fg;6�ɑ��{�O�ʓ)nR`�B��lh�@���/zG��˶��S+<����?1���?Y����$�OL�c���C�ҳ2��,1��Yn�q��ih�KU��
J � |��"��K�ʐ$rT�K�;�,]Y��}���qE v�RԸAY��0<a��h7�����(G�NH�v�#J���Iܟ�&� ��]��<�**y��a�G
�<p)|��g�e�<�%��%?nԪc�P$V��d�C�	a̓)n���'��ɱo��my��Z���<�D4�& �����qW��nL�D�Oz�:2��O ��h>y�G���D$pfM" ���C
�L�ȩ�剽\�4�$���;��̱�IQS�'�� ���z&hŢq�90?>����\��|����!(r9����\K��I�._"��ʦyѨO	�����<��ʪUd4I@��Ox��Lp0�)cᇲiy���ɜ^�!���I*$`���L�nH�D�+w�r���''�\� �x�&���O�'0�6h���\L���-�:�� p#�S���?�f9C��1�C�8Z-�A�
���)�|��˜ c���#nK�qt86�R�$�#G
�p��}>�j炧ym	�4��yO�������Pp����,:^�'j�����?Q��?���
�L�{1J�:�X��f��'��'<\X�#ׇ]�X��ѭ�8V�pA��bF��P(W'�}�R���	=��tg�M+��?��X�` �6)	�?���?	������+LJ:���E�N����m��Hn��'"M�h��61sx��p�|�ň0(�\I�K0[���Q� ;�8�YF�C7Ô����㮑[�'F���	^DbQ�Ǿ:-(a�R�}�
����i-��'!�Xje�����',��'���'��IP��)8݌$�w�R�d��D˲O¬@W��H�v�	��؎)��X晟c��d�Y}bQ���a�V?�(�ӄ��.e7���⌓�4Mqc�'��'0���~R���4⅒Y�l� �H�!��P�$��H�����9��a��'�JM� ��F��"i�@���!�bE*'�A(F@���P)��5�<b��'��T ]�\IP��.��jq쌦�?Q���?�������OJ�8Sw�ϤH��'�����*2D�@y"�Uڮ�B ��Z���@�3����$�<�)�;6Ǜ��'l��4[d��cG�i���Hwn��GaB�'��M�v�'�0�|��ф� D�%HD so�7��%x�"��פ,��Pb�X:iv�x"��e���� �A�W�B} �i���G	&T�H!׉_�ZP��"
�'�P�I՟`���,S�:�.�J�e޿aQV(1�e���	�\�?E��$ڲ|� �&��4Ik���t�H?�xB�e�\��$d�%���{��G�S��� T1O�ʓ5���b�i�B�'o哠(�0��I�<�՚��F�.��h�� �&;.��I���r��#-��� '~Ӳ�㚖��i�|�d�]�9�Y��dN���9�d�X`��FG�-3�̬t�,=�#A�#\H�����{:���SL(_Рs�e���P�d��O��lΟD�O���O�x ��h�pQ��l\� ��y"�'�yBg5C&��� k	�o�p�slQ�0<�6�i^�6m5��K`��R,��u+���������Bx��{t���g��S2얾+;� ��&,D�Z1�O�6��Z��3��,A�>D��D +	�F�Q֊�kp����7D�����VX�����e�z��w�"D�p�f�X�^�l)RFb��_L����$D������r��&�^� ����.D���g̀�|�LbG��D|�|b�n1D��b�%XzP�#A�,j��2D����@͐��#w�޵.���q(/D��CGP+b������;>���+D�D*2K�.(2��M���0k-D�X0/�	6FY���YՔ,kr�,D�$��oT���BO7Z�D���?D��Z�"�39~�84�`����;D�4�tNۚ;�Ȃ�! fp��Ī6D�����.O6P I𫇠j!p�8cE4D� 2mۡJ�(	��eK��64[R�%D��@b��04�XJ��"`GK8D�X'X�I�RyHGY:fF"��N7D��5��X��p�fļ.CPzq*D� !����;�� �.��eRD+D� 'C��|�IRd�KZ�ƙj�#)D�x�PD@��r�p�>	ؤ�Z��#D�8c(��(�`T�� ��L����� D��0�{�^�)WK�r?�(��:D��[S�L-2�門�q|v�1��5D��� �V�2�Rl9��'D�̑�ΦT���I��L�ziz	��3��Ao�8���'��z�@(��i1������h�R)�C�z6��	3]�Bp2�a#��#5��"]������O�p��.�a��xr���ڤ���P���(�w�@�"r	h���'%��h�%C�Ӡ����-âՋ�O�@��O	 ۆD����\��e����O'Ή"AL���|S#��Z��J�'�ryH��<�((:V�e{�x��%��$�~9�G����?Y��'��O�P0�O�p��S�-�l5�w%�+LJ
�'���fg&Z��\���1lϤ�r����b��a���ݕ�h��D�W�,م�-1�����Q�hT���ϭG����D`�D�f玏�n<�Ȇ�$�ȁ#�C�{�n����q�sԉ�PxBiR��n��WM-ZMx��-�����64��:3K�W8(L��)��X����Eͨ�f���,<S�����?�Մ��0?!U,-.y0���p%|��q���Ж�'S=�i�ɸY7�1�O���O�^��٢d�+H"51�OM�I��n1��ۦl.\_A*��R	S�|�H��R�M&���m�B�.�0���~2	�<)e�/R��XHR��?�@���U)(X��XI�A�' O^�HE�КeE�I(�Z�x�~!h� fGmY�/Q��re�	|r̠<�V�ڵm�l���)��y��$_\��$iۂ#】��-�!��DE�� !G�K�vr����WJ?�I� �������t�,U8&���:M�	�d^=@�H����m�,�`%��T:�ͳj�w�j��.ނI֒IJ���O�x��v>�O�^�� ��"�� �Ca ��LɅO���&��c��03�<F���bAeW!{j�b5n�,sC�'��I8����ڎ����f�(�ِZ1\Q��e��axB�ݦl`�ш��4o#~�`��'(��:� ax�UҰ��"^6����s�qO��A��'��>��5m�<�.9!�f�p��E~�#M.2�~̺�,�J�0a��ݹ�?�{�I�h|5X��5v���+�'MB���G�n(��	���x�V����pm�w�ȄD"����$��+��Y�T�O��=�����2��h�`K��3���	�"!D�C�	3r.ȵX!훒T ����,��a�2��J4�-VI��,(#�� 	� ���O
Q��2(��a@��J!�D)�0i��0<	��'��	[#BѤ	Kȵr	4Y��h���3�4�Z�O��s+������;wBS�|�)8�ʚ.�iӍ�$�	K�$�!���Oz���`�Ҧ����C�AE�D��t9eጄ~���D/�V��A�3O]�F!��0PN΍�.�b�	�zs��k�=���KN��@�h۹"堁Ї���81�5�h�ꟜE{�O��S�LY�u+qh������뗀��xҥԁ9^uJV�ʏ��֡O�l/�����^ֵ T∘�8H���d�O�Ūc畷5� �:&.�NR�jFX9���d̔�P(�`WaS_���u!P)`Ŧ҆z>j�)cH��<���?yEG��d��ro҇*��� iH�?Y�mw&|���Z�H���MW�ud�Fy�Ź%XP��)F�Lj8�H���Wg�aC�iEH��?�)��T�ZE/� q瑷B�v\;��$�tS��!R�x��i����N0d����C�7�
V�)|O�}����O������)Qr^Ya��D�e@s7��ȁ6���[�L����HK�!*t.�>��<��n�=kw^�ӫ�8!�(!��Dd�v7���w��{(_�b��S>�M�$��,�rmY�EP�} I�P��(b�̀5 Ƕ%���	�ty��O\m�w�͚_o���Pgz���0Oڭ��N^�1���s�W��p<��Œ6��X�AޘO*"8��k�Syh]'9�a|2C	,�0��m�w"|��-_8�t�n�3&���FzZw,v݋�%J�<aT�79?d���*��0�
�o�D��$Ƞy�"���_2�,�ID�[i�����e.� ��к%�.�"���2D���_�Aq�i����2B܍�Z�1o��'���㞌�ݴBT�$�͸hL�4��
ئU��'4�!r��E1Y�Ԉ5)G#T~�#�c	W�\��aQ�r5@��<q����;������e�Sb��]��DP;I0�T����!������fxR@�Oǒv�ʤr.��W��	��HO��H�N��Ye�;�ِ&\i��V�I[�m�QnK�1�k�-!\O�.YA�@8k���3�L��jוp�'B�bǵD��O�	^�r�x�U*R�ǌ()� ��xL �S� :O:�:bLY�E)�a	��DP��(�[''.�|��&�5�\�hW�T0f��Le�����N�Z%#��]�P.�)q��}�`#���Ĉ��� O�I>$PIt�ƽ��$P�t|I���^�;��3����s#����&n����k�3'�Z;WB2	�����I�_������'�� ��JY*��u�Qǝ(Z9��O�X��B%d�1C����B�鞵~�,U D.�:3�t�a�/�,@��y���SF�Zw�H��O�@�&�H��g_I%�!:`� B����j���.[� � �!A�q"�(��Z<[z�����F�X'!�O���!�>§|����a��3ָ$d�N.kܢ%�K;6�y�剽V�DI�<6��$�r�
�$y.T�	�� "��+cEG�)�(�P�C'�p�I��ع6^d$�*OTM��.�*#g�y��d[
�T���A��I?8�˵N��^� bJ�+0!
O���Ē*�B�0��89ֈP���)Y�\�2�.UnQJt�F�
����OM�<��p�byªuu�=�W��s\����(O�	P�&7]*��S��U#����ch� 5�rqѡʝUIL�V�U.�F(S.���0�O�
�+)�>~�!+�_dD����2R��#)�yx�D��wX�����1x��]*aj�	��(!�\�V�=§�ܧ�yҊ�����N�4Ѫ�����^��)e���"��峍�d�?7,zpd��-��@��F�*i�F�"�2P��c΃e���g�*N<��.
7[wv䠞���06Ѹظ��� GuT�b^t��#L�j {�I^�v'���̜��ɃrZ�9UǇ>8��U����1��6EG��zؑ�ծn���R�"^�i<�b�)�����ٔ�?��ɓ�a�l����Ȼ8�L��*Ng�'�hջ��ſ/V� ��QDZp��F�KX��f�y�&k L<:=,��� �;�����9���{U�X�q ���/��x�
=�@����=�s0���b�+�q�\8�E�,syZ�,1������*V&�����|e�8���'rl���k���5$Q@����>��OD9Z7���a	��VMV^n�  �i�� :p)Eg��pZ`5#����g_��1���AvqsJ���g`�-*����B=�~m�0M b��w ���i������P6l���@��,�2J�P���Ώ?� 9�4e��fYV)��C�7�d��NE�p��Æ�Z5ߘ'������J�D�G}����MQ0��hġ�C݌Pm�y8�V��QNRQ{ҕ�e�љd["|��ՁRb�e�0dD&~���:��A�h�Z*!.-O���7�F9�D;p�j�k�jL	1�A�g[��4��r�V�*%�'= �86�~��J}� �udZ9yvU�# �kQj��%@�3�n6:F�̨2O>tW��"�I
����<� �{�çP(ʜz��A��\�S�OߺC' �(�'g̃W�>�@U�ģT�R��㪮>a`F�o�J��3I\!*�4�D�1v�f%�Ҧ�y���
\�d��g������m�YK�U@|TD��Q�'���Ӗ)��P&Zd�OUp]tz��	�ae2D�*�b��靷��R.C R��>ɬ���q� �9��D'k�0%o��Htb�/
�Ju���'�:0�	��yW��H��}�D�̸$L��WA����sc��O ��t'�$c��Z�
ī�]��j�᧥
H����bFׂ\nPpGy��Bej�㣭*#���f��d���2c��R�9� ��|ޜq+ѝxr�	y��ҪJ8fb�RBR��'G�� 2"G),V&1s@�ݫr@4I��k�8���E`�P:�,�g]fxy
�5�����x!Zz�e��g @yRb�=O�]�����O��ٔŚH�x�CiR�S���"X����	�N�ɞz�Y��u�y2��!}��黦I��8��<�p�K�xc8Г�'8���+�:�5���  �]�7"�M�"`�$�y��a��|����'�&�Iа	
�3���t�6,�p��I�Q$�$@P�� �ւЪM�*]��T�,i��Q�. �d�$�`MC�h�I���Op�##� ��!rɊ�p�Ђ����nثz����(k�F {��x��,9��#w��!a%�(�~Zw/� d.�<y��	 a��f!UR����	P�6�Y�B�!/�R%"ǋ�8���f����D�'�JdMkW-Ķji�u�v#(���ϓr�RL��IW�(����	#tfvQ��&BwL,C5����p<��펹<��s5��|D�5��*^I��rS��'������d'ʓ�v���ɗ�1F F��~׎i����7�l�I� 9��_��	36��\9�R8G_�M��.]"$��#��O����+��� C ��3� O��(O�����_�[?��)��� ���1�X��1#A�jN�3&�L|��ʖ��>w��R$�#����/��,Y��3'I�+A�N��?�!�[�25���Á;[�B���ËB��+W��|����'Ԯ0�<�����ZvY��	�hsz8�4cΐ)$z@� e��U��@ʶ�&ғ��'�V�y�(Kg��a֊\00�f�'	�xBͥ�b���(���)@��7u�P`
s�V9?�P��j �	j�'����� b����Х1�f1��.��a'�xB�)\��,d�שZ/&�F�`v�M$WCNa��C$x���""�ې`rP�!o:H��R�Q�HO�1�e� p��̒��J�b��P��{�� .8W��c�._|5[0,]����-�;;������G�ECҤy��x����}b�MV�uaC* �-F@��n�'�y��L7v$�f��Jl�x b�]y�'�P�PA�I3|�\�v�1 "�ĩE�(Ut�5����mo��<يy�o�/N�t�b!ʘ�f}����bz����XGx�|�'��&��������ʲW�`��V
@��⟠E|�@�p�0�PR��(.��"����?B�d��bY5�HO��h�g5BPT�AF�?a�2�Z��
�RwFpElوV0>��RjF�i�>���ln�'"�,��'P�J�J0�§��{�,(���O�qG�L#�h�Z|�l�%A�Hݫ��i�H=���?b��԰������7��!�h8�"��
*mjy%	�vj󄖳oB��֮F���c���Oݘ�	�=`Zģ��׋Q���iG���	�����D>^dn����<扰���B6�FT���`�)�z)z	��#�$��y�!�#>�j(�ݴz$���J+6�АH��r�8��?Q����v���V3!~l�r����K���H��d�#��T�&����	H���P Q&d5b�%�ڧ��%���pB����N,("�P���D4ּ�
^�V�XՋ�'��C
�y9N��3�A	2���2�4?`R�Q�'��<)�ʙ���4<���:5�߀F��ay�ؠ8~���R�ۨ$Ĩ�6�שe9�Aid�)�ɉ%��@k`�Y=nQ���R��E�@�X�D�	�@�My#���O7m����r7�-g�1uI� 5��E�|"���OXH:B�H=!j|��J�f��s���c�Յ�I�{��{BBc��ȱ4*�M�d�� ې�2s"Ϫ`` �6hI�7m��N�]�I�� �f�dC��OH��i�>qR�=�`=tB��"�
�.AX'�O� �'�_*uӛv�.����SF�=]��J�I�7N�Tp↤�~�`���mȉ�y� G5O�@q�0`�:�A0�?4JN�h�7O�,C��\}��G�;�j��o(�!��:e�n5�נ�{1��A�(�y�(�BD�Fx����}(<i!�Z�n��SC��5�n}Y���r�����t������%��P���-8�jc?AB�'���� R�/1��f�,D�$!"�P>+<��B��n�tXɢG%D����کv ��/'4�`�!s�#D�Ա���sB�	�L���<D��Pi�9����% Q�X�ޙ�g<D��S�,��;�.T��b�m��I,D�<#�HZ,A6mROG(t�xI�V&*D�q�Ë(��m�e�ؖ��9��;D�\ÒhƁ\���k��:R��!"�/8D�4��cW/\V(ؐ��^�Ή��&6D�D��M�lX�#�"�fU��!"D�� ���c��D���x�h�;O`LH�"O `t���l.�	��@�	@��"O�0��;��=k��݀[�pe"OL�җ�5��8���������"O���"j�$ER���S�"�*k "O����)��4���@Yq{�9z"OV�A���J�b�s��,/G��f"O�y�I��`���9�Q$G��˱"O�u��i��!���G$�I5"O��(��	&(��i��(��H�"Op�j���p, ��`Z\��|�T"O�P{"C���W��:�h���GP�<Y��	�l��U���I�L�h#FF[N�<q�ӡd]}�1KJ%ovL�N�<���I'0�1Y�'��K�d�H�<����Â�K��3o���3�H�<�B�L�Y�	��e2P,T��m�B�<��ɍ�D@ţ2خlƾ9�AL�B�<em�>
}�y�FI�iP,9�5�Xf�<��� ?6�80�&�a���a��K�<yu�ʓKr��N�����I�<i��ժ�H��c1h��r���H�<���MO|E 6��Y��l� ��F�<)eՏN��\򖢅�� )�&Jj�<�6l�s�x�b�%yF��v�i�<a�I)h��A+��� f�a�<����(mB���ޯt�L��k�Q�<�&gs�P$�NH�e�8]Z�NJ�<Y�LU3��SE���5�\Z�<A �k ��O2
6��V#YS�<qbH
�HƉC$��
:+� =����@���J4P��¶����Uc�=	A���ƅ�k��tA^q��%�������9��A���C��5�ȓ�T1��33���:6�ɴ<a�|��f 0x����M�Xr��.E4d�����-r*R�>��ȉt��.'�N���O�`�ǫَK����ȫA���ȓV��)�P-$O%��V�SzX1��JT��v�ɻ'��XS"��c�4��hA�]z�ەӚ�xv�M�n�옆�T��	���G��`�T(ρOu�لȓv�� �\$<�B��ӻu�@Մ�<��УA�ɪ �F-6>�$��>�������5v�r�(�F����A��2���K�Is��0'� �^�Tq�ȓU�L؛5���`I���E(ڻ7��<��\��Se@�L&�4ڂ�4G�I�ȓI�h��e<S���T��.��L��P�p؀���v�蓀�K5x�ȓI[��0#��"A��C TG��A��I�Lx�lS�
���ЌL�r��ȓD�4�a$i��p���5�	�Zn�Ʉ��B8�O�0L�f2e��m&�%��m�X�f�+�t���(�&�b�ȓK	��Ȧ��mNZ��ӆ�-�v���r� PP�m��a�tġ4j�	�>���N�&�a# j\������1t��ȓ>�,�yT�ϖFv����'�
��G|2�=6Lfp�aD�NG� �N�=PW�%��#�8 M�=�8�P ���JRd�ȓA�p��C�3�T��Γ0kI�T�ȓ@#F����$%��l�f�- �����SӞ5 ����耠�/��)�݆�S�? 8��A��@�x�dnN,B.{�"O$��r��l��l��F?��B"OT��������Iksa�~���ȳ"O�=aɝ�O��	;E ��I���"O�傶�%u�����e�\�F4�"O�y��i��ःt��#H�6���"O�Lk�0���#�A�J%ֈ�"O�D�u��9N ���\��c"O�鑀�$R��ZpʖR�L��r"O��I�d��pP|<Ѐ	�^�<���"O,��b ز@8��H�����p�"O�k���HH� iU.��DkS"O��BI���j&վ]Q�Ā'"O4�Z���nZ�(����_^XM�"O�uI��dm]P� �aP�P�C"OL��28¼�sc��eD�S�"O&	S��^>�P3�A��}l�##"Op]#��X�R}z�"���pԼ��"O�Eq�M�'i�� K���}c(��"O�m��nӺe�z�	dΕ����2"OD��ѮE�}(���P�'��X��"ODQ��W�ki�-��&�B��=��"O���UgП9Sh�Cu%ع���g�'�
�V�9bC%�'���F�ѣ|!�D�+/�4�:g��3Z�:��?Jt!���X�>��B	9!��IGh<A!��u&Ҭ9W�˗��I�
�;�!���SzR�jb�E�H��y��.\!�DQ�m�t4�0ȁ�>� U	!,��G@!���"�ة�g"����K�q=!�D�5p��y#���r�b��RAG!��4�����̨$eؐ@��!��!+<|"%�֋0����ԍ�>!�$��X� @J{���l�X�!��F�>h ����5¼L�'̜=1�!��U���Ȗ�\6u��M����:�!�$��s��=ɃM��t����n�b�!���!p<��bf�6+R��qD�;)}!��̏B�n4aC���+vT
���n!��ʹ/J�(�b	�4<H82�ĝ^m!�dHG\����@�8�;g��9�!�N��flU]�i�7�Γ�!�$�8l2��[e�W�F ���%
4y:����K2n̐F͇�3��}��
�U�D�<��T>�Q��K�l��R�ܛZ���3�%D�\�ԩ_�@. �c���gv��AD"D�`�Pk�y̮) �	]�`XH� ?D�0ʳ��f��n�*,�I�0#;D�H{�<��HAg�p-�N8D��a��1

�Fl��y&nU��%6D���"���V�b�	E��-@9�y�#�/D�l�gꀡ,��Ƌ.y\��8D�d��Ȉ'W"���J��]�5��*D��i��h�@�'��&y��qʆ�'D�(��E�}#B9�'%R�>��)�J!D�\p�'�<��Ŏ?62��?OD"=iQ�"X���g��_���#&�{�<��ON!L��:Q�ٔ,t|)��r�<�"M�h*]�]*�=)��w�<�g�ϯc�%���i���H~�)�'Y�����^�Q|H��
і"a��1{B1�Ч�-]��T�P!]s��1�ȓj�> 	@�7�X=k� Z1u2Y��M�bʛ�a�s�-g�����k�P�<� �Jv�<8�� wcK�pP��'v��� �nh8�Z�a�(%�pI©$D�< �c	�q�@y3%J��'�t�"LOJ� s@�ծC�n�"(خHl�hG"D�LB�m����px��,y��)a�����1{�>� O�!!Z�i�� '=�C�I�/AE�J�qv�Ti�oѬ=�B�I��c�/Ĩ�e(�2x��O\���C�D���ף�e���Se	Εd�!��^�@�
�+��#"�ő(h!�]�q�k��s��S.P!�ĖSp���nX�*��648!�$R�#�:�z�L��G��0�dC='%!�S�+<�`��P�:���a�i!�v��HfNX
@��IӲ`O'vz!��Q�?-S��W17�6)ۧ��u!�ا0���� G\I�BaE�3ph!�$ǉ�ĕ�5)��t��9r��Pf!򤋄J)sÍ۱Vp&(j�ʔS!�*d=��zu`>)�*�zFǄ�wQ!��=mbbp��Շ$�6��D��P����щ�<��%�$��;�� �&}��O�=��@A����zdd�+�*������"Or��0��5-��D�1���r4��B�#�蟀�8B��sW.��G�`��0�"O"�!TMA�i�J�Ǟ/?_��Y�"O
�p#A��t�VIډ2hy
"O��k�%��5̝y tjW"����'2}�vGͰj��5�Ci^�	JY�,OZ�=E�dl	<OgnY��<���跢���yȌ'e��T3`�]�\�uW@K��y2�Z-!��t���+0p5�Un1�yo1(�q��Ĺ.��@O�yr��a���H��.��e���E �O���SD1l����Jͤ����o�<��#�g�A���9yr���!	Qc�ĉ��0>���o��tP%�mm��+CV�<�p�2;��p �P�NMb�s�M�|�<�!"�/\���b��\����R�<�Vp��s��R\�E��MH�yBe]�[�`�J��4K�� 
��و�y��)m I���^BR�=�J5�y�f֩i-�1���] 0�fP�j���y�m2rb����%|Ub��$Y��y"�+�<Kֆ�'v
\X�t�σ�yB��5;*���  ��$h��P<�y���&z��i2��Jd �:�?�yǨ{��|����& �Ģ��yLo��	1)"~ءÔ ����'�az�b�`���"��-���w��2�y�c�N���cP�ҙ�����:�ybF?z�X�7�Su���#�iS��y2oA6�-���D\��<���c߰�y�*�1m:�ca�a\�Ic�
R;�yb/��sq�0[tNԍ,� 5�bZ�y�O�Y���hV$z�9@L���y��/��C�ߤ��X������y�K�v9
�ⱨ�-��G���yrK�k6�Y8�e�{;&iK����yrHʹ2X��ĺ}G��CN���y�oɢ
�Ԍb���`���<�yB��F  �3�G�\/��ЃA�	�y��P{X)" 	D7Y� �c���y��/p����ďX T���:�y
� >�Ʌ��;6��xITK@����"O��q�U1����S�c1�I"�"O� ����$������*@B1�"On�sd͂9��C��V2=��š�"O�@K�/��Dݚ�T)�B��}�"O�e�L�-.EV[��x�\�ʔ"O`��ǫC:f���cB�.�&iY�"Ol��2�M���`�7j8�$�b6"O����e��yM�`z 鋷Z�́�"O�U�0�D!&�@(V�N�~����P"O�Ңg����!���^s��"O�U����Ia νorIAp"O:�#`':V��y叆56�$���"O؀I��5q:�)R�I�D`1�"Oy�.ERu$�Q����<�3"O��c-LD����:q�N @"ORh�Á�O�/�^��S�"ON��֫��)~�H��Ύ-���sv"Oz�Jq��vr�Z�F�i�Ĵ(4"OR�1��cI�w�¹^1 �"OAC$�3lI�!r�F�:{<8%"O ��fÖ́i�L��B����x�"O��RĨ��
���Am@P��"O�XquD��n���=`l�)�"O
��rd����gmŧe��"O��nC�=�bI�e�ZYn˷"O�l�����f�t��$9#U�)�""O���4�J�QT⧃ǫ�$��"O�`��H�:M(��ö"	�^��4ل"Ov%2'�U���W8c9��
4�M��y�i^�7�֌C��h�6�1Λ��yf�	]Q$��;]���g唕�ybኧu�l`�0���ZT���u.U��y2������i  ��d�F)�yR��oм�6��TT8��b����y�OP����惔�H��sU+V:�y"+��@ �Xs�KW'P�i��/�y"(��0㚸�F!Y�Qݰ������yRM�J/�,z­�*Mv��9�F�yB��,֮!srM8Y^�TL=�yb���O�}��ћL`��:�yb��+x�e+��'�V�E��yrF"d��K7uBz�r^��y� ��nI��'�¶p7� ���y�K	�@�R"�V����LY&�yr�H&Z�2S`��(�4�I��y"(�{�ܛ�&_�RE4��h��y�C� �@�CčF���Ca�ª�yB-L<v�����(<��c �D0�yMF�_���a�N��:r}��M1�y$��Cp� $ Ϋ�Q������yשRzZ����0d�>�cB�߆�y2+�7m%\�#�!�\Į`:!+V$�y�$ֻ&��!�(��&�0���HM �y�k�/a�t@;�
��JrJ�C��ls!�DLW545���V�Tc�m���ʋ-!�d�y��[��&)�v�Q�G�Q�!�dJA,dX�wK�3$��]�OȖ*�!��#wy��f��5�b
�֍94!��<��o�u�{c$�R1!��3�����2eq���ʍg!�Y�&�Da�H�kJ��� )$�!�d��ysh�!ԣݝ�|���G\�!�䖚}P�=�RǅA<�G�:�!�� 0���?v�	�#M��r��"Or<�F�Y�!� `��e��ZR"O����O��m�u!�=*M�YZ�"O����e܂�&�#�D�/L���"O�����ܞY�^x��"O�5Aa�\�a�ZI��mܠm�dl�1"O*�CL��~~=S�%_�4���	�"O����EE��0�ԬYs���`"Oh0�e�Ei��ˢ�� �"O��/�?:�lz�Է��Ds�"O\U:#`H�;g!Y�3݈e��"OX���w,fܱ���'Ō-!2"O"�Ju$�*U��9��ԅ$��T�"O,p��"�?-�+�V�@�<�B�^�<Y�眊���㑭O�<d�R�mEe�<quJܺu��]#H�W�0��BK�<�ƊP�@�.q�Ѝ��lѡ@O�D�<��웅_LNu����
��]9*Ev�<�u�P1����G�,\��s�<�bh>_<S���z��ׯ�I�<ys ]����PLQ=l��(c�KG�<9�	�"I�SB��Q���c��O�<Yvσ���D���6���Sv��J�<Al�+@�B�aS8F{���΋P�<90���<<�}��K�5X�\'�I�<��0���+"T��`�09��y�ȓ!�\�c�G�y�$)s5C�-�lɇ� F }�Lݵ���B�!�zʀ��ȓ(Y�BTm̥d��y
�c=,ɀ�ȓ*j�c�
�3����d̚�>�*I�ȓ �R	2N��evƹôb#wD��Ū�su`ӹW�u�Ac��T����� '<P��E�`7"�!�n�9�����hg��r, �u�n�!#�NOj�y�ȓ#�pH���G�O�pء��E�^� �ȓ>�@L���o���TD	�iĴ���!�x�n�TVt�߷mڠ��J��y���ǻ[�`	'bF�UԐ$�ȓ p9AC�V�	�T@X�!�`��ȓg�� �_%�x�.̶
6pM�ȓD��	��(�)q��9����ZцȓG%��t��W���4)��)�>A��
������Cdv���O�6!ed��ȓm'<��$#ĠT��Y��$Ι�ȓtz���@�<d�����c�"��ȓ3��6���0�"`��.אS���ȓC���[�A/$�D��m�4_xu��/1z,�tF�Dt�Q�"A4H���� J����КG8�"$
�0dڐ��ȓ|�ă�숗s�p��æd���>��B#��
�|�� 
DD�I�ȓq-��é)�db�'F�{�����[� ��� ,� ��3�M�mȢx�ȓ	�����c�1L �3�+�`�@T��"��Xq�d- �q
�<~sȩ��f��b��d$�B��5�n-��:��)�ˈ�7�c�ɜ4b�b�ȓw�"Pc�OTs=� �UL@�JP���ZP��˝K�
:��\I��q�ȓ\�T��DK�oX:��C�SPA�ȓv^�Q��d F��Cs�8�ȓ.�㳌��+J��af��9�ȓp�ڠh�N].babA��R
F�i��|�]cRn�5b�L� �Q��|��S�? \u��
�?�RL��`����<1�"O��CG�3KHܴ�D������"O����OC�&��\Bc^�<����"O�����A(<�#"L�M�ڤh�"O���)G �&Ł@�;gp@UY�"O����E�$da$0��U{�8�5"OLD[��¬:���GFΡbY:�#"Ol�فJQ�!�l��Ŋ/pL�<R"O~Ȁ"P1a-�\Ȳą,CN}9�"O�W�R,Qa6���yY|.�yR+T>N���FK�	p�Θ8�y��N�����^(��u�
�yd��>w���f��9Lܤġ�
���y"�Aq� Qx��U'=H��Q*I��y2��3vUz��0B�#Z2�;B.���yR��@��f�]��DYPaT�y�m|�V@�6�5���a�M��y�Hȡ!F:|u��&���%cI�y2��.��M-J+@l��G)���y�`�1��m�Ǥ��p��ȶ�һ�y��L}|�� z�1�-ת�y�O�$�栻U`��]5����B���y����3�P�*1 ����y�B˥l�&��8�ֵk
���y�D���V.�0䑣l��yb�*D�jP
����$l�)x�`Ѵ�y2j͙+Jd8��2?��pcCφ�y�"K�)����������b$���y�j��SӪ��bŒ�z$���U��y«۹%��T�sN֋�"��` �y2��l�H	�0r]��$ *�y��S�������Y�<�A�<�yrj�;t�Z�� IS�K�7�y�Ƌ8q�z�Zo�
�3f^�y�J�7,����S�_�,�� ��y�K-l�d��J�j܄+�  �yR�� Q(N�2�kհ�F��щ��y�M
� �3�Jcs�&!\��y2K�&�$$����a���&'N!�yR�Jk�$�+�F@",j��'-�y�ΗIzu�G�o@�Q����yB�L2K�d�%C�w����	@�yBÏ�l�v	�f�(t�"�"�ʕ��yr��D�E���� ���	s����yB@���BPB��z�L`?�y�҈$����>;��&���y��Ҋ,&fxi�eY<=o��z���y��^�b $�` �4;.��!"O��y�B�HJJm֥�1.������ �y��~��#w�'&LL�vӾ�y�h_��ȍ:alX�m�h�qi���yRƜ�c�^�C�D�3
n�f�G��y�b�39����`�5u�2��v�Ȳ�y�Dն@��`�@���t\E�u�;�y"hF�g%��2C'��x$�L�P$��yr�*B0��4��3@�@830g�d�<G&ɮj��iMR�I~�H
�Έr�<!ǈߠ\�U�6 M�r#�y�%�
m�<��	
7VM�����>rZ��
��i�<)�C��>k���t��4l���"���o�<q�-ʷ?\j�h���0cT� 1Ɠa�<)#�O�K�����Z$j9~,��.]�<Ѥ��2fj� ���3�!�@MC�<�c>w"`� �V#�q
t@�{�<� ��:���j��RV�^��f��"O��S��/&xD��G�~�Ĉ�"O(���P���SNUt����"O�y�AD�]� C�L̀�S"O�A�n�O0(jtJIh4x�"O�h;�����-rħQ>�n=�"OX0��ӑPD��De>� ��"O�l�0F
O,L���Z�i��hC�"O�<��x�5J�	]�$ذ1*�"OP��5G�\q�����d�:���"O���/M��!D*�T�x��"O���"&
X@�I�HX*nQ�IC"O.��#� $Ȉ��e��]����"OA�5M�$ A����6p `�!"Oh�3�dҲ_l�P�¥zJL�"O��cW{���*�!k2t!�"O��b�*J2.��P8��B�fP6"OT��I3ޢ� ��МO�쐹P"O1;��[=|��� �G�3*�A	q"O
:�G�*��QDǂ4N�p�"O=�Uh�.j�v����V�<��iK6"OV�b���I��gE��JY�c"O dq�%�3H�՛�A܄_���@"O�L��&���D��"�F�f���"O���˞!iVh���kצ$��yC2"O>��Ş`NU��闢.n��k"O2�COV.>���H�^5cm�=�"O���i�0�a�E�Ι���ӄ"O|�c��0(�Z3�皂�j�( "O�1���8�zu��#<yw��"O,��5cM�cU�(����1`&�)t"O�Uˀ/?B�����%"LP�!"O, �̒<O��m#�S�;dr,W"O�d8Ì*.8��af`��HH���"O�8�5""(���@ �8(R؊�"O�	���9N�NX� n���"OlH�c[+�`�D���O��ѡ�"O�0��I#��E!���-&\���"OD�hcM*|<�)VmU�]%	q�"O	��m�6O.�@'��1,�xS�"O0�1�D�~�9��!~'�!"O(�����lM�C3'.eI7"OP4`fA
<>	:��r�BJ�z�3�"O� x6 �'Z���.T9Ѽ��"O�̻ff�U�r0�U���"%9"O�u��Ȑtt5	�M7dD��0"O̜��`E_��9���=Vdt�b"O��߃_��`�"Eθ��"O�Tk �K� ����pO�*+R��e"OhB�T$M�R��D;vyrr"O��p�˴<�� A.KcJ��T"O�P ���`�����A18I�9�u"O��Z���G@���#&.N��"ObeP�'\l��D<�,�Y�"O̝	����#���#��"i�40�F"O�9�C������\|A""O�9�V%W�w���*T;^|��"O,�����
�~��W��F���W"O��[T��ZX����(�sݞ�ɠ"Ol���E�+��$C!*,9&x
�"O� ��jG!m?
\K�Yx��U�"O.%k��� d5�����R"OR������0`���n�(I�"O��"��+! ̌�%�L��īc"O� ����(M j��YTNN
g�d��B"Oj<�ԣ�`a��bG�J�,(�i�"OJ����*vi2!A%�MJ ��SB"O��a�/N.wv�`򇒕%��2e"ON��D	 �����f7����"O���WcU�7����fŔ<��D"O2��t@�2ٌ5r���u�V"O�
f,��r�0Y�E��Y�=��"O� sI�T&詰*�o`�"O��*@�=iVAY�i�<{g�LJ�"O��2��`�V��7��%�hC"O�� �L>Wx5�V���<�\��r"O�=�Tc�����ω;���V"OҨ����!T�TE9%�s�js�"O>q��`��(q��w��	�"O�5��@Ϯ"��\�0#��.��H#"O�I�AF����1 Q�-'�j݊�"Ov���P�CD�s�Ȋ}�j��&"O>(z��J,c ���i\?g�6U�"O��1B��5�hpJPh�S�.D��"O�=8� "��(V&�C�n��E"O����܇k|����G�0��"Otu���"zO謁�)Гh��)�&"Of�8��ZC���!���
t�"O�E�63� X#P��^��u*O�8����o�`��>C�6U��'��d4�ڞ+�R-;c��D1�' �	�V�'#��`�(�6��'���[���2Di�`YP��-�\d�	�'����C\.2���2�Y�x�Ze��'P�͓i�E��X���p
r��'4Hx���8���+�쐛hm��c�'_l ��,��V5j��+ �\W�P��'4�i��)�1^�� �ڕV. ���'&�i��WITl�R��� E���B�'����\y��[X(-�1-MB�<��--��:��X�"�R��#�G�<����2�p% �+��&��})H�D�<ɑJ̜z�a�$�!Vڭ#� �B�<���#oߜ������V�n���+A@�<	E��#gŔH�%ǌ$bukFd
}�<�)����yԊ�<		4Q!iUv�<�%���[@ uf!x-�Xc$�LN�<!�K�"N��uЁ�[�zt����O�<)��T�nbn����+]�PP�J�<���^4X �����i�֤���
r�<��A
r���#�͖M����j�<���´tBօ�D�ɸ'��K�_�<�w��/�z�u��Ԟ!��
[^�<��o�`Pja����|�*!��b�Z�<��G��B�ҕ Ǘb��B�D�X�<��C_;xȦ��B�`��H1׬�n�<�siy{d|I��*8��8�"O�{&���-��(��)TN��"O=!��ΥY��|(���6����"O\�3( G�"���_��p�"O$9����M��Mk�l^G����"O�H�"+jʮ`rP�K&��AQ�"OL��$�[�21��Q�`�
Lj "O8iA`cm7q𰊝��I�!"OZ� 3O�Y��@�F�i�p��"O�4i�j�:�rh�tb��k���"O�ыѣ�0H�j��nD����@�"O3�K wp�z�^B��)#"O� .-����5*����:r����w"O��ZTL�=[��}[�)M�X��T�U"O
]إǖ�����i\ l���aC"Oā+@��C��(Bi��X��"O��ze��!N�I�5Gޜ�q"O6�:�HņF�8P�
��8�K�"O�8��J�TѢ��S�B��b"O��X� �%0b��g�ƍr5+t"O�9�0�T%D�Nx+�FJ�*���i�"O��3�Q�L�D��ʛ`3\��`"O��[�ϒ;��)��-����c"O4L�FN�u�������\V����"Ojxz�HS:J)��XlA�^�s�"O��P���:I|(;v
ͭPE��e"O�� ]b(0s��$B ͢%"O����%_�Ӳ�����.���5"O�(���Tu���w�	F���D*Oh��cՒD��D�P�5��0�'7p�"P�=EЮ�I@�N�t��8J�'�(���4A�N�g�]>:���'� �)��Є5�<D ���d�(�'$X���pUiBF���{�
��'��������8�u���p��A�
�'�%��4� ��u�mD��"�'��k"$�@{F�V��fi<	�	�'��LS��5z�xb��ێY0(���'a�$�-�>B�b�Q�>^x"
�'Q&� *	(V�rD��ぃ� 0�	�'�$��)\y��h�2�T�u���;�'���ڷ���X�h:��-p�<���'�hA3���0uc��,<`6<C�'�� 0���W2���HZ.q�)�'�������h��1Jw@O�"_8�q�'^�I�/[�\iz���%�H[�']HI�$�˩ ;|41���.5���	�'�B��E���q�����)�&)	�'W|���i7P�݁�
����'�����M�]��B���Ra�'?$3�l�t�*�@��|���'��au�� ?Nɡ���x�Z�Q�'�|x�����En(�$/R�nF\��'�X�8�+� �݂�K�bk��b�'�nmÀ�t88�c�7nXN�"
�'ᠵQqEBnn�BƓ,aOV�[	�'�j�Y��� �~p �f<���'O �X��3T6���9^�X��'���sņ�G�U0���N��4@�'��Y��\�������M�J$[�'\jŹ�h�#G� `%"�F5��q�'�:}�3șN���%&�8Ŋ̆ȓo^ŉ�k�d(��I��*P����[�nlA��	�q��t��"��q(sD@N=.Ô��#^w��ȓ#g�-���**B�0�e`��^�Lt��-��IG�҂-C�m�G&�lTl��6�l�;�&P6j���ө�ZUPՇ�xP�9j�J���,�Yf�L;��ȓv�"s��j���� �"y\����=�����W�~��p	WOK"����ȓxLN,�1 (l
H�� �E$:���l7��$�b.`�Q���G�~i��J��hж���L�Tb�ӽ&�Q��-�6}!@H��"��cˇ�h��ȓ_�qqc�N�\貤c��X�C�)� X�6.\�=���9�#s� ��V"O� �C$�5˾ S�"I�Լ�"O��h�
��JK6��8��ʷT�<��d�8G�@f�	��w��K�<�"�$VP�s��M�t����H�<��ყ�<�[Q/��:"|ٵ�JG�<)��^�켈3	�FN,�ࣼ�B�	��xQ�
���CqI��8,B�I�v}�����+[�p�2�G�rj*B䉼{8��0��Syd��G��0ZB䉡 LB����C3�д�_#g~~C䉪}���1�ʦ��=�R�%�B�I�jITy���
SU����J	�1]pB�M�ֈ��&@�Tը��U`��"tB�)�2��C�Ѣ4��X��/���C� +��5I�k��Z+�\9�ʡG�!�������U	)@XyQ�-X�l!��ʀ^����LdG`�tcA!6!�G8L�Ѡ���-�\D��W�!�DW��%��b���ZѤ��Ha�}:�'�BŨ',بf��}�`LN�3V�X�'T���򃟠��d�!I�8R��I�'�F,sa�×%@��#�L�1��p��'����f������Q�T��
�'i����Y5%ꈩ��	"���9	�'��SsL�""<�%iujF��@��'����4��0r�B�U�ޓ�Ѕ�'m:a��!��y���_�s@2I��':N��2�E�L�4�N�3n*���',��C�kO�Fj��HO.]`>�K�'0����N�s��Ҥ�G��ʀ�
�'tH��B$@Ay�^3k*���
�'P�<b��L�N����@�g�셢�'Y�4�|D�w!��_�ຄ&̯�y�#(�dh��մV�Nm	w͉ �y2%T�SfTp���,U��u`v%�y"��cg�1��)�R����/O�y��Z��6�X��u�DM���_��yb`A�k�L�	�8��p��H��y2\?�.�(q��;`�|���y�D� SE4}�D�ٳo+�h��)���ybL�G�|�ӄηj��" ���y�I�%h�Y�&�ɺj��=����y�L���hy��<^0����bG��y��tv%������lR7�y�A��|X��!E��q���1��!�yң
8���W�¹��A^�y�OW�Gtt��R�w��zT�ʞ�y"-Q�d4}�%oJ5}�RԠsj���yb�P%3J @�3�I�q�@�f��y��
PC�-�'�@���S����y�JĮ�x��D��E�$��CP��y� �(X��Ir�6sy8��1&]��y��<'�b��D "�$Z�?�y��@�jM�,�A�.T� OK/�y�d�	3xQ��+@�"T��7KT��y���&fpm3��3��$��Ѧ�y����$�L���)�pڽ��Ø��yB�BS-��Z�0t/�MR�Iң�yb�v�~A  �g`��ӡ	��yEM<�R�ᐲL�cSJK�yB��,l,0�P퉍[i�Pr�-�y҅��]@��BI�Y�L)�*
*�y���(C�}#� G��X��	<�y
� ���Gυ't��tO��C�Z�"O,� gҨn����B�"���2 "OfPG�ÿ[���������"OB��ׅȱfB2DxKɪh� xz"OF9k�_`�x�֪�)5F�h7"O�e"R�R�VX)�cT2`��"Oz��"!�Sm*Y�1��A�&�kV"O���bj�rX���S��/7�v��"Ob!"� R�%�]#��ܒ/rV�)�"O���ݩi����ԯ�*m2"�j�"OR�qdM�e������_�P2U"OZԸb�<uonx���2M�0�"Oph@�,P3����ꋍ2����#"O`��u�<���")�5XJ��Ҧ"ObD(�#W*p��T���28 RR"O�E�s�̲.�|�'<.��#"O�d��nY^mZ��% E�1��'�T2�K	�K�$����f��	�'	�����:�����,5gn���'�|Z���r	�5���Q0'� ��'�p�*�A�-M�"�ai�&��':d����ȁ@T9�G�^�}*X�yR�ԧX���u�V�x�3,U�y��� �� �q��q���� �yr��V,�]��O�w2i�c�V��y���}�,y�Mf�r�Q���yR���0Ebw'\�`:��*'
��y�K<���LX�`(��-�y�	EF�(RF��:܀���x<�ʓT@��ҁy6~�K&헕��B�I&VŪ�A�D��n�	gD("��B䉁޲�Y7�^�&@�쓧#�B�	)@<�po�7n
�QBa�e�B�I�5y@i����'qÄ�c��C�I)W�^dh���
��\Y�A
Sz�C�	�Z�, �r�p����Ԩ�9..C�I%1����-��>�q���SZB�I�@k�e36$?�@��o�8K
C�I1G�� ��m�2�WJU;I��C�S��jc��ujڝ;�!�4��B�	�%��"G�9�^4�k&hH�B�ɥa �=�Ѧ,O�����t�B�	)6�^�Y
�z�޽��!�v��C�I�M��X��2Bι�0�ц+�C��4��Q��ۓ+�����Ђ+�C�	B�p�D��+5�a��
��"QfC��&Z'�(W��0Bp�Y[6�ȼ&�xB�ɞ �nْ� ^I�e��(Čr�C�	�n�dtr �!��8�j�Ec"B䉪'�J-��)R~�%34�աe8B�Ig�Na��kǑ
8�<��G#;ZB�I�.Qਢ�l�'+K��+��D�8��B��4uҎ�IծuͨT�c�=gE�B�I�|hٰ �.0w������
?GXB�I�R�
�`�/F
����E)�"m�8B��:~�����۾'�,R�*^�� B䉖+>�CA-�}/�I�c�FC�	�Zj���b�Y��ɡ�!Ȯm�B�	4)����5I����C�ɀ��d�a�5A bDʐ
e�C�I�Ҙ��+8$̲���EʔFӆC䉓e�f �֨[-�hSwKȪ��C�I,|�Xx��&�[v@�!>XB�	�H0X!ׂ��R�1�T	D�-��B�)� �"��]�X�6j�m��hX"O8�'C�v�I�F°\�r=�"O��jBcU��P�u�K�z{j̹S"O�82uӯ}�-�fʴ<p­��"OF�6l/2�JTҀ˄c
�]p"O�q���W5�l`��׬n��p"O�Y`(á;&y"��6U˄�x�"O� 3�T(`�xD[�H� � ��"O8�j��	r���/E�KC"O�l	˴B�T�%g'W�h��U"O^���~�l�a _T�Qk�"O�ԃ'���`�� oS ,Q��2�"O�,�A�߮M�08z� M4P���"O8���{�yбnH#4�
A+p"O��J�,F�x�v8qX��t��"O�$�5�3�Z��+���[�"O�T�bCӅ;.���I
sb8:�"O�k��ӊg�$d�CΗ�5@h�"OXA�񃐤k4l�@Bm��E���kG"O�-)��8
 a���ne�"O&��ׇ(!C���L�x���w"O�@:�l� \���Ō�W��uc%"O�@H���k��� j�����'r��S�Ua�\��ɃGs�mh�'���3�ڍa�D@ʁ	�F����'��<����	�$pQ��)m��5
�'�ѩv6ϼ��U��hj�9q�'B�� 4iO��� �K:u���' F�.&+<<�@i]�^f�1
�'4�k�\�I���.�Q#tl��'|�I"6�\!S�j���&�\��l��'n��R�@K;���+GI5ZKF<��'P�5�
O#�B��Vj��J�<u �'���IF�0>FmhQ!�Ia>��'h��go�5oӘE���7H����'�J����O_:�'nV+	�"i��'���*��F!�e9H�Y�'(6,K���c^�����̠R���'��+#�(h|f�#��W1,�)�'c>�Q��Ʃ\"�A	6��_�Q�'=������.������B�$�y��(�^\*$��`�YK����y�ـh،���Q��z�υ�yr�ȿL��[�H��RT�P,��y"�D;��"����o�L¦Ƅ��yB"��
{�d��+jK�����܄�y2�_�~�Tx�C�Β^,8±�V�y���L�F��C�QXH�r�� +�y�g�=u��g�3P��`��A���y�Qd-��jeIٶ��HPt��'�yrD��K�!��bN!r��X"
��y�BԈ�Ψ#�~��Ы�b֗�y�iՈ
R}36��G������y¡�Oł�ɷhҿ=\<�A���y��]4-�ly���W2G� ��@�И�yB�+q�tU���ׁ�J��u���y&���pk��5���Qg��yr��-��0C'+{��e��h<�y�GO#
�q�3�׿y���@
���y"�J$E䶤�Vi�1l/��ܟ�y�V9�} D�q����7��y� C�v��tg��9xfu�7���yR�E�s�z�����&@���!��y��/=���� �9$�-AR�F��y
� �<�-[�2L��h�;PB3�"ON���%H(^����E�L}��"OT�2���jD�˴F�1�^��5"O���tK�1�\c4c�=��4�P"O �K����o��tG��B�{D"O� � �V�����;Li���#"O��[0e�y$rt�2�F:E:ʄQ�"O���կR�B�Du�e$066v�a�"O�a�@b����O�_�I�"OX̳'Ųg��t��f���H��"ORP��	��kb囕F�8�g"O�8�t���km����a
�Qn��a"Op�	�&--D�)�����ؚ�"O����%�7���P��� h�
�ڵ"O��6i�+�4��qF��DP8�"OF�	#��MzT�Y?5���B"O8H��Ѷs��Y�c0��1"O�0EO�O��曕D�[v"O<X! ��nqD� f�N_�`g"O��Q���
�Q���w\�pc�"O{0p�VN<��@`R�o����ȓ#�$شQ&�\�p��YBd�H�ȓO�r���*�.(�P�@%A�U+݆ȓF�Z�A���m�$���:=�=��jq��z��X�MZ�q� 5J���ȓ�NU#��B�y��8�'@ X�@����=��� ��HE�9\����ȓe�X|��eR|d���X�Ň� �zA8�D��I���d�diր��4���U� �vu{�l�	E�����I���4|d����ׅ����ȓV�����B�dU���b��r`�E�ȓ\�T���҇mhh�Tm��JC@̆�8O����$@.&@��L�BbJh�<1�d�Kx���C�B�Ȕ(b�N�<1U������̔�
�1�n�<����+Ӏ�27�J�����I�b�<�@�B� R��5�*����G`�<Q`F�������L���࣪�[�<I҆Z��x}9��P-R��Ejeh	a�<Yr�ĮaJ��Ie �m�UI��Hc�<�U`�g�L#��
"	���g�[�<���V��1�E�\�Zyp�
�M�<Y�ح{�x��ѫ7"���c#�d�<Q7큏�h��7��/gK��:�	^�<it����x��
�a+D��P	�^�<�n�<i��m)7㐊mw`�rc�X�<����\lp ���ۈS  �BCJ|�<%�\7]��;�m�S�I�@E{�<�`C->D�mɄ.�(p`��Qq�
C�<9�H��^4�ɑ7*�V�N��f�]�<�A�6t�� �A�i`\�s�a�<�gc�� ׀�җe�\`�HK`�<Qo��L���rF����І�a�<9�i��>}�Ɣ�9��(�#�^�<Y0�t��T1*�<x���]�<�2��B��Dp����1 <фk�n�<�7�ݶ6y:��E=G���c�m�<Q��H�"݋r�,�D�x���c�<aW̆#zal9
�aA}����AI�<A��B#$`%#���&1i\8Б��@�<A�oR�L�B� ׬!;^�H��E�<�2f�M�ʨ@�g�MP@���-�f�<9�͋�Z젩��*Y����#`�<� ƉxV*�?P�zf�1G"O�[��!��+5�4Y;< k�"O�����
�
��<��������"O �� �(�� ���T�&hH�"O P�%�P1UbM8�*���J�"O�ݨ��J����!Lv"OZ��@�%�>4I�'Ⱦ����"O$E��ʁ�37Ne��˱rYn��"O�4 c�ȇr�\� �D�/bD�*�"O<�E#�!JQ
�n�oD�)9�"O4��h*r\l(��D�F�"On����)�jT���FG��d��"O��
�D���Њ��:z���"O�P8j]jH\1 j���0�"O��+AΆ�o�R	��o�+ �it"O����!6OL�K��9y�x��"O)�t� ���{�͇��""OTa�"�7��<P'K�w�TlqB"O"����ϩ<h�1�gB&��;""O�`���J�N����� ���B"OruB�&+�&���FXR"O�-�@�Y O����ph�K�d5�S"O�����2��ufF�Vq�-Q"O��kD�˦V�@�s%T����"O�D9���u�^#NZ*UG�mQ�"O:U@�h��z/����^W?V ��"O�}h��L{h�y2FZ�Ap�"O69�T"�d4�st�K�mY6�rc"O=9U��9@��p�K��M(��g"O���4�Lr �a1el��d"O�Ɋ%l׍������
o:�г"Oڨq��$@T	4&R�_SVuI#"O��;��:W-���0��l"���"O��Z&K̂t%d9���?Lc�8�"O88A��U���� �  �b,D*O��F���!�/]�7����'t�p���ҝ	p�ҋXe
�H�'=�ZC��m�����I�V�^9c�'�u����y��*H��i`	�'�QQ��7>܂Q�B5o�!a�'��L�V!L:R������~���K�'����ݜ6x��Z�)��|��U�'X*)HG���$T0�1�fE`Ѹ��
�'YD�CF�P �s���7e�8I
�'�h26k� �-H��G�.M�T+�'�h�9��=�t�a\�;�R
�'k��Aj@p>�Y���bjM�	�'^��qA�1"��r�R�
Y�	�';��97n�{�2͚qO�!V�$E�'N�=YЀ��-8e�3 HK�|`�
�'�8�
���ôT�%5�8c�'#V�P�9���k�Z�^���'a�p�'f�%!3���l]�mF����'�`���j�c�6AT���}��< �'������w8^DsS��m��h�'dX�I2�΀2ll`Z��B%as�q��'�R���6��Ͳ���P��h��'�R(�p�USXz2,� C[����'�<�I]�<���ʍ q!8�*	�'� Xt.Iy��*P�p.
�	�'� �8��M-Y�j������e�#�'qT���m@�z�l��wd�h�vQ�
�'�lz�ɬs2q7�T+�jܘ
�'L��U�?p��}(�Dĭ��%3��� �P�E��b9$��L����X�"O�4Ц�$hU��'��)�s"O�m3d��,G�)l�Bl\pY""O�l��# ͢�����W�Rty�"O�1Y����Q��\�B�[�)F���"O0Hu�+ �N5x�O�~>&��7"O��u��2&����u��`=~i0"O�1ʗ�=x�Sv��h:���"O��R���O�P,ysπ�$�Tr&"O�H[��Wf2�ℍ�(5> �"O����Ke�°�����y�"OX @�jE�+؃d,�k�&�#�"ON43�P3j"|�J�q����"O��tA�U	fu"	�)���R"O������E��D#��R�B�y�"Op	��g�(��C�&e�@a"On�[&��Rk�-q��'Dr<d��"Oi�m n���rka]t,h#"O��a�a:u4��y�I�{��J�"O�|�w�R�/���H1n��N�<h!"OF�%��*'�ԁ����7DdH��'�P ����1M�d=t���X }��'K��'�&(���-EO7`���'��0)��
& �Z����V9|�@R�'{"4`����B���E�x�8���'��0����r�p [��Z�oY�t�
�'
�A�ˌ�!�8���<T�<��'d,jv�Ž_�Ks�$0�6�Y^�<IaȞv�.���5h�`|��P\�<�&��R�Q�����b���W��}�<9��h>����?p�b�!���x�<��kҙb�.�# �ǃ}���Uo�z�<���
Z���sm�>Q�B0�7��j�<�`c��3���/�"YP�Ih�<��oI;I ��k����W/o�<9�F��D�ԭ�n,��%R�Cj�<�iF�/���Ae�$�-{p|�<I�d�!2����7	Y���X6��y�<Y3DɧH�!��̗U�|u��
Ha�<Aw��m�ǎES�]p��Z�<)��*b�FS"��K/H5���k�<��oH8O�.y8�m�>g�b��g�o�<���_'W*(|KbI�=� �r�m�<A��8�x���@/L𠥅�f�<9�8Y�%k��-6�,� ��d�<�e�;v��++�)~
�ʖFE�<����lOԌ��'�+DV`4Z�$@�<	��
U�)�%m�1`�P���o�E�<i�ó{�����09�F��t��l�<1!�Q'_����+Q0butmx3�Qi�<� O�#�j����*R	 ��P�<1�)��=d0�[e��z(f@�u�J�<��g�+86zp�G�E��h�D]�<i҇�_�`-S��rtfu�sE�d�<���ݰo��qg"1j�$ܸJ�^�<�����xp�c�0# <5���[�^ɒ�02�,Q�E'��B�ɳ*!���w,-{� `D< � B�I"P �b�Z?r�i�B���FB��6X��	�@z�x��ؒ&��B�4T�H@��ƴ4�4���ˌ+#}B�	�w�'���y��I��E�v4B�I(N�h	&�ūr3�((�·�p�C��}K
!Xl��D� �(��_:T��C�)� F�a��xd �#�L _$%��"OFtj��0�j��yl>�
B"O0��E#Y���qB%*YY(���"O�yS'�*:r��ʲ"�W��ȹ1"O6��&�&:���ҀݘJ�V��%"O$"�DY�"����\�*1"Oht�냇
v�E�EnӏW���&"Ot!���t{�8�5N��vz(�"O�}b�n����,I�A��a�"O� ��H�u^)�� >5l� �"O��!���"u�����$+�ԙ�"O��v�W�/�VY 1�(<G"OL�x�� �r1��
�`)zA"O�Ay�(�͐Lxr�A� 0�"O8̻#��6e�m��aX����"O�i+e�τ=X�b��0s� �"O �2V�S=�����NY�L%�V"Ov6c)Mz�鄋N(&~���G�(D�+��J�p� �:�%�w�$=�v�2D� Ba��6M�V��3Fʠ#��/D��	DH�7kD�*�Ǉq*�a��,-D����HEX��ڀ�
�B	�3�=D�P�H;+���3��do��k:D�$Ӗ�D�9���a��P�(@�U 5D����,�uFB�z�aގjNd8�f%D��	W�	�m�Z�D/ʯ`,���>D�����*;�eᶏHܸ}�RM=D�ԣ�
�Y N�3"/���=1��:D� Y��ɊNJ��@�;�<]���<D��:�	"?H(�p[�3Q�HG�-D���l_/X�HڢJ�7+d���$�*D�����OT����S&��l��+-D�H��I%��c0'֧E�"8��*,D�gG�a�0��t�T!g�"t�$*)D�����&��I*��E�#{� =D�� ��T�n3��;���9^ 0H/;D���͐,AP�s�`� o�����7D�PA��'�f��R��7����3G4D����fH��y�韫��[5�3D�(�����GW�TR��	[Øɳ!�#D�\�"��Ԓ��_�69�	X �>mn!�$Ļ޲i�@�!`.<Q �J� 3_!�@ �2y��m�/:u�D�R�&�!��Y Cc�hla���@"OT5�B�#����FBJ�l��"Oҽ�CΩ�de��
�<u��"O~�3ODad���D�_]P��"O��3��o�V͢�dC�X1Aj�"O$|�f-�-��Pr#V>3x�z�"O(�����FM*�,�*��	�"OL苠��$a�ƽk��A�j/
8�"O`5j7a�<� �q�� :�Z�"OpPA��lX͸�i��~#ޘ�"O��*a�aP�	�ŝr��e(R"OĴ�%ߊ3^�@�锬=��=k�"O"��Ǧд>"�:3��mi����"O�!R�(�;?]D����:h�9Ѓ"Oj��`�L��懞UHbŉp"OL�(&�.?�:R��>L�"O��*Ѯ�/x�"r%6U��$Q"O�  A`\�c� P��X�g����7"O�}�E����HI���	)vt[2"O���aÁ�uH�%\)_w8p3"O��҄%!wа���20e�` "O� ��p��&{�<"�41F��r3"O ���ɝ��L�� ��7_9P)[ "O��i$A�X����Ğ	Xz8+�"OJ�ÒǬ[x^��"�B Z�+�'�h�Ԡ[a� A���ӕq}\�X�'���@���5r� }��]/h���p�'�0M�S1=��4j���a��'
NP9�향yp����<cؔ��'RD�baB;�X��!�
3Z��'9��P�+��X����Ǟ2�X�(�hO?�I-G�.=)&kP�^�v8�@���'�lC�� -�@=��`Y���Z@�®XRC�ɌfmH�I7H
�4����q��Zl�C�ɛB_2���+P�C-0t��^h�O���I�73f%� h
4^�%�b�;(���ß�i��
!
�\�H햭'^:����+D���E���6NVM��d�C��9�R�(�d�OX�~D�����(�C�˓M���1��=(⊸+�O`xq�h�';,|�S
�<~c��r�G쓄p=i��»$��h�� $���@�QE�<�F׉e�!M#�� ���J�<1&��!��kAՅ:���K�EC�'q��E�tF��H��\���On신E���y�oĳRv���~���I�#]��M�U�N����<�|&�d���R�K�e0!bRJ����$ D�D�$'��XBR�b�+�'���c�Ŀ>����D(�S���Y�l-�  ����5���Q*�y�?i��Dy�!Z����c��?�y��:VL�s3½P�B���*�1�yd�*|���C$ �C"E��aЍ�y��T�{�|�C�n]�)�f��f̤�'�ў &� C�ǡG�d$k�KSиj��7D��2�N�ft�bʉ���xX`�5�IU���O6NP(֋�*r�$�����()��:�'*�LX�eG�@)A��3� )����;<O ��LQ���aۻ3{X�Kt�|R�)�ӝvm�Y�d� �(\�P��S��B�	9R�8$۠��G�ZA��U��C�	��Lٙ���  B��uE�>$C�	�m�L#� ҙ%�Z���H!88
z��$6�S�`޲_
�P�O�|�`,.�f�b�T��O|uY��`���2� >�F�p�ϗJ�����=C�>�k��0��c����p?)�O�q���	�KB�bŃ^�f$�Й"O}�ՏF,P�C�X �`�Ȓ��{�O���)VGR1?���'��Gܺa�
�'}����!w$ �(WnJ�?���N�XG{��4J�z��5h3��k� Q���y�@A(O<t��i2_��A.!��5��
���(�A���TSA�D�	rz���IS�'�`M�@��5��ճ%��+
C��#�'+�Y���V<{�f}U��.��X
�',�{Gc*v��3Ԧ%ph�I�	�'�����Mذh�N�5fx��b	�'���I�/T'L�&ɢV�A�d�&8��'<�M�1$ԥUeB�e��\�����8D�xs3cŒO.��q3
�/-�2mД;ړ�~�/ʓ!�i���VY`e;�c��Us�Ɇȓb���#4ٮ��󤩙�7�\�O�=���cQ-�|��fn���jOm�<	o/���+���2Ж`BP~b�|���+4T���q��~n���G B�"B�P�<�gG�-bЕej�,rQ��鉢Bs~  V�������b��C�)� ���G�v̆I�eOU�q���4?O0��Ė�����ٖT�L�-�<��ɾ�HO�<�
�~񩖤��W��3s-Kp�<Q�M<?6.a3�I�o�XH+v%��<��� �Ԣ<1���8&2��E� � ���eA��y�N�>���(Д ��:�m��y����MX�J�瓉ACT��dC��y�����C4k�?<q�}�J
��y��}kt4�"d��8����O��y��MJ}(��7�����D܁�yb%�7u��ϟ,A�
��� �S�O�Ҩ14��7$DI*�$R�@R	�'�z��l� �z���εc
 K۴�Px�ތ(� �ÅB���J$�w����y�i[�4��݆ ��+��U��y�i��p�i���0G��]����~B�'�b� ^�54�s��Y� ��
��ē=\�c!��$a��$���� ����Qh��0H�*�z�.Q(��ȓ{���G��h�8@��J��j-�ȓZL��� xw0Y*�"�\oZQ��sב>�F*��DF�����s�œ�{¨�ȓA"�@:���5n���A��@[�`oZ@(<�ʝVy���!_(�$��s�<���N6$��Ub��AXgd�n�<y�Y�#%�����#VJ&]��.�p̓�hO1�|��W���a�!
eJ�"b tZ�"O~�c�E���
�tOf`+'O&u���q�Z��S,Q�i���8r�+$�d���1��[���%F3���O�*�y�ƀS%�� v�J�l�&C��y���w;�Li �N��ĉ&��'�y�C�Bz�����<R>~��F�ɴ�yB"�3-J��K�d��B?��� � 4�y�ȷc������ H�hD����0>�7+�G�e�`�ջ��#A�]W����'���EG�id��� 	�k1�0�'�ބs7��;]VL���o@찌�6��
���!͇[�jA�#V�����	g������Q �Q�q�����*�� ���r��hG{��	��/j4�V�ݶ)>e���Z!��3q2#p �:w�
W_&����dH�v���G �u���!�ʊ�^��~P�PԢ�$L�M�`+g8�pq(�<i��哷3*�1s�Oל7^�`5�E<l �C�	4L�Hl	�KҤ7%!��IISnt7�(�	B}��L�$�P��<�e�a�/�Q��4?ُy��ӆVx �r� �Gf�Ŋ�.��p?�0��7>?�hq�ѩj�$��#o�c?���)ڧz˦	�@I�Tꩩ׭�/(T��ȓ�H��#˛_�>��
���եO�Q��'}9@���[�d�28q�ǌ/,r�?	�������!����P�՚Y���'Ѡ09w��_*h\�P��7Q�>���'���{��ВK�,P��)�v:(%�'"F�h�J����0"��A���9�"p"EQ+�e�#FC���sV�'��Ɋ=z��{�JO( _���b���?�:B�I*mkv��w C6"0��h���2B��	m¡��e�D41�B�!W��C�I�46�8�	��k�J���k��B�����! U5Os��7�.eF{��9O�iAo�0�6Գf�f�i�%"O��*sk�5 א�;GC��#�v� %�in��)� �`�rÐ�\-���"�q� �0"O�M#h��EV��cĂZ�2��3��'���t(�a�w
	2"L�id!���!�$� d��m�������)4}�Ȩ��)�� �'l�[gM2Q�>  ���Z�<Q�m�5̐P7B],&��K���<!Pê�H$��F�Ĥ��Yt���#Q�Rͨ���y��
��QZ��I.x�:��G���,�S�O$ *^�g��r�l�= �R
�'��3�G�9t@��g�`�
�'{���&��@:a�a��\VNM�	�'�{��@�"���0o�*%����'��p@塞�:�n���D�)vqP�'&��@����y��4�*�'��u"�c5d�dD�ƃ)��Lq�'+`�1�O��)�)��C�6+�	�	�'��I��܏-Z�c�P�y��� 	�'?��#΅�_��c$�`�NUP�'��2q)�*o���i��@�XDL���& ���Y���:qg�i��\�ȓZY ����������Y����$_Hɺ�I>���a�;Z@��d�����*�����ڂ��hj�|3!��+=l��֋xt���:d��ХS�n�@h䂌/m�V���'��qX�G�
kf��-4q���y��f,K�s��`�InD!�ȓs��
�N�=%jjuq��J$�؇ȓ�rȨ�@�{R&9i�%N	N�
���Iu����oޠ]i�<�+I�p�N1�ȓrhި�#�X�x4 ���+���b�@ ��dJL�$_;$�ц�
���/L�XKn]��/�5$�X̆�v���D�I���W@ǩ���ȓ1]���P�
 ږ�
 �%mz�ȓ4���a�i����㕦U�p��ȓNF�1�DL֧M��@�%G�J���J0�}AC�;[���ࠁޤ3$�4�ȓ|�Ӄӌ��m�ծ[�'�rć�T�,�p����#�^�ɀ�	;�4��ȓCل���쀄>�<��O �G�TD��i�`LҐm@�i�,䠷͎�V�l��gO��v�;y\�!T�ы1��)�ȓ6� ��d��5`������*����*L� \ �FΏ`��I��L�;��oj� C*B���"5�-L�k�h��t-�B�.�v�Ф�$eC��@f߬v��C�ɔ��U�iԶcX9@�>��ȓy���;2���x8��$ҵr5�H�ȓ5&~�[���2b
L`qj7!��ȓ	�D�#t�Y�Z� �V"��ȓqW�ȡQ"�I��1���A�%��1��rH��@�
�/���4�O�~4�ȓ0�>�Z5E�7�����7\��,�ȓt�Q0r��
[I��� ��	����ȓ-��}Q�c�2�^�0&�S ~��ȓ!�ʬ�2-�.���6΁�&���ȓe�Й�V��$ox������	ె�H`�A%MWg�l��˂o�&U�ȓS�z�j�Dé�츛bME�
j��ȓs�@ᶊ�0}.���Y5X���ȓ ��Yʧ�M�+�v}�I�%>���ȓM���3p/��TɊ���A���-�ȓO@��cŏ��JpRd�Y�n$����S�? � �IF�	5��`ӫP<���"O<10���&
B�`�j�- R��v"O$(�A	�,[�� ��/"(d$9�"O�2G`��R��u�_�#\��a"O�,Ӡ��"����$�K�B��M�T"O�H�BVqgH4�'G¤����`"O���5�̀l�Ry��B"O�yQMBp��;��X�%fHh�"O�0��ˎn��0���w�u�$"O����Rp���i  M
Z0 �Q"O�@���ٞ�ح�Av�x.��'����m	�Q�l�?Xa&���雼T������l��*�."|��Ђ������ri%D�,�o1X "��R���A#"������c�$�ːIȃkX�|�q"O���V�y*��r�� &�d�V^��G{��[%!��ѥ׉T��C�ݶP�!�D�}��iq���s��h�%
5։'��|R�U�-�+ "tj��	!�8Lp��~�j)'��Gc��s̍�ae��y��M)t�T�Hs���b1:�Q�?k�ؘb���������8]�őV'��f��1q�ݼ�y�����ee��X�l���)�%�yR����'� ���љ^��<�0�4v�Ѹߓ��`���x�$6��*�\Ȃ#D�=� zQ���K�!�dׂ^S���fiѠK��M��R�\�O�LZdb
,��P1��	U���a�`(��\�'�[-�!��	Br�X�i�}�x�b�A${�r��d��X]�O��}��P�0��zC&0K�D�SGF��ȓf�,��e��9�&%c�"Î��0��xZ�E�s���u/a{���eL]�d��L�xr�)���=��I%"�6����c�<��BQ
nKD`;�gX5F�4"O��(���361�ٔe½<��@
��DP�K���!�A��H��,{�#����1�B���|yr�"ON�r��GR��y���q�lQ)��*e�x�E�=��s�81�%��R��PPB�H s�bM(�>D��F-��&ДT��Ȇ]�F�� <D�|�0+�*-��p��B��x�<�$,	�L��@h`܊X'��b�C�<����*8"F�K�o�XI���EB�<��J�N^��{�Ɛ$\�%cG}�<�Ď_�.K8��v�+� 0"W\�<ɵf�|�X ��D��L�F�_�<�qȌ �y@�.YqT��SA�<�����PP���%�R��1��x�<����1m݄��6M��g�a`J�R�<�'�+�L<Z"��QX�R�<��.^k�-�-݃q��M�IL�<�AF�?��X㠂A�{�v�!��O�<�bd�I�* ydܜ!Z����B�<�ǉ�*}b^1S獞5X�ܹQ+B�<��KW5.D|��#��J��y���<�P��4�Ը���+����q�y�<y#�FDz�Q�y��0�$\�<Q��U�p����6�3_�V�a�ςF�<isl�|�.��`"!�>�Ya �i�'����w��h?�ՁO
�L�1~V���C	%���ZW`�U+�B�I#
0��tMڲJ��Tj�BM��I�LӮ9�dj埄9���!4�F����ڎmZ��T24�������yW�z��L�e�Q	 ����9H�OW�z��i���L��(��	{�}"B�X� ��l�-!j:\��  ���>���`3P`�sk�/a��pɒ�*B@ �  �cI��2�M��(���@��`؞<��@��bn���wOF	` *�#&�S3
v ;�&�>���N�b�a,*��ū!☊������f�m�rbأ9�(�`۬9���x�/D�� �0∓"|�����솃:�2�;����"�8!�g�Νz�l(�i��6��{S#~�����l��i����`͏S�Z����9<����ϓS�P�����>���҃�R$
�m"`�� k�(	�N�@�Xpc�\$J$�6��h�D8��򉚱��'!~\pT�E�r�xԒ��t�x�J>����q�l�!��FBmT$;/�օ�Ɋ�
����?�xD��+��e��˔(��e�C �D�����^�TJ �H�"Q��-^����!�����1�4�r����\���ّ�K����4k�g�����_k�ڷ\�4h16�^.���@�jy����.\2��6��L�zE��AQ�O�ڭ�����kY�,�D�}����ܨ<6���eK�O�by�g����Z�H����器Ij�� �@[2C����_�.�NQ3N:݆)��e��Ql4!�Ęg��5`�旍ɸ�8'��QI��`�̜`f�h�,[�`v�Ss�'���$+
�Bp�n	pT��OB��$��(����19ʒ<CeQ>A@�������@����'�9I0`���Ԍ�6�PDjH���>��KY�z~�q�o�:_	���t���y)��D�B���@X�KNՠ���}r�a���[����4�y�[Q��`���v���������?i�%�U���$��X�$�eo%Z���@a��K�<x赫^�X�aO����\�0�%/Ke�I�9|U�ƏQ�:�� ���8/џX(�=C��軳`A$��v�� �(��T?W+��tMX,q�5�G� <J牡HՀ͢ �i����'eX�`�ш:�R�J6��(8
��(O��b�*X�H��H�4\ c"ή��OWҙb�`�� �H`�'�6 ����'��
�fm����G�bO,��Q0
�ff�)�zl8�$°=OQS�1>J�'�@�	��3;�v	�4�Xm�8y`��v�J�I�J��\&�P�A�N7���@�� g�`ZR�K����!S� O���TȂ��d��:J���T��3QtZ=KBcɐ O�4y�B�e+c�f����+����|K3��iB�I�2�	�)�l�n�C冚�oV�:ۘ�p�7	�*��� � �$i��m9� ]�-kr�B�8�~8h2F�>a��B��#B`�i҇懟J��ĺ�) k*D TY&|i~���)�-x�j�֢$��z��x����4b@Ux�ɒ�P��I�\�] �^��m@���i,���O��`M�1��Y��?9�F���<	��:Xt���I�Y�E�\rX��0!gS�19�q�T[�d�C�G�h�܀�F���e �L0D����$E<N*ՀP)X�E���q�%�	G���a��)_�V�v`���[.KQ�@�l�bv!�d 9�:H7���u4Ā�q*�?7�!��ַ3Pf���oD	Fh�:둞�IW�[)��>!��,�|����f�"9�#,D��%cP#�,9[1�ƌ9�62ԅ��X0!�AO3��S��?�E��m2�)�!�ص9��xQ�Si�<�saĞc�R�;�ȷ9�y�'!��<16�U8 ��d��@<\OX��3�ǟb�d� W*�%s�X-���'s$�g*��*f��lR�<9E���U�,���(�yBj�	#H��k��\j5ӯH7�O���Ճ<H����iY�~[�� ��B���M0�K�5*!�T(D�h<iA��g/`	�j�:T.L�zt�nv�iN�"~�Mn�� ƮO�_# ,��椇ȓD� I�#M�/D���0�'|[��ϓ8�*�"Di�	F,����<`����H�-�0�Q�]�?fa|�Ɍ���q�鞰F�>��c�Z;'����k]UX ��
�'n,3Ԁ:�����r�y҉��@�M<8�`Rƚ(�(�n�k1�܀�F@+2-ڠ���� "O��:$�����p��͈�:���ɭBv�$A�
HK�)���u��h�L}G_�BD��)D�dx��6�"�z�a�3cB�[s��>�5�U;�j���΁6��DqQ�ʳM�(�u@[d!�R�X�Xi��� 9l\�`.�a|!�Z����tEđ!I�F#�!�>.K"MX¢��]��X��O�M��D"�S�O��qJ���t��@�j�X
�'�8��(�g���"��ј>�L�R4�<��'|�����~�?�gR�`����@�^�	��U\���z��H�,IJ�W�V�<�� �=����CF�%&�x}`��Z|�يP�&�`�!M�F)��D}ҧ|��黠��o4��+ʟ��a�� �[s0����lH�l�T�'��ic�D��"������
T'[]�I�BKƭ[f"����M����6+�p��%f"�� �(a���;.Ox�(��W�p�B���׹r�H�:�'��M{祉/G�c>���i��d�%��jY8	��G#�<��I��M���(x8����'PL %DK�8@����ώJ℉w%�SD���d����h�����O��		�4��E�9]è;d�	�0�|��6 ©XH���'Zp+!��?x��ӆ�Ͳ<�|l14oŶ�\��w �;o��8��+@�Rh�ɽ ���f�L2=���#U�z�X��n����D�ɇV�����\�mʊ���
HU��-b�?�(q�t��'4z!ć� �!�sK��?Q�`Dv�,R��0}���	!Fk��!�ޓ�21ҷA�����<�G�]��Nr�f�+����h3��
Z��� rh�^�)�V�Aec2����>Y��-���>�O]Ѱ��V;�����
s��!؆D�G�4I�c@���`�]�hD񟴵{�'��[�A�w�ډ�E(_��TX�GN�=g�=`��'݈X���ڴ+攑ZE�� �՘�׸e��N��W����^��@��v�@��'� ��H�aZ���K�c�f`c���?��y��`�h|[^���IȎeP�������F�ߠP�EB�� �+�X���I��e��5@t>�P�D9:!~c��@��E�8$t% PI޶��D;$GӋ��'���E��pb���Se���`��2Jި@�F�7�j�0t��(�R�1��
@��&R���A!eՊ�(��I1f?��%y����.���R�'o�d�G@EX�<��0f�.-Tm��{��ŗ�2܇ቝI�z1�cP�L��r�mI4m��C��-W`D]tJ\�$&X,dJ�C�I�j2�X����1�PL�t�RʤC��?3�r��L�B,��ϒ1/��B䉨C���� .�%�7GE"#ٲB�	b�z� 1&~W�0���&Q6$B�I49�j��S�R�2�YR��éN fB�I���h�˳8��)��G�!^^B�ɔmښ�%O͐vv�I:���3�@C�	.<G؁"&�J�b]��bT�[�*C䉜H*���&Ⱦy<�1FF!*TC��]P�͐�ߢHw��8�*C�ɡ9����oK8͂,��
D��vC�Icd�\�S�O.?~��a ~^C�	_�̵�#ALZ�4T��Şc
C䉏n�x��L8�R��2'A�L��B䉔|�R|��/��$مB�C���D�? �|p�y"O�y&)6��/S@m J���yšeQR�%`	nz�@p��L��y�n�V��)��S�?f�pY�-P��y�O�:][��3�!^�����C��yB���YƖ ��c�8J�f��a�<�y�ʭT�f���F�|y�q���y£S�s�ԙ@��8t�9��y��xs|җ�i=�" kY��y������q�S:X��09��T�y��ʵ��L��Z�_
��@PH��yr��z��r��7Oü�`��X�PyR��5s�P��󄎴B�p��E�<a�%�-(�|ݠ�Ŏ
���9��t�<���äJ9N�&�W�ER�Dq2"�Z�<�2+g�$�5��=7�p�2��L�<�m̙FFpm��g��80D�I�<1��ih>8Y4ǘ0/����rbO�<)d��-WW��zP��]�`a:#O�O�<I#�p
��[e%�'T2��Gna�<ɄHЗ6����dޖX4�Ap�<�jKNsR�yg�ɛKU0��R#o�<��HB6�LK�hǜxm�1�",�j�<)u H8>���¬�N:	�6�f�<����&6è	9r	�BtA9�G]�<�j%&î�qCfA� ��%�� 
@�<	3nŻD�6ة���v��<���H�<��r�J�Z��K Đ#)D�<鑣�Ff��S�V5Lh���@�DN�<� ���0KC |F8x:���94w���"O�����]�fb�dT�U��h�"O��)S�"U��a
bY���s"O�����v�VL �0��z�"O��s�Ўgwb1a��W�Ī8�"O*�E���"D+T,`(��rO���yr��&U���j⦚�K��)���yR�Y�fa�	���A��2�l��y�ˈ6�&-�ѯ��8��d��yBe4���0�W9, ��P-�yR��`���;�cC<7�6�C�̝��y�LD7�Uæ��ϼ�y�( �y'=64p8�ە<9�@C��yR��v�R��WB�5fJ!�a�@��yKǤK�$� j�6�Z�	�b��y�o�%N0}y%"��L�k��A��y�(�d�vۙj^n��nO�ylj����
*g}���ТY:�y2�Xr��W�)P�nm!^1��C��*V�����dp�3���D��C��P��q���1D
N	Cg�-l	�C�ɄX=x	�!��q�"Y0�&A0C�zC�[0lD;��_�i�(ZWn���`C�	 -���22�,1����C�:v�V�aE΢'7��bE�'Do��s��E(U��"~��*uP��iU�B	�!z�K�,;(C��0a�]b�m@
&�.(���j9��I���X�MBA��ĉ�B�P|�ʓ @Y���P�";|O���Ɉ�P �љݴ5�:s�T�q<�̃��v$��ȓx��3��6F���g��20�?)���A�S�(�'$������Y;�WԽa\��Iq"O8�� ˘�)�P��b4�p��i���5�b��I��3�g?!�˘Ob4!G(�X�.�R��e�<v��WP,օNrj\`�W��㟰@�E �bV���'�>1k��վ:��9��b�D����pE)5�87�� aFx��0+xZ�k�%Ax!�D��i��a��A� mh)So��~��{v蔑w.�|�"}zU�Hd�i��Z����4jy�<����".�Ҁc���v�	wnԞ4 ���8��S��y"��A���`�^�Q��P�s�Ԡ�y�oτ�,E�U�~8=d��yR#S���Ap���=,�5���˓�yj�+�Lت�ɔ��<�5��y�^�/nu���
�|Xe W��y2�J*m��!ƨ�'�V��DC��y�d�Aй�U�pU�a+��R��yrb���-r@"	��m��yr��D���ሸn �@C�+H%�y��	�  ��.X�t�X�e��y�-�7{*8a�(/]���e	I��y�߃,�6���ݺx����!���y"i�+Ah4)�̍�-���CcL��y$�������^�	+(��s#Ɔ�y��N'XFdbFg��Ȳs�Ÿ�yb��E�%"�B�)+��ɳb����y�'8���Ӣ���$�BM1BM�1�y��ɧA�Z؄g��di��	M��y��?D���7#�-�8�
����yR�J�]Vj�@�,֍ ��
D��$�y2'�6<ك�����-i�ǖ0��O��q�#��~R/�<��m�'�FP��0.�&�����v����ȓ ��U� *^צ䪷#��k�T��^���%��.�?��͕"����/.>pڂ�*�����#���!�A$E"�yU�[�^��,�"H�eLPbTB_&S��u�eH*$��I�T>����� �H�t�>8W�X ��P��a e�'��y@��H� �p�)d�f�9���Bx��9d�R1�
�v/�G
���	�I;��X2��}J�P��SK��9��c�$���/O.QꗀR+&�䊓�-��m��e�'|	"���j4�&O8 h�%(�/��[��C�	:`�&bG�4��AX����Z����R!w~x}��_�'���L�9g�"ZG46��QH�?YZя�3It8Y���zV��Bx�I��5yZ�;��փ�8�'U�OG�!�a��A1�R1J\>xuF5���[�qB){ԣЬ��՗O
�u�>����<7���!�+`64CR�A|�I+b&���u#����ZJ����ҍ��KA�3BVe���\�7�H(���!�(i�T
�ܽ;3	�@؞�C���=w��v��%� ݘ7b�8B�6I�����b���D�z)
�{�;}��*�*�&�
՘�B ��5Ƈܝ(�t��J�v�h�)Čڂ��x2�ǂU��وѪǌ�*����p0u�^��p̐�LS	��ɱ�G�R���ء���>�рY>�[�j /˸]I�o� +	X���Cx�Ta�/�#-L	Jn��P��* �!�0�Ѷm�@3>(�@+F5q�	�JÝo�b	`��B��nH�Ov��Dn��T�Z8���WO�PCD-���TG�� Ä�,L��HxE�|���0�0�+3�I�9Xt�Q&��"�C�?<������d�}B��_
�!���ΟC��xP��*�� ޣjI���W���b�!\�9���N�A��x��y�o�`vp�!�2"��-�7Nر�y�B�1��}x�,Q�k��x��̳(0 0#��t�A�6� H�d޻�1�$M6�������X�r�&͈Uh��]F�z���H1f�C*_ɛ֪�%4�L�GJ:{��!bD��&���u�mS��'3 	��2UƠQ$�3*��k�'4 �B�/πc�F ��5-�ɉ�'�$a�rMәy[eB3LQ6P@�'u�@ӥ��2ѱ��\��-�'�9����]�NU���Waxb�'XL�"���0A�������Os�'��z��� �H���B7�P8
�'2�e[EaQ�bê��#�]j���0	�'hx��qiS�!@.�Ct��0K"��	�'x���6�.|�*�9���~u.(�'�`��F�N&	N��H��]
9*&LQ�'N�_[j��i���0ڌ �'�0����,�|zq	���"O��p&:D�J$�R��5�1"O��Qc`ƳZ`��c����(�P�"O �U�$*\n ��@^��� u"O^���G���H��e�Q��	)�"O��E��3�
 �e�Q�s��t���ɕ-��2S��M��E�'�8�P��#]��B�	�IH4��ևӬ��*��y	l ���S�lx0��I>E��&�Y���ʭ*j�34@ˣ:����w& �@D�6w������֠T+�̓D�fxKwJ��yHn���� l��DO�N@�B�茟K�a|"�@m�t��-��S�e��$�e���K�j�	�'�`�y�#�&���9@U+$<,*����F��hSb�(�*��VO�/:�Z)q�@J_�PBs"O8��!��H�^��Ӏ��O�hX8 �ӠZ��Tŋ��)��<0�Еw�Ttk���<�Msf��`�<�Ռ�WN�ţ��M kT����
��<a��>D�,�E,\O(�I�ۄ,]��P/�p ��'��`9ł�;��j�iK�\F�3�)W��а�e���y"c!l8%2���+��0󵫓W�'���W��e����vJa��g��/��Q���^C�ɩ9^0��G��%z�ˑmS�HΞ��Å�:{a���I>E���O	����G�A��5�$�#5�T��
���"���#z�̄ �g��  ��'\�#FfDI����`�ҭWT-xb�E�VJ<u)%D���	�-��COU�=��ƅ%D�L;0MD1�6��Ǐx|0 6D�t����l��m냡���6�J��"D��bG.g�`x�	])C�:PQ�>D��3�gM�YI�p�`-$P�l��(Y��'�ui���>�#���s�����'��<�\X��mH<9B� pH����/7�\�T%��Ӧ��a�ǥ��z�g[�Ѣ+V�k$��!DA0AC ���ɮY`.�������ɢ'Ȱe3�,��Xz��%�J�����_>|dP%�>ق)�2
�T�ѓ �<HX�SJ�m�d9A;l���g�5�0|Zv�3zr@��� c�l@�q��o̓c�dT�!ۮge�6m�5�8
��T��"u��X��mR*;�HY�J��_8BO���rj�	9q��'�~�Q�f�:0�j�!���WELYaםvo��薘 ��ce$A��O���I�:��� /j��*ܐpu��*qN��v%�X��''�qd��q �Y��q�K��&D�����w�n� a瞺w��i�ɀ|����t����ԅiC�,9,`�4LV ;���Q�34P���ע8��(��L� m���LW8tb�CW�2ߎ`���з�?�4EC%30`���(}��D�ǲ��5���A�i�T��	����h�|�d�[�Gnp8�a��!�ܣ֎(�b�$�?F!:p��Ù"r$��$��1���3D�DVa�g�	�>_�-� ��K�<u�q�W��2A�3Y��̀�M�4�r���2��/P �ċ16F(g[?fN�	rg��&=�8P�8���{�&U5v��\��Ћ@�ZXr��\
YkF}3gO�$:t �h4/�t���9z@"ٱ�x�(�"d��aoW:� �I@���<A�׻� +����b�N����9��zrjT!�1� &;Q̩��!�O�� T�ĝ��)���@�v����$B�|�����BTHș_�Y�$M%>��T�פWSl�v�V.P��P�s�=D���1 �>B�,{!��Y�Ӧ��(����4e-�`�`k��c�P�D�,O �+'���J@x��hQ"t�0�"O.�B���r���0Ӈ�,羱c��d�r��9��&P-J��?3&b�"I^�E�>��ȓH�4��"�Д���hv��0g��$��"��x%B�w��@��L����q4j�pv��*��V�܁<lX���<�XD��#R����(L%I+N�ȓ,"ƭ�$��r��t��"C���ȓt� }QF끴
�u9C�dZ���Oz����ɝy�F��B�'��t��u�f���, ���% B&c�~�ȓ	�j$�A���d�^��(�`��}��yLF����?V�Mٖ�f���kNn�����`�����\�Y�ȓ@�L$�b���p���7�țjb$��ȓ\�H�j�$OLf8�AL��$TՆ�$��	�(�wr:	���q D��A)*U��H�[��[��eꎑ��5}��Hr�|Sp��n�y ]��'ؾ�ɃMs��5j�fвp�*���'�<�s� �-G(*0�i��A8�'J��3Ԅ[�'l��Ȁo�>��I!�'ǜ,*Vș5��C��-G�*�'�>@�ע���r#G�
 c8���'7�X�*>��WE�ȍ3�'�����$E.�i�d�����	�'�r�(&O5I=���iW���,��'�`mB��i���D.�BT�'R����lL��^yIfOG�{)��Y	�'a0��
�xժ"�q���'A	��H̘<in���IJ�t�>�DP|�ڰ�c&�,��\8��� O�\�\�b�<R7�����uV�-����_{?��Ō,{��hA���8���������@-4�#�� G�����]h����^y?�ç<�84��9ِ-���v�h@���C����=O�,a����L�f�VH{��o�^5��bF��j�j!��'��K�物*ga�H6�Dp&�M����(�eё�F4i�kT�g���b_��T]>��K >J�OJ3G2�2B*ʭpN�'�4`@u�T�S�'/4�wm;6���v�,�-�'B�#=E����"{gX������M��'�S[f6�L�<��{���O��Wp��� 	T�l�� AWO?z&���;	�'N�`�(vJ\�����׍�	 dp���,6���� erɆ� LFP�IP��2���D�dO`aR��EI�S�'�֙Z� �v�-2��ޯF��|�'8���H1�)�g�? ΅À,¨��!��M��=��nZ�dD���}�����C��۲Unp���2���w�����'��4
ç"��	�u��?t^B�Z��%C�Xm�'���ّJ�ɧ���V 	�[�Z���I��bV�	�1O�6mr�6-&�$�d��'R�r�{UH[:jx�;����I^�yn.�mCW��|iϟ�Ope�r�T
e�)��㙠P�XC�#�/vL� ���V$j�Mй�2�01j#��㟨hp��v>M�F���k@��PA��V*0�CE>��2V("<ͧfx�I[�ʜ0§V߼L�s���p����}���54M��`�dGY�P ���5>�~�	�fL$�y�}��	H�L��ra���tE� Vg�8'� ��dl?!�O�O��%?���V74n����F�xg��baD/�y�&��I�b��g��WB�Z���S��7>I�i���.�qC`��<.x�y��'-ZA#�(�oQ�Q`E=~��<�	�'�	ە-�L�n<���>u���	�'&b�Ó��<A�s˗�a��-		�'�8�T�C��`1 G,I�T�F�@�''��!cǰ2,�(����[P��p�'���dF71�a
4�S�c��q�'����	i��X�嗨[� aS�'$\��ƾ!�aY&#��S!��*�'�1��B�G��@��bJ�E,f5j
�'0��ُ_����F̉<
ޱ��'�N�KD�"��]�F/5�|iA�'@R�bb���%�l���=>����	�'�<Iه&�t��)���J!�-;�'��I�䉱* hY��E�!?Z���'�� KV��<m�u�'KL��!
�'�ʬ��� �h�R@)��O�A�	�'p$)�!���Ό#���W�<���'>�Q:��P, ЉP��N.�ɰ����oMp��c�)t�<�C!�g�<9���"X�ڤP�٨gHp��Wjb�<�a�) 3��Bj� Oؔ�����_�<)w���xQr'�V�$(�;�-Gw�<1%]�f5���폽ly��:�lQu�<��mO��9Y�bݲ@����p�<�Ԁ �xh|�vï!�`u�G�c�<A�M=�
Lz�CQ7!W�}!�'`�<��Eŕ#��Y	��{�H�w!v�<QEÉ�HM��xxaW��w�<�A 01�r%M
�)���1�w�<�C@�iw\q��$�
aHB� e��w�<Q7)�"����ԃo5�`XDG�v�<��W,�څб�)���zq\p�<�6;�<����n���2%�o�<�#"��"x���Ğ�h��U����k�<�$�f����G0Az@ʠ'�j�<A��Aqh�"D琬.�t�A��}�<��#N:W�:,`��������;�y��X� �ڝB�a2X�xň����y� ��p+�/[�\m�e�0�yb�މW��|C�!�N^��p���ybiM ��{�f��OTP
 C��y"w�Tm7m�r,��G'��yrIB�zs�i��OI��Ț�q=C�	��h�WO
��UI$9GjC�I�q/��eR��5�@�B�|�ZC䉳hO$����B
Ȱs�L���>D��s���=�z��/G)\�`%�:D�H��Y�nZ�����ɺ6p5�c7D��q1�X���Z�e	,����(D�D�c��O���4MF�.�����%D����GG�F;���'䂬~��#a( D�� �HX���s��B1A�6"uh	��"Ǫ�
�#p�2����1�D"O`I�sWz�����"ֺ�s"O�9�T鎶pd�i��/�tՊ$""O0]CǮ��hV�}b����nPy�"Oڹ�Ԗ~�-[ -�C �	�"O�4��Ȝ/w���:f�S F4��%"O��D��3p�pQEK�"�$�"O�T�c��E��X2�*[%v�5�"O���!!�
Ϟ1��Ǔ*O� �6"OR�2���4R �x╌�"`W��� "O�dZ�c�2S�L�9�˗%\H��;�"O�D*��;kP<���i�2AvD�"Op�"��L���d����(62�:p"OnՉ$J2wԱ�'�.2F��"O�+�,�>O^����$$S'���"O~��U�
e˚��䴊��W�y��.���p�\Iɘ��D��y2��4��hB烑X�l�H��L�y�iY7���%�9A�H�E��y��K (�D��&�4Vܱ��H=�yb��Lcl�4�U5Pt0���yr�@5<�v��7He�``[炆8�y�C�C'�)�W��4d��ӁeS�y�Ã�mB���
�[�ґ!��Џ�y�E��2]Dp���L�A��.���y��=�2!
&�,Aތ"D��y���=e�ɑ��:p��2�:�yB���F ��I�B�NԈ��ݫdH!�d��"�(����g�VQY���Z!������f.U� �PS��
k!��5mYh���Ŗ�襂R�Wq�!�[;J��"c��^����#�!��B�A��(p�G�%Ѭ]�$ʥkm!�$M+��,Y�F�xel��f�;S�!���Bi��M�$ >��P��	[�!�Xd̐�ʮ;=`� ah~�!�$�Z��ic�	�j�53�C�z!�ڢ*D��A�i;���.i>!�$	�d
 �/2Wt`����4)!�Ǹq�B���b{�iY_���
�'�d;�i�Mv�q�-��O:��s�'�8A����,������;EQ�I�'�B`Q�}�DP��@�>��-j	�'��X����Cn���,Ha�a��'Q2��a��ꐄ  	�F����'�`i񌚀�����$T����'V����Fn�$St�Y�B-`���'T~%I*2NM�t�#ˊ-E�� �'DT
#& �	T�6̐�Q�'.����.R2�Ԉj4�9-"�a��'2�9[T��"^K<���J+JL�
�'��퀇�U''W*��*Ŕ%4L�K
�'�^L1A��9��pzEgAԠ	�'C*��  J?>̖���)q����'��p���J��jÆ�#����'ah�Qb
9BܠB����Đ�'�\��֍�Y
�ة�h�\�B�'����cL�H�M+Rsw6���'�:��O��`�n�(EJ�{���@�'ad�3�_�v�l�3�h�p�Xy��'ڶ|#�KU<`�i���<g~(��'g�P f]��BKg���boZ(b�'I���%Ɂr����g��)��� PqgAM�5ƸٴLU�q���A"O�q0�D	�{L�k�<�pi�s"O�&ҟ#���cfj�'q#�"O�|����Re��H]�c,츣"O����V{.J�C�gʿx��d`�"Ouj��۩p���p��o�NLZe"O:�����g	��s`�H&u���3"O@�c��47Z`���ذ,	��'"Ova@.,�*���>/
ȹ$"O�C��[N��3p+�/9 ��W"Ot%Z�j؞BG,��"�ڐ�i0�"O��B��B�EP����.?q8���"O�x�u*�*��a�5��A���W"O�y�֎	-n�0�{Q-�J#.H!a"O�l�a.Dt��3Ma�$�r�"O��&ѥ8B<*ѬP%��)�T"O��J�ܞ"���
��g�\)@"OTa����ܩa��p����"O��I�F��C�P�R�N�0cPiiU"O����� {�ܼ���q���y�"O"}�ߔx@���J����"OoV°��/��"��u
�nC�~!�Dj���V	�T�b�XP�̺�!��©��j6���wu>����<�!��'Pd�x���Qv�=H$a�%W!�D
�6f��@�	�3\Y2qs =C!��̘j��Q(��(���Bԯ�>@�!��2�r\Q3g<z"�v��m!���������,8��NZԅ�kކ��Ň4fK��;wm�8����R�d�
p�S�rw2�s��E�xR�Y�ȓ���0�*�)D��T�_�U�ȓUb乊fO�\OR5���pi���ȓ	��]�dg@��F� )2��X��Qe|���b�5v�|9�P�z��ȓ'u�ۀ��"gj��*��g�p�ȓ՜���I����)<�~T�ȓ�^�ԇ"1~p��`��J���ȓf��9 �^�7�
��Pk�.M�L��&a��	�JMJ'��X�д��)L������Jţ�1'(�y�pc1D���J�q�p��c�
"<����#=D��ybD�94�u��	O�(�����7D�JB�Ɂjh"v#�6�h�Sg"D��R'�%����!CX�t��*D�@I��U�����%$�DMp���(D�B�N�2[��u*pO��9�f�qu�<D��◣9dKz��
שS�T&D�DKg�F-'.v���˃yA��r�h.D���*C���ʶ�S,�xsQ�,D�L�$��%�~鉱J8N��$��6D�Hj��U�3���'!@��U��3D����ڰoL�	��[ ޙӦ3D�,�B"Q94��I�!�-��"҇3D��hF?z�޹�UM�A�n3D� ڃ�ǁ6�̹�C���rA�a�B-D�(�-3n�x�BA)�6A�r�b��,D�H��ǅ�	�2!�ʒLp>��O,D��R�%�b4ЌP�&1	�,D��K��X+ ����!εW���*D�d����]�����N�cjr5�k&D�l�ש�_Q��`O�, Иty�L9D���EW�E�-�GZ#c�( �O*D�0ڄUj;p��n��_��)��)D�� :EI��.�~���	I�M�Č��"O��ʔ�K�[%�?c��p1"Ol4z��0�`�g -��Ŋ�"O�,���K +X���Gϵl��@҅"O��N�72��!�i��(��M:5"O�P۶�U�'��!	#4tٳ@"O���c��TH�$�q&"O����/a�>U0��[-�`("O���"��,K���/0����"On1x'�8��A���R$��HT"O2�P��Ks��M�em<DCt��g"O���g�h��x��썛@WV��"O�LIp���x�|좳˗�2�NI@�"O�ɛ7nD=KtI�?b�y�"O�%Fŏ���ɚg�-8E���"ODI"d�L0J�~���HoZ���e"O&��E�G�L� �� fsp��'"O��PD   �8�=�c��RFG��4��D�Å�(��U(1�}>���i��>��=�š��vT�i�eM�^�$ �s)Z]H!{g��_԰��I2^Q�Q"��P�```(�E�G�f`7
>K&�%ľ$���x��l��M�6 ��J�@���Z|d u#k�<��S%V�b���	���kŸ��M (@#o�.��3�j�օ�a-Đ%�8d�@�0&�L�ȓsO�e��d �Z���	f	�()�pL��D�y��q\���`��!sَ��ȓt*t��E*͏?dB��eU+}ۂI��7?4=[D���b�O��la,���]9t}��B�{�xU�M�"����4���qO��/�\�I����/�p�ȓMt3��ֱ|�F�C��� �����/L�Ha��E�	EN#��P�48� ��2PZ1���Z�*��ڳ<̄���gK�}�k��V���j"b�16i�d��G)"S��׎3W2�aP�.6��ȓg�J�S��_�Z��"'���	,P��E��U��o��NuH#�کG�ֹ�ȓy�J!j���.���;�H
=RR�0�ȓ_���c5,�5s����S�:��Ȅ�?���6`LlΠq8�ع��y�ױXG�T@����R�0C`��y򈝌��`ztA��A������� �y��5�:�K	'����FFN��y�$�?"��$�q��p�ba���Y�yݥr����I͋k��x�T����y���,���Ԯ�8`SP���,�y"������gg��FN���	�7�y"��eu���p̊3t��dn�:�yRN�"f������>Qx���FI�y"��2Ȑ��M�31��#���y���m�l���њF���1c�$�y��ӔG�ɢ'.�&"LEJSnы�y��2� ��
�����JN��y�h�y�hL`���&iN��5���yr�@@�-r�)����$P��K,�y�.�7n�m��i�ZE�u��$�yb��-r��!G�/R���2�Դ�y2��5b��`iv(ޜA�x�IBdO��yҀ��* |��(�a6�	��.�y�B�v�z��a�-���p��!�y�O�8qx�јvĄ;4`�a�n��y��ɭ`z�;���+*L#����y���hyR����t��� @L�yB΁���<���C�=ö�8��4�yR�X�@��d�̪��u{�h��y��\&]��\A%��~Wd���%9�yB�����A�� ��0�c�3�yBaX>+��p�b�x�s��yB���,|��)�ՙO�|���ݡ�y���]���B���Gi���R`��y�IM�2h(!0�<��l�5�y
� 6�j�f "����;f���"O����20.�iH�C� �xy�u"O��*�B#"�T`��d�\i�"O�����S>�p\�a��P�f"O���P��6i<�u���V*=�Є:C"O���M�W�컶�:|�t�cu"O�u��
֋L4��1��W�{��̹q"O�i��O�>��P�%��:K{�j"O���H��c.�9(�ڬ M Y�"O�aS%m[ �5��C��K6<�"O�u2�2%�A;�"R�xk�"O G�J_�Rdp��Y8"O(��k�79�EB�C
"���"O4
#J�F���ː��,>~M;v"Oj�H1�҄T�|�	�&�*M
��"OB���!Z�>�M�T�5�x|��"O��vL��]�\�s���,�nq�"O����I��S d0�bh\�t�nt3�"O�t"4�D;Py(tbɠt�pt)U"O�키c/_P\�A�O�P��`i�"OZ���恚A�~%1�Ínܜ��"Oa�&�I3+��M���ж���v"O4�B.��Ν
�V�q��T�V"O���ǟ�S¡З@��@��t�A�	P�����(j�)��R+q#R���dR�t>�B�I�v�B�-��<��ЉbԾ�D��6�*�H>E��2||9��Ӗ9���R-C�R���ȓ5�������=��i�eF����̓Y�� �s
^d��ď�	��9���Y�4����'��"a|"M�9`�P�GW�}�ΕKb�R7@�e+��>f]�9
�'R���P��.���lH�W#zD��$kJ�4;�A��(��2�#�|~�l�2Ύ�n���"OhP�6���7b~��%�@�<��"��F�m�0����)��<ycG��5���̀FT��� �PW�<�����P �+�♉���<�!i���z�j>\O�p����*yi�D� �_��Z��'�����Q b���įC�A
�t!�D�|�ʍy����y�OA1NEYCO��Z���A��O"`S �_!d>����:9�v�9%�K0.D(��17�!��,TFAXe�۲0àR�F�,�J�� �TWҸ)'�"~�I�-�m(0��8K�j����H:P����$��`�Z�(Ǡ֫^)ر��]����	gh�I����U�'n���J�NA|�	dަ8�^���� zv^=���O;�`��bC���LD���G ��	�'ڈdx�AJ5jA<\� �	�<��b�w�L�f$����+O?�˓�6D��Se��o��{��^�<���Ҏ\Z����L��:��6��Gy��R�7Bt�@�Z=ax¢�?qU�ؙ�C�1�b�������>�WG�. ��s�k
�i�lE��/~6��k�͇�q��T��'��Akb��)&0��w)�`4�������#oڂdI�
�~��c>igË=�#Hޒ;N�}_�!��c�T�Єu��QS�l������APa1�M޴w��)�'^���B(K&X�Ez*\< UƱ2�'���M.鄔��NҔa�,O��#��?gXhc�M2OR��5�[�F|��EK�(?�0���'>�$ʴ�ը^��p�Ң���p�����f�I�6hO6,,!���_��d��`)E�Ȍ��`��R���Q��N|�3��	��']���� �K[ ���X�!��R*2�'�O'�" i!	S�g���8X}>Q�7!(��S%7s�	'k��&T¹b�œ�nzB�I$]B5��֥"�`��3�R�1�`B��8i�	{`�O�d~����lN+jB䉩'81��K��asP�;B䉛I��1	A�ʋK�%b�cH��C�)� ��6�V�G"Z)P㫝+=�,�"OX(Cː27��U�Á'b4r�"O0��ٰf���*6CU�1����
O�X�ǍD�=) ��$K�!d^�p�J«�L��'}��d�X�}���;��I�OA�L�ÓK�2�S�\��]�����+��"XR�`�l�5���ȓ(�XЁ�Bs�MH��O$��'�ezD��=|��OQ>�	2-� Iꈛ%�Z7���¨*D���n)X��a�� kh�y�˚���
�"��SV�3�I Z���(ũ�4)m�P�Y�f~�����Y���zB��0^IBӣH�%�|��(��!>fc	��$��,Y�d_�%�M��(�6J�<F��]�xq�l;D�Wc�K�<���?H�Y��a�=��B�	"�\��W�S"`Q
�jR)����@����U(J�$ҧ(����)���
�& B��G�Ѱ8�ْ
�3��[C�)ǘ��ǂe��,�>yUO		�n�i*�N)�L<&&�0)2�*Ĩq�t�G��5�I���1,  e*D9�՘�#�4!���FƫR�N�Q�3O`�isX�rmn�"M�b?�hpoQQt,m��O�EB�}A�1O���3��Z}��O"��ê���K�c�80R���f�=���'rh��q�,�3�)���CS�",	�vm��C�\G4P��:�)��N�>�[�-+��K��;��h���3�6�R�'T�a��D�x��p.�i\�˓U�4�Y�`�:�ʓR���(���6Җ��u��`���ȓN_��Iw_!_Xh e��]�u%��*0n�+'�8����'��59�Jz�	��E�fB�	�P5T�!�⟼K}j3IKO�hpX%��\�$��z��~&���� ]�l;7吵`p�i#^�!�$��?���qe	�X����e*A��SQ#�?]����G�~���@\�.,A��Q�f��a��	�[H҂�Z��剶&�����(Zi��y`� �\C䉉�XX��1m��2�L�8HO|�dY�r�:��Iu
��3��Ѩ1�q1��F�o�!�(R�rT���R�� xa��Cz�2%�|rE�A��l+g&�p���#�\N�����$���[34�.E˦�Cx#@�IҌ��i�����#	�P�����?@͒�,q�`j
�'�t$����OKl����#C��ٱ	�'�JA�D甯ɾ�� {[Jh0"O����#U���8��mp\$i�!"O,�R�@-[���U�	.1�`"O�Dʖ$T���Q�ȁ�
1p�R�"O�p��o��J3V�	A�1h�&���"O��D�C��d#�C>Ap��XF"ODic畚P���f_�Vܤp�"O�ty2�ӡ�R��7��L����"O��9bI�D������G�*�Z�"O��i�B�|��� f�M�op��s"O����A=�E�	גpY�h�"O*p"�Y�>��p2�8�3"O8 1��NuT�M�A�
��x�u"OZ9�!l����0)Ǯ��k�$��"O�Mˣ��~H(dXAlč5��kD"O��KPb� �����3R��li"O�1�D�	|��k��Y���8�"O�uoK�Rnqs��9u��1"Op�!-��
*60h��cFl�F"O�a*�eY/J�F�ya��zJ:}�"OڵɷG�A� �PE **Ȉ0"O6$�Q��{��m��N�B�����"O�ň7�F�c
 q����"O�9�Sc�B8YP*��n�B-�P"O�͊���Pm�,J։N�7̂�H�˝�)[~a�V�4�b�.v��`�ɛ ��}��\>�.D%�p8���+r�d�8����!�� ����a���G�;v�n��	�8oUD@16��y�K�o^��Ʉ�c���g�?��Kk�d���.rd�G����d��	�ya��sA+	'Jj���� ����J�%�V�ʇJ��A,�=��lsR��jϮ`���]���O�5�qb�;C��]�&#�!S؊T8��D[�	��;0#ĉ�?���F�F��5�0�1Z�K��z���N8o����F����Đ�+���0?��$ ?%FA@+�d�B7"U�<H��"ե����/q/J=����>)^qR��(�n���м��-!=Q�@L�rtA:�V�<�Z ���QeY�N"�C�,ΖH;]y���U�9��=��x�Ӗ���%� L����<�� J02��Ð��#4�!��B�W��40C�)% e��iOF���� O8(�F��S�f�3U��;��8�$c��k�P��9UOB���D٣&����	�}���yrh	c�O
]��!�BEޥ�w�B!�S��6�+td��y�HX����t(�Q'��(�g΅^z����W� 5)2VU(��8��ېf^�	A�钒!FdA�	�R��Q�%�V�,)BĖ�V/��(��O_��¶�dJ�?5*���GÔc!�d��X��i�7�&(�Q���\	%��ͣU���y�m��JQ�kP�:��a�g��'*���R?Iu*@mf�}�6��B�ژQ#�d8�{C1��DD�x�9��Κj,�9�wڙh�@Љ� �訩�B�xE�����ϨO��siK8/�q����K8FL�e"O8�/#�Xт��_�(��)��*"�y�ɝ=K��9��O�h�K�`���yBF�*b�b���D9'�h�뵡)�y�iЬ|I�*�b��hBd��tE��yB��TZ�9#�#�2z+������yR���$�aV�˙t|�0��[9�yb(�-�.DYS	�-]�؄�W���y�� �G�< �F�J:C�����)\/�y�Y�a>� �&�ۇU�z��Q�y�A�;Y�*�AŌ�@8�v똾�y�"̟MQ�d�Q!� @�����9�yR�ٸ+�H+v�4C�Llru$��y�b��GĀz��FiIJ��y��@�7v$���ج��*ق�y"�V�C���a�+ܝsj�\��&�y���^��$�@H
��	�����y"H,t�NY񆌌7M������y��%
�BY��"�0@Ju��'���y2 �tY��K�D�C#��y��)'mԔ��m�9EL�Q슯�yBL¯t�� �>�h��+���y�"��P#ʱR���
~婕�N�yb��<|�i!��D�R�@�����y�	�vt��J�g�<1H�Х'���yR�F�F��m#1�� ��A�����y�`C+u�x�q��")��i3�J�y�> ��i�`�,���#gݰ�yI�&'~�=���^�sdk�+ -�yrM\��ʡc����`�ނ�y�VY\�#7H�4��8�lZ��yr�Q��\P� �����@dY��yR%��
;ƽb�_:vTR<[`iY��y����Nf4�$U�`��ja����y���@ؐd�_̠�)���y�d��BL̍R�IJU9,�� ��y� <����Ur~�k~��'�A1b�-(�A� <�"�b�'ɺ�6MO!C�XVF�%%��(�'l�q�蚎i��0��>(ͼ ��'�f�3������H1I"0t)
�'>���
�U�V��G�U
#�&��	�'F�څJȯ��D�C�V�tE
�'[ld4�%@�u���%	�'�X� ��ڜYZ���G	Јp�	�'3ց��=PY������0ʚ�H�'ul�su���PmqSlH�c=ʹ�E�>��x��{+4V���vL��P��	+@�F)ZPʓ	@=��'�jE��3� 
��'�۠B<����!b��e�$��1����z��;')>����DSaBU���xr��I���O�j��aVb���F�0%8�OZ������"C��`c�08����5�T7M:m��	:p����S��M��5����)�~U�`AߍH�L�'S�)�p)+�i\�D,�)�����p�
Ѩp�i�0�c��>!T��M>�y�M��w��q�]%n��q��Wg���O(u�T�K�W��SF�Y�֝/�D�9���bE�m���(t8�%ň�<E���Ɖ/�^�8�*
&b�~qrK�yR͕O�����T�ŧ��DP�J��m4���m��(O���!T�t���� ~�9�g�>m��#<ٷ�)�3�E�~��5�C�9S6p:��w�9R��b>ѩ�M�6v��Ņ	U���'-?9v����O>u8�fI�.`����)�)���l� ��"�>AI�"~"$E�t���ڭK���r����BSv��'�lYTL�#D$��Ӎ:\Q>�!E��- ���9ʇ/]c"�Va|��ݳ䔟;fB���K�|�(�3S�鈟�\('k�'dT�1�#��_�]�E�'�|�QfŘ:���u`�e?E����Yˎ\��+ԯJ��l�gAQSK�=��̈��@��d�F?�ᓫ_$\��GG~E*)��Гb���R�e��Z}vp�G��8!V�/���"�ԓ*(�!Ӎ�7c��9-���2��*)�����c��=9�~
����ݚQT�)��.��g�����ׯ/ܩU%ۂ�p�r�ܮ+~��
çKu$5YǮ��(j�i2k����@�DgRu�����ۖ ��1�iH�?1Q�� T����fؚHɄ\��Eŋ�HEkKj����l��L_V��A-�����e�R���f�TxdʩO
h	Yv
|X����I� �ͺé�-Ix��I��0D�8��Oԕc�L�kV��-]�|T@��/D� peO�7ֺ R�Ƃ,��I��,D�đU��Nl��§��P���;uG,D�غ3*�>,��
f��!8 ��r(D�H�Ŧ\Q�YQ7�I�A��]d('D�P[�,�<��=�䍗0"����&D�VD�>�9i�k\+�Ĩ��'�5�y�F�8du0�@2jƋ�̌�a���y��Q� ZJ���g[�a��S�����yҎ��cZ@���N�V̢�$�y�;�8a�Ш�C0>�R@c��y�� ��1Z�H�=��M�7/L��y�Z�%"l(�W�G�6�\4J���yBk��p�A/v��AN��y����~�\@���=���ܜ�y㔟���Q׃Yp��	�'߲�y�n�
8����V'�p�����y���?'<�f�U�d���Y�eƠ�yώ�m�X�ҡT��d�ʅ�y�*J,j�0���<F\$5�y���)_3�P�EZ�@��%���ɏ�y �kV�왃bϦ4������y� ͯ4e4A�'&}�``�$X3�y�Π<+2�b0dC�&\�P�t�`q��_'&�RE��'Y��Ф��'�m�ȓ9p�"��%J�с���&y荄ȓg��<)�`���)UB�&�~q�ȓ r 5�3�15����1ܢ^hr�ȓ:��ږ��h�Qb�	¡xМ�ȓ" ��O 2�$t��I���M�ȓ0�ޙ{�/]DC�xz�$�Q����ȓ[ p�憼:��YRp?�nA�ȓ``RRC:'�J(��o�J���ȓ<�|A�`%�Cﰘ�� L)�0��ȓ��H۶���6�44{5'�G{ұ��1�d���!�����g��6��ԇȓ@�|HKU�Jw�v�YWC�#@�<܆ȓR�n|8�ծn7�]	q�M���ȓs_��@�H'| Ɣ:���k��؆�S�? `�цc�R����Ӹ��{�"O��C+�}��󖬃g�}��"O�!��J�/�Ь��+�[IΘrP"O<�ieƚS�5���1�6Q�E"O����e��}�Fe�$r�4���"Oh	Č#}�9
7dڤˈ,��"O�	��	 G��҄�I�MR�"O�.)�t��3� ��T�T��yBł�Fȼ`�3̕�w<
j�Z �yB
j@,1��a�Y.��䆍%�y����3v��&Iӟnt��rN�
�y�A�!i?�h�',ȟ q�ykr����yrN^~�F��7�F&K�b���ݹ�y�(
,��������&.���yH��$���*�Iҫ5 	F)��y��/�8�I+���P�����y"��dv��pu.F�R��N��y�䏟 �h	�H�&(���p���y��F*%�L�@�S�GR�(��y��]��]�TfL|Fp�����y�k,Q�����C������y�����)�R�KKFt���ߑ�y"e��b4MC�O��;��I�C���y���@ψqn�#Rf��`�k!�ؽNԆq���z�X�Xv�O!򤅐��t���j���ȇ��:�!��&7�6�+����e�(�qć%3�!��.?�Pr2��4>{&��WBWUu!�dCl Lpw��<\��`����\c!�D�@�a9�ʏ{��D�#��3Ba!�$��MX���us��Aփ��>�!�Dʄe�������HO^BB�
9�!�D\c条фV�IKz �3N�!򄒛*�TJ�ϐt665�*J�#�!�B:B0(b7䌗V.ȭ���P�E�!�d�1"#ĭ�хR�XT]�5��*[�!�$�![�!�+́=�,�,8�!�D�NU(�	L�+`�>�f �,L�!�d
H��b�*F�l�/� N�!��JO�U��oʿ?�|D��.�>G!�DB�o�BE�G[7FFEô��=q,!�:p�:�`�%T�.�"|P���y!�K+#v�ʁ�D'f�@09b��`�!�$���8��jWz�x���͐��!�dH�>op3�ʏ�>��Lf�!�d�42Tu�6��5H'���,\0(#!�Dބa��yW��*42DK�> !�q��,�ë�!&'"ę"KU&'�!򄜾Ґ��t�0w"� s�еj�!��;��y�aD�	i� ��C�`�!�ZU�I���8Z�$�v��!��ͫ9����[�@Z���]f!��jl�Q�ɉ(�0}���C="H!�dI/iޖ��6	J�L�,i����V8!�O.���dH�3f��es�5!�D�L�
D����1���3T� $/!򄂬
6����L٪`y6 Rшˠ!!�D	�K�ʙHB��&�<���׮V!��5{��Y�2�� (�7���w!�	�)_D��F#�]�^-�&噣Rg!�R����+�:l�͉��UI!��>e��\r3K�>go�s&�Ħ6[!�L';��*�K̶3g�hHd�
zH!�9,�n}��`�KԮ�.\A!�� vM�6`�l:��'��dֈ�E"O~DWKS�m���Ud�!�H]q6"O6I����V����J�n��9{E"O�iRҍ�>�#� ���HQ"O0dZƉص^
9���ۤ��A"O>=s�0.��᥮ŕz(L8�D"OY�u�����ճsZ0 n-��"O�mp뛡SW((��>v�`4��"O�����+G"�� �b�������"O�t94h��yT��2�`*}��zg"Ofm�%iX|��E)��+�����"O�\��Жw�:q�(�.cw���"O�:B��!���у��Tj���R"O
��7�ǐ�!d$��$�� ��"O���d'~�(�X�B]*�K%"O�RP��bh��P� +F��0�"Ol�"���#S~�y��[
�z!J�"OaK1��<��ӑ.�Q�=p�"O�1���1L��xX���5W��9�"OB!�3�U#4+�����ߞ� �@6"O6xA�Q�^����&����}C�"OA�/������ �Ť~d�"O��seA^7T���w��+ԙ"O����(.�����6�t�A��'�Q��h"i$o��x�LP
g��A2�&D��R/_�d�d�#�$��6j��0�!D���)�G=�QTC��
0X	I+D�`Z c�U$(`U��:tų1*$D�,��/J
$���7�Ւ��ybC!D���G�������rl=K��2D�����C�O�vMZ<(p�`�4D��(r)+9�t����JRa+�J3D��k&Ez�����GXJ���c0D�T;!m*tj�0���աHS^ĳv�/D�\Ju倂WF:D3�mߢ~��L��+D��##���B�abe���,��*D�`�دR�}�� �"4��9��#D��{3��Y��1�L\ ��X�t�>D��ڂ�P	�D2e��j����I;D�0��MR�X��0f��3h�sŢ3D��1IU�9St3P��p��!�k,D�$��G�'m�2��v��1Y}x�+D�4 ���t ,�r�	�9��Ĩ��(D�����}��s�T�������9D���槐�"?Z�b��rz�]�;D����P69BܔKc���t�zi�Pl;D���"n<�����T)���8D���%H�9�t�5I�%H�Y��a$D����m��6�`J�iE�H�&	�g� D�8"��D
���f�G�`	P��!� D��7�ݓqW�-Ȱj@�Oi:|@ա4D�� ��d����K�2�X\��'D�0�s&سq1�h+�B_�}_
`�*D���t�̷;�x�Ц�[&%�&�)D���$��{��1i���?Q�ea�a3D�Њ'�Z9\F����~ȴ�
�B2D�H���Q�8`2�c ^�I2�e0D��
��	6?�ʝ���-2H0�Xר.D�4)bn�=G��5+W�^�d�Q(8D�d	��]-h`.t�pbˋu��ؠ2�5D�@)�\/^�1p�\�L�����2D���� 8���ہÇ�V%;@�.D�d�$�Q����sR+�S�>M��+D�l����3f��(���"=�jx��.&D�� d�I���r�!i3�W'��@�'"O�� �a�-6[�� ���R���i�"OZ1h��D�J�2%*ĮܱjG�Z�"O��נQ2(�|��gD�-=?ġS�"O�X9��͆J
��jW*! 5C�"O��e���j��5��"�)|$�7"O�|{r�ѹI]jH!c�W�:T��"O�-8��Rr�p�bZX����"O $�v��:B���R"�t<p&"O�-�R��<9��U)�j��"O�I�Ն\I��{"a@�t�
�
2"O�U!E�z4�<0pI�#/�f��"O�$���/p~E�p��qiD��"O�J�-wP�ۃ!�$<X�=��"O�ɀ��3b��d3ЅT �t���"Oޝ�bmH��~!#��O�Ș(�"OR���W�`6.pP�I�B�R3"O�Q2��6Z����%ꁌL��t"O��ɧ�	/X�^a��蜚Tb�x��"O��C��L����FD8SD��p�"OL!�NI�U�F������O�~L`6"Oެ ��<<�끎 �"YHf"Ol<�C�M=:�t�b���5�!��"O���µ`E�Y�1�̄w�vp*�"O��w�_�D��,ʄB-�8�R5"Op��
����{%,�%ǚ�0�"O�����	�~1c��?*n�p"OF|:�b��/~�YW)\��Z�"OT�'   ��̂d��� le��I��`�t��(�O��.}�~Px�� r�Py�m�0�~��B�6ܔ'�ȉ��*5Ѐ[���tNȊ|�����C&1J6HC�0>9�3Ch0�����G�Ut+�Z�hó8!՗'ص�*@�	�ꌤOQ>�a!	�0����D� �D�0o=�ɨc�c��RQ`�>���O�,�������o@0�x��[-��kؔP�1v�3�I6{N�� �bۖ]����BV��u�+44T���%7}���xD��: ��~��m�GR��`�׬X>���}��xY�JLA�a
e�7S����	��Tpd��'"S�S�O��=�qLH�%!1�S�X�H�J�<0TH�U	�/��7m *%�NQG��:M���0��*O�剽Y���vB)m��S�OH�%�8Yɪp��?K�8���Bi�5� ����O�Xi�vZ1+=�KPAO;F:����5}��u�z,¥���{�'G��[2�~�
p��oX���P��Dν&��''�>��GSy�� �׷7a�̲�fM�p�Y�w�̀��?�t�\�s�`��̦|&$`8!Q���*'h��8;�x�w�|2(A�99�|�<�'�_�I��-��b��p�+pG�C�8��  9���ɼ~(4��a�iP�E��+ٳss�B�ɃBwrf\�6���y�&�&���<i�Z�Cu�#~"���^(�I�A�.%�ܪ#+�s�<Ѳ�A#	(��C�/��m�'km�<'�Y_�Jf�7g�Bq�Fnh�<1�,W�b��T۠fR)M��eȶLi�<yjߴz\TȀ��+b �&G`�<��#�>�+'�X&;�{�+�^�<���^*Dt�����Ҭ�WF�[�<�6�'lJ@m�)�z��E-�}�<Y�#��t�p�y�!~�8�C�x�<#��4�8�&�L�������z�<��eNA���4Id��!B{�<AӠ��0�{��%ξ���u�<1����v���	�j݀E���k�<�q�jv�MsCY��M���c�<QEB��X>�憇�Lm���W�<����8H�xc��� h�i�<� e�} ֐�*�$w8@xa�Gg�<)'ֳo��8��e��#h�)�oZ�<� �=h��82v����톝p�6�H�"OB��cל}
�XB+Y/.��:U"Oz�(���>Z��3I_w�jDx%"OV��Wb�_'�Y����'@��t��"O�8q��?|�)Ip/���t�p�"O��s1.��P��C �R�a|H�*�"Oh��c�8z��Y����l��4�"O�E+1�<vTĸ���Z�\��,Ї"OLꖀ�P7�h�'�1U�����"O+)Z,
�Ρ�b�f��EbV�Py�<��P1P�j��#Vp捲�!]R�<��@�LlB�u�V�{/�/�E�<���!u�Z�I��݇2v<�MX�<y`��>$ꊁ���R��as�U�<��"ғC���HR	��-�ꭲ�OV�<��U73��A�4aо4ztݠA.	Y�<�3d~�ur�µ+bz�@���^�<��\T`.��e��_�����c�<q0�J"w�hy�B��#ZZ���F�<iR�_�7@�eX@k�r�Ƥ��GJG�<ɂ��*�Ԩ����#!C�}cgj�~�<A� /Z��=��BKB�C��r@p$䆁z� R�J�/nC�	4)$
��@iG�R��A\4.B�	�w)&\	�^�`�����ܳB2B�	�xt��
ֹ+F ���]�G��C�	x(�|+ÛbxNx[#�նe��C�(4�*�c[,(N���Hӏ}��C�I�Twv�'ǱM�(`R1�S�QLC��]?��eֱGk�-j$O<E�C�A�~��G��mI�$���8@�!򄇥T��/�4q�B��LB��Q"Ol���@̸e^|T���,��-0�"Of���[!�@4���&����"OX�ee��y�`i�Ӆu�P�Х"O� a�倪`&xYS#���AR�"OJPW�
=-�N���b?Y���"OĔ�A�&K�Nd�PO@xL =r�"O��A%jU\A��/�!n[�(6"O D�e�ӳ?�t×-3lO�0�0"OجK�
4xU�74>h�"O��"���R���,Ǧ&H��f"O�X ����"��J��{v���s"Oh�1��'F1^��eFM�{2�Ipa"O��
���*�6l�V�: 5�u�c"Or��R�)�$T#!@���Z:�\��^�b�����ąYs�ܨ��	9w�Ʌ�ů �X��-Xjv�{7��\)\�ҭe��5�k�N>e���UVj6ዧĳC�,�֍m�\��!��@7n���$�p�����0R&�]PEG
��~� ��5d��:��ª:S
��i޷@���(K�EI�=i0��c��H�wca!��<'d��S�O\�R0T�W;|5"�٠
`h�!Յ��RBQp���!�	��F��(�j�i�Y�W�"ŐDM� �ug�~���(���I�f4��'v����(@Q�X�F��+@\I�J��L��̵h��t�Tӎ�h
�'8����ȧ�G('��m���^����U>@=�%N#��Eqg�GY��4g
�>U�S�T?��F&�?a牊���O�L	�b/�,��i��j��~[�D�H>��J�%~Z���>	cǅ�0i>&ei�F�Q��ՠ��fӺ�m�IX��H~}Ҿ�MG�Tf1|�NT�
ԝC��P����dd�ˇ�1�B��'�!��S��v���-�j��/�?n!L�:���,x@��y`�OJ^�P��Li�;p�H$:I ��n}�L@*�iB`>	��N�V9��zR|s�<��訟���Ζz֎ᓳǉEGa�t ���:�l[�ne�LPSI�:�M��ӝW&�i�Í����L����Ǣs�Ј�O�/R�T����=�x(2g/�A�铎0|n�@H����(PYe���_��54%P��Ce�����3� v< �ңtl��ڷiE�y60,���x�O�
&�nd�=�~"'b��ow�LI#$\$"�ب� �{}D
�!� �=E�4������#!B:�}���5�M���>���ȟ�D)#.� +�v��!�g�ܙD��'����Iއn�eKԢ�8�)�Ҏ\ K9�O��+�2�)���?.R"�9���f�L9�$��'�,�b����$�vࡧ�W�M��C4c��_�I�]�Xh�?E�4O�A��Ւ��AZ�6���SQ�<�F.ɻF��c��7�$�#�LO�<ae+�XȒ����ߢy�,)*�	U�<�-|y�9� E�ʼ1��M�<���9 ���:�(�e���[0�]A�<M��X�d�ʛf�1!ӥ�|�<��)��� "h�RPȌ�Thy�<�UE� 3���#���Pf����@�<��-D���Q%�Z(<+,Ip0&�z�<y2K��-0���ǎ� �|���s�<�@Ř&7<Đ{P,�4�V	;�Tr�<���S�S���É0��:3��b�<i��[��Q8n�� T &�]�<�`�3f��DssD?E�
! ��`�<�G��[�&���C�82B1ⴣ\\�<A��d�0p��2Q�bX�BΣgD�򤋹n��dS�&Y�>4DBa��C!���t|�C�ɖ$t�b���5o$!�$�$P�D)���e^�2G�!��B�kt��A�d��@B(XYDIX�Py��L�.��(ˣȑqxP����y2��.L��]Y�D��4�֭ҍ�y2m�U�iz�I�' �������y J��(<8��r��<qvʅ��y2ۡoq��5LX�P�%�yf�6��Jd�E�Uy$���fC+�y�͘�HiJ]��f���E�qˏ>�y� C�YJ�4���"��B EA��y�͚s3(�2w͚G�|�@0�S%�yBc	�-+���<��`r�E��yrG��R(i҃��)3��]�f��y�eO%&�8p�ߢ@i���� �y�#ՔF̌���۹OD�٫t����y���9�h��r�ZP���y��ܤuɼ����!�8��h���yA�,����d�~N����G��y���t`��yD�v��DAb��y��ڿK����a͕m �����y�%0��a�H�SL��`�g��y�N��)��gG�1_Tu��Z�yr��6st���fɃ>�`�g`��y�iZ�zU��z��ڈ �N9ɷBC?�y�+5t�8�+�*����ch�+�y��?c��n
n�l`C��'�yf+x��x��f�%;��BH��yɓyھu��#�f���
q3�y��	$x���Y .���X��DX�<�U㔋bd��',�<sb�N�<IDK>e��������K�D��G��b�<YT��%o�2���ɹ/W�2�,�Y�<Q�*Kp �G׌1�Ғ%So�<A�c޾ V��"5f�w��TMV�<	 l_�F_�\���3p�޴��[�<�D
���%�F
6&<z��r�~�<���1���@�,�*�13A�@�<bF�m�PQ�u�)sn�T���S�<���
7��a��������Cj�<� �)R��;\�zǦP�~�X��"O���'�Y:
���葦��0��!"O:�w�ϊO[��Q������"OP4��'�Fߚ=qA�S-����"O0�8SFG�3��QֈT�	���D"O����I
�:>�]�FBN[4�I�"Oj%�e��*u�J(H.�S�"O��7��U�0�!7�^�#(�K�"O��`�L�M�p���7�R��"OJ5��{��[dl�����#"O\1���40����?�lJ�"ON�rR*G�K:pM�G �P�^iR�"O�=S�^��� q��Rj(Q�q"O�	�m
�yU�'�ڟk[^�j�"O��[�G0�`����$h>��W"O$�	Ջo��:Vɂ�nW��P�"O���S#�${t���([9fj.�u*O$�p5���5/��@A+G�QS
�'!�yjЪ�5<���� ���	y	�'��QTL�"Q=���@k��c��-�	�'*,uX�A��YV�)�lK�:\�J�'*��r�H�ux��;�bҪO�v9��'���n�0:@���H0F�)�'iL����U��	�%FڅM骡��'�����;Ym�л�H��X�٢	�'8|�"�Eh� 6�2�@�"Oz���8["Bd:4��_A�U`&"O��q��-�BMRr��(]��"O��#J�q����Aū_F�xI�"Ob�"�A�^�Py+�`X�f�� ��"O���
�jBB|��ʉҼ�*�"OF��T�M532]� �F<���A�"O�=�d�#NC>���IR(�6���"O�uഊԯH\Dg�$p�"�"O����9f -�Bo�UxTQp"O�[7��-HQ�TG�,G��9�"O����O"t�<�����{�Y �"O����B��L)�r�Ɇx<���"O�A�R@U�"5Q��
o^Ƭc#"OZ���цLz��t/�5a��E�6"ORtI��Q�! �����-Zq��Y�"O����#�]�`���~X��It"O���%,[�j��� ƍi=:�[�"O�0j��H�T-�u:s��$'&�=�"O�xy��0<���l�#	%p�"OȐ2#��8"�P��D�!R��!5"O��b�'��#�YCE�٦yZdE"O2�ҐEҘ\pD蠵n	�.vp�8�"OȻ�b>o\jI��E�
Ԗ�1a"O��2���$�G,�i�"YA�"O�4��Z5i�Ա{�a������"OVT���F�9�E��čw����W"O�uӧ%�-�v4@�"�:<z�Сc"O���k'*�� �9G`4 "OF�6����ŪB	�R4��� "O� �͟�^o���k�?PfTy�"Oֈ�R�[�In�@�ɂj��D��"O����S���a��N$\���j�"OjX�����<��E[���Q�"O D�VF:-2Ȉg%��>��m9�"O\�0!�����Xt�לzq��p"O�����}�N�s4���RH"W"Odp%2�JpBn�Q`��t"Ob��U.A7i�$esAn��m���R"O� L�ʐMк�Cb���k�r��"OL�H�FF��y�� {� �G"O�0*2�3F���UN�;�13`"O ��"Lù�\�RgF1��"ONA���!,��`@�ӵ8sR�h"O���P��^aKT�O�!E��:a"OJ�bu���a/@ 8�bB�V�؊ "O��1�ؼdrb�sA�_�hbB"OdH)���0 )�腀��`ۤ0�0"Od��AH	�_����ȏ0˨��P"O��)�@"h},�Ô��i�.�� "O�Bh?�2$��U�b�]�&"O�Ec��$m4��Ԏ#rð� "O�c�cD�N@�Zଈ{����"Oq� M�0+��9���C��P0"O %h�)S\_v�ӆ��9v�>,j3"OX�r��O# %�$X���� 8,�X"O��HBbW2g�i���l���Y6"O���$��N����ר��e��"O�[�a�Jx(A��"�49բ1w"O�D��!��"��-[�! h�zf"OF���a_h�-2� ց#9X���"O���&�T8t�`�b�`T9o����"O�)��C*z�T��(�
&�H�!�"O��ز�΅GL��CpM�"o:@=J�"O(�`�`ۺ%�<��a�-# D"f"O�G�֍�( ��ꍰW�D��"Oyj�H�v	��J��Cv�ts�"O�9aցJ�l���Gh���,9��"O l�f ۃ=B�X�w�ֶD�n�Xc"O���Ŧ�$��)6�
�S�6���"O*}
���0��ѻ��)lhTP%"O�xi#&G6m�0(��A/rq��'B�x�I�8>����5���':v@ �o�a��9����C��;�'��!�SʧZ� �լ�Sв̛�'�P(����5��rT&JV~���'�
����ي X�5��HC Bo�1�	�'u���4��ZL[ �Y�H��ѻ�'�yr��cv�[q���A# ���'���a��*Kl�AN<���
�'0>�ɱ��|!P5� �7����'��(i⇂>7db�/ږ7>.<P�'R�):C�.QD��S���g)���'�б��1kX	qB�b�� ��'�P�p&�9����$͕Z��X�'	�l0a�O)L0�&�#R���'��H�u^j�|��`�Q&���'\��B��'!��M �ݵ9�a�'���w%A�=!����+
��]i�' ���!�eA�H4�Y8줸��'��9A󨗊[������)1����'#*t��^�@���Ǧɾ<ׂ�2�'�f��b,�"^ew̕<g�y�'�"�I���d�4���[:��J�'��jf�,A��8��+C>]a���'�8\�����h۾ �u��C)4�'�rQ2��>#��l����*��'>=�T$V��j����7�2�'�ri��X�.�XD�FC��,+ll�'�4�%H1#j)ض/M [���'��1�P*�5�ݫa��66p �'��Ĳt��g�@h�u��rޑ�	�'岄�C�ԣ?~E9E����	��� �<b6/]�6 U����"�P�"Oڥ��@ G�\�X�O��l˃"O�<{��΍3H îY `A"OJ԰�`�)i���i�l��<W.H�"O~��(�!#@�1���,�N!��"O"	�'�W/�����אwlH�r"O�Ѹ�L��������c"O|���nɔR�u�횇b�ܙY�"O4����3n<��� O��Z�"O��3�ɤC��h�Q>9�qK"O��Z�,���K�	�\	�J=D���3B   ��   �  	  �"  �,  �6  -A  �J  �R  $Z  �`  [i  �q  �w  ~  ]�  ��  ߐ  !�  `�  ��  �  )�  l�  ��  ��  4�  v�  ��  ��  @�  ��  ��  r�  ��   E �  � �$ - �3 .: �A H JN �V �X  `� u�	����ZviC�'lj\�0BHz+<�D��g�2���	#���=�?Y�� ��y��%+�4y4��%Ӓ�Y���|c��P�d^v(��q�T�ٰ��w�
�	뎑��,�	"���	�
�Π�Q�'��B$y�T)t��8���S��3Iˬ<3#"�2V�Ŭ�G@�]��G͛V,J�Y�jp�@gP-#�<H�0�@�6N����
�=�n<x@~�rdo�o_�m��ޟ�	ڟX�I
b��'ӝx��	�c�7ܾ�I��h`O��M{,O�L<N�����O�����mQ���T�
�2���Π"�|���O��mFy��'��kQ>�M��)��"�zE�6�5"F
�1ւ��:��UDN)eT�x+B�Ob��'ɾ�f�A�T���@C�&Ţ���ŉW�����7������?��ň�Vs�m�p��.�y���wm ����q��H����#�?��?y���?Y���?9����)aޕj$�ϔk�ơ�v%�٘��O�O��m��M��iN6-�O�m�6c{�,��4&-���u�X"�Xt�/!T�0�XP�==�pE\� ��֟,�ɫb-qO�'8K�q�!Q�>�XU��6�ZM����x�u;I$U �L�Ɋ�M��i}�Bu>��Ǻ�!Ŏ���������롋���M��:���p�W:L<>���n�@@[B�CX�,6@Ϧy��4e_0�� a��<��A ڙ\X�p��%�l)� X �%k��xm�( �tpgE� ��$���0/�@hӖ��N:����;�xC���mP ��4��H�]��4��G{�Dp�fP�9���(�*L5 m�"�հC�8�B�^�;��h�Hѓ;&�	o/Z�$��o.-R�r�oE�a���II�P�F��ג=��H�!�;:F�H�����hy���?�p�i�4�Ozܱ1H��q�X���'�vii��˰A͒%f��%I�4�';���� �����P`J]�t&H-#�E��M���F�ߢ�(�#k���TȒ
F����C�����j�(k➤s�4<�zp)�(ۄr��)t��:��#�k���0<��ty�+�<IG�Z�N*e�7�F��%�J�䟬�I韈%�\���x�'��퍴mw u��͵�, ��k��y�R�''$�@��ݭ6��'�������O�AKA��Gั3eFT�h~��P�'��I�H����4�?����=��� ��4�J��B۳	���'����3��J�b��-�6�^-3��?}��F�t��EK�m6�h�h��'%x��AĂ	AOQ�6ǉ+����`��D�O��=���]+�v���MҐq�����O��1�'D7��S�O���9LE(�M�UaA&J2n��'��'�2T���|���&!��c���N(��~�'�R�j�d�l�����4���
6N��� c�u$z$Q-\����'��I�^�8���0���p�'��!�LH��n�dKȍu��P���\6M��J�nA�Rȏ#(x�˧��=1�%��/�u�f),\�p�㟾J0�%��R'Y�rU[dhƃ8S2i�|R�J��d� -���XW���G�
�+r��k�7�GUy�\��?������|b�4[5����.N���b$г�ўT���>J�$����G�lΙ��Er�Z���O��nZ)�M{I>�'��-O��"A��l�Q��L�����Cod-�'���'	�Iy��?�x�b㭓m�	@)�5��MJ��D4��YЦʛ�2�*7m٫��x��-n˰�;M�7?����n�"px ,Y)�^������Z�"��ʝb�TGy�*�qD�p$�	�����X7����F��5ғ��/?I���Y�$i� ��P�(�9 F
֟l��	k̓]��tz��Բ,��hZ����hX�I?�M{�'>�VEdӔ�'E"(!��iP5O8������37��ό�Ԡן`�'���'=�	էx�C��|��ҿiU�)8�,�0��D�4�� w0����W6ax�N=�f���� �j���	��n���е�+ID���լ� @���)ĕmE�%GyB�X��?��\Q�&�'����`�Z�*A�$0*�M�h T���I`������mP�L�D��b�M!{gJ4�W�$,��|RչiP�E	�cŏ=t�����7��qB��x�t�d�Z�p5�iH�S�`��?�	��X�;R
�.6=h�c�j�/Ì���䟨Z!ȣ����jT��M�'"���O������ݛ^�x�s�MU+Q�R{����Ct�V6a̬�ye�U.-��2�6}psv�~����?K$�YHvc�34��Sj�p~��Ɗ�?� �i����c>=���&X.�U	�Kъd�R�8���O��O�#<��ϑ��>�h�ǚ�Y�gER�'O��x�f�lS�s$����g�:~����s�ז)�b�8�4�?1-O\�z�l�����O���<	��Rl�NX�E�'v��x�2��;�Ⅹ�ω�Z��k���Ӛ��(�j���1d���Ǌ�^�(1��0���AK�8͢*U��x(;��\)&hʧcm�|���L�+�����#Q�2"�X��4�M[� �>1b�����|��埰�I�B�):%�xj��@eG�w���&�l�IJ����� eJB0c���,?Wr�kb��O��������4�?��i��OT��W>�J�M݃(+5k�� �V8�FNH"`�r-��4�?���?�,O1�MR��L�G����Qf��ep�3���Cl�w��,�l�!ڃ��<���wɤ%D�:��<s��J�G,�`7L�W���m�)� 	����A��0&f����B�䩨Gi
*r��%��=6���F.N��0��͟��?�����n.,� `엑'��08!�� �{��$E���u돎G�F�j�Ӓk��'[�6��Oz� 8�TZҵi���=�hXC�L�	�X��IQ-̜�Ģ<����?y�OHh	��p~\{ǆ�c��3� <�#d�͗MM�0�U		�2V0���' |�#���;~&f���DL*bx��ʙ�n�c�˂N`���c��L�tZ@M�~�I7�|B M��?	 �iB�O6ꭙ/CDp3A�V�{{>�'���I�5#�f[�;j����^+b��<�d>��|b&�i@@���cY�&`2
��}�.����u�N�v Pf�i��S����y�#�GC!�-��e�x@fXh�"�'����/ۭ JɄ�[}J����i��bًG�P��qHebI
���W��C�L�4UJIh��6H������9�� �ŗ��b����e��t�oS�k�x�0�d~�g�&�?qe�iv�#}B�O~��9s�7R����d��� r���dG�BbҐ�`�U�}�)0����ў��	�M�E�i��'bF\���Q�8�0�صG�*�`�A�'P�W���b��D�	ޟl��Ty��-0�(�<|{����Tv��\����(ـ$§gەh(HU`�X>��3�� ��q��G����J���1`e���*��hf�a#�%�"l3tᑚ>�t��O���@��y���=u�������|�VY u���<��������|�L>Q�G�:v��:���	�M#�@���$�O���O��I�>'�:��D^+&˥��U���'F�7��e�I2�M,����|��"՚R���T� ��"${ң�M��,��i���'/�X�p�ON󩙆2���H�჆����el@=3
��4&i����D!I�^�A	�%H(�ɤ�&ũ�
�8w:D0F�:UhP3@
S	�BUZDeO46r�+�@Ŭ7��E�K>�@ů[+j%Jrƕ;u���)�i�5���I�M�4�a�6��U@U��!�v�s���nLF	����?y���hO�b� ��?�8	�C	�@�4q�C6��ަM;�4��D	�d�|���O��DG�*Hf���+6,��X�m�{���d�O�)��O����Ode׸18�K�ȦQλ8ƌ��E,Y�ڽ���Kh��>T�
H
U�H�aypDiA	�S��@�We��ee�D�@��3��U���~=��:A"�_�"�I��M��W�ĳ2�:� �аj@�9H�>�?����?I���)\?wD8`;���1�!J5�;�Bk�	�O��?�ߴQ��B(ՑO��R��	�.лE�ir�'�*< �}�z�D�O�����X���O���RM[#����r��
[�Zp�f�Ot�$�[���%�|�Ot8D��<V��#�c�.S(D�B��L��+�S�OU���D,G�چ)�1Z�<C�O����'��O>���LF��tP��b9�5:`�0D��(5�T�)T^b����5��5
�2��,��>E�d��&4gB��F�	)5l���/Ԧ�&��R������OX���<qL�\t�ԩ#��u�"uI��
�R��b�!@�T�S��RD P.�����_"B��M�E�ްp��d��l�5)�z��w�љX�.�4��'c�2]
 �:u�2�'�j��/Dq�1��h)�1��V�NO< ������+Oyz2�' �ĝ?�O���!�M�֕�FS/p}�"N#��`V�>a� �	 g �����<LA�B��O��$F���Qߴ���|�����Y�0��H$�NuS�=�W���8�V��Q�^����	�����ny���j�C���*�k�Tw��C���A0��ʳH�B���7�$N���I�W�~��`��!$���T��Ӗ��hSJ�C ��\x��ЬQ9�`���1Q�|&�|���+�x�3冕f<NP�P=Ia~��O��D$�	r�OC�hXE�B�=&�`,��A�������'�TBq�#��y�P��(�:��N>y��iX���H����i�O�٦��/��q)�|4d���O,��[7F���D�ON�ӻ1�j���1���(�ş�1�)^�u��B��^J�)Da>O�Y	P`Mr��t:p9
�
�����X�4<"�Y�6I��d�axҁ��?i�����_H�0���M�}��뷅��'�a|R���JFT9��n��B��hz�����?q��'����K��`*�Ps�
�rvB0#���D"x���m�ß���c��mV�`R�L�?�3��|]�)��	4�r�'󢡡��\�"�T��o�?�,1�0_>��O����m�h�0��2�@s�L���O2�3�c��<��ځ-�81�d�aQ�U8)��Y�)�1�H�i�j�i"��=<��p��=E��I,xx`�$MY�)�'L�dH�T3~�FtZ�_/�ԭ�ȓh���d�ǌh r8��H�T��D{��'��"=q�S.�8��1 �D
1�����]�	ɟ$�	�4�\9RCԟ��	�� ��¼���]X>�k�c&8���a���zD���*vUd��Յ$��՗O���{2���rGek��-�������<���tD]67*��A��ubJ�2��H4�=B(2 &ig��� @�;��	�d�޹���{ҧ[��y ڴ�?�g΀+�?)��,O�����pC؍p���_+�%I�ݕE��˓�0?)TM�Qj��@1�L�2���D���͓�MC����(Z�h������+x<q���|��q�vk�~k`(�+a���$�O����O8�;�?!�����ؔ1߾`S��!d.�8�`��
D
|q7k�2ǮL;�%�'�j���	8(�� �Q��ķ}���&kȈI;�� e��~��{��P�}�XD9�E �X��A��޷r�R���A;y�P��o��\�Iɟ��?�����l�pc�܁G=�]X��Ԗ5�!�$F�7�́��N�6l�H�K�@���':�6m�O�ʓ����i��'����d&�8�Hd�N�-Ш���-6�S:�4���OV�D�pK>��b��0�$0����ߡp��%^�Da'.��9�H<!4�4OR���Ň"ap�I��dG�QȞ�Οt��0IǍ�'{��|h�+��<ax�I:�?ɑ�i�
7�O��;�L!oV\̞: �q{Eʥ<�����(��M%�ӭ>�L�[2�)%�`	ۑ��F�'�7M���.�S�c�N��*��>n�2�d�<y�	�@����'��Q>�bH^ş`��t,�a'ԓu��E���
ş��$;�� tL)
:(�i�΃DB�L�O��S7𵻷�j�n�[�
��k-���ze��l��b�Hz��H$D���S1KڅI�J�k��|ҕ�G�̌ѓ�͆w� �����~~���?1�i7T7m�O�"|
K�-:����n�*g�F�zk��Ԗ'�rX��g�}*&��g����I�'��!Ti��G{<O6�ͦA����M���Q�-]7�~��R�n N%Ith%�?���?a�"@[C.eZ���?���?Qd�� �Q�C{��H;q� j�V�(Ppg�(�� a�1Q��6i/�3�Iz+�����߆$ǘ\���
�b��}�fFV����A*�(f���q��^�JENa�O�j	�AaU;�yg&/P~^KL��d�! ��`w�'�l�����Ϙ'���	P�-0��PL1_׸x��'J��ˀ�ۋBo�<�@ꌖR|�����?��i>Y$�Ђ�"Z�x2.|����=�^��r.P�a�Bi1�E�ğ��	��D��7����Oj�X w�t�*wΙ& `L"e��3l�~�����r�B��☻bļ���'�.�z�+@�91MX�d�䊑Q�h����F%�BO�.l:\�v�
,.��|b�����1M����Үm���������4����'j���@�'k�S�H�s�"�$'�4�+RB��@c����3�	2x��A�M���k�FM��O����O˓!{tbó����OrL8u�Q--�����"?l``	���O>�$O�]"����O�瓹�,��&`�&|(��hd!ݟ��ʨ=(´�"*YD$�S@=O�a�O�U(�щp6��Tzâ�8a�x���q�aJ� D�B�ax���/�?)�����Ӑ8�tUr֊�2e�&ͻ��O��'���':"�� �!����`�C�p�+�=�fR�(�ܚ�(�H�J=k��^��?1(Ol����9��ޟh�O�T����'A<�	F΅&�,�BG��F��r��'�� 	�`k5-�)s��@�.�O�o�o�
~,�4;�ǋ]A�@�AP1��ו-�\�q��F� ]"i)�'G�fĀ�h��L��P[UN߽G��'�T����?����x�tw�D�B�}�୘S�l�2�5D�,�͑�/�P}he�׮B�L����>��8I�>QӥfK������+�eaE[��i�Iџ��	=�d��u�ҟ@��矐�	��Kկ�'?�l���ϋ?	"���g�V��`ς�d� � ߺ��|r��x ��J��E�bꆶ/�¡9�Fđ_jJ� �V�ìز1)g �������1�D7M2�K� �;:�����R%���������OL��)ړ&Pn�ӴdT�K� ��d�;͚��	�'�0Q�f�l�#ɛ_����)ON�Dz�Oe_�8h��^i'@�X& �;�-*����+.v1����̟\�	��	��u'�'GB:�y�#�Tz#���gZ���4	K))�;��)�V�yF�'<ON��pɗ!<�NQ�DY�v<х�E�u���.: H�)�!�j�axbm�c���ц�[�'��Q�U�$}��۟���^�'}���C�;s���,�N��XK/D���U(�(p�Ĥ���XZg�.��Rʦ���[y�HF�X�P6��Oz���=�pq� �#~bz ��)E�
6��OJ-���OF�$l>m`&�Onb�xP��6W�HȀ����-�c�)O �!�	Uƪ��\�e(T8�\����\!(�"�#�Dف2�n�G�['A�3�U8[�!���P"8�8H�Xƈ��KR�J��2�O���-�*$�Z��UjA���!S�|"�K&-��7��O����|����?�&	6
�8s��QS�k�	M�?���;��`;�Ƙ��>a%�ܲ>���t"�0%.L���P~"I��O>�X�N����!A�]�Tu�b3?���퟈pN>E�
��j�b�y�ӞR�9+&g͛�y�K��j)dr�j�����9eN�*��OTXG���Jgn�7�^)C�u�v�S3j���'���'�vl��`Y)"�'���'g�=17�W˔�V�}Z����r4�QS!e]�Dۂ�d�/�p)���$ԽŔ`��m8hz@lU�;[�]+j=y�d��I�=��=�B��� �!�S��)�,P�kM�)a@�'���!�����O�=�g'ʇ6�(,B�'�+ĸ�����y�N`o�� bR؈Z������w���t�'��L�d�(�"	"!���X�!4�觮]?Z��h������	͟�[w���'�U�L���3���`�<�yCC
�c���`��.ĉ`�NA؞,)���0!ɘ��kk},�����}ܱb�nDj���ۓU/���
Z!6)F�a�(e'.4ju������}�'��X�QM��J\)�
.�̬���'D�t�tA��L���0��^��H��9�d�����`y�,�9!r��'�?i���6Ӛ��ud�tqNT
�N!�?q��Ҽ9����?��O�D b��ۚ90� �� $��
љQ<h� S���ʇA�-rNHC� Q��B��;d�M����R�Q��x�
��lN�ż1@���4�j�,NF�Q�yDJ�O9l�9���ʷ"MD��&IMq�8�ۀ�1k��'�a|�տ2��%r�d�,X�4���O<��?i��')�H����"	�����C۲tC���$ĄR�ioZ⟤�	A�4�	h�"�O��F-� b�71�੢G¢/m��'2��Ѐ��:�ʀB�݌� C��EL\ر�?��6A	$��
O��Z0��e,?)�М
k��9�	L�d�f "��/h�"����&�4�����AU�Ԅ�3K���B�+�"v��E��4�H�"d�0�b(���	ci���u"O����l�#Uk�a�H�W9��3�I�h����^",lr,���T*I+�@a�Hp�����O��d�4y�n)�*�Oh�D�OF�dq���*�*8��yF'N��j%k.�ɕ"d���M#(@�3���:Xs�g�50c1O����'�����f�-,�pP� @_qz8��|��@�?y���y�+0y�����?_�\�2a��yRmB�5��Z
 x�rf����W����|���3v��X�`?)��Xч��m$�H���c
��'VB�'r��]������|�ᤄ�
��H�
7s-؈�����aP��P�Ŕ	�b�Eá?̀m`e��mAn������	��lÕq��pe+
�r'&$�"�Җ5���d� `�~���L�ơ$����/"*��K6���,,}�W	D	cx�D+�� ��2VT��Å��k@�0b?|O�c��а��W���`�y�"G�;�$\Ŧ�'� y��ø��	�Ol�Ã�<A���Z�K���9@��O���Y#�����O��Өv�N@1�[�}0CW�;]�5�ϔS(
��Q ڶ'��I�WM$O ��&���z��D���jLTy���C�4��(2K[�(��T��^���Js�F�ʴ��E �D�����'G�I�v�hT�O=X���kA�X'��O���$�a��)AC��� ��M�Oj�=�'Y_�k�3����@J;"xx��t���?�+O�
�������	֟�O�i��'k��i �|�r�`�A8{�:���'����X���ް.EP�k�n��˧���3@^��3E�ŕO�`��bg�9F*B��,u{ I�H���i��YE���L�1Y�̑���8|�\Iw���$:2�'2>��b>�$��G:��7����쩀��8�d�O���
9�r��%�'l)VT��.�����?��O��lZ8�MKI>ф��+1�x@@/�"ӆ��G���V)���'��']�
Y0Q4b�'$B�'��ǣׂHv��6V���ƞ�A*��r2�ě^��l�-M hR1�(�3执KֲQ���׃m)4� T�O6.�����W,8;����O��X�bM�'{�Z��Of�]�P��~�ŀ%3��9�3�Ɂz�
T{̔՟��'�&���?����'�F�x����@�h�ߝ�Ȭ�E"O"��c��u��]CUȔ�w},��r���K���D�'$�>C��X�J7ou�a�� t��@�tH��4��ݟ�I`yʟ��$2tN�a8p�_0��j���	>(�� ��Н4 �l;&x���''�����*�PY��L�t�� b�A1,8�qі/��D�U8�بः +Ȝ #k
8s���X ��<�����O΢=	���fkL��lFw��+���t!���j^Ȅ�Ÿ���
�,˼#��'g<���?�x$?��2G_ [~�ٶ%	 L�v�z���O�˓�?���?�%�7j�a��m؜$0V�ƅ}�̬��˞���QLɖS,I"Ów�t����Qj,CsOR3R
�����;�������9db�4`�,�OX��+?Ap���R����7*��F>֘�R.Fb�	`�|@����h�� �x�D�/1�O��I�+9�Ri�K���8r2���<	�����?��O���<1�]��Yc���e�C6W#�'���1���"MY��'$I$8b���)J=e��SNV����ׅa��*w�� � ߵ8�H�ٴ*@�H�|ڲJ�1W��QkD�V4l��D`	|~��@-�?A��h���)� ܵ�5���#`U�A��G+N�ؒ"O����e��c#�s3`��^q����	(�h�>I�F�pw�ـ� �u�2���{� <3���<y3�@$���I;Jt���I�7�,�a�i��T�B-�u��'����s�B��=�&�9�3�� �~9�@��-�E���7U���H�=4��u{!�5M����ƍ,�3�	"k�&-�g���E�b��B`I���mn����o�O��3�d���<4���"�rtd��B�I�8U <b�$UQ��q��&���+ґ���$C�~ItUf��3�fG�;��0�@�8�o/\O��Q��,��I�K�J"�k�Ȑ�tr���V$ND���$�p<�C!$O�t1i��i��`i��
#b��`�WJӈU fyQ��
RX^���)Mb1�į�	�ܐ��Ks�.��'tL7-K_�'U���d��'b`3%Q�<�� &D����9n�ȱ�SM��;��q#�"��\t}T�xPa����M�3)RGE�^�2)p�R�c�V9��lk�'��D߱zn>I�a��@���!��*��e(ŉ-O>�c��I�!1��r���}>׌�	C�f��DM�3��7�$ۭ
�R]B��Z?n��Af��'#v!���,� 9�@k̴Dz����i��B�O|�Ϝ 
�F$ w����X`�|`$'�6-I0<Q?)��-�!A����2��I�j�j G1?y!C�/�zi�ւ�;YKv-qg�=�'"�8�����"`����&)'B��'b���/Mz4�s�[>&�X�E�d�[2�Da!����$V���䝅��kӆ�G�t<��=���͈5Xh$�5��C"O� �A�8�����]WnD�T���h�H�ᵦ� 
�|���薫.�8��5�t�()�n�<a�'֮���	�7��]{t�Ef`����I�y�4c���W�%LO�ԛ��U���񳄁�>5�F�dI�yaz�n�+��%q��ĹEܘ�#�>p��'ې����Ϙ'ըa+�[S�E�T	��q�H�;�'a��Q�eŽ����A�b�*Tz/O�MEz���,������B�.�`d��_"n6�.X��i���x�jy��d��S`�y��q��//]ܛ��w�*i8�E7#��U�N
�!�0�'���Z��'h��'�ՙ���5�$�`��I}�OGX��q��Gsh����3ZGz4"����0/V�����~W��&>-[�h�8Y�f)�'�"�z0h��8�fHq�I����|B�䛗���!i׺s�H@�bkDEy��'Q����I�!���5��M�	�J	�I�{E0}k�FI@��#wN��v]��E��Y���?I�����]�D�v���O�B�&��a"����Żg�@�*�&�Ob)�S��_�$z7+4rk��3� �|z��=U��	���~3��yR � t��I듣s>�0i�Hۥ7'\ٙ���/׼��7R>e����~,�}���ظz�y�D��b�O���+?%?��'i�a�7��6��x��V�**XYp�'��@�A/v)��*Rn�����'�#=ͧ`y�8�.Y*_n%+�O�2�F�����?��?j�E	C�	��?q��?q�����?�����M����c��!EX�r5*iN�K��\�
�D��2������/Z潐���ncf��`�^Z����� �ҸZv�����GXY��M�-��X�4��:�yW � MM��!Wd >9�|�8�˻��D |UR�'�ў�Γt�aG/F �3�ҙy;0-���U�I�br��q�$��22�@���o���S�ܗ'	�h�M��6{B���N'�f�h�F�IT��'�"�'y�)�S}4��(��	�qop�Cf�"k;�1�$A�I�ؽ*��3ֈ�u�6O���dL]�*���	�꒑4亴�B'�E�<=8���F��H�G��p<����ן�SB��FY޹P����R�fן�D{"��9��!�7�P7!�(�_3J�B��F�� ��ń\yV�z�Jj��ʓl����'���&j�N\���ľwQ^�X
��b!r�QǨ�;nD�	쟀�	��P�Ci Y�}��	Q�+�7�|b�)�;��m�Ec_(�P��6��l�'<��94��5Z�(آ���G� ��|����J%���2��k\(E|�o�#�?9���O��T��4e�؍���F|8**O�����2n�T1�^�]����"y3�}2e�<q���7Ĕsg�1���&_Iy
r�R�'<�	y�T�'=ذ@�FY�5�C<,����˟r�bm^c
�|�cLD�6�dx(�ԫr�?eC�f��.��xpL_|紘�U#q���AL�0�*]��j"l5��"���{�#k�2о��
�}��	�0�X���O��S�Q~
� T�sbF4S��<�Ӭ�,�ZR"O��ʐ�>F�0�I3�+)�CT퉦�ȟ�[�TNCh�	4J���8XF`�Or˓i������?���?.O�	�= �$��7�Tc�t�����=��\��^�J��ɐիʁz�����?#<��$���Q 4����q���N�8+�q��j|�T���ܼ9v���OP���s<� H��;rݜ��"�����O���4��yA��T�zu���'f�Z�h/�3�ybMB
I�HHF�J�-�4�R��$�?i��i>��Py2L�1��q{�HU�zOƼqR¡y=��p�'���'5�R�b>�h��E���;�nM5!�Ix�+W�,}�Y����@�LЮ�n{D�Ǔb�q'���-S���ɦ}�L���P��@,�1�Y�	a���tM(O���'c�@s�)Ƹ^0����x^|l���'�ў�F|rh�p�^Y1dG։��4!g)��y�h
� m$�Ȅ��/	w�DA��������M�ILy��;;d�맅?A�O���'��>wX�� ��fp����r�8M`��?i��f�l�jDM��Y�&�>ͧx.h�$�jBH��tm�H-G|JϘ^��!KL:'�l�t�
��$4#ATr�P+��I��$�O@b>�0�l H����_� ��9Ö�<��BL0Pp���k����=���ɂ��DO1T�hh�+�o�ޙ��N�2d�	���	⟬��џ��O��	�xaAEO´+�N,:�&3���I�IGxD$N�|uP�L��BD�|&ώ��'���iM<	��D�'��%X��/[��I`j��F7�Or��e#u�h��H�O��D�V�$t�0��䊶�hi	�M>��*d�	_+nZ��Xc�ɕ�\̓E�-��ם!����&u�@ȟ(EkI�hf��p��R��?9��S�� ��'���O������i�,����Y�<HfL��NAa�
~�����O��J�$j�0�U��?7��T��O�ܸ�5�ɌXP��TJ��"#����Y4�d����*B⪟���O����J��-�`4� 	�i��U�u��g��T��������O��0�G�Ob�ɇm�
�s�������4�J�b#DK�� 7�ӦeΓ_f�(�IٟtsR/)���?1�'M:��땏Y��+�!e�6�߱}*�Γk�<������Yw��3O��Ytߟ��0^nHԸCC��D�\\;p#�F�0���d�j�	m��n�#�Ms#T�$�O��Tń�,�<��bH�Z3�|�7-�Ȁ�\j����O�I�O��	���'Z?������$ ��ĕ�Ѳ0o�;R�����Dy�r7�?���Fj�#,�I�C�	2Y �s��x�!��\'*������6EE�����;�6�'���ߟ`0��l�����2vqFP�kn��x�>>���'��'`��T?��E [�^>���(����% )��`��W�'�Q��Dnڅ0�K!>���'S��g�1=�d���± r� �'�<��aKԣITl���@��6���':���
E8YxҴk�

6y�'n�́C�VU�I	V�zL12�'�����埆o��m�e�յ?�p*�'Ox	0��YLv��i�N��FzEB�'jt �F�/	����7I^-��'�q��Aσ5ᔀ�0�J�.r�3�'Q�(�qh �	�h����}E�Y���d�O��$�O���O��I#�D���:��@���Ϧ1��ߟ�Iߟ�������柘��ß`cT��M�T�@8fwx$�����M���?1��?���?����?���?�)
t�d�  OӢo����l�>s2���'b�'���'���'���'�b���d�B��6�b�xm���Q�6��OL�D�O0�d�O�$�O�d�O���P:xY��BZ#KT��	Sy�0�o��\�I��t������	�����I++w.8�$�/^i���D �Z� ߴ�?����?I���?���?1��?���_�`��#%\4hH�50e��L8V��5�i{R�'���'�b�'���'��'a��Xj�;O ��lZ�S��$�no�T�D�O��D�O"���Oj�d�O����O��9R�ײB�	Q�Eǘ5Sj�Y"��֦������	�X�	�@�	ȟ���䟼Z�aR�@n���$A2pcD��M���?����?y���?���?��?!���)kNH+&�C�rF�<&��ٴ�?��?���?���?���?i��c\�4��5x������
>�5���i�R�'Q�')2�'���'k��'���(Q/§gr�����IǢDI��j�d��?�*O "~����$H¥�e�ҾGR�P�Ζ��M��D�x̓��Of�6Mm�pa!���m�$� ^�X�� �_צ5;�4�y2V��$?q�d�����rm��2�NR�h49xv���>E���	$#J:u�FA�d�(E{�O��]�wN��A�lU�R��)��\f��T�H'��Q�4|���<q
� *���@(>� 𨒌��!i� "��ET}�`�Hl�<�*�ƴ�'�yM2e�s
�r����4[��ɔ�1y���3?ͧ_�>D2^w�d�	�6�X�B���?IX����˓�2˓����O0�}��r^� �Kudd���!R���I��M#c�L~�#c�(���D�MrǂD�:E`�ɖ+ؚ$3���ɔ�M�E�ifW-V�&��0ɖ�ل 9�yT��}�c�b'����� M[¸1`��џ��'^1�4i����~��"C%T�X�`@KU���42�F��<������*m��#p�\Y��QG�1ga��+����{���Ix�O+�|8�G)2���c�,s�)s1!�WN|��O��Sb��JQ� Y�	 �|��Ove������	����pe��Bn�r6Ì�h[!��>�HI��Fd	'CL�<J1O�`��?M�ģgՇONl`���{%�`EN9p���-�H �M��q�4Їk�4%Κ�a�a�t<āq4F@G�^��!+� |h~� �Mw<��m�.����B��Xc a��"d~�[���
u6�YZ���8H�e�G�,��|���Ծk�Ic�C�!��æ�I�iJ�Z�ad.�l�`�Ai��?��4n8�����?I���<�]u��Ap�F)�T�H(��c��nZ=
<牆�M�S�ʧw$hm`6/!d . �$P��6%�O�����'�z=[G�|u���놠.�����'��Q�E&&h�L�5Fj���I�pW�BAP�L��%�r踔��g��7 l�PN�!n:@�FN�lJ܌�7�#�@[2��'4B��eC§EW���S�٫ǰ(��I�T",���5(��m����- j���@ũY�6A:�E� ����Ƀ�ھ�T�8~#\q��/��'�@�L��K���c��V0-�N�sXw�t��+w�����e�D
JK戬1D/�<ѷ���?��4{�����O��	�O(���u���#@m��P�RE��1�Ų��d�O(�l�K�ȟ�)J>!�*�c���X�"��C�Lt�<�p�³(ɮ)�t�H������E�	;��9����d��رM�hH��BZ��`�Q` KwCxu;�Q�nd$�J[�p�D�yuU�-D(%H��D�.�l�T�ʀi+��z\�Rb��H�MT�D��\8�X�1�������ж`��Z�Ɯ�W��q�����o�[ex�"�	�4AS�<؄턀K��Oh%@�$�2/��u)�����hR"O|�g9�:�r�?I�"��e�>y��y�yR�+I H�r�Y7`�d��Dr�|iRC+m-T)R"{�F��ȓ0��y�@�F#9v��@ fp��ȓ �j1a��A�h����%��i�����ruf����+ 8�IVo�	>���ȓ��2҇Q�FP�iWl[?��wP�	��K�Ɗ|��d��Ԉ��e�6 �Ȩ
~��5N�".'JІ� H$��G�mՄ	�S�љ`b���ȓ)�P��"�	+^�۔Ė�JJ�$��9�dp���Th}��ɞ�0�Vȅ�]��Cs�V(^W`Y���F#�M�ȓ���i�낤'��,׀�7Z��I��[�ޱhEʏ8b$����߭S��!��\=��w��3cƜ��w	��G���ȓ/����ː)c�P��� �$���ȓ��,jeG�3yW�T�LD�A7�ȓ �̨:a�[�Q'�T�P?�N5��A;�$"���j�@ ��O�zXd���.ђ�
t��@P�H�K,V|��8�^�oɝ>OT�I�m�)oG��ȓkpq��� ��Z6**̬h��U'�<H��ĵv��A,��I��i�ȓu1�D�e�[���
�.ƥp08��	�w3*�Ӑ�q��{t�Y�mj�	a�.6�zt�E�;D�P���Pf��;�j�7�r�:�'6��ZD�ԂTۡ�h�ś�$�2�|CDLK�z�p�"O�L��,%�p�CR,��
�����r�zRkG~~��;�g}BJO{5>�CP�Ԓ^}��S�#ؓ�y�WZ~�:�k�lp����OYti��gI!P���`��w��(P#��g�ܺ��߯N� ��"LOl���W��z$���x}��%���f��H3��ʻ7`�0у"O	�E0Y>�iZ���X�άX���1Z�ބ v,ГA^��O��%M}8����V�JYf��m�h�<����(VEL!8q�Ⱥ��4��kR����
��U 1����̓;�*�|�<	"h�3 �UC���#t�hU�I����Ĳ^�]���ߥq9x�`�ǋy��u�e�4_��abG�F�p���)� ����/*�$	U�F1y��ɒp�ɇ'AtI	u��)I=�����W	�dp2b��J�ٚa���J��,��h��y��1�����S�腺�)�*�~,C��
6��HZN} ��̉E�T�͈S��U��[z�T��K��y�e�rH�4����W~���iQ��Yw$�y4�P��,E�-�Οp��������Y����P�VE;7�E�(Qa~��+rY��m�|�0�3�[�ݚ"I�q�0M�gaJ�:��}���٬�0=���ޕ U�Հ�
\&�zD9E�n�'�8ă��;�B���/����e�ü*<�mۂJ�"��Е�v!�B�'��*u�� [���0��׎oOq��S�����ȎT�`р��v ��b+���O���3���,`�*X>�6���"O�2&�&WW�d�
J�)���P�d��\"�EIX�2=Ȕ�P�I���+*M>�B�yR��8X�fD�}}�C�H��>	�JQ
�\�0"�R0:4�M�g�h]a�� b�*�!�51w� �j�Q�
� �-a��� ��7 v,�EzBI)p�n�"�)W3K{�M�6/ڃ=�Δ
ȗ�b4"���%F�r5�T�Xo�|B�	/$\��b�R�.A*e�8y�H6���&L`h�j�O�V�z��^�XD
��qbED������*8�p��!?��*�D�<�b/HP
���+ۨ�`a c�h*p�ڴ�-���B1�ׅ5K�\�O�x��5�ɘt��(S�
-KJ{�pq�'�> �rD�r����I�k����a,A�hH�i�c�89����֪��<��D?LOX��VJZR~V�b�jw�%3��Ɂm��Y{�M«:��(qw��48Ĝ����RV�e�'�\� PTUS�6G�}`�'E�I��n�� �0��D��Pݴ	���86@@�$4�C�(���� �]N��5D��^���C����[S(C�	�p��\�GA�(�rL"�@�?U��+�oδ|p�b��Q��kU/�|B��dI;�z\QB�X�3L ��#F�/a~��ϖM�1���]���P2˚&~x�,��h��!�A��$���i
��<$�v"S4^����Z3�UG}���i#:U�����r�N���8游���Q<>���ȓPrY��޽p�����I�e�L�'��k���]I�O�>5���=G@M�DJT~Ɗ�Q.2D��"�+�%�41{�ѳVؒ��6�5D��B��`�R��O�HrAC��6D��#DE�+	���k�J�s}V���;D�| �㚺z���F�6��<�F/9D��!�j�nʞ�[�"U>�8I��*D�0y �.wn���WWf�Q��=D��$�J�+��8V���v!��;D��k�.����X��J;G���h57D��
bWp�@sM5ؠ)x�/!D�d�D��b�`�3%�7z�Y�!�$E9r��3O��ks`��bB1~�!�d��*�J*U$
&�ƌ`Aj��p
!��_�@T}P��I��`ab�iQ�p�!�D
�a���U�gx2\`�+�g�!�Aw2��"/�3-x��� �h�!�$թk��שDTi^��2��^J!��2#O�I���3Ejڡ�mV�!���r���5I��S��s!��.^��9R�h	SM>=:�.�W!���
5N1�0�W�0h�!�#O�5a!�@�����&$���
��B�}n!�DX0���YFH�\�V������f!!��\%��x&�G�G�Ԑ�c��{*!�d& l%R�.�n��i��:!���#���VI��/�KU]� �!��_�^,z���%��!]M|!�d�;6xH�I�*&Z�Zւ�6rV!�d�����!؆@d�IrသZW!򄕘q�"��P�D�a���3=!�Ԃ�PbKӴ_�J�w�ޅp!�Đ3ot���L�:�H8є���y�!�$�:IG�@S��%�4X3��&�!�� ��Ӄ�M2 �b�JG +\�q�"Oz��&��U���jf΋�}�ظ�1"OnuQ.�lqB,b� 茭�"O���CҴt��4,�o�|��s"OXQ�"�5t�yRI �&��]H"O��[�N�֘xΆR�"�(�"O��X��\"s�M�mF�V��6"O�9VmF�"�-+�J�7� P{�"O�����V �,KR��z���c"O� I#�3R��e�3E8U�J�("O���fO��A��N�e�2�B�"O��8�G�8\�
�9Į�*>˸�Y�"OiS� MZ�]�ej˶���ʱ"O��;1�+%���3ˈ;`Eh��""O��Ѡ��$k>�T�TmH!N�>qH�"OB`s�W��٧,�8Z�"O���WN72�1w�^*\���R"Oh5�#��l�@�K2�288\�3"O�}!g�E&	26Lj�,^��ܨRG"Oh;�ă)i��(djǮl��Q�u"O|)BT�H�r�R����ͯ��#�"O�u2S�}yv9�f@;t��Q "O�|C�m@T,У��%��M��"O�,���ҕT:ZP��#��2��c�"O4@ŃP�x�.�`�ܫw�Qɑ"O��T���4.��d�;5Ũa��"OZy��ěgW��ȕ�P��Q��"O����,�!z r�"v��%X @X�!��8+�f�' i�'����a�AKAY1 �r���kq���#M�e�dqsk��l�a�,<��{�N��6��ҧ��B@Eښ@󖉰��L^&�Ȱ"O~��&���}z�+L=D5�9I$Z����i�/2��P�d�h�0�c�/9�X@bU�?��,H0�5�Ozy��P�z���W`L�x�6����� ݶ���.�
} �l���wז��dĎs˄�iWB�@��Ez�-��h�^yz�GJ�fG�'?yӒ	_�2�DU�1�͛X��H+D� �%��$LS�p��΍lS�x g� YTQ��%�bb���V���?E��Jc�DVL�7 ��)RK�X-4���)Ͼ��SS��!1�Vs�`����'�f%�n�U�p�x7ΖHF{bs%�1#	C.8�`\�R��5W����!\�LK�䒴���XP�MI��q��MH�0�
������'"�������pP��/&F�Q�hz�O�%'���Ά�vX'>u��E�����uA������4m0D� � ������*^>g�l�,Qj�QA
	��}���?E��8�N}��I�i��=A6�T�cB����0Lz��b�6P
���JFkb�����%曩d�e��Ƿ2o`�3ړ?��T
Ǭ�
SD.��V��+����	��E� SvF�4�����z�n�L�L��q��W�FZ��?�O��j�!t���1��=�\��s�	B�@q5�ڒ9�B��r��tm�>а�����'&����R��y'0(ф���jR.�ucr�Ӛ�?�"�(�*�b!�7���>�j1�Ҥ[��n�n�,�Z-��I���0�Ͱt��A�g$lz�(�'���F����!��'�J���bF)l�R�D͗0�X��	��mr�2�+?$h^(����^�����g=(�K
�'����aY>gt<�r�L'1���DƑd��#|B��[n D���Q%&���hb�G�<Iw��j���[�k��D�>pëC~�<Y�A�S� s䂠X�h����<�c�L~Ƃ�pVD�bPS�+J~�<A��D;3�����q(��Bֈ�]�<1�h֥b� ��Qf	= �}
`�Y}�<�2L��>*0pd�³G�v�� Mp�<��EM�p[>�C��G$i��hQ��z�<� `p���`� �!���"Oz�J��ݩb�@���R6���!"OJt!�MY8F��gC�Ѯ �s"O���@�r��|��V�.h��"Oh�Ҕ��O��z�嚕'�p���"O*�P��#��d��$,S�<�9""O��+�
�?@��;Х�����[r"O��Zg�G�AHv}Q6d],�z�"O� 1o�D'�����}���"O %`���)PE��d
*[���a�"O��e+�&c@`���^	��"O��,F�~b�R�"�<Z$.Y��"O�=�@���'�n����<0�lP�"O�9�5 �u�ԇV�p@ڇ"OvɸEس h�$K���*����"Of���l��|?�1��	����g"Ox<2��Y T�~�0��K
��"OX)v�ՈEnVz��Eb��؁"O|ٱ�G!=Ɍ�f�v��B"O\��	��a�}´ N<$��"O�` ���e�$8x��V�U'�q��"O�S���7� \Xdӛv*�)��"O6����P=l9<rv��9:��"O���$J���/x˂ ��&D!��.Z����a��$d �m��-�!��ۣ(�IG�&��L�O\!�Ď
yf<�0dS�r Z8#m!��WE�}��O��~�$M�%I�!�d�(t��#v�ɬf�`��K�|�!�$Q':�!��͢�R�)�ِ�!���
��Ad-΋?��=ːkN:�!��	2z�+@	O*E��`8�k\���S��	���;!>�eX񡇌s
6��?�#-��&�!#��ø}��=��a�<����7Hi������k0�PGI�A�<9�a�#L�@y��k�
��e��<�Հ5P�K�A��`K¼yvUg�<f%D�B�i�ug�1(������Ze�<u�.C؜�D.9s���5 �`�<���Υu�����i��J�0@2��Z[�<Q�D�Q��,�"#܋d.��!��]�<Y�"0�p���*�$���ϓY�<�@n�Y�qe� 	ո8�w�M�<auȟ61��D�w�
�Nj@�cM�<���� k�&�iS�ՂEC:@�ዏn�<��D5>�)��A���^-ꔌ�g�<)⦅�x�v�@�P$
�!���Y�<٣��'xkB��bm� 	������]k�<	�G�%�5	%d^4���c��f�<IRқS8��QcX.��MSOT`�<�FMLU>$�q��K�M��@w�<a�M2��
`	7S��Z�M�r�<��-5ki���T)��A���p�<9ҩ��@��X#v�@( �g�m�<�@E8t�������c�j���o�<����8'(�"�"�N��8�ʟi�<a��&v��˱h��0����\]�<	�\("x��M�� �Yԯ�m�<!�Gҵc�\5X0�,G�)�W��B�<�!��%
���&� E�T��{�<��$�.2��-���R�8l�1S ��{�<��&O�ff�9&��;��@�<1J�&I`J�ж
M�h~@Ȣ�D��$�<a���{Yy��Еcb�i��I�D�<�lP�U	U��\��Z[�S^�]���� r���a�Z��բq�A�O�����"O��i6�B�$�7CȘ�q�tAM���'��p�p��>a&�Z�9�,��l�~�L��P$�eH<�RF1g��E�3m����M�`qB��0԰:�NK@؞��hP[{.X��얻] �*E�<Ol�dA˓nv ZW��3B�$$��A8�z1���#��dh���9�y2-�c.��0�SX���r����	-j&���G�=nզ��fҥP�>��䦄k�ڍ��j�(�>-�J&D�Ԡ��8�8Y����^���U-*I���w�����I����:
�Zb?O�d4��!d6�A���]�$�QR
O��fN��7'p|�� : ~�R�H�Sft9{w
ׇ[�b��o] 	�y2�75�(AAĠ�P����Y�p<� ��B賋�
'�����E��Ȥ��%m:"��&��� �Ɠ�T�f�U�c�!B�P�6���O�@A�.��J�l!7�F�*Y���u����zyJ�[��@�F�B��F�	n!�ʈA�5�D�O0du~a�u
I����d@	d�AR�'�;E��|��+z��,+u�$ON����Pxb��&~h��A��~��5b��/%1\)h�Ɲ^���S�M6������6�(�牉?�P騐k�a�x2�D�g���A��R�m\�h��bU�7�����iܼ8�z�[f�1Y�D��\�N�Zs��a
F<�B�W"�x�O�zN�:&/D��#�)�.TF���^��3�˕b�$i�*�yb���4g���M<jWp5)�)�IIwn�>Y��m�f<��e��|r`%X@�qE!�fo��w���Px���"�D�A���Lk�dܻp�d(�i\4X4�9��ڔ�����Z�e�:��T͋�?9l�Q��ȳ9�x��Bo
��!OcO�]�R�ig98�`ױvX�����`�N��'0Pu+V΄R��3�i�I�th��O�U�c�:DF��b	6�'l�%��/
JRp#�(U�x���\����.ۯ+��%.<�@�A��iyRć�Dp )E���{2���x�)���Nh��"����?�6��/T��m��DS C�x dn��`�V(<�BL�֜K�.)�f�H�A�|�'�xYqF$�Z�=������#%�	8�.5��8�ȓH�j�������'���2��ky2�J�
t�OQ>% ���1;"ѱ�->(YA�F5D����G�*z�I���2X�y�H1���r���牲-R���+�*q24�s��lN������mҎ�:R哝P�p�"bkY�P��،�x�H\�<�6�p���1j
���Op��`�ʌV�q�r(�6��"�ޅ���txvi��"O���D$�"
���83�I
�D
wV���W��`&(&��|b�c@�|2tqK�GT�\n~���R�<Yǯ�Ud��4���ȥ�T����PWȤ�P�R�g�C�k�A	v�%�@k L� ��	�d�h�'d�q M�"g��,�ѠOHƐ���AR4��d��t2���dȶ!�|�U-8�qO����|~bؖa�ܓ��\JRNّt��h �Nʬ�a@"O���4Y"@�Nh��2^��URbd�����%<t੠�8�gy��-~�a(q)�x�����,�=�y"��՚T���ҵt��4[uEH#E �[T�YE~�⚰
��?It�C�5�9��ѫ�:����WD��`b��і��S�S >11$�)��X��;��E:�3��?AP/Y��q��R$<`�æ�Dx�p��`�w���s��B��'��Y�%��#Ȍ�s�8r4���v�Rв��ϯ7�r��6	���9a�&5?�e#�*�q����?�;V,"�������(pD'X/��p�~�0J�B�|k�
-�d� ��g��*�OPi�#����2ƀ:�OH4 5��S�^�����1}3�(v�'{6��qD�<!1�O��`��T����a*��u�N�@�{eN�P&az�$P~��	a	�o��)9�	�'V��c��>9/�l�l�'f��� "Q-h�P�f�C����2��M�`�B�ə3c���bM�@�`�/X�HJ��;7�'��Y�_y��=>r�T>U���x��#V瓀m�UR��mm-qE64�|� T� r�ܧT��������@�P0T�$��'�,�J�0���1�!e݅���&�D�\��q`�3uW|�%�Y��yh�5�}
�4}2V���C�fD��rt���*���f��R��	1?5�च�u2�Pcr�'��Za��jUn��e#O�"�N>�m<"�d��U�ja�R��yy�gǟXs@CJ,ep(s7M�J �" �Uh<)TA��	��A0v��ARC����yBH� i�� a�O*�!q8O�u$J��;��
�))
��!��4__&ԇ�T?f=R��K7ddQ��-�`ȳ�'ݛF>OnӞ'�f<P�5�dP��|�	�2R��A#�҂A�p���ۀ��<A'�¢o�ˠ���)SeA�7�ܱ�6�	jue��Ϙ��'Y��� x�pE�$'��!��:�O�#���<q��+񟛶�:I�\���DW~)0!��B[���M/��xS�� �����C\�~����
��wŘ��'���X?�T?�'��DćȸT�f��W�U]@�mQ�'�m+5�W�LNt}Sw��	b�YF�Ζ3z4��L�ןy���O��5I0�0b#�"�H�Z�Kט��$�YH�X �7W�\є�8rD����>w�l-rl�&8p 㟬�ϓ?.`�g��a�EzA�ٿ%�jq&�DxE�ɟe3jp����:�`�|2�	ɒ�f�pPe�?��C��a�<�B�gۖ��0DZ�+�n��LV��Tpy�eI�Oä扎QMd���O���Ć,F~fL��E�9�e�P"O�eДË&E־
ef�I4~�!��N�yӠ��!�-"6�'�y$�*q�Ƥ�S(� P�	�?Ј
5(�"F�J��5�	)Se�u�x��'���j2�<-s�l�[H�3W��<׈O਩�l �9���?1ʶH��t`P�(�-�A[ra;w�7D�h�I[׈�25�XM�V�U�t��q��
3�t&�"~f��2p�T(W	~,�����`�<�&�Ʊ1:��a*ϸ���,��'�`��7���+�:���ϓ��MUR!��s'��bh�}"��"�~=���\�T���C�/q�y!D��T{�C�I? ҆��3��fB��C����i��">�H������Eʾ�ZE�a�6�Hp�W��y�&��y2Q���*9v���	����$ܾ&kd��>E�K�(}�yx���"7Pq��B��y�1,�Y��^�I�c4`	���)*>`2�'�Hy��j?WDR4�pB!��;��ca�x�#.ѡN��E��OS>}�0)Q�8}"���L���sU���3�J��W
Y�Iџ\S��M5��OE���dY�&��k�A K#�a�
�'f8Ӆ��a���PDٯ@ް;)Ot���[!���(�fIxᯇ�,��HKvF��tT���"OVh��ϥ7�b�:�\�j�d��B�|�D�
<���Ǔ*��M X�D���V�x����bꖌ���68X�]�''��1�����M�J�(B�ɾxV�e� ��9�X�քߖD�?ё�<n�fc?Q��oQT�ƥ�W��N;�eY�h#D�H&�3u)�EW�P�����<Y��_&=E�OQ>}3�
�6�Dr�J�; �"D�8IQ ��T��h��Ƀ8<L��#�ěcļM���6cz���F���F�����5�`����zU�҂՚u��\ �C�3/`�A��QUh<q󭜜	��iB抾0#�m�5�\�'����0�S�oB�ai¼k1�5S��	�B�I�~�Z�IE�FѾM��� ��˓{͸E�0��S�q�q��?�bS^�@�'D���E*�('�P�B��5�j�;�I&�%u&����Ѷf���A�M�����	e�X�W!�$��:?j����S���mI?�!�$f�v3�c<m�����62�!�<<^��Aቹ@Q���#H'w*!�DM�o�(`��Z;VB��c�`ڜ !�dI�4���Y�( e�Tʐ��$Y�!�d:�α�+
�7� Rm�(�!�� 8�Btf� �d�rɝ
���b�"O^5�3m�+#���U�N���� "O�����\��@�&+J�"O��C+љ-y�1ACJ�~���"O���6�6�r�c�H�
k�� "O,1�vO�`S�^�W��t0t"O�P�	�5r�x�3�%\��4{#"OJ�!WD���`z���.�+"ODhKT�ӄnn� �
��mR�"O�!A�ԈF�`��!�8,��tk�"O��l��!� 1�$ �3�T���"O�%(�Իp�Z��4�%kd]3�"Oj��r	<J�y�I�<��K�"Ot�r��<[t���h�L-Μ��"O�HQ�c.t�͡ �P�-1r���"O
t���+R�P����W�Rts�"O|a0���d�4�C���;K�x"�"O���I4������M�=��w"O��sHQ8<A�U��*M!��x�"O��,�h�`���3E�^I��yR��?_�aC򃕭jXh9) ���y��(��ZE���w���+�JA�y2'�V7L� rE���&�(��G�y�!�Υ ��ҮuźyU숪�yk�S�<� �NB%�H�#�Ǻ�y�����xd:ע:=�y��Ί��y��.�%�T Ǳx��Rm\�y�.7OT�X���ك�����N��y�"�&$��T��U�0���yrJ?Hz��A!�R�[&a��y� z�r1A��Żl��h�E	��yr@�����S,�3U��$B$P��y"�R8s�L�M��h4���y�e�[�@`0T� ��H��y"�G��E���=G�\zc�Bi�<�CH(����������^i�<Iw��E���D�Hi��p�$f�<1��m2�Z Ɉ+o�qb�^_�<)����\�A��� ���A�_�<�r���vv�5c��~2M�PJ�[�<g���gUly	$�U�v:="d#�Y�<1��!rQ.G�MĭXP��S�<p$����k��W�s"� F�KY�<qr,K#5�uaoL,ODh��D�IR�<��)�m��p�'[C0�����O�<����8\@�zAI F�蘑H�H�<a`
�v��Ң
�s��@ m�]�<����;L^�:�@R9��q�Y�<q��N�IN�Y�"@&w����X_�<�3DO�7Pr$�d"�P|>$�ɝc�<9!�3�6���
_���p� ��b�<)��B<u�&|��NX�����a�<9�.�5T�8y�cI�c�z�� �]�<�u!Lc�0��dֺFm��Sv�p�<�%bߑ)��q���J�)���X�o�<0J�["�вB&ZU��@�,Rb�<�%m��B����f�73\�� ̗[�<��J���ܲ��̅G�kF#EV�<I���Z�\Zgl�8Z���� @�}�<����|�z��G��?&0.���n�y�<�n�>Y^.i�@M�&L�cIHt�<���Ƨ:����o_pk��\�<��MɏX
�%�֮���pP!�n�<!�`Z4}XPhY��H�(M�@��q�<� � �F� ?_M`h�U��y�"O:ذ��s=ti�b)L,�
��"O�!8���А���)�=pc"O�m�V#�',��;s��;FE|�k�"O8����V�}��G�s7�]��"O�P(�F�j/�m 1G�	$x�(T"O�t���Y�HK�QG� '��]��"O	��.7{�@�� �Ț�"�:�"O��{rIb��u"��&Jˌ���"Od�H�A7_,H��Xd� "O�*qFS)#�TM3�%_��X"O�eC�Ño�܅񵯙7&���� "O��)��ܔ^�.��7�D�Z���C�"O�lD#M9#� �N�&��(�p"OL 	�b[��@f�1gz��f"O� &A�.g�-qEĈn]��rE"O�!K�H�>\�D�
��:x"p�"O�Ђ�e�~L\S1鍵0�<M%"O*Q3f	"?e��&�<!s@��r"O,qCJD���@(�,#bz%�V"O؄�D���@S�J���C��I��"Ox�+�n�_��mش&N�Vu|ذ�"OFpaE�Q�Mⲅ��V�WD���"O��QQ�/j�=�rĊ�oqP\$"O(��E�G:�h��ɍ�Qq��: "O�	�f �}����Q	�$m���C"O�!��Z;���ڃ���C����"OR������,;L��E0\��0"O�SD�X�1Z���Ņ�$RtV�`�"Oz(����mB28�U������"OVչ ��m��񓶩�~Yݛ�"OTA���߿x}���)��`< �� "OK��T�%�\�!�G�=4�Z�"O���R�w�`R�ǑX'PT�"O��6��8(L��Ŏ���J�"O����䒩ybd�S�ŋ�!��5HP"O>a���*X�CD#c�L�KB"O���AĀbĠ]��BQ�PpV"O��ȃlxV<���R�{�P	�S"O��2ˍ�O:�����D�����f"Oh�	�aۊ0S�K%o\q��e��"OBB�j&j�`��?:�^�z!"O�H����#aà$��[/&��"O����YU.��Ifa�F�.x9"O6P���5Ms�()2�!z�.p��"O
�`㧛Z�0� $�15� %r�"O�5�Wo}���'�	^�&bU"O�����,�f�r��M� � "O*�TE��w���!oA
d��w"O��! �
A�b��MЂ"O���L԰���2�']	.�zȻ"O��Sj����HD��s%#�"O�m3�@�2 =�c#�JP��"O��q�U�KP�Z�ߋ��""O6uUA
%��T���$��)8�"O��آ���2%�=�`G�P��Lpf*O�Q�%�ȩ��d�wE�'�~�J�'Ӕ�1g@��B� G
\)����']"�pA命w gm����S�'��U�T�#�nu	��Q�(�H:�'b�	��ќJ�[��:����'���AC��8`���i��Y6�x�'��0�2��stk���y��'@&T�� _�<�r��N���[��� z8&��|Jx�)��J�k�l R�"O�4���H��hE*O�q�v"O漺��ͿY$�3�8����"OJ��F�{4���'���	��"O�81 G��+�:�)DW#�P@��"OrȻ� �&f��6�Q�O��9�W"O�	 �F�ap
!*���<��Ah�"O.�*�o'jD�`���7�<�"O6Hy掄����aJֹT���I�"Oބi�hڲp �$� j�@H�%�"O�H�P`]�|���U�m0"�:g"O�`��8zX5@���&�Q"O��P�P��Bd�k�=�e�"O�ͳg�&^�� S
n		�>�y�`�2i��V��;Y2uYGZ��y2�X�i�>A �GI�p)�g=�yR��E��	2T�9d���&O�y"��Ѕ�(=�
Kvᜭpjܐ�'2��۰@��9r-�2f��c�p��'�,�2	��I�IEȌX��3	�'���題˹~��!#'ܐ��[�'�$hb�T)d aS���������'�N1�@K�Jköib�\��'��!�cD�Rp���&��`�
���'6ԝ�+��'bX���äY,Jx�'�6�!@l�� 9�H�г0���y2菶rn��M���j�
���yL��$P�!rIA�nz�l	�y�@�Hފ����o�����C�	�y�
�x��	B�h�V�B��L5�y�B�*KD`��B�Y��Px���
�y����5z$mP���9�hڝ�y��GOo0!`���.ְqz�����y򂐄X�A3�"���A R��y�mY�urC�j�:lƢ����0�y��"~�	��1�B�Iw���yb��<l�~t�	��1J|@X�X��yKŷbh]��+Y>DRI�����yR$[Q��L��I�="����ҧ�yҬ�$Z�����B�#��A*����y���0mP���SN�1��ժ�y"�E�]`N��f.8+���CMX:�y���%@N�gbV����A��
�y"$ǽ�r�L><P,z��Z� bB�I�	�:Q�3eU
U�U	 לt�^B�I�D�Xs�F�88�x9d�GDB�	��D�[���	��!�5�ȯ ��C�	5oP`q�F�ru#�aB�L�&C�IȦ�j�́�\=�9� ��(�fE0D�l2ƥ�x[~uۤ� >k� ��B�:O�#=9b�׺E��Cs.Y>5��h1aOY�<�/W�a�,u�!�H�x� lxÌ_�<���:q>@*��.ޝ)�@�R�<��,i��5&N
�0�9�m�x�<��("]<�k��� �s�DAL�<YF��.RV wF^�&��PPP \A�<Q��D�&��]Z���?��u���Jz�<1��F/ ]̴�-�*���	Q��u�<	����=�hx�ꋛQ�r��r�<�M�f��@� ї|Fv� �͝r�<���@M ��J�c����1�Sk�<9�-�%]�p|Z��m��%K0 �K�<�6� �6��or����s��b�<�E��(0��R;�mq5�d�<� �����R1jb&�gH�P@"O���ܡi��az�D�;d_�e{�"O�XZ�J $`���焉�'H�(��"Or�����$O�)3��Q{;�`��"Oj� �I��A��\�T��u.J�r�"O��A�hE�q���
���z#�Q�"O���kF/�Ҹ�P
U7iLb�"O:-��-3Ac�a��II���͢�"Ob��c���w��y	���6c���U"O�Գ�AR�:b��@5F��}�BE�r"O��)\1,	Sk�,��:D���ċE�4�qbi
�7�!)�L%D���3�-܉7)I8�(Ea>D�HvF,�l�@�[;^�[Ä:D��qK
�8��\P�mك�pw�<D���3�O6>� �	�`V2\���u&D��"��M� x�%�1�Ը7�%D�8:�`�Y�*��4Nš/�Ā�q� D��	�jW	,)^(�� ����֤>D��B��F
0��rՋ��3����3,?D�����C�j @�$�cŒ�g>D���V��R���!_(����Q,;D�X�&Fa �|k#5`,Y��9D��C$o�q AM^7�䩀��2D��I�Ǯ3������UH����)=D��������б˞�|Y'�(D����<��@�a��Oڶ�چm�V�<����6Ɍ�����
�8�j��~�<qEN�
��0�L�Vb�]"1��{�<��	� ����Uc�(�ɂ@�_�<qT�Ք 2��Ą|I<���a�<�-Ƃ /\�QX���+t�^\�<I�o�#/p�bӇ�;9�F�Ҍ<T�ȳ dO8 K�JxAaq�Н-�!�$��G)� �t"&�Ȑ �=!�$Li�XI�D�TZ4����C�!��ُ\����2ÝbP���g<�!�$��%����jK�d��=�DE_�`~!��*0�D`vM|t���eI	WH!�d� *l�x�B�!el�;��?:!�X<$%Hӏ��ޙ{ӂ/P!��VY���
�
�7e��x�'_.h!�$��|���ħ[��+��ݮ�!�$��V����oלʐ��"T�q|!�F�W��-KTçZb~5֮Kq!�� ��}�׉V,Aw�,eMڜ3T!�%aBt�Qң�)vv�r¬ȝ)D!�$^�i�c�N�(æ�1$)��^9!�O���q	ȖE\X�p$�z!�$
[��)u�:9VX�Qp��c!�$�Q����^:
�
��ƥ�Py��H� 4ۀ�C�k"� �n�-�y��:wz���`�Mc�����n�*�yBl��(u!��YJ1�R���y��>{�&�9�����*ҋ��yR*N7�u�"hI-
�"Dc���2�y'�8BH�l	�H�mhͣ0n��yBB�;x������/f��8�H���yR.��P%T���Y�d����F��y��K!Z��C���W��8X�M��y)�N�n�c�.��L,�@�)�y�m�T�8C��2EȰ�i5!��y�3SPy�J�?#�aY�Ě��y�N
ڽ& ͛:���BR�E�y
� �)�� <A�<�C�	a@|9�"O @��`� ��8@¹E:B�(�"O��2��I�"::]�b(QZ*��H�"ODds�hE�?  ;�̇d��z�"O
1���,Vz��U��َy"O�|��ş-V���T��.�"OF��i^.��p�R�V�y����"Oޅ���7r�&�
� ��`��)2D�@�gG�)՞�*��].'�5J#�.D�\ZM�[J�1o�8&�ɋ�.!D��0 AJ]e6��t�MZ>�z�d#D��ISOŵb��tˎ5 X3L D�t��_<s�щ�؝^��Y*=D��t�)
����%��iuvꆍ9D�\���ń$�n��2�EY{�0�G�7D�xX��@?:�hi���FL �҈6D��3��K15��9Z��ͽ~��-Qc�!D���d���NTP�)�L�]K��:D�بG�M�Y�f�R푻|�A�E�$D�
r�_����U%�"R�B"D����7|��P, /���s�?D������� �+��Z"�����=D���!N�$a�l��.�d�v��/;D��@v �q Ӣ���Z���7D�|�F,}���UdM�J��Q"�9D���Ph�.n]y��e�d�u�8D��Y�c�;4�ΌcV'h�8��W<D��a�b�[����gP�{���N&D��q��	Ls����5m��L"��8D���b&$!��d	��<��P�d�7D��QAK?`�
A`��� >��|�E6D� at��
-����p��m�lk��5D�4����|�����u�=��2D�\�����3�~�6t�ڠ0
1D���j�8˸#�+�]��i-D���&�<[��HhrI�#2��\�B�?D��@��=��cv��`_�0hԅ>D�ع�!P�6?�{ej	1lafC"�;D���4
�-s�	���2�0��%D���gȎ>0ͤ�Z�ê,ܬ�B�>D��#�3HNDY��T�s��(�k;D��S���_'4�k�M�9	����.D�8��)�Z�r0�T,Q3S��h+D�#���;[��hSC� %g���/$D�DJajF�A��!�#_s��sn-D����IM�H����VJ�%�b�HS$*D�(g+�%%,n(���ӗi���g&D�P���;�0��T>'�^%�tm9D����!ŌLՎ��G z+Dݣ`d9D� �a�7� pC��5!��U�<�4 ��8ҡ&H/[좤0�˄O�<q6�@$s�(�n�*K9`�NQ�<I#@ȅ[1��.@=�"�[��IX�<-=�� �n�?nX��%�!��B�-��4�@�(h��Ǘ,s�
C�	�e��G☪a��eat��G"�B䉐gպ��tē
 f�+�V fC��4���ڧ&�X��A���X�V4�B�9�Ph��I�)p��b&��"p�,B�	�l� �z�ǿ1�4�g�W �ZB�*(C� �gა��D���>B�I�i�@ ��-}��e*��C�$B�I�J�����)&�,��L7Y�C��9h�d�R�� 6x���ʊm&lB�)� ΰ�u(��2��|�0�J	fJ����"O�xX��1�����&T I>�(9�"O���#eZ�a�����I "O��AW)-K��A�P� X��"OƕtF<Z��0Z#$�zJA"Oz���7$!��1v7�"q "O�X���FD��5��d]uoD|��*O
�q�R+w�����⍬�Ի�'*P�C�/U#+��]zBLҷx>��
�'Н��iV�iH���q�E�	f��	�'Vj��d�	��ы�.���t)p	�'��iZ,�J��3�c�5c.��'(��xd����^<j�zb�'pĕa䢔�lB��� �b�6p��'�v��g��6 ��M�A�;F��e�'Xv��N�[�hY���g����'��}��i�zW�5�W�#�
�+�' ��4�[�'MP!a�j	E:�x�'�.h��B4?���@B�)�}��'x�9���Y665���U�]ThEi�'��QS�J��z6H,B��:�'H�� nQ�
%N�`�
���yr˂<&�\S`�G\tH@A�	�y"�
��c��:ʼ����y�U+eH�Y��I�:�� ;����y���n�f�����&�HR�P��y�BF�H�4Zc&ȟD�4,۱�� �y�
1*���H�k����`/��y��[4Ȇ(��h?ⵈ0�B�yr��?&|�Y�D=5���w�@3�yB/V�Μ�C��ϧ�F=`��y�ɓsid�X �q� ׯ��yr�])N���k$�H�p"�#i���yB�	�`��0*g#�q������֤�y�E�*.>`�cB�X��}�wGĳ�y�i٥d՜$i"��9U��P��2�y��
Z>��s#� OΠ�����y��&�8IM�8Oܢ�Ʉ����y¦��x0Ӑ�<L\�a&N!�y��qL^l���K�9� ��d���yR�Q�	`�af�X�<o��d�O
�yr�ȡd��(@!F�!��L��
��y�d٧t�xE�w�[-�\!;�Ż�y��&<jDA#3L��#�~Pw�"�y�<?��5�V� �\D�O>�y�X�(
��Y?;K")1�%���yr��6�8r�$I����m�	�yE:-�����Do �j�����yBO^2h�Υ[��,g�й��E9�y ��&���_Q���8�y�$�^O�A�Z�Wcd�aD	Y��yb��=�����U�M�����y��',���cj��R"��k��y%��#�*�#gC�D�>99rʆ��yb�J�GQ<�b0�]�n�^\KA��y��ȕ ^,��b�2j��x�!F4�y�d9�^m:���c���E/�y���:O���X���Z�N!�@����yRMZ�w��B��CT;Z��G�^3�y>���p�ެKҊdY��N��y�eX�^<��[�H?:ȳw�ڴ�y��ו;�X�86��vF虪ƁQ�y"IA�_��P�#���glxE���
�y�C�~���q�ι5���H��ʂ�y
� j��q��bh2��N�SѨQ�"O�aʴ�/tv�:�&� ���"O"!�	�;~�ּ��n �T�(#"O\)QV�
g�����-��N� }*�'q�A�h̯#@�'.��TX���
�':@a�
��oL�TLا@�T��'[$(*�ЗZ���� &�L���'�DUK	κ7��aB��m*Qx�'
*T*��t�q)��m`�'
�؃�^��� @�z��"O�%��E7N�x���I$Y�f��"O
�
�ՊnlpQ����R�is"O��x�-��)v�T�Ԟ��1r"O:T�UO�>X�Z�jӵo�T��$"O�	(�iL�g,�@�Q^�(��"O,0;s��"/�m!�댷9�11"O�8j��Ҿuj��A��ԧv���K�"Oְ� m�8kZ��bd�	�~��C"O(9X�hR8����^�5trk#"O��1��Sn���:U�ۊy<K�"O��t��38�`�alX	g�R)sQ"O"U{�lÃK�R����*��X2g"O2���uZ����H�0�Y��"O�e)��ޤ"Y\q��K�Na2�"O\t���I8L���[rG̶S���7"O8R�·Z���E8==z-a0"O&�@#��'�dA8�MB�7�屔"O0 X3C	M^d��qM۽[�"\�5"OZ�{d���{�U�c��/]���k"OV���J,S��H�!F��Z� �"O(�if]�zFN�u������"Oލ�Ѝ��dw�����b��-x�"O����"�`�����wF��"Or�	�'̄7�C��(� I@�"Ou+â]�H2r������}��Գ7"O�Ȥ擞�ԑ��	�5wf�`��"O&�(�-�b��%��'/b�$��"O�A�aXzND��q��G�I��"O�������`R��f����"O�M���,w>�]���,l$�s�"O֙ Q&=a65����Z�� "O����GU�QV9G�d �a�"Ot�(2.O�N�:Q�1�����$�t"O�<SKہ:_fi0�T>����"O,y�����j��#�������$"O�}�hh.%j��e���J�"O<t�`�=]HF݊��z�v 	"O>M8ш�
PFq�w$�Uh�h�"O,�R���NR ӤB �BB��"O����5�T4�ޝ9�	�*OVd{!��?Lr��-�dx蕢�'~�p���F�qɄ�۱���\�2�q�'��h�7��5�ll�d[��H}0�'�vM�""Nx��<��	_�Fي 2	�'�p!�Ď��X����l٩A_V9��'�]�֬�<e�lLA`����3�' ���F��3@S(Ĩ��,~���q�'�~���(�20�v@ �${�y �'Fƭ�EN8��9X��G�u'D��'��!��.X��nԺ�+׀_qnt9�'s0��P��`��8㮇�U���'�2t"��̑gCfe��@�6Otd��'�A2A��?$�!RnT9E�5��'a:4�&�<��1��C �MG���	��� qS`
=D
qsr� n��xʃ"O�]�%��C����L�5�.��"OnB��#'��2��+fv�P�"OL�d虍-`���dH�;1h:D�"O���G=�:�P���gP��U"O(�j��ժF �o�(T���7"O6�p3�^�\W$���ڔ)��U"O��8�K�@�ە�/��TP�"O�I8``4��ũ��5Y�n�0t"OZ���N�|�*�0��$�����"OJ��rDT1e8R�!�@�+\����U"O^8#奙��@��切�d�dH�"O©���
L���Ŏ
;
K���"O�(����� �LB�MDKE�q�"O�i�&I,b��BW�Q�r\��4"O`�p�e�z�HTM�,JL�p"O���S�VH:�	��B:����"OT9c���<�A��A�$C�~��"O��	�ɑ#N��E� h:
�ه"O�Y
 � b
����ՊM3��ѡ"O��e֘jS>����#��'�y≙�]�0YӴU9r�K�.�+�y�A�k���1#�μ 	̽aaK��yr��XGpQ
碘5^�����y�.�i�`�c\�NhQa@���y!X)�A�|N��Bh��y��\�*�Ƥ�$�~��A��y�%�8
_�$�#�43̒��0��.�y� �(!�R�	.9` �Q IA�y���󠉕�9�^�I��9�y"&��w��z`F/f�ƀp  U�y���{��R��[.3"����ny��\�!���UQj�#S�����dXC��Dk�E�)�p5��Lʘx��/]!}��⒣��4H�݆ȓO����޳C$,a*4%��t�ȓ,%&L
$���"BR�:���$D�4���`��Ú>��tpA�"D��0�(�+jH� ��X.W�D	Ʉ, D��umY���i��ׄN̨�r�=D�@���V�f't@��H�5��xr�+:D����O�k����W,� $O��	pD,D�P�ehZ%���@�OY�h��Y�#�/D�x;mC6�\�9�e�ފ5c�1D��Pǌ<b+@��n��fH*��`�<D�8�s��V��y -V!|�fh b�9D����d�1F��Q�WB��2��3D�8�gɼ3�Rd*��V
<ʜ�C2D���V��+J�Ҡ2dJ�QZ�@�=D�<
d� �1z�Q���
64la�� D�\s�C�� 
lQ uF�/a��tv�9D��a㮗,a��uB bH7Xh�xzЉ:D��p%�JJtdZ�nE;���p$9D��S���T�(C�Р�6$��!D�,��-�2�mE*`������=D�p�Gڃ@��҉��
Q�-��O0D���Ʉxֶ����1��Y8�F)D��a_?����iQ�-�V�2��3D���� �|�8���Z	`�|m0��/D���5Oʩcж���C�X�)��8D���cܒ9��\å���_�V��7�5D�|��EϚ#��m�'"�����s0N>D� QEf��~��u���5��(q1=D�|Q��� Vz�����a�ʼ��:D�� X�B��4'����fL��~*&��"O\�;�"Y�!��rJ� W��z�"O�Б��5@��0��"8y�D"OX��G. Q����6 ��"O>̘vH_H�b�)�2��� "O>�1�U
bL��Ċ�P�r	I4"O�)A�����]��'YN²���"O"�:QfD�(�P�HC��#"O���&ɏ �`���G��8;V �"O�z����JXq���)t2bE�"OrE�v�ƴ��Ҕm' ���"Ob�؁JO�N�Hab�+]�v����"O�Tz�A�7NB�Ǡ�)��b�"O�8���8]������G�O�<%÷"O$�;��V�H��S�܊��u!"O�����"Op,�2䉪^Lt]bs"O��xq��d���Z�d�)V-��*F"O����nD�K�R��*�$��@�"OV����ͱ4��IB�W�7��A��"OL���N��Z[��A镭E��L�`"O�$
@o�2��VB�4�ȃ!"O�S��<_��r��aUl�+s"OpC��X5q'O�S�Ȅ�R"O�ݳ[!���"�ԑG�콻�"O�� #	Q<�����C�}��ɵ"O.��Q��! ��G�Qa�iJ�"O�I���͉G&�41g��%A���"O��� �Y7�X0� ��o�r���"Oh�vn�+�z���0��-��"OJ퀁�!\��&��t��i`"O�A�sA�$l�PZM�f�b}�"OBMse��(g�S)G���l�"O���G�4�i(D��+R\P���"O�k�dB����'Xs@�<��"O���M�)2l|��&	�y$�"O��&��TN &/�k��k�"Oذ����G�I��O�X�Ң"O�#d�"-�V	:�-L	(��P��"O>�I� H_��s���_u�q"O$03%J�>p`�%��(��q"O2���J��c"pj��7���s"OBMI"D�R�~��O��n�ʽ�V"O�p(&����(5 ���]�Z5b�"O.ܱj��{0초�NM�,��8�"O��Y`�Д���
;����"O��r�+4��52%��XH���"O}:�㓽:����@�#i�0��&"Ovi1`�'��2���h�A��"OD�{%��+\X�2�ܚY��!ٱ"O��;��H�Hu�	��j�
SL�}��"O�:�KR�g?Z��)�0A�85"O��@�˖GήxJ��`��A�"Olܑ���J��3!J�K���""O`pA��J:T���"SE����"Op0@�@�=n6���p��*o��,��"O�1����R�b�'V�ڈ�u"O����m��̱��M��x�03"O,,)É�*Q��$@�ikxr"O�$��%)��b*ċV�X�3�"OJ�1C�N
	�>�)UIS�[�R���"O�}�]�6�E��g�(�:���"O���@B?��@^�F�xղ6"Oʔå.�V-��dL*b`��@�"OV���G�ed����,U޴�A"O� t�ɒ�	��8�Q��ƞpqz8"O� (F��0�T(���Vq��"O����=FOtĚ�&kM���"Oh  ��	[|������E>�x˵"O�Ћr)�~��;Q�^�F<��J`"O�U���*o;��(0@ܳ>)�ɪb"O�)���O������Bq�d�V"O:���%KA����g�%o-�ͲP"O� �Ed8\��1����NP��"O���U���t׍T�/]`I�@"Oh�`g�4+4r��ǌUkCt��"O(��@��E�E�P�y'"O������?�v��c@�!�Du��"O���V��=W����/S�0���"O�Q!�'���"�(�F���["O����I�Uȃ.#�yS"OR��ѧߓF�����	��M�`"OV!��DX�zp�%������"Ob��R��s�\`c��D��}�"O6=
tg�2wG,4q��?n�rq"O*TQ �D��yP�/�6t�ZQ�"O@��c�NB~ّ	/�`0"ONqC!��!Tk�Ģ��	H�)�"O���ť�"/��U�3.şB����"O�-��;ȑ�AM�6p���	a"O�)�L]�"�P�4,(0s"O�-�0�=ر,�7�(�q"O�`�!E9w
��D�o���0"O�Hs�Y�<%|<y��] +�ԴT"O�iS�7 �T���50��P�"O2u���8)�lA]9QU�1��"O��{@��^sh訴"� A;4]�`"O��;� *��V��/���t"O~�97&הĐ�xT��A��q"O����#ú5��e�F�Ҁ�"O�Ѱ���OG�I�t��]�D)�"O��c�:)a8y�f�;)�z7@:D���섧8��u�$̈������7D�r�բ+|(�!�t��t� �7D�\��\�y��p���*db��+4"5D��*GeS�y����aD
�1�ѫ3D�  �A:.є�Z�.%*�ziR�2D��gA�
  \b$��q:�k��.D���4�>%���'��Vn��p�E"D�$�f��o�����L�PD��ڡ
&D�hZ��U���B¯�	.�\���A$D�И��ɮ(m�]��H�><�#$D�8��$mQ����K=$�����B!D����h¶(���+
)�����J9D�̂�E�6��y:I�k�(b"K$D�ة�Mm�Ĩ�@� �H�ar�-D�|X��q? �YE,\�q!T��4�/D���dO�>z!�C�&$<kq,9D��#�<)
�e�$t�ⱻm5D�z��є��Q������e�o7D��#BN���a�%��w~���+D�88��M�1���I% M,n��;D����OK�校c#c4v�H�4)9D��Ób00�9ѮJ����Ў2D�\#c	X�)�Y����B��I���$D��ң�0���'Z!�rѱ$�'D�P�f��R���;�>r^HX+%D���&/�=���R�EQT\��0D�h��ƜV� ���%Z��@��*D�� F��nqR`Q��/�B7x}��"O� �'�/U�$n�)T0`�@�"OP���XZ#6�*R�����G"O�����S�tT;�+]� �p�3"O���À�9�v����"�\	 �"OH�"rE��<��@HĲnA��I�"O��۴
O�t��!8vǑ���`"O~a`���ld��F��2#�Y+�"O���E)d�z����O�3�P�S"Ov�B��-}� �@�T�ޑ� "O�Mv��P����u(H�_֨��"O(0��ðO��D*HVke|`�"O
�sMO ��ѕ&˪%[���"O�An�6<Y P��Ĉv ��3�"OH9*!J[> ��e��d��{u"O촃��I.m&���	'��p�"O`EyecƝ|�L���--�v��A"O�1��	cXLR�E	0�v	��"O@��l�8�,x����*T�d@��"O\�r�����R݃����u�xۧ"O��Y��8H����]n�X�"O��Z�!�	<$y���x�((�p"O�,�'��4z�"d��J�+����"O΁qĆ[1 ��d#�E�~�j"Oj<��bU������g���#"O��ӅP�y� �Sr�B�L�ç"O��1M�<�P��o����۔"OT��l�i�\�.��*ܠЇ"O�1!#B҈h�}ɶ�Byʥ���y���iM��*cM!)H6�:�O��yO2c�$� 5�ݞ(0��HAL��yR�	/��x���otU�F�2�yr�фT�I��'jᘒ�#�y�Ϟ�d�2#��| dL�fΌ�y��L�Ez0�����j�>ٰ�����y�E�&O@����7MK��gbZ%�y�K%��x)Ӊ�7X׸=y���yBCF$D��$���@�R��q&Ď�y����h���H��X�B�0�N*�y�ƀ7I�
0+b,N�:�C�[��y��_�HŪ�!�J6n妰�2�O�yBE8R	�}8D�ۓr�P�2��V?�y����ջpA�"\��	�Ř>�y�A���0$H �=1��U���y2�H�t�E�'���_*��j壑��y� �� �ђ.��h�~(R�i�1�y҅^)M���hE��oF�=U�A1�y�"�~��舰.�ijNYx����yb���d|-��@��_�t+�F��y⨑&��sÌO�^����$��)�y�A݆|�TX�m�&]X�UK��P��y��8"JZ��D�a�M����y���d��y10�\�)'���޿�y���+b��p��
-`1�R�\��y�_�M���V���nN�9�	���y���.84���B�f���
�<�y���<i���$f�F
u"Ԥ�y2�Y�a�p!�
�%p���*�':����I'YxLpH��
v%[�'�H�1��a�,��G��Т+�'c~��lȷp�`4rÎ(L�h�'Z�%) C�	c{^���E�1 �D��'�t,�� uW��d�сL�T�r�'�aIp�6+�ҥkT�E6Hp&�x��� (X�	A�@9�ӈA�K��Q�a"OR�w�H�5Pr��a'|��Qv"O�4���p"(�`؆��AP0"O����׸d_����%@+I�6u"Ot͙d��ukZ��DLe�����"O8�8�e��)P41�Se��u�V=Z2"O��F�A[��!�$��v{�\��"OY�����P@�CDq�"O�f��% ��TYt�J�KB\�f"OЄ�I�����e�
:�H�"O�d o�`�L7�	--
�A8�"Oz�Όm����Gͱgy �"O�]�WE\�T�����uq
���"O�I��`�"d� �òG� I7"O�+ů�0a�4Hr�í	FLA��"O���&mՍ+ŪM�?,T�at"O�0[5���\�-��e�4*E��b�"Ol<�HP{��@���Y��D�A"O�ݠ�)�<��q��
�x��|�"O�95aO- �	���G�h	�Q"O�т����{Q瘿&�,�"O�I�¢	=���1�]O�ҥ�3"O@��s�0�dL��HS�R�jI�"OXeh��7ᐈ#sh�k���"O�Q ��[6yZ�ɳFM?�.� �"O|L#d�?�`P@S\�>�-(�"OF��+эj��ZR.�.�\��"O�5��q&�p�&�	3Nz^�[e"O�=y� �,.��ъ�Ej��t"O�l�R�U�-^��j�\%D/�A�"O�D��ȝJ�*���������"O�H;F�xg�\Cʂ�x�!H�"O�
�ڥ15��b§�J_�X #"O�����!`9xq��	~�l��5"OA!(M'(�z䁗���uv��"O6=8���6}���S���7b���"O��G�To���#EY�DA��"O��C��QE&�X#�_�b�xB�"O�-ـb�:>�$�q��׆�%�B=�yR���
���P]��@��: �jՅȓo찭SuK��~��H�;ui�i�ȓ t�8�s�7[�=�P@V�x��x��r���֕j�2p��hŅTH��ADL�%"RP���Mg�݄ȓH����-�}7�'K����L�)s
+�.��2�N�M>8�ȓ8i���f��5h0�r⥒��ꈄȓ:��5�3ģW,�5��c����ȓ<��!�B�v�I[�e�~�)��m�r�"�Po��kAnڢ���ȓ<w����F�Pj�1�a�"d��B��@�x��0 ! ϐq�ԓ8��B�	�%�Z1e�M�T�b��'��~B䉑#��ѧ/U8`a*��ð. �B�ɧ�~� ���(6D͸���i�B�I�cC���d�;��$����$�JB�I�T��d�QF"ld��랄`4B�	�[Y�
�(ۺv� 5��u�B�I�Q@�AG?��x����,JeC�I�*>m�C�1��c�k_,G$B��.k�b��'	f���K�j�l]�C�IXi�fgܿ&	�q�l��	��C�ɔdSd15M�JJ���t-=\�C�46�hei�..�<�θ4sB�)� B��g̊�f��x�Yl$��"O�Ey���eR(��uD�X� �Cb"O�$��o�����@�
� ���"Orh����g�H�Ba�h���3!"O�xBAR9}�8;�JUYh����"O�Y�p	��bd��� C��`b0�"O�7-�<"�"@h��Dn��2"O>Dr��m8�Q$a܍d�p"OTtS.��N��mz&�G�o}L}�"O��p��&Fp��;H��-��"Ob�8�Ɂ�b�<}j��Lw�"O��'`9t��$�poT��UȢ"O|�,솄�E�-� �fH�!!�DI�Θ���<@,���F�("(!�d<��k��M>nI���+��X�!�$M� �����g��v:��Љ�!�d�.Bd�c,O��;����!�?m,V5��f�7,��J�T�!�$��eX�a$A���Q���U!�� %Ô%����$8~�a�� �!��	s�U!1$ �{a,�9�bUn!�$��d�r�θ	F�j�Aݕp�!�	�.��c�DJ���P��!�$�iN�ekrtC8e��`l!��I�gb����o��<J�a)Cb��!�d�D,�D�aIT= m 0�x�!�nв�fD��H�/�:
�!�䗠�>�4� Mn
�j��,x!�$��s�K�Ĝ���a��\�uL!�� R+Ĺ���5}��ʣ��.$!�Dk8�����$ZtN��%T��!�$Ɍ ����%��OY��A�I !�dP�rR��0�T�]Pb|9W)��!�]�d/*0H@ud�a�䮔^�!�I�wM\���!�/Zء�� \�R�!���	�L��郷SMd8aB�ͅ �!��܏����ʸl5�1K�
��_V!�ċ�N�؊%`� k0�ȉ5��#Tr!�DH'����R����v�P�>l!��Ż0��w�@O�}�e��[d!򄏁YP��􎊨7����\�bZ!�d°�T���m��hÃ��70N!�d]!E{���D��f�D�Ha��a!�$�,��<�!��fI�P ��%!�N0-j����u��	� �$'!�H]�7�U�l6YK5`�5!�d3A��*Dfȭqt}�򨕅N!���&aR1�EgB�Gʠ��2�,�!�d��G�OD��X����5/!��M�bͤ�귣�+c��=���*\!!�=�b��g#�*4m��� ��A�!���Y*CE	z�DYk�!��TȦA+��ݷ|�t ���Ƨp!�dìN@�h�[�i���^"I����"O����E�%t�A#"aĔJ�"O�e�T�N�4X��(�j��"O丘CO�4R�LqЫd�@A6"O�=��M9h)���A��,� X1�"O�[T%L�^��l@�i_��2��W"OX��2� �t\�����G�$��ԙ#"O> ����N�8�a�*vv�sg"O.���+Û]��#VoZ�g�{�"O��jӠW�����-K6|a�1y�"O��"W�`�Vi�2��OP���b"O� �d�M.��X���jT0��"O��PnH�0�6�A��29=�!`�"O�f�.`ʹ%`-ŧb$��"O��1��a�(��K]�2t�"Opx�Iː~�H�1Tʍ�`�܈8 "O*�r-[�7E���@�Һs��DRE"O�l��l��8�����й yP�`�"O ,��B&s<�Y�чK;�	��"O���pG���`�CH�(�*y:�"O��CF?��ɻM�lt�Qb�"O��g�cR�����N�����"O� 
���l���ö�S�tU��	�"Onm;F�W�z-�X�5ֻ��R"O��a�o�b�l�0�m�&Uµ"Oz]�CM�
�A����>[���J�"O�����&�X	q��Ј0"O��e+P�5C��FJ�K"OH�y�H���D'�~�i�@"O8 �D�M�~���뗚�h�kc"ON�)���w%�1��)D!;/�ya""O��!㒍^���zu�6p�`��"O��ÇAT�-�*}�� P#@8��sf"O*m�dL�*:���d�\ %Ҡ)'"O�9K V�^��A���+�tٱr"O�	���ՅR�*�`��
�H�B�"O���K���a�� ����S�"O�8�`+Ѽ(��0
f'O$^��)�R"O�mj�)ئ'/��El�\�����"O��,�$�RBE��g~"��"O�@�.ޭ\�1D���"O��J&A�="�%�G �p
`"ODmR!�^`�#Rm�0V^�AB�"OT��ɽiZ���UX~��"OX����a� �����>9P@�"OP8ӂ: �P��A+�N'���'"O�iIF�W|��E��H))��"O���F��<�yi���3�T1��"O�"��J�Y{$�x#Ϛ3|����"O|Q4�[ "WHlж�E�l�=I�"O�A�I�*ȉ���ߏ�B6�=D�,�V ��:i�Xr���u�"�8D���A�;x�б�&U�+&vEyS�4D�\;��3e�HHH�NTc�"$�T�.D�p�!%�" �a��ε74��� D�L���װ
�!�6	�C*�AIh>D����Ǝ{���'Ǜ%
w�8D��Xc�JA� <·j��s3�%�@�7D��Ӑ�^�1�  �놽::r]�Q#D� ��,9Y�r8��h��J��"D�x���/�&�J�%X9�R�q�	 D���@OK	(�&dQGֱX9���F1D�t�S�גj�:���cɃ/�W�#D� ��b�;�@ H���	)����#D�h ��Zb�]8���7:ך���&D�p�lӺct,�� PW�>��e D��*&k�>Q0��l� yځB��?D���V�S�ِ�a�ta
�H��?D�8H����o6b0�BR2%F��<D��1͜ [Ֆ@� ���0R9t+?D�ԋ��\=�lt�`l��o����;D��)��	�J�NrFm��4f}���9D�@��
HAd|�x	��b1�m��<D�D	��6Ǩ�(�0]�|�Еc;D�� q��Z��z��ht�Mc�-8D�� ��3qHN.
jFi�4�Y4ycҬ�"O����(�G�Ii�OW")Mf�Y�"OX�x��<͐�$N��b��D��'��D.ib|�
�,^x�@*���B�<��g-P�񔋃,�t�a�M�Y�<� f
.�8��Ί��.p�3`^j�<�p�>Ĭ����y�i�b�b�<�a��;{Vء��� ���h�@H�<�Z�4-2׀V���+��
�!��B�"q(�p�iZ�4'�x!!	�6}��B�	'SV��h�oSh��y"� ;^�B�ɇ4>�J�)ĘE������:��C�	�'�����J��N �#H��_9�C�	�"��X��\�EYLP8s�Q�y��C�	�)@�9Oܭ~7L�i�P6�B��R�p���57j��T��,�C�I]���� �hN�1�v��rޢC�	>C�Qt'J4r�t�X6���0C�ɬ{�F��B著b��c��x�C��3����@ɞ���]kQ��Fh
C��#�:dJ0N��V���R$$��]	�B��'.�U:W�?�qA�J]�mo4C�I�GA"aqP�D4.@8�Zej[�y�DC䉚	%������8z��3s��jC�(:U0�xU�L�X��V�>�&C�I�|Ǥ��Ѐƫ��&F��v��B�	������&a���ڐ�֣L��C�ɨUL�Sb�3 ��l*�(��C��(	j��l�2�s/U-�4C�	�*����a��0[a ��soƈv(C��B�k�����|�����2��B��ZUz������c��yv.C�o
&C䉺|�v�4"�!��3 !�.7�.B䉆xt��ZD�{��}�D�=%1�C�I1F,��(1��w�aG��q�C�	!��օN�?��RR%�~|XC䉧BF�Cr�W�Q�������44��B�	:1��+7G	/_�I���
��B�ɑT�@� � �8y�"��d*��y-�B��?��T�2�R#�.���m�;
�B�ImF9B @��P��I��A�4�B�ɦ TǩA� R��A��E4fC�1z�:$2���)�\,p�_��HC�) &5�e�J�>����)��M�(C�=Y�\��m׸3d�����#�B��"^�J��r"ƞrϐ��e��C�IQ����pN�&ت�"G�Xl�~C��>@��uv�S=���Z֌�b!�B�Ɋ%�l���c~�jr�׎YC�"༴��˄$DCW� �|�C��/�Lj�Ϟ*P� �h7'�Y[�B�(5\BA��a@'xY>٘e`�SY�B�I�l0����L^ >D<�1�+]�B�Ix�8�`�dA0$(�U�ў<Z�B�I"I���4C@�.Y�r�љCC�B�	ah�dfHʟ|� ŋc�N:p�B�ə)�� p��P�%D��1�/�-�B��n���ip��/.zL�qM\�q,>B��g{�Pr��-f�QJdŌ�`�B�;Bǀ+%�Q+6���Aɍ*��B�	?�4ɷ�	.�h}�Rjϕ $�B䉮|h��$,Y�t�\Eq��M�9�C�R=�aj#���m����T��C�	�%[t����.��А��E�pC�)� <L�uΜ3P��6�H�@}�"O���F��-)8���E�,j�st"O��t�M*���
�1>r�"r"Oha�6 �29q�NP#��T�F"O�@ga�lo�;0��b�Td�5"O�2�d�;: ����%a�"OĀ��d�*D�rm٤�t�^�"O*�N�%,f�K�&Y.b�JYAA"O��`��@�q��$��U�0�
�"O�1U�ܴ?���k���Y��0�P"ObA�	�vN��#�q����"O~ԑ&� p�T�P�A�3}(���"O�uz�B�#��1˧�T3}kd[�"O��YC �+�Ve{�M7|��"O��	F2OH�l�a��x�$���"O��j`�>!i�}� D8�kv"O��3���j���;5�i�"O�t��ř���A�D+ .TAD"O�s�m�>g� ����?V+:Q�"O�8�b ��Pb�;!�*LsRɃ�"O�U�BlR*��R'ebd�8c"O�%�w N��F� oG��"Op���
�4z4�
�C7�T*�"O��{�\�v!�\h��_s��)�"O�0abȀr��-A�458��"O�吠̚��&(�p�ۑa޼�A"O:����@�vgPm���	�&��"O �"��W�NY��ڡV�t��"OT�����y��9�Ă�7Z�&Q��"O��`�	�$8�@�j�&�7v,� "O��P�[6pΘ�"u�@6|\F-��"OB8QJ��&� �g�#G��"O�T�DB�� 4�ea��r� @"OȈ��$8��z��UkT�Q"OA���y��j�[R���"Oj������qH����l�6P��:�"O-�E�Y<2�� #���*|;\��$"O�a��胄jyޔjW��j��b�"O�%B�4[��A�����.�z"O̙�"b�Q��=b�B�����"Op� �F��t��%�T'Q;ӎ�SE"O�d;�H�$b�=�g�	+�L`R�"OTݳG�V2ŀ��ጒ�p�xH�4"OD9soפ��J�Lߧ~J�-�y"�=���t�
�V���@���yrd	�F"����ظ`g�C ����y�c����:B�?*yRQhV�?�y�����]Y���2M�� d�7�y���f��|i#Fش%5d尢��y��ږwS�����F�vP���y�Đ�e��H 1�$`p�0Rę��y���2G�8�#RěXÖ�Z�`��y�`�%[u,� �@N�(]�.��y���-P-!A�R�Ry�hS���yb�6Q�,=��fV�QZT�⃎��yrT1D�L�#E�H7�<�K��y䍷&��@�����hG
ފ�y򫓅g��\!UG��u����O��y2�R�{� Й�h��oT����N��y�Δ+5T9��g�c�̙��`ǣ�y���(_k�Fn��Z���y��#�yBk��t���G-�N
J5˥��y���Gv��K��C.} �uau���y�&��[�r��W�_#n鈹C����y
� H �`��q� m�D矘;��y� "O@�3��C�*��5����67�b�"O�� �I�t�T�9��[�+:�ux"O��Z$I�(Q
	8LX1&9(�S"On ��(g�.���ѧ2���"O �a¦[�'_��� Đ�EFr�ҵ"O�U��9&L=�A�}=\���"OZ����:2�ж�R�l�R8If"O��!�L/[�lە�̢.�|��"Op-`��èZUPT��N^�5H4 P"O���a�͂`�h��' ��"O��;G�1K -Iff���%�"O���b�3Y󤁺�@R�^M�"O 	r���j@ntyB��;cԌu0"O�̻�`�)8�$|r��(�f�A�"O0��a'H+,�n�+�����"O�B~.���Z7y�fuKu"O(���.�"j��%�������"O�5Y��� :��]�����*A"OfW�B
0]�\�jV+w�@e�&"O�@���
�I9��Qg*?w ��"O��I$�69s����hD�v��"O<�@7(]-C?��p��E��"O��3�,Þ\���a@��Pv���"O�d���Q�\ܞ��s.J�}����s"O�؀aA�0C�YB��PJ�ճ�"O�)�k�����N<�y��"O��ȶ�L';f�sW�ͭo6���*O���UOȑ	�����]��&tz�'��4�w��>C���ʨ%dej�'d� JrLT�
�tI�l�0��%�
�'(Zm�r힬5~<}Jq�G ���
�'U>�A�䘭=4lp�ˍ�u��\�	�']d�(�.ʗM���#P/po��	�'$&%3��� II�L�GM�m�=��'-j��g�Ѳ_g��1'D�
}��|��'8�[�+�=}L�(�̔&n/��'gz8��i>�J-���>\I 0 �'H�3cj��4�h�gR
��A�'i*�j�]�z�JA��ܓQhv}�'A�Z0 �/q(#7�K�\1;�'�������!L�0A[��H��Z�')�!�����}i��� h��5y�
�'ӾU�Q
_��� y%�H&���
�'�P�ˍ�%��9S��_MF	i
�'�NUS�M��R)!�[�N��i	�'_�`�@)��)�X��K�!"�'@qJc��=���7Ҵ}K>�y�'���R�!@4�)�-t�z		�'��	�% w�y3��o�(y�'��%�6�R�i��8#�)�.l����'�93q'��=6�6*H?Lڙq�'3jz#��B�θ���M<�v���'K���[�|s�`�`��`�$���'�\=�o��b���#D�*�x��'wfU��1||AE P�k�@�'�@M��Z/'к���F1Or)��'bМ���į7u*�/���q{�'��-�b�~+L�"�_\B���'~U)����d߄�х�@f�݊�'ep�i�� -S��i H_�"��݃�'ݼ9eG�,	�؈��رkI�@�
�'�TL���4и��Ɉ�ڤ	�' D*4,�Y���oIѸ�3��� ȨJ�'M���]�B܉+lI�"O��ö ���b��f�h�"O�gA�
p3��7(05yP"O$�
��0Z݈�vM�fz8x�"O6̃"�T!_ -�� Q��A�"O�`���)�lT��?�(E"O�(��F�t^�l�AL�N"X`"v"Ot�)"o�Sj5�&���s�=�%"O���HEn� �>:(�"O�M���YO:��%@�"*��7"O
4��dX�z��G,j��q7"OȤ8Q@59:��8�͑�f*<	Q�"Ov�� ���l�B�JuKw"O���$�h�v�7"�>l��Y��"O�7�$)�� �X�c�L��@"ODuH�	�g��0X��ПV�`Tx7"O
8㢧ʥ8|6X���[��"OV-Ѧ�_���HӮH<h��9"7"O��*Ů>3���F�D�|�}�Q"O�| �
�d�j͊$g�jY��9e"OZ�IS F�i�֤*F�X7Zi.�S�"Ob]Z6 �&i����Rg*T���S"O���"j�!v�>5J� ��WI�X��"O�
6�Ŵ��%���2&AH��"O�lH3���R���G
�{"Ĕk�"OD4�ab��9�yR�	[c�eC�"O�zN+I,�$��M@��=�T"O�Y����~� Pvd�R�"O4s剂-hhT�V횓&�����"O6i�N�hdJ�ѱk[�Vj�hٓ"O$��GT�l����/D^�T�7"O�-�~Z|�&�I	cQ�4c%"On��$���v�^g�a��"O �{��W�t��]�sË
�j���"O+m]�&�� # S��db@nGy�<�u��I�]�V`	�I� �ӣJw�<�����aF"�@IK
�n\���o�<!�a�:My�
��eY20+rm�m�<�D���Z#s� u^L��f�f�<���B)h<�;��
%m[x0� �_F�<QB�=�T\�2�
7["xx�An�\�<9��M
;k�tbԭ��u�����`�<'m'P��b�ۖ+e��tJ	\�<)���N��9��"= �<�'a�U�<�I�4�.�K��ּnv� f�	O�<!�i�
Dtx$AD퇏Y�̖�JB�	;b�!� !F� # �S1Ɍ3jV^B�	�n�
�Q����N�����#J*O��C䉦I�1
��W�0�`� ��C�I8?~� �Cc�|��Ȓ�C�	&��9�&S�Ro@�+�C�x�hC�I�B�|R�c�a*Y;'ŖI��B�I�N�H�KL8�^9[�/M�p�C��tU����`ֻq�\���2A��B䉟zTX0j1��1D�N��Sቋ}��B�ɞAj��5gˎ[14(UI)q�B�I7!��)F�\(q�堉,aC��C �=;���!��H/�;P�B�ɛSf�=:�"\� XJ��H�f�B��U��YR3�D�$6�{���B�)i�L�ڶNF�[V���w#߉T[�C�I�Ղ��˓#[��[6G��|�XC�>�~�93e�!O�}J#�)n6C�I�C���cu�A�[-��)䄫V�2C�)�  (9'�c^)�쑤Q�Z�"O� pAB߂A#�qP+Ʀ��U�"O���#��1*5,��ނj��AB"OBq��?~���s�눦8�0y��"OF�q���9�2P W Be�<Ъ�"O�L�!/V\��h�~�X���"Ox�y���Q�R��f���e�`���"O��Ec��.���0��\�~�	�"O��"Q��]Z�x���٘��3"O���3��r����[��"\��"O4��e ��a(�@M�8r��l�"OJ��R�W��c��[��Yz3"O",xF�R�l8�7A��\�2�It"OBihb�:i�⠺��C�n�"OfIbG�J93�恊ݞ��xW"O���AAº-+]!�fY��a�p"O:A(d�ܔ}?�B�eI/__Rz@"O�u �{@�q�5ņ�j[��"Op�3��1���d3�d`w"OfMc�jC��)��W���"Os�_�"3��a"�%�(�&"O��D-"K$E�Hѝ��т�"O2����C,NZ�p�sd�(��""O�@ɠ�#&t��f�G�O>���"OTa��� 8;h�:��L&a
ѡW"OD=�ĎܟO��Pf��\�ل"O� {�
CZf�q��s�Id"O�Dp׈
�4����h�8�"O��9��/u�¤@c,�2�̔:$"OB|�էK)��H��^�T����"O&�Ĉ�u@z�j̉\o�$�""O,�����Z
j���25BHR5"OT�{b�Q���,���a�"]1�"OppQ�	<n���L 
~���b"O��#r�@5B*bTq��[���Z3"O�����g���	g��*Q¢@��"O��Qd� V����%��!�̰��"Op1����0�^%P��!2�&E�V"O:P��ϟ,E �����\h��"O���-o���!m�A2��-L�<	Ջ�135��{W� � ���Q�m L�<	$煩+�`(��l�ѹ$E�<����!���t&J�q�N����D�<���Z�W�0��,���4ԈS��u�<a�lH���l�7�C/J{��`�͇Z�<��sYŢ�/&f���C SO�<�P蘺�]x��L(/�5�vn�L�<��b��q+�]i$�]�5����f�C�<��h�Q��Y��4|x��'�F|�<I��D2Xp-�/ �x�3�Np�<��r ����
��/��+�Fl�<��i�U�\���T�u]���B�C�<��mFJvPaD�{��b��~�<�%áy�̤�
�=;A�0 2+�D�<�qL	+ r&i���X�>���rcD�K�<)�拤Ψ�x� .&H��bJl�<���ĩcb�����ژe� y22�^i�<��d�h -���)���Eb�<�F`T�$Ţ0(�e��E,UٔKSF�<1�O��Qc�$dڄ_��T)��@�<	�C���Y��3Z�E���P�<��!�|yb��q�ð	�>�󖂐g�<����,��0�MJ�w� h���Hd�<Ѵ�ݨ:B��'�&<U��Ì�T�<� ��§�0����7)6=̎���"O⌒"�C2�
��3G�^-�3"O\��n��>�jmR&L�a�@yj�"O���BK	.y�8蕄��u6z� 5"O�1�k0p葖��� P�!�"O��� �8(кd�H�f
\�Cv"OBj'�^�AR6X9a�,v�`A��"O�!s�#K5�"�a��p�d\��"Oh`j�@��
w�Yr��O.?e�a�s"O�q{���tV�+E�F>(�.���"O��a��5-���)2�����|�"O�\˶n��F��a���W!*�>XQ�"O"U�Cd�;Ԅ-�6/�W�@D�#"Ox�X��_�P�"eZ/՚iJ	B�"O��6 Z�V3�� b.K02���7"O�ɩf-^�L�k֌U�`��r"Oz4�v���":fl���ùDժ��"O�1y�eԩ#�
|1�@�&:�ּ��"O޸8�C�u,�"�eíU����F"O$ �0 �Y�̥��X�@OV�ئ"O(Ȳ�����#3�2c�]9�"Or�bG#A ��śrC	~v��"O�x�GU�"-UI%�7:^����"O��S&�[2V�z�� ��_o�X��"O2�e]�P�R�җ��f�A�"O�����?W�Xʄ�T�(�4��"OPܢ#�[�:�6�(g�O��.)�"O��	 ,	<O���4�CP��,�P"OL�{�"��y���D#;8��"O���'��I0�{Pꟸ;��x�f"OF���fгg��<@�o���� �"O<Q����7k5��ۓo��,����""Oȹ��JG!x�(Y�ŕN�"�"O��p�L� @�c�Ӣi�-p1"O�1�C��s4m����&�j�"O�X��c:N���V�_%�ي�"Odt`�I��=�H�I�ҟw+d=�U"�S��y,X�� ��ݸ.��!���y"� M�Hk��2 hF� Vk>�y27��RR'ڟu (q�5�y�A�L��$��B(z0\�p��y� ȶ�9�@�$׮���W��O�"~za��h��q�T�U�V5��^�<���Q�$!�EO�.nv|a�\�<�&mzV��U�'���{B�[�<QV!P	;{�u���H�It���І�|�<�Ƈ[���%"@�� �b$��Aw�<Q�Ή���s�J	`)�A�v�<�&Gd����,�Dc��h��A�HGxJ?�i�H9#�"ș�
,x�naC�*%D��{�g]�CU�J�0nd9Ȃ�$T���W�D�Oy���p�߻E��1S�"O"0�D�x��h�vl� \zr,B�!BbH<�6E��y�tj�"�-Z�as���E����>�Yu���x�ME&
$)�@�B�<Q�\<bl��w��.N� 3��f�<����<��i��(�^�JHd�<��em�e�'�ہF�N4C�ʃu�<���	����#s~����p(<y�4l����Nբȁ��2j�
�'~��Pj��;��@�7'G.L���'��`�}"��(!C�,�
�'!����4#4Xc��q,��	�'���ZP�%_�*ta�Am�t�	��� I&-�61�&d�ѯj�>���"O0��#�3x�>9[�bE�b&�!a�"Oz�B3�����b'�K�h#"O*@3ƀ��n���5�����'ܤ#<�T-�I�L$��.��(#�T�Ǉ�g�<i%n�]�TqՂR9sV��iŃb�%�(O�0k���!C� <!K����"O��(5g��"�b�k 'hɬ��"O���.J��p����|�r"O�|�㭉q���㏞?6.|�G"O:	cf�ݪ5�d��t`�+���"O����Ǩk�rH����8 ^���"O����cC�S>�5#��b�"O���p+�Y��b1��-/�nQ�t"Ox�c�;bH�Ea�g۠t���jS7O@��d�s�p��O��Uk��h��� u!�d��J��S���&o ��BE�at!�۳m_t�ţU##j�d�d�38!�DSwDzUB��\�0a�,�F��,1!�dV�$�����KX��a���(�ў��ɐ�����<g�0c��G��,B�	�K�����[�\��Rm+|e�C�	?}�D�P
F��mʣ��s��B�I���i"�Q1Vyf�i��^�z��B�I;?�69�o� �b�ڢ��x&���E{�C�<��!3�9�v��&*����e�U�<Q���5@j*��*�!ts��C��R�'�ў��h�p��.K�TH�C7I��I���~��./}�$ �o5r�N�l�v�����&'Q�P٤gO�9����)^���xr�L�@�ݲp����JsF?an1O���dI�����!���E��hm��pD�d���4H��Ȃ62�R�����B�I��vX(��ʽ2�p�r
��x�Dʓ�hOQ>��=*"�����C��<�F� D���� P��1��@�,ƨ20�=�$3�S�'sb:���̛
��;ņZ�2U�y��Iy?�m.GW҅`�@�$;X�� w@q�<a���l��Aq쉣]F�� 6I�a��hO�O<�]s�`�.=f�:U"M']dyq�'���C$N@<�RTl��3�=��'��٩�V!�$p���4#���
�'"�AZ�Ɉ�@�kroO�.|���ٴ:�!�(���C�`Hq�8���� ,azb���+<�se���eǘ0h��;!�T�W�&i�aH|2f�Y�7!�B�L�@�$g�2FgP�`aʙx!��ZI?��tn>ak%�EK�3�kz����~�نP�'m��a��I!O��dC�-D��Ҵ��#��P�f��&J�"+&D��X���:@���j��Q�,�~t ��$�O �	 "$<0�t�I�҉��БR��C�$%�l��BX/)���ed�1g
�?y��������
uA&G�.�Cg#��Z!�D�27�P-D@
�.����Hי5!��V�0a��B/2u�b�Z2�̤gH!�$�
�3'US��ŠR�!0<!�dء(x�<K��{b��	�AA?/O!�!Ŝ��"eϣU�@	ǩBr�y��=g^8�pHG"0~�$�3@CU�@�ȓ�`sU$1�ZbٌJB���:mƆN��t5xp���nFz�����8 �,Q�7��ԓ%�M�4���ȓWy4d��cרMCp��`R�M��}�=i	�S�? .����8x��IX��=b���SA"O�#�k��.'z(��EƗ`�b	�"ON��7�.�=R��m��h�"O&m85jKHۦ��G	^��$8�"O�:w��{�N�@,�:U���搟F{���ǭ�V]�#I�3|�\ԣcNV�!��+��$8WdG1qbݢ��?V;�O"��׻ro@(��c��-�^bA� F�!�ʗhZ�y cl��G���P�v!��]2�t�X4N"V�9��,�5��x��I�eh0�
��YE��ؠ"��&j�C�	�	+R��#iT�P.���J�9@�C�I,_���WʂP�����	�:|ĬC��2&,��f-S����f��C�I�c���7��F���
�K�;@�B䉝z+<с杍��x@d�9 �bB�	/6��i#�hϝ sHQ�AA�0`��C�	=���pE��,����u,�B�I�Y�l8�U�	�- 
͘Љ���B�I 	D�r�+7$��0Q���&�"B�	¦��JC�t��I7n���p���~)h��ֺ<Ӳ`�P#^��Մȓf���1��L�I��!�<����,� t"#!ϟrh60C��x����41�����	BrAp�c	�{�$=��~>N`�3��d�,�%��	X�^ԇȓ;R,Z��2V�`Ļ�
<c�&Յ�FL�2��#J X�*����n��i�ȓ��2E�/Z�@<�tރh��Z�'�N-�֏��upE)d��2N���H�'
L���ݒ^t���s���6϶d��'�}���;A�����Z� Z��'�ܔ{�I_	|�lbH��x�^3�'�
(�ƈ��Z���G�G B�F�S
�'��LЇ��'�5ن�Ln̢ԉ	�'�j�r�>m���3v�h&�@�'4\�A�ji�dB��T,g���'�,|�@T��A���l���fm�<)k�jl��{TL:��hf!�j�<I�N�	��EA���fo��s0N�m�<�g�J>]���D�	1Dd�tJ�i�<��j�+O���3ʝ�֐`�6�SA�<I !ˑav�@Q���t��ī�q�<l�#�`���9V��0�GU�<i�ע10:!y��Ļ]��y�-)D��qS��fb�Ȁ@q渡��	3D�L`��Y 2C���K'`Z��U+=D��;uJ��w�a#%�4���ɁK>D�Ti�K�;zt:�H�$ZN1�V�9D�X�SO��l���s��c�>�A�8D���ƣ�+]v�jW�[I*���7D�`� �L����Nz ��A�6D���A�Q*a8\��#D�RJ�I2�2D��8'�N$Q.�9h�m+I':�i��$D�P�eX]Y<��ek}�m�©!D� ��A��M��6b�ȂԆ!D�����!}�&u)gǅ����ҁM5D��H32g��K�L	-iu�H�Ea8D��HC�8uW@�"��[
ؘ��e5D���� ��Vќ�F�Y7Dv��ґI7D���F�I�^��hQW�ӓTFh�SЈ(D� �&FـV���q�ҸF��	k@!D�d�A/O�"�A�פ��%E��9R�=D�y� 
78�)B1��4C��LqC.D�� :�0��HF\AA��+ .���"O���jɔ#���zGN?�Ω��"O�5�gl��M��kϘ���P"O���w*D�������"Oii��S,V���*�́�}��@4"O,���O��N���Q�*�H��"O�E�gg�s\|ؓ��^�-�d�6"O��� ���b�[V�x�&�H�"O޴C�C�@��pA�Х\G2�(R"O�J��H>1���)�\;�i�V"O���$!
��J0'I���pK�"Ona�ƅ�{� ��� `g&�"1"Oʅ�������cPœ4W��q��"O� �7#�8��Ĝ&*��!h"O����ۆ��@+g�@z�>�e"O<�B���!f��� 3�F�3UޭБ"O�䠃�A�24��1��^Jڄ�E"OP��֏z���9 @�2~*�0X�"O�{�AM�+�B`���Ŗ]�D�0C"O�U[t#ۡ.���k
� #"OL�
�b[>E�zTFFNP9v"O���V�T�J<�Ͱ��F�3�ʁ"Ox���O��	c�+rBt<�#"O�5x�.��:�൲$��48L�h�"Ox���F/B;��0D�[���"O�`H$�J%yD~c C	2TwE2�"O����^�w�](uLK�1af	�"O���D�"5q��*��R&?Lb]h�"O�L��*bvM���E�`96��g"O�p酫g�dU�C��M/��"O�Is%,��Rb%Q`8i �H�b"O� �s�^ uTr�����z�<:�"O�AswZ�y��	��P����"O��+��JApP�c�K.��"O��H�`ͻY��Y��є�$���"OH��i۟8y0�˨c�^Mv"O�q�����H}��-ȸM��@�"Oڸ�T�P7K$�hP��q���$"O��ؖ�X3s3Q��ѐp�n�"O�d�rJ��'N͞d�ܡ9F"O��JP�� U���*fG^<D�,�5"O����i�Y�Fq�R�ޚYs��"O�����O,'B�����(I�LtZ�"O��d�ň����deB��4D�"O�\(�N�Z�yRߴ[E�Ek�"O���Rmt�YIGAK�*8��"OZ�a�+�Pv�k� B�%6t�3�"O�=s3g�:\ ��H�)R5|m�f"O�)����llDU6(�:^$�T��"OV������4�Wh�3ՊS"O�� �C�0��RgG��,�8��"O�I�un�BK"�E�d~(���"O���a��>�^��#$��#jv�"O*=��� ќ���	_ D^�h��"Od-�e☟l�M��J͢kE���"O�uHC�^7@����+~*䰊w"O��s��ΕA����e�@,��"O8���H4u��w��i	�<��"OH5�4➮���I���y��܃�"O<�)����tb8A� N�2H@:�"O�hi�./t�8`�F˜�v�	�3"O�L맡׳(�`���aNl��"O���A�$]�����ǁ�]$�ʗ"O���v���U��Ý�X���"O� �̱�ɖY{���B"��b�(�bF"O��˗Y�Di����7P�Zِ�"O�H�cў[�<,���\&�>���"O�Q���Y5�)h��W�`�l�"O�HH)��Lx2��T�V��"O�I���&��\�2e��<H��"O&U�ƃ·?�
L0���R\"O�̚�d�-���V.��~��7"O���D*_3F�I���6�:l)�"O�ţA�[�&�90���4��(�"OF �Q��z	���a��R[����"O��11コ3�d��щW.WX���"O�Q 
�p�z���NI�VB �"OX��l��MU�	#��}Mn�pW"O�e�soْ}�|C,ő+X`��p"O�ykň@d&b�b@6���"OP��ʢ<�i����/�)��"O�7���(/�\yŉZ�C�NX�"O<-�fQr�(V���"���"O���c��%6�[PGJ0^�~hR"O�exA�0+$z��T$<E�2�"O0���)3@�sE$���T�s"O�0��n8&�pcT�;��@�"Ox�AE�1zB�u�F! �k��7"O��bVOۤ9�>��4��������"O�$jvd�&|Y ��zQsV"O" ���@�g�jТ�bv��r3"O. ���݌gMn���O�Sb�|�"O��
FN�*{��9�A�$_tͲs"O5NA�F�@��e���M��s�"O~�Y��V �%Ñg�^E�s�"O���j> �b�����p�ިRC"O��9��Č��V�ɂ
�<h�"O��`IʡI1�0�$ܻ?m��`�"O~	���*8���ף�67Dձv"O��j��؃(=��L
�O.��'"O(��P�u��iAk�(-�v՛�"Ox����8)��׉��]Fx�k�"OtȷB�:��K�F-r��`��"OQ�F(�,JX�6��1���p"O������H��9H��
	����"O<���Bl�1�TDO�=�h��"OF�Qh�f�rdI&#D�e?^�2�"O��dū#8J0!F+Ț==�Q�B"O�uY�	�TbL� mEU; ��0"O	�f���*�`���I��K��I��"OJ�R'kL/A� P!�C����e"O.9a�$�e+>�����:k��q "O�0Al�E���	�u�p�"Ov��g��M ��cp�͞H��"O��င�n�Y��&���� "O�؛c�C+�@��ֆ��a��IiS"O`"�G�H���n��r����A"O~j� :�"\{U�G�3�(� W"OJ|D���m<(��T25�9k�"Oa��hʪt4y��+�ܘ�a"Of�Y� =L~H|��k����{�"O4�@���'�8%��A���s�"O�%��Щ
�a�v�Q  {��1"O~JAjI�63�ـ�i
vbh��"O�A�8E{�H[w*Z�'M��"O��*���2
���؃� :8y�c"Ovu���ܐݦ!K�CZ8�%[""O0�x���$��y7!J�e�4�"O� 0m�u�ԇx�`��H&dT��"O�uj�D�RrN�Bq���r��L��"O>�+կ��*��p�S�¤DD�"O�0�a	6��x`4�A�i���	�"O�u��-��/�8�bG�=���S�"O�b�%do����ڎ/��0"O̼[Ď��Y���9��J7FH��"O��A��;I�DÁ.; ��"O\9�PME=Hoĵ�VBO�+�q��"O���ץ;ni�|�V�46���"O�i�e쁾l�����.'�捊s"OBL��";m��jX��
�:@H!�� ���A�� �LzW���!��FI�cU�H#��R'�
�I�!��Gt�L�)wt���<�!򄞔Wxv�S��1g��-��|l!�g���eL�"IS�I�K��=`!�3~*�p�f瀙	F�H�w�&HQ!�LE� Y�q��u�#�E�8!�d�H�,�eƀ �0!F<!���X`����2��[��($!��1	���cú>�����EY8�!�*~O��X��ېg�*�8֏S�R�!���s����q�=HSp4��S�!�ĞEe�y)��K
�N�Ѐj�/�!�J�Rtd�1�0=��HW�ً?-!�]�!-��Шł(��A��R)!�ėu_�̳���/h�j�^2S!���d,���f�� �����G<!�$��(F`�#�O	LF��f��=i�!��s�\��aBO
$,�ВDLޫc�!�$P��BL��dC�6���� X!����\��Q������W�B�+!��	=,Vh���ʰ���WKDL!�D�sz1����.�Ѝ�/Wf.!򄒨4m�X��F:҈��M:�!�$K�f�����Ǖ7��$�dˏ�cu!��*Y]����T�Q����M!�䔱o2H!�n6n�6��F]�Xe!��""����Dc�)�\=���ִW!�D�%�:%Pp�^�x�z�w��2|:!�?%����@B�,�F�S�ЀJ!��3� b�LT=*�^�2��X.!�D\ ��e`�,��O�� ��!�+L!��Go�U�q"Z�?��t@��ݎH�!���"O��Q� ˤ8Բ��'�{�!�dܸ-�X�bB���q>����O�D�!�䆁vz�QG
��oR�*�C^�9�!���(�(�I��Y�N���F�&5�!�$�"��`���{и�[w���!�$ŬL4
�r�I�?��!*��H>W!�d��B�0q�׻��Rl��OC!��[ �����;���P�C�N�!�dE0��D�U7>������q!�^�=�y���P�I�p�Q��
q�!��&��!B�0�Q���,N�!���a�L�Q�'܄03��Q&Х(�!���/GL��!��i��W9F7!�D�R��HІ֮Ux��h��I5h'!��j���Q�.s!+��X	F!��:$"����Ɩ3c�X�D&]�ef!��Մ�l�r�	�O�u�6�˪lJ!�$�,Ĭ��blR$8�p�� �{H!��V�'�J�vn�,8�6�����$2!�� �<b��"V�XA��=�
��"Oz�uF�9��@A�プs�ؓ2"O6Щ��S�EP�#P�L1��iQ"OHd�fe�7�Rh;�F��F��Rc�>���L�b�x"U&�
ܲ�ƜI��X�J����:�~( ��+r������K�F7�5�� ��A@~Ʉȓ,���Q��q�H9&/ҝK� M�ȓ]4ru�Ȋ;��@�cN'@��ȓ	�h�y� j����wA��3���ȓX�����׸Qr�$1���h�8Շȓ�fT*�䖋RK`�A��7�&q��\�$�`��<�0y��J`�����h�Aʋ�d�� 1�@Lvq�ȓD��2*�.g�Y��K�9hF^|���DՉ��'>��T��̎�F�4\�ȓl���B#*��C��̢p$�X�ȓ%q�x���[�!fݒ��	�S�d<��xt�85$�: ��1���� �ȓ�8����k��P:6�A�#�洇�q>��Y�թb�8dj7�Vxb�\�ȓ{��9��O��Mz����^�{���x���PV�7}BȔ��!"Q ̘��'���UE˼|e�X��ҥ!�Ѕ�]��\��]��0���9Wt,���>��A.5P8��� 9=�=�ȓf�ba鶤��Y��4�G��2-�rD��]��\0�i�=�ij�䜀3�}��	�'� Ԉ!�{�\Xo�A5$��$�GZ��3ӂ7D���k˨j�fUX@��N`��HG� �ɷ� ����h���`d��ѲD�(KU�YY"O��J��N�J���2���@$�޽"�X����Ty~�("�g}hث#�U��B�[�X}�f�'�y��!��Z�@�# HT�F-��~y��0��/
�!2���E��kFEM�_�pR��ݵ#�����.LO:%В�F�t +X�+k��j� �T�&��`�Ğo�B�
�"O@�Y�AK�>�v���y����0� Q�gfE�  ��ᓀ����Af�9Y��)��䐳��C�	=Y�q��ۧ;ȉ�u O�N��kQ�Yf@�a�C�ܸZ�I�$>�3�	�3�d�x`eGN�����\B���d�2�lyy���t�����ϊ�R �	����u�R$W+M�	���u@ LO��j�&\ ��=Qp�\��H���+7����/	��Ԃ���d�`�z�J�\���`6$���`gE��y��7h����&��9&����F
ڤ�~2E5Z��-��V�<�Z6yW^LG�d��'7 |b%D��u�}�%FZ�y�ʛ�v��[���VI�%��Um��i�����o�V%�S�tj��'���6o�v)���alk��ɺ
�T�nA�@�7
��tÐ�<XI�P����,�Z���+��	����EDO'2|P0��ɶ(hp2F�N���#�5H�T">���ŌJH�<��TF�z8����n/X�� 9H�!ذ�Ϛ]�<�b�n�\�<�F�BU�9���^��iJ�͙ş�0�[2Ng��5JX%sЂe��&NAS�1�"�GY<LP���ǫKn0�ѕ@F0�y2&�\Ybh)dfŘ~�n�:��ϙslܭ�e��GeV�����($'�A���ӂL}�o@ds���J_�|�oĀv������ �8U�5�Lk\�͸��/��Py��ȯ�=(5LB=�o�s؂�jӓ5Z�IABCJ���hk�k	1\*$@Fz�R�.���ŎZ|�	�Ed٭2��J�H('�j6����JS�h�xC��:hzơ��mI'
���e,�-X;~7��¨H,Ya�k�]�l�2�-��7U�%�~�����E���E��$I�b�2O�m��9����
YZȵ��a�&o#TM����d�؜����	}P��"v�d��.�Lb���4��O^8�tK�&c�4=`��9�O�yJ� �1v�,�T��*L���fEZ�9=�e����K���!m_�٪�CF���Ə�5}�`���������3ғG�d��[�	]�|Cjʊ{�~}H�i�0ļ-����4��`Cv��	z��ҵ"O��Q�S�N���C�+a�.����i�f�BJ�R�`�:�L^$2R���)��k� �4�͎�3B8�HW"�C�ެ�"O��z"IF�&��yh�߂�����ج%�lpB̟���1p0.�9:���1��'����.[?��݊7�ոE-~ y
�<�(T,�}�h��c#�$8�>ѣ�lb���)Ʈ>4FE�3�S}�jS�S�=�qI]���h�'�7�8E �ޒ�ҽ&?-3��M�/�Dq��ۺ"/�5��#T������;^���b�Ǆ�?�~��P��bt喛>$ ��N<E����Lo��8��50`]�5����yR(	2%b�
4�):|�	�!��y�@V0PPx�0�� �y��F
0�y2f@�A�đ��sOpX1�A)�ybͪ,��Ǚ�h(����i 2�yB��qx )�CF�k��u�`� �y�,L��.���Ǔ�lѨ	dǊ�yAX�~�hX�u�X��p��yR%T�G�&|���?Dψ@;����y���.L&>��Aυ 97
��n[��y����j׬�.ϐ��_�yR���O�z!�"Ǜ� 8
4��kC �y"� �@��I��#н"���2v�A<�yB�%9"yX�
�m��2��ٴ�y���"}>��BR6�� S�-_2�y�Ϟ2 #��` �<.����˖�yB*C)2�"AYjο.��e3+ղ�y"cTI�&䲃���$�j��^��y���
<�w��+��$)��^�y�C��Va"�aV�P2����q���y��ք5H�i1@���.��ck��y��-)26�C�� �]˶�9�%��yB�e� ДdϢ-����i�#�yrBף}�S2Lޜxp�B�L<�yR��_�p�B�|�~%�b�I��y���;��̢��X�}K3�o���y�k�([&Zȑ���p�.�飌ʝ�yҢR?��GT?s�����yb�V�.�H⤨C;,1���ӭ�yr�W�E8�t�q%Ϫ='��)�猾�yBE��L��b�n�(�)�2`Է�y"���,' ��$�+[P4�A�X�yBhV�:o��)�L�%���6�y���4zM�x��!'/��Pǡ8�y��E�pᾨ�ǫ�;��RF��y�锓k�������xLX�����y�bƘ"����C!�"S>dK�ˍ��y��Q@|`���AI���l���yr�݂{0ڥ��ꔞE� ���ڴ�y�K8\F�yu��<�BIk��=�yBoY�En@X	��ч7j*�B1���y�͞�������$���Ճ�&�y�.�?V��Q�P(ټ4#Ef@��y҉ހS_bU�bb;��)��y��ߺ�`ܡ��v�Tm
��[��y�GO�N�P{����6hl�҈_-�yB�#��hR����p�z���y�*�>>�ْ�=z��BDBҫ�y�Q�T�HR-�j���ЎR��y�b)_ �(��֍4@�(8*��yc��|eld@��=7�E"�$Ň�y��ݟ%��hRB��&� h "͇�y�&�h�k$�n����˹�yb�F�,[��T�3a,80Ywd�y�,M9o��ܱa��R��������y��2z����s�%��M�$�ҝ�y"`�GU�=�D8�|�Ҭ�y
� ���gטS��8��#��&H�"O�=9хE!㖄�C�@�����"O�L�f��)jq]��Ƅ��I	Q"O<S��B-|5X��8SU�B��� 1�:��C�'�FpySEّ���`�bG(/T@ �ȓi9���o<kt�Q����1D<(�̓O��͓�؅+�ҧ����z��ӱw�xi!a �E��h$"O�,�ҋ�|zmWψ)L*Q��^������![�$�t��z���&��{GP8���;a8d�Yt�:�Or���(�4x�J$(�fL�1��5RRa��g����E�qk���Xx�eQ�V����W�;�&�Dz�Ć`+,U�"(��@j�&?yr!Х� !�2�Szr�k0�"D���w�S�f���c%���R6 �"��C�y4]S��8SnH�B��?E���}?�mؕ�Z*�F�:f���dY��N��%��Р|��#�.���z0�d�'0
�gm?t᪔�mGrF{�h��0^z<sA�(pB�, 4�ݴ�p>1��)s٨�C��3�е#'F h�鳦�Q�.�*�{���;�?��XP��$�o�����f�Y�'c��!P�Y�V����W6 ��Op}�ÚX[b�	�ԇ+����'��%��CFZ����3$��4��	Y֊�2O9t���8I0c3��O?�d�!6�B����&W��8X�� A�!�U�c�Zu�B��A��r�#R� NV!�	�?,��S�o��250�:�ԟў	�f�{(���} Pd��G:�O�	�:Yv�9YRFR�m$8`P7F\C7&B6L�Z������?9$���5m�ڥ)M�A�^��ց�b�':3-Ø2� ���F�`�]�(��&]&��(� �']��B�I6jhZX����
��ԓq�� ����E�~�љ I<D��S�O-t<h7C($���B!�� ��$��"On�+����x�������4�@��W�@�ǃ�h-�\"�\����գjfA-�j��hR� �O��2�/W���`$��ҥ%U�1�A�gi?4����.�q*��W)P�KD8q*���;h�UD����ZiȔ�&J:��9����y��S�ӦA�q"�z���[��$�yB�	<7�
�Sd"aGv=@��ڛ�y2�� �*\�AJ�$4yD�6�V!�y�E�5U �(cw�"��%���R0�yR�O�l�(չG�
��5�e��y�J��ZEg���4��L<�y�AL�O~�M������*�-�<�y"m��>*�E�T�)�f��蜢�y2���,��%!�*{�v��E�I��y�>����^�-�P�T����ybn�*ar�#��J�#� �Y$��y�#��[+�u�r�[#K�6��V��y��e��!��Ν@��t�B��1�yb���l�$��2�C��J��Q(���y�횓3�=���R�i0��CQb,�y�kߨ8V�eZ�#Bf���X��0�y2�6!�ظ1�Z��A�5���yB�S�2�;�  ��"%+ט�y���[�@��������(Θ!�y�R�M7��9�,��nD>|��	,�y攁�T�(#�H�T\�h��	��y"IBGw��"���:��*�%��y��L��dy����MR��Ճ�y�,�K�`��BkR�q�̒B�<�y�Q�z���q��s��z��^?�y��Y5ܕk�nָ0j�14�&�y2�6H��RW��&x��g��y"�
G�B$o�|H<��Q�Ğ�y��U�k���� �(�c�����y,�d<��1�$�,\�×�ĩ�y��"���u�W�v|�0$
R��y
� j)� ��.qE6�xu@�{�m�"OR4��9S�(����a�0�;�"O|5�0�]�S�	�N�+^����"O:�a��ol`���ْ*��mhB"O,�X3	�O��0�����7��XX�"O��5��1���"%�`��P"O�ى�h�2\ ����L����e"O I
�O��*���"L�0H�"O��A�fA [�e�)A��@a"O"=�D�A�R�օ�5�2vf�8!"O~`(����Wd�%�!�t���q"O�%b�N��Y��:���`�6(�"O�M��h/1��g�FkN���"Ot�z��V�&���ۖ&NuK�ة�"O>��6��`����h��*�.$zd"O(��B�ù)-^]�u� �l���Q*OTa�rاD���[C�ޗB�Ȫ
�'/F���"X+,r��GE��8n�L8�'��z�kߢL��R��;C9F���'}d0��ɇ*�"&E #�j
�'o� !��W���B�!�i�	�'�|��ٓqXT[B�'"$`	�'����͓(}Z�D�5V�'� X֨G!_�~�:&fW�ȅ�
�'�������1�T�bVKنBHƅ��'3�2� �s�ba"���	ަ� �' �
I�}�Z )�ȑ�'�4yS$2����GƬxIN\2	�'w^��r�D�?��qj�N�<t�$)�'����s/������ H�o��#�'ͺ�&nM�!L� ���\6̨�5���@�<�a�Z~�y�v"���`�k�<҆�q�V�CtFC)�F���l�|�W����w$���>u(B@ �z�2��q���3W\Q���?D�h�f��H��ecJ>���'���lf��+�����y���d�!�4����_��ҧ(�?<!�$[�f�� ��'��N���EƗy�-pf�+,��o��p=ِ�� ~�輪�̟�R:�����D���Q��(e`��`�B������Jn�*G}�U{l#D��Zb�H��lQ3ʖ�{r��� ��~|��5�A)0+64��	/�'OZ���H0`����*�ƌ���@PX�d��O^�@�W�'����EA��dա�zm�0bx�g�}��8��`� F`�d��V.�b!����|��(���� 8�T�M,>�tiC(�� �I�!ҋFx���c��W���b�*P�|�.�J&P���S5n4�U���#��3zp��eD�)t�T)i5��x�����Oi~,�M�"�!�䕷8�0���j�!t  ��*�)��䟤U]��s�'U��y9j�L��Uj��I�	Tظ��*�!d�)YgCUF`!�D^�v ��c�?$jn�s"��%��݉�Fi5z�C��c)@�R�?��Ǆ-�	"f.ذ
`b�)tɰ�󀌁�=4���d�� +q��u�)c��҇w����9
��g�Q� �6I ��ڨmaz�I_�s1��H�㝒G�������O2����d�;"h�39_������,�h`p�I ��bGE�+�fE05"O\Փ�!��;Y ��7�Ԣo;:���'4���%ѪLP�FC�XRB��'��9[�6,��܂�
m�p��b ��b#(D�����12>����Y�3ix0�׀�9�lr��R�JڎaCf� yf���L�V��{�2%�f%�/-аtJ�АE*a}�� "�@X9�o�<&,��fF�r����S[�|WD��"��ki��I���
>a���$Ԛ����mƤ�� "�� w�����w���YB�D�ƃu�<��Q9y����`�Q3u�m�j���A��y���0S�I�W�-U�k�K���(S���:zE���C�@ȫ¯�5n1�Pyg�?�s��;�!��~�0�q�T�uW�9�8D��T%�y�>y��
XP %��O^���'i�'HVĔxq���T)Z�'L�0�7�$�F�)������%ų<a}2�dp�s(!� >����6�h �q��1^~�(�ARE^I���G���}��'���%��7�xqA�������]�Ҙ��aC=R��� �BP�Б�g�خd�44�`4:V�!�ʌ_a*���p��=��B��	@޵���Q@X�l4;V4ѣ!�92N�Pʈ��Q[��%��[E
�ʈ=��愞��� ��}�<�!�Z�T"���J)o�}����梅ie���H�X�����6d�O2�j��[�%ːI�`��x��0n*�O�U8ge�:۞А��ϰdv��҄�
ĵQ%����/9�`a
�\�<�RmRCP�� 5ʸa�iE}r��-W�.�D�\��U�ɂ��K�ʉ�`�BmV��*������`��Y@S΀5 ���'D����s�O�>�q��,^ "�bU$W5^���9�M2D���v��w5�զ)*��`��"D�$�f¬z\y�"l�f����D,D�P�D�Y1�Z] F��B� ]���!D���#�L�
�8D�ހ�:M`��=D��ag�,J��#�P ~1� �>D��yu��!N�y�0$K�}/��)S?D��b�lPy6DH���M&�ܝa�=D��C�OҁpYJ%�	�\�-W�;D�D�r�Af�"����;���@$7D�X���Sk ޕH�,�C����$�4D��3���,�qP`�0PE�b�5D�@�W���,���Bu���1�-Y' ,D��)6�%TԸ�JQ�v���SQ�-D��B�03w�ģ=��P�jC�gY�B�	�8��}#q͍�;���;��b5�B�	�E��{�R�Q� �0��/t��B�I9S�v$���/AF�ĪB�!'�B��(E��9QA�^�3���j��B�I�#NQ���1g�$�"G.���B�	�
@H	T�UB����ͧ�~B�ɅO�V�b�A�/,��qzB葮�8B�I&A\fo��U�y�A�M��C����M E��)H�d-�Ui7��C�I	/���2�@�$E�DX�B�ɝ6 ��iF��=�^]BХ3��B�I2!2�`!a��}��fE�{�NB�(K�LR�O�B��h� ��=D B�I?L��A���e,�x�kȘx��C�	�+��ˑ#�6rP!a�ZO��C�	�}'�=�����!4���K"\B�I UqxUBᴍ���xa�C�$B�	8}>�툦�V�Y��!���&�jB�ə}��Dd�5����Ar\B�	�DGR�4mԑ)$�B�6%� B�ɆQ}��B�4z6���ѥm�B䉫
�걣��.y�����/d[�C䉡M��hPRn��ݠ5 DW�$�dB�	%W��MRì߀ �����z;&B�N�0ɣ�E)}������/j`B�-&���ǅߥ�Ti��Ǉ!B�I�_�Pa�  E�c���Sa��;2s0C�ɭ&f �@F�ŵfI�$��v�2C�6(zĜ�Ƥ��Y�n�!R(FAzB��?=�@��nP5]4J���:?~B䉙D�&�0�m�M�K�,��~@XB�	"l�i��LZ&��Y��M�H}B�I�|��bǟ@�MlǏ��C�kϜ�tNLy�j��1�F�2{�B�	7.�bH\�2�x�B��?JDB��6��`�m�hu�dLU�z^B�I� ��)3$�=FNQ�c��/
B�I�@zr4Y*Ǖ	������ֳ~�B�)� @u؂p$Z!��3��y�"O T�$H�Q�b�2��|gT�*O2-ק=r�e�H09�� �'6n�S��A��!�d�Y�!�n���'����� �6��i���5�r��	�'Bl�u�N�s�Ԍ*�۲+�B�'�4��E�U�u\p�"�G^�#( ���'3!�f��J娑D�j���J�'�eXg�F�77���B�7\c�D��'��@�#B/+D�U��
O=P�x,	�'��`�G�.�aJ$e�>J��}@�'��3�#��fp�0
��@��x2�'��p	rI�� �MXX �[�'@i(�K��pv�yx0�@� =|��
�'��K��Q�I-t9XB	� ����
�'�z��ꊪB�T��H�x��`�'M��������ҁg�h �Q�'���vDG�\�b�K1nĽ(�^l��'P��k��i{�	���>���
�'q}�� �j�{���!�%j�'���d��<R�<-2& M"�Ld��'���{&�ί K1 � ��	s	�'\*�8�I��b@0�
@F?s��)�'1�H � ���!P�
m\�h�'
���a@�q�*$i 
�=T^B�J�'��Q��ĉ
B��E��Byj� �'�<5�s)�5*�pY���Df �
�'`�k\�Ao�� �%�<�4��'���p�D݂P���r��{���S	�'f�Q�g ��o��%R��Ѱt����'�v���K�-N��tA��)>����'�$��"��<���ٶ�ʎb֘���'�@̩�̯2Ln}9F)Ψc��8�'AB(j�/�G="�����"$�p��'���W��3[Ȓ���O��5b�'S������ iӈ4��X�]L�k�'�`4I���bH���'	.kꠐ

�'������_%��с�g��h��'�퉖�����yr�ؚ^�hJ�'�@g��N|.�I�#U����'���p�d!Z���Z`��W��#�'�n<�# ��l�Qb@�Yl��'��%��uv��TLV���\h�'�MZ�C�ik�e����:q�8�c�';>Ds7ˍi�NP��:oP@�C�'��|)A���hA�	"b~^
�'�V�9��T�F����X�O�Tus�'�|`�c�g�~�r6�GSM�Z�'�pc � �nY�ehh��'�tq�C�;G�F})�)F�D�Ĳ�'@,�RU��
�&8�1'[�E�H�@�'��8�L�>08E��T����I�'H��'SDA�"I�N����'�X$:���$�Ĝh��9�Д�'�@���)dXREhgK��6h��'?Z��7N��6�.PA3Jx�Z��'ɞ���<�,L���QL�Tt�
�'(�!�l\ �H���e�B®��
�'�:����
�2\�Q��]�!-h��'�%@���l�D-�L�#%HT�
�'Rp�+�g�pSP[eC�+�18
�'1��c�h�,M������6ڌ H
�'�.P
��dOm�c+ڟ|�<�y
�'�jA�a�
�r��ZTf��}b�b��� ���3"�w�t�T'Z f�����"O$h��O�%��ǉ�)y6i��"OD-�!`$@	D� Y�HQd�#%"ODD�3���#�R|R��!g"O.1����]�]!c���p0^�	�"O(𐠣��><�,r��+1Vt"O�2$��T$~�;�eȳm5���"Ov����	��y	(:H`��"ODT �]�`��-�6��0!���"O��B����v��@��/=6��"OlQ��	A�d�s�ږ8�D��"O�'��hπ00����� �#}��W�O4*����^����ؓ��DC/	�R*�q���X#*���`sF&�S��'��d{VE Ө��6�_8Dq�h�O&X�Z���#�����N�⥢�JF�S�O�x��ː�9�|t�۟+�<�s�'�F�!�S ;��O�>-@J�m���í�@�2�����6uY�.����S>ɚP��*sR� [��A�5��,	�
��I���TKG>i��.#���i�NT�g�9C�$�d8f�1S�ԟ��4���0j U�8Y��Δ&%��}yPEx��)���\�'n��4���Xyb�ծz�'� �i>i��&&_�K@I0��$wX�CN=hc�A�L�<����O�?9p�,�|� ��E�Z�Jָ��s/�C��B5&�r�4o�aD��'�B��x��E�[�T�ƪ�/M���'�\6J�Z1�ٟ��9��'1�49b��@�)��*�_u�kGӣV/0���ۑa��M�EG8qa��on�0K�R�Jd*Q���т8����F�I34�"��T�RŦ=R ��zB�𩖙Q[ԅ`�,��gxL�E�sFh��'��9o��[��58w�O��xC׉��z���5I�>�9�'���n|�@0�6I�g~������`ȈC�x�S��gT��BDj��0��?��O|调���gQa�#
$2g��B�O8��(�_�S�O���'�0@!T,�{z�$
�47��X���S(<"���s+�*{<����݃���3�V�O���ҍ�041�I�	e��`qF��ܜ,�J���L%	���R�(d�ؙ͔N��'e�ܑ����Y�Q��0��JO�a`H������=���t�Q�"|BD)Z�,v��qWo����� /�j�<9�I�2���Gl��0fn]��M�j�<i`NݲWr�$��o[��
�2V�[�<���K������K��y"�bJV�<Q�D�Z��U�� =:��bg�R�<A��ĎV#���)�8jd`�s�
M�<9��,C�̜kC�4W7Ɯc� GL�<)p�Y�$�8�W�M<>�`P{�+�E�<IGA�-p�N��Z:Mo>��@�Nz�<Y����o�v���]7f�����~�<���4Ӳ����K�&c�ģ�$�a�<i�Fеi��C�(-6P!�D�DB�<9·F�\��nJ"X��֍@�<��e��t���V�T{�)�D�y�<�&��.!zQ����/:!h�����y�<���[(�e���*Wq���׏v�<q�jϤQ���������A�J�<ѐ(� �h�#��;P�FqPgNE�<�A���ޡXWnǴ}6$�yA+KE�<�2��6}{�AyM���T�Q NK�<��6�&�xC�N�䌽�C�MD�<��&0A�`0v!ߋ�^��`I�z�<�qm��5�� ��W�z�}	���w�<��HP�\�|�1�� A'���w�r�<!T���| z�c���/Vh�r�a�c�<�F�Nkuę�rC4Od�:�!�]�<Ag��;��k�-a`@��`Z�<���N�p�t��-� J���cb�S�<Q���5\V����!H�G�� %
�M�<y�N5Wa���O��hT`z�kF�<� �u�∂�6��`qo�K��m�F"O	I��Z(6Y�@��Hz�x��"O�+G�2`Af��	ϴ Q���d"OV�"6m[[�|�;�h �5�ց�%"O:m�fƗ43�r�D��sa9�!"O$Š�A�WҐ���>9FQ��"O\yq�cZ/3,�ba�M� �r�"O@|
�T(k�hI�e�Y�7�Fx3"O� @dX� �"
�d�)҂"O�x�&l�dF���G:���s"O�����w�9�'�[��PJ�"O&Y�c<�칐&R-�.1Sw"O�d�v`�;Fd갹�e��*#n*�!��C+[�8����կ����6�T�!�ۼG�~�0�HܛJ�L;�o�&�!��(`$��!�J����A��S�Io!�D3��͘F�]�(��q��G>p�!�d��O��D1c.B;+*�@��X�i�!��n��̸���2���o�+4�!�0o��s*�\��*3D��H�!��?Q�Щ0T̀�u>NH.�D���"OL�[C�ř2�`rH�#��H�4"O��顄�;r�Jq�'*#y�A�1"OH�x�@�1E%N�j�(�� ���P�"OX*�nI?=0p��8x|�c�*OP��W�Zqa̵4+�.�Xh��'ɂ�y2��D�:�kD�P��i�
�'���ㅩ�_�l��2�^�s;��s�'9��`�?I��!�Q�U.eȆ��'�����|6R$�#[4\��'�j���"�sG��2��a�p"�'�,�(�
�=�<lK��ȓp �p��'t�Ek�&��HD��'��w��|��'ز�am��:=XW*�k����'���m_�K��fhc�(e��r�<��-��o�����[�#�eȔaGq�<�EC=EPU�Q+��@�@Un�<���0uN��&�%Y�ڄ� �i�<匕�w�24�3��%$�T��U�g�<��	4ϖq!�� #�f$+U�d�<��.A+}>�t������w�`�<Q"k'!Ә�#AU�2
hU�(�X�<���c���R'*�J�!!čo�<��X�68(�]�Sh�Cv�Sl�<9�ыR��8������� �_o�<�rIJ�3��-����9�X�A2�i�<�DoB>6� �pg�|�	��DNp�<�Rn�Ŕ��&�R8͹&hQ� �!�d�@j�� ۮP;x���^�/�!�$�����Ta�L5�Y��ݛ!�DW�HQLArC
�,�P�!�.[�I6,0l
c�ˠ�!�D	/uǾ��w)�4I��q�g!�O���1�CO4� ��BXf!�D�2��A
�a�N5j��]?�!򤈐
;@)R%�T9��8���3|�!�D�}�L4S������D��rG!�D�:D���ѧ%I����Ă]7!�J-qƕ��!zcj�ŊC�[�!��)�j�z�H�6kX�;���!�$�R��w�
a	����U�PF!�dͶA7܁���O� �pD	X?'!��T1zjxt�p ��^� EZ�G�$�!��[ Y2ĂV	��s��U���F�!�� �ñ�߉CPvMk�&ʩ0s5 �"Oĭ��!�!f�ܐ���Ǐ~`T��"O�؆��O�М*f��
rh��g"O��2.�03�H��4>Z��3"O���!O�s�fl�iT N��3"O���f��;Z���i	F��R"O���,I�Ҩ��@524��*�"OX�PV��8T���O��Y�I�e"O`=1 ��'6V0��2����h�d"O�<:a ��[��5B�K@�h�\T�T"O U�"�ͤ*费Ї��
l1��"O���DDgt�#I߸	!P�S�"O��6�B2�HX�RN���4�"O����&X�Ơ�桔F/b"O�����3D�Fe�ЋF4u)p8J�"O�ģ�Ү��M ���2�T�"O��Ǎ 7>I�i���+���b"O&� '�={FCR���H��I�"O�h�2�^�sr�%��� ͎���"O����k����aŮW)�p��"O�I�ϾNU0�x5O�~����a"ON蠅�ۊ|�ʝ��-�t��#�"O��  ��Y�j����|0�u"O�e���͗w����M�<S�0��"O�z�U��U#e_r��a`"O�,0�ڼpd �n?]���"O�`�r��?R|a��LX@׺=	'"O���6m�z��s̆�4�6D��"O�m Bȇ�E��� �(T�:]tdQ�"O����6z�QJ����9V���"OLh�F�؍9Y^�዗���Dd"O܌Q�J (�q��ă���"O|L�d��I�����6Z�4|��')�u+���
�� ��@�l�Jp��'jBi9b�U�xb��΁e_ LP�'|2�S�d�14<������/b�P�'%�5�B<Rb$1���,��ę�'.�³�Ρ~VtRq�Lr/(��'~�\+�GW�i|��sC+�)l���a�'�T���o�le!�`��S�'=�j�Ȍ��"��dL��S�V���'
�ؤ$�bp���i����X�'�9)�l�7k�=3�(�+8h�� �'��)Y�B��(ӆ+ٮ'�Ԍ��'�hm;��]�X���T#4
��
�',H�rL��Dj-�F�N�B��	�'�عRS �X	��E��=��	�'�zti�eɷ�L�#tF�;:�a{�'n*uB��G���dҔfC�2�0�'�( a�N"h�ܤ��d><�jyi�'ج.��� Jׄ�����ԙ�p<9���[��8�@� _�)X�ӪN�+�!��g�rfϑB�4����Lj(IH�'p�	�VԬ5��y�Gj�O��0��'>�����a�b\��+4I�xE��'��Yp�TJ���'��8�(q0�'g@Q0�7���ڎt�4@�1D��%�ƨ������C�`g8p%/D��gg��!�)(SE�|��-D�H#@]2{0��@ݠ&P P%,D������8t5�����M�b� h���*D�(�r��")�����5C�] o#D�@o�&�1�6H��Tg�A��,D�L1���{Y�A��B�|J|���L&D�� 6y�`V���tZ�
3l�\I*�"O�Jg,1`rvE[CJ ?>�ҠS�"Ou�m�&~P�k��>3�8ih7"O&�C#�U�2q>��g� ^3��t"O�1�`�&��}9��B�R�Ҝ:"O��V���R�4�"��	�{�PY�""O�=���
�čI��?�N�"O�P����}��Jj��*��( �"OR�ӡ-�3u��!re�K{�� �v"O��Z�L�Yld��SLT+)����e"O2�koA�4t����,��%�"O�[��%Upԅ��W�����"O�2F�U,<0hE{�c�:%�Z�S�"O��wm��&��(P����#P"OR�b��ow��@5f�Dc!"O� '�.79����} ��RQ"O�Q#� )���?�Qpf"Oj�3u�p�
�)0�ߢU���@�"O�i6a��F�u�PG ���"O��q��)�t�s�2p��"Ov�b��b�J�"��/Uz�X�g"O��q��ُ�  �w)�$kґ�"O��"�N�+�X���� V�q�"Ox��`�͕Q��q:`��	KE�R�"O��	%�g(��"2f�H#"O
�%��'��x���E< &D��"O^�C�g�<��]��`��^f45�q"OL�� ��;�\y�n�=N@�2`"O�P1a^�P�U$��;/�P��"O��{ʈ 	��4��Kp�t�"O���ÇІg>��(�.�,G\N�Ҁ"O�|�Ņ$4j�� �LL�:t@�w"O�q��]T���+�=g�lQ:W"O%��DV�>�re�!�	�#K�<��"OԸ@�-�eD����@+.C��B�"O�]�3��0h� �"�&֧%���7"O��م��#����KݜZ�d�q�"O`i���Q0hMJ@Bea��`ys�"O�}At�QQѲ�*�ϋ�s�@U�"On��'��/���"'�M~���"Ot��c�P�pT�ЪV'ڒ)?�1�p���O���&*�M+�����^q �2�#f�J�qt�٣{���?����(s�PU��ߦ}�'n��h��y��Ӭ�jd/�86�HU坈Y^����k^�MɲU[ra��r��h���N"&����ڲ5X�e�g)��c H@�Ӌq�C���*n�O4�`�'T�7��x�Sp�t!�1k�0@�#9y��!�逌. ��)�gy��\1t�p���� f)�s#�2�~�6�D�eu� �zG*�����!~-��p$�Y*�!��H/�7��O���|��'��'`���-*zL$� c,c^r �E��`��uágH�?Y\3�"�Z�)x�?����n��^���`e)��.^�	��@(���-WF���#d�Ԅ����^�(A&��$�vޝ����v�DȂ�%> H]�ߩ�?� �i<���'l����������͒}).�4�"n�jH;{�"�'kҔ��D�5]6I�g��|�D�rAdȢ��'cx7�Ҧ9%���S�?	l� 0rbC�B�]-���W���W���	�d���*ٴ��<	۴%�6�W$	<hP�H��m����ıDT��) ȕrU-��mW�%螤Jb���'4`̓*Ǵ?�u���̰>�zM�C!�1A��Lk��ے��ՆQ��P��P�����.��'w��&�4K�A�pr��ߴ5݄�����MF�x��'%x���R��"�8��S��2p(��=E��������F�a�q�
��􋑀p���dH����	�Mk�'��I�.u}$�m�⦡��,|�N��`�	xB��6+O��$L�LI�0�C׃�xA�	��4̺��G]�Sy�Ԙ���!�|�I���47<!Bv�I�_r0h���<���I�#�&��3*LW��j�ʂ�v(@q`̃���BiY�OX骰�'�&7�#OqP�
�e"�� ��C���Ɵ��H�Ib�'���7�ǲ8h*�#"��0\i����d�b�p��M(t��+0�'08��@f�i��mZLy�T�D�6�O����=� �IP"`;\e�`�B����)�2�>���p}�9�ac��9#�lI�+�{2�`H$��;:�D��}뺥X���D��`ЗI22c�@��sWr-�,U7�ƴ	�Oԅko��)�9J�R�� ��� $���p*�.2�	)���dI����K|R����@��N�m(6�s�5aH’$hK]���?E�,O�T�gJ�C\��@���*M������O�%F~r�~�4�n�K}" H� ]���U�
h���h4A�2tk�'N馽��cy�Oo�����,M�8�SD�֪k-��H��\a��Y��+$��e���C3��)����y���'���(v޽�󤀱gh��h�C2D��hH���<��z�bVa�8�JǊ��mldu� �1Pj���ϻV%~5bU@��'�`�#ڲ3?
 h��'��6�Fyb@A+���;DнaT Ҭv`�m�3�X���CT�'-�'�ay���n�4Ȅ�	���ҡ+��'e�6-�ަM���'�Ms�7Sx�p�#D�7rL�`�r��!�O,A�q�  ��   �  s  �    �%  2.  s4  �:  �@  7G  yM  �S  �Y  B`  �f  �l  	s  Jy  �  х  �  W�  ��  ݞ   �  ��  �  ��  ��  �  ��  D�  ��  ��  ��   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ��N~��\	?Cv@ӎҿF��(8`����y�DG�|�mYDG1E�>-��'��y"	�*]�MYԤG,Czr��v���y�M��ۗU�~L�S�Q���(�'j6�!�j�Sy���(�GD�A�'�l�`���!AnU1���GH���}��',�(�N�B�=��JG��<S�'(jE�fT#en,}�Gm�<?Y 	�'��`�i�t7��f�5�hu	�'�}un�D�fl�
���'A�
Ū*��a��������')�V/���	�e��rWZaC�'�̅��)R�B��Q'�Xԩ�O8�U�'�X �q���д!�A�5Y���I
�'����� b���9RBX7"?��(�'S>]
�!'c$I���-�d����:�S������Уu�Z�IF�KE`]��y�
5	���@�i�&>�T8D".dў"~�k�<�#��Hf$�7�jP��'J��w	�+y���2�`�`�А�'1b�RB����'퀶�:4�'�VmFK�H��}���C6U��]��'w���Cg� :ܜxA.��J�����y�)�3� ��3a�88��}��a�>���H�"O
��� �	�ؔ�PQ���A"O�L�0 �B�rX��N�>z@@"O0�IѮE�bd��W&6k�"O��i��|�b����B��Z�"Of��$`�6=�Y�@��,F�昩�"OnX�㨐���4�%���X�2ёV"O�����G'j�D9V��R�� �Q"O*8���ť%٘ )���X�� 剘�p<���A ��S���r���3�LEK�<���ڋ
l�@��ڎ)xNI��E�m�bB�I�e��;'�.Xv\x���h2>B�ɣ~�C��:!R0P�HJJI6B��(*�j���I?(�0PF9'��B��+th��W�._N��7[{@B䉎
 xQb�ON��J�z$��A=�C�	�vj|	#���` P+$�[>Qi�C�	�9�;dŀn�$��)(�jB�I?$�j�*�"����BN�XXH�=ç,�hD �u���]/PT�a�"Ol9��ц"�L��0l�e6Z�b@"O\�`2�%T?�� �W�*&d���"O>,���6Q�a���$Et¨��"Ot=�vM�<ʤ�j���!i|&$Z%�'��N�v��jݧ��)�Q�В_�r����`=�N�'|l �iׄB2�9�ȓc��ge��%�:�3f��Fz�ȓ{b������<�el?^}���ȓ$/80R-)1�0l҃)Z89�L̇ȓOt.�7BM?)�̣Ԁ�3=�y�')0�=E�t���C� ���]�d.r���V'�y-�Pؚy�Ak�6a%|,�$GO��$;�O`�S�[��s�e?�j�"�'��I�	I@�I ��p
rn�0X��B䉪,@=�fO�E�j`�g߀1�Zc�t�<���iˈ\�Qb�B��X�Q�$O��!�<8����<�հ���j�Eܓ��=�5+�:+s�0��n�G��E�}H<)��D�`A���<�\t�@�;!�$;2P� �M�:�y�Ԛ[�!�d�Ba��7/	&3ar��<再�ē d����_p�]�qNI~�*��O��=�����&Yeb������}�E-Zw�<�w$�]]�ċ�����x:��<��I5��j�\�R*&P	�"�bި�ȓ=Ji�a��uNr���dB��R̄���@�oA)�8�W�T�S��YDy�g>�S�Hɫt
 H�D�Yx�*���+=�yrB�[�p	��1%=4	rՊ�3�hO���8Z�����H:4��1�=!�Dѝi@$S�@и-9T}q���%l�!�$Mh�W�L�(9��b�%2=a�۟�%�`�F��FI/OWZ�Vb$D�4Z i+�3�C�K�S��"D����!RR�P���>��I�w*?D�$; ��z!O© ��Q4+;��:�S�'}���c�&@�M�7��6m`�4���6�ad�$~H�"A����>�	�X1X���ؖ>T�3Xj�����|$��㍾Q?�e{&��eZ��ȓiJF� �j��x��
�X���A�� � ,!���,f�@k��M�[Q�@�ȓ\a�Ԋ���?*X�!�'Lα�BE�=9����4Ή�����äc�d�s%fM�y
� ����@��m�Phˇj(s\x��"O��a��΅J�HD��o̬Yg9��"OX$��-�,d@=���h�Za��"Of5��_�m�@q8a�I0	�HK��'��O̜���
�Y��lܯV��x�"O҈�U���b��#d������7"O��صBS�g�F<A�L2���;�"O��*�EB�'����"V1i�t��7"O��t��?�D����jc}��Od(������"�&��F�=D���aՇ{�����ϊ�;$�, � \Ohc��KVV�=���`��\�M���*EM=D��a�
	g�<��ڿ�Ak m9D�d��AU�_����«x�|��Q�$D�T�DnI�Uk0� 0kA�F�x�X��!���<YBί}�����@��n�dM���}�<Y�S�k�\iv� �v���$�|�<�0-��{vTH�2�Z�e4)cF�Q�<�A��m��*��2t�հ(x�<��(� d؂Y
S�
Q�P�c�v�<iBꈉfFFTU%��`�Ȕi�X�<qЂI
`�0�)���;<WV9H�EQ�<QE*��[N�YAŪ8ʒ40���I�<٠�?y���㋅(h(� �Ҋ�C�<�o8v��l٣	���{焊z�<�U XQx�5C�`4Oh�����@�<���J�SΥ���EZ�u��@|�<IP�� Nj銳 � m�!��z�<qQ�ȅs7l���O����!�S��M�<��NE��pc�ܹ%]��ZC�`�<��F�W����섪gҴ EΚR�<��٣?�P��@�F*9K^�;i�<��%N�ԑ7�����O�`�<�&� �K��i�eS�P�r�Hu�<)V��?'m��"#"N�X�=
��Dk�<	#h�c+&�򫑞"0������b�<�3T=��"&_��	�,\�<��֪$��T��H��2���A��W�<9%e@ C@xqu�P�E���0w��z�<A��D���B�V����~	�a*���4Au���=&���ȓ((Xj��C�Bap��J6U~���ȓ?M<�z��]�pqv�P�ņ9��%�Dd�b#�g��Y��0Z�b(��4�J�%Z2#2��BƗX���H�\��X�w?h��6+�FG�Q��s	 u;���^�XT1!�`���3E�aHǓ��������,/�ć�7U�p�@P�l������.r��ȓ4ų��ĕW�$���+v�|���,��)�mX�G< x�g�Y�g���GE��R�PJu^P*�"H	w⼅�eE,-x�kܪf3�p�ab�N�\��i����uk�&FXx�B�;j����|2t�s���~��s3���S�J+D��y`�L70��b��:P�@��5)7D�Djp/R�^˼Pb0�����t�(D�������xu��9� ���b)D�`u�B�T�p@���pV�(D�p�D!&�>A0�YO�\(�4D�4�a�_F��,PJι6$9ˁ�-D�x���m]:Y�MK�o� �2C6D�<0a��#*�����d� Z�E��9D���u�D�Y��)A1���uL��2U�+D�� �9���ϼ�D�
�A��I�tJ�"OPI��F�G���Q
	�,52���"O0�T��?/t�p�����$"O@�A/9@��I˜B�(躧"O�Ѻi��{��8"�d	w,��BU�'���'M��'`��'��''��'����d�*T\� VMDl3�Ѓ�'W��'���'.��'LB�'>b�'Rt C"A<t �"�R�1Z��4�'��'���'�'FR�'��'6��!�`�0�$��i�<�`E�'���'�R�'���'vB�'���'�"yJ1�Y��4��jÆX�r��a�'���'�"�'���'���'���'�,$ⱃ�.mE|�؀�S:ծt�3�'$��'��'�'S��'���'*8�7��)�X"�ް��Y��'��'	��'���'�B�'"�'d=�&˙8TQ$`z��x z�s��'���'qR�'���'G��'*�'�\ ǯ�2;�(Èl���u�'���'q��'���'2��'���'�5c���S%���G�ݯR�ސ*'�'$��'ob�'��'3"�'���'*,]���S%i�&q���� �x�!��'#2�'R��'�b�'���'�2�'-4���2J�y)��ڽ%J�A4�'�r�'@�'���'\��'��'�~���߳F������EP��k0�'%�'�R�'��'r�x� �D�O�%K���G��@S��H�=�l�u
ry�'��)�3?���i�|���	!d���
��q�q ʇ��������?��<�i��U�ˆ�u��aE���J��A��~�J�$Ƈz�t6M6?ydC9r�`��8����Be�y
�Ü2�DѫA���'�[��E����Y�����+8��x0�S�~6홼/�1OV�?ř���c�˶[p`2�ǘn����d@f��vbӦ�ID}��Dj*��f0O��X�ʅ�D�*�B�(
ZlB�1O8 �J��7U�8��%��|��r��]s,5C#�����gD`�ϓ��D<�$���H'�I~�n3`��:!
ى�\9>��?9dS�8�4ht�66Oh�Uc^�Zv��6@Ԝ�Iv�S�z�HD�'���)cO_sձ����cu������aƓ�"�� ��5�>$*5UNybP� �)��<�����d���	GC�2�H�
�O��<�6�iѨ�9�O�n�u��|������<�� ��Q�q���<��i��6��Oq��v���N\��eN��Lh��IYP���@���ٲ%��~�<)�g��@C���QK�=X�6Q�E�S�<)�j�:�6�#�~	�iv� ��S��%	�&��m�7P�ޑ�G���*�p�2��7�.��kj�P)`��Q^z��q��(��g��h��@� � A��r��һ~j��!&�\r"*ٰu�"�VmK��t��Eh�İ5D}*u��7NT�"�CL���$�8l	������F�tjO�K��t	Q�T�4B��|Ѱ z��� S����мo��1���ʣ�A�r��t�2�[&Ol��Z�	4{���v�նs޼�aF΍8
(1ei	�|�����<_�(y"��e�N�jgN�>�`�S�"$R�x��l�hڼQK"� 6C�X��b��b���L��@5C,Y�e0�n	1����G� z���j�Y��\H�Cݛ]�!�N�@>���,vBq� �(�!�$'|� �(<S~ix��({�!�$�]冝z6�+61Du�N !���aa�ű�F��鈒��%
�!�$J/3��r�
\�:�f�9P��a�!���6R�qf��G��Ĉ�؆�!���^���q�Z r��ku�^�ji!�dX�!F@�ڙ�T�5�߬�!��H#AP`mߗO��Y�l�q�!�$��hE1W�2��ѧ��%y!�dM�K�<	�C&4��X�j-Zr!��4�`����t��Sf!�D6"v�As�&ʂ��wc��!򤁪���JQC���}��,5�!���g�z�PD�I4��	�B��!�d�Y��A�1���*� D���Iw�!�d�2.B��`�ӷ=����kH�**!�D�%u�H	���ߐz�@�D F�j!�?e���#���\�����o�!�W�ڬ@�E�<ݚ�V%ЖS�!�� |��Eh�A�
p<���nS��!��ɮ	25"D�+xa�r���=f�!򤝪[9`��BO8@e ��d��:�!�tnLy2X�.�VD�S��!�� �t�Ukݲh�8� �A�,<��ex�"OT5�H�;0^P��/�<�����"O��Xw��!T��q����&{�Y1"OvI�ÎU�
��ّ�J�}b ��"O<;�L�s+n ��DyF"8ĝx�)��b�(9)gF��ց��F)�:B�	�/Vꔈt�ϟpg�\1��A� �O�]3�Q~x�t������HHp���J���� D!�O�)�Fm�7M�8=9-��=9���4�ZeD���POf-�v���Ĩ��ϭH�����2(�P9�EA��>���X�l�|� ڳ/e�T�׋"n�m2�s�<�!��:��ȣ�K	�`�"���<���|���b5B�lr��%���ZЂM@�.
1~!y֣L'3RC�	"�
xR�(L@Ң7>:�"���gu�x���$d��p�1Fxr�Z*Y����,�+n�Rq�q���p?�Ghý*)d�*7��Wی�Q�B	l�f����2�<`z��X?e����$��"�6��/�`����b�vM��PW���dX�HZ^�YǦy>A�uD�~h���V���Z�n"D��"���
l0��q�O=����#b���ӫZg���%g�I�"� �?�'�Ie�$H>T�#�ۊC���ȓ ������V8w^)���/|dtDg_�L/n4�w�"o����CIVW���ĉ�x`��֢D�(z
e����6&a~rP;SΔ��쇒7v5��%�s,L�A!N~)�skG3^�2m���3c�9��f�Pd,��֩E-K�#>Yfn�G7�m����3[:���]?=�d[��@��� @����!D�l��lH�a���J����$b�t��	�
N�E�4!�B mӏ���22��-�%dV,O�xx�o�=�!���7ڀ�7�K���ȋv��q�N��M�Si� 4{���Q���d�)/��]�r
�-,K��q�+N�O=a~/Ӈ^[Nx��E�:1��(���8��(5(��1Z��뚩R~,��������1��0!���f�V�����+!��0�.Աt_������!��Ӻ(��i{����m��$"O��X �ݶPB�1��A$.{��	�6O�l	!�
�-�E���p츢�R�@�p�� -� `8���+�l�<�p����<*����̂�E��Fy�'V^21	2=�axB�����Pj��Zl��!u/Eɰ>G�N�hh�c���Q��P:��Z�r��	Xbbz0	�'	�ѓ�/ʎe��[�Ē�C�:��$��DL�H���x��E��X�i�res���O!DB�)��AS6)ܯ98D}�F��-1, 6O(J&���{���i��])�HA�2|������{e�)�'�z��D�ܑ^�
�`5Ú�B�,�s�O���P�6�O~)���M�tb�Y'�����'�$A�}�d�U��3&�. �e)R` ^x:F@-D�lj@�A#����Ei� <7�8b"h0�64"��!ڧcx�[��&)�v��3 U�D�ȓl�r��DE�kռ��"c�.S��oZ�
v�*�)���f�T�>u��j�EJ)f�ti�C� D���P���5P���o9^�ۖ��>at��G'&y��K��Ia��՞u���!�
ه�	2a
ر��4m_� #4��s^��ADX�e���ȓ$�1���\WT]��
����O���֗>�¤'�>%	s �s�b�"b�Ɂ@�Hs�?D�P��ޜ:��CΉ�q�8�ӯ�>�E��=2�<\����|~��1O��"� :Xt�`
�	{�>�O��&��>qsL���Hq��X���2[��'b:݉��3LO�!J��-Lp��`�4Y�~hH��'Dh`���&?I�L�dfd�e�h9d���/���[p"Ox���Q�41#a�څp��`A��&?aB��Ka�:��Ai��g��<�r�ǻ����M��C�I;�nuP>hӚ]i�c����� �@���Z�_kd-���ѢC��Z1
�G��Z%
�Hj!����7>�����Rv�i��Q�W�č��i��IE����(��g�RR�a M�=KBֹ	T o9�!��	#(��X�O� �$-z�? |h��NK��m�U�ȏ2>PlAR�i��keA#�O�Tss��{2��4E��RG�뀒�d��a�:�򤊻k�dٹ�OJ#4��?�{��3N�r��T�/$%r��'D�XP�ț0^������m�X���e���X�8ш�0�,)h��?�٢�U��	�K�6�C!��<UP��V*R1�2	�$@���6(Ï�^ā�lL+B29���iUd�ɫx��kA�S'w�]S��_��"<yӃ�o@м�u)�p;��Rc�A�'L6y����M��J�n�6z׻i�H��Ս^  ���X��ߴ9�>�"g�ĸ]��Dϫ�0>ч�!_�� ���|�TYR�QO}��%Ĭ�Aܴe�҃�	"a�����y�OTl!�eB޹^�dHA� �8"�,E��'�8���fQ!O�Z����+Y0�x00�C//�𐤥<���p���{!���O3���"+_?�J]���ش`a��&��ҨXg�a#����w|)�ڻi��	6�C�AͧPNDx���b�S�� �hI������O�)���<�L[����G�@#(��!��A��;\jp�u��!�M34����0>	`��Xx4Ũ�c�?b�["-W}�!V�\����2)�������|�NX$ad�*�d��<g.(���L�<��̈́�m�h�@�a^�j`�(dLZ�([L��23O攫2	V�<��S�L>��:l�s3"��A��e�e�N2;����B�5�>�8ug��i�[֨��8�|�Џ��VH(��%�O��3��U�}!��(C�^3"�B��񪂪`#���	�lW9Jt�kG��T��\	���vl�;Hm<E)�� }®@z��S�ԥ4L>�3wݻ �,�CQ��>a�I��{h�c��*m�(G���|�6'؆g�`;P�]�}���Y�-�s�<���7���"p��@K��&# ��(�r70OX��,��&>c�l�*w������D�*��1N5�Oƨ�4�	�:��DQ�鍼_{�rr� R�蜪GBZ4E�����'�؄�$KD7$*��0l�t�b����̦�#U�F�!���[?�P��;Qk�8Q�O�;F����A�5D�2Ǎ	$l�^9��H'p3���(4��,y�~<Q�W�O���S�h�)��9���P)+<�D[�'ݴ0x��L`�d� +� ��A��E�'�.��H>���O��q6I� s���!aQ�N��`�"O�B�.�2D(\�v�۟M��q�'k2(�E��5(�a|������h�IT �0��[��=!6��W&Ru�6O�
�/L�TRP� i&}p
�[4"O�A�hV�r�d��݈L`�8g�$8���؟`H"~r��xy��сi��u5!c�\S�<	�aS2S�-���F9A��p�a˱ �6$1���R��Q��~�خD��V�
(,?��(!�4�y��\���T�YbFb9�DL����D�"O���I�M��H����_\�mį�(o����O^��i���@�1�T�ӷ�RmT��<�X�v
G8��I��"�EzI�#^�,"~���	wO��C`����ҧ�Z�<Qw��	!�*�)�,o���R���Y9%�@��ا�����H���[�4�Q(�)Y��yR��$5��E'��m �·���Ĉz9<mߓ��P1�3h4���9}FՅ�	2:���5,m��0��	|p���D��Q"O�dhw#	����qI���Ƒ0��	}�����4ҧJ��a�t��au�0B���iܪI�ȓ3��Q4�[�P3hD�$�#�B)mZ]JFu(��sӂUڇ���k!�H�&Αnj���"O<�Ǘ�N+�a�c�Ђv��R�tX�,�0>y(�%7�}z(�
�n����FX��	p'��yrB[8\UـnI4���ui@�y2�߯0z���4&A�x��9eO��HO�����Oh�O��9�2�6<X�Uk ꚿP��3�'+�y��@��Y9���+_�K)�PA�4Oג�07��sӚ���D6R^�a.�R�*�D�4!�T�K��-rrPpC&˕O����S�dq��
E,����OF@��r10��	���Io�dr��W8R��ƀ �B�)� `� FDXpo�l`���YN��`"O�a�S�!Bi;�kG�y1Y��"O�r�GPV �{��z3<IA�"O�A�`A-Uƀ�@�i1+�r�"O԰�Zh�-
��˯-
�I��"O��I�+���&�SE�΅j�!��"O -9���FpV�D�J&)����"O����A�@r5��Ɍ��0"O:M1����_���j�l��%P"O�ґ�R+��9�-U�p�Ӆ"O8<��K�c��-��
"H�h���"O��cN��f@��+�'����"O�T�"��=-��H!j�0�Jhj�"O��'�߇3�-bW�ͫ��I{�"O~�yj��\~� F���q��1D"O Y��#&-"s*�%S�"O��s��Fnž�Ks�L,e��<�"O�B#MЎ��q��{��z'"Ob(��&�Ӧ�1$��n2�L�d"O�!Z׭Ԡm��p��倣�b�s�"O�a���Ӳ�1��A,g���Y�"OD�����^޼�C�ڷ<5����"O"�KsE#�i냉^�})��j""O�d9��<OІ0�c��L$Fdj�"O�E�Q70Q\hrF�>)��(��"O>���a^:6=F k�G�	Z����"O�z���)�ڬ�̖5:�n�sP"O�8QF�-�(�3�ʅ�Z��i$"O��b�D�w�Ҝ���:^�2�P�"ON!p��*�^a*cS�fGB`"OT�!+��3�`�RrAӬ]&�y�"O:�q"oO"SAL�p@g��3T"OX!$�Q�<A�[�	Y�Q�|��c"O&Ek�[id��sC�;s�riڃ"O��@��%l:Yꗆ<w�p�&"Ot�z���~��L�!%pၴ"O�<:'T�^h��NC�ɰV"O$�hsa�:D�L�$�>~}¦"O0��%ש,�6�q��09?�œ	�'.s�W,���6�x�Tq�'@ax��^*�%���5~5�
�'�(Ժ��&rɐ��'e�La�'�x�ؕF��~kS$R�v#��Q�'.N08�c�2�:UЂo�����'�
��eO3� 4�R�\���'���KS��v�xDC!ڽmΜ|��-b����Y����2��
���t��Ci�i��J�7z,�����-����ȓ _uj�_%|L��Q�&d����ȓkF���._�h�H#u��7d���OA�2��D"I�>kL�p���B�{�o����]�#愠�ȓ�E����ag(,�2��|K�Ї�lN�JD#���"d����&��	�ȓC�n��!+
�RH)&%A�����ȓx��HB��C�N]�v�:/�ְ�ȓc�4�Ri��*�D�dOG-R��܇ȓ_�Ju&� l,1�e���5�.)�����d�h�L�pG��=]^ �ȓt�2)B�	�R�d�0�*�5*p�؇�~����4�ϗ	� Re�gIX���]␼S"�V���X6�ۯ����ȓ<��y� B�]G`�H5(�p��8�ȓs��i%c�\cθ؆��B��,��S�? $�x�H�VHEg�2k:����"O.)9w �
QpF�b��)t7�T�A"O2XiS�^��)���_�X?���1"Ox�{��ԲW������h7Dd� "O���,�������1.A+A"OR�1IFq��9[��@?Bͬ�y�.V�K!n��t�_���)���)�y��b\P�b��L�d��"0D�?�y�f�;i���5-�u�TTJ7���yB��U��(W�G�o�Q�v����y����J0�b�k�=tSܨ�L�y��!�����o{Htْ�yr�J-�Y���s��]�6�)�!�$��gx�d� ޒ���Pj9~�`�'�0e�
$j��H��L�d��a8�'"����j`����G>p��'HxȻ��R�f�U8�e�Pn<	c�'u0� ����P���H��u��'�6���ċ�bR��ja�X�9y*!�'3t�
�EE�/��u󑆎�)�"���'��0��C��=u�zQ�,
��'���ҎM#]��u�e�+�v���'tĽI�`��5bp�*�(9�'ޠH��o( T����c�m�(;�'�ƀC6��Gf�;"'
�|����'ZܩFfK�u�hPRI�5u��=��3/�Qe^0J����hf��ȓQؤ0k�䂤:n��j��O0�`��ȓ\���yqo�A�~�"a�QQ����)}�PΈk���	��U�j
���ȓ;AhiY�`YQ�\A���fq�ЄȓY��yC� ��?� \8��_p8̄�9�����U�r#��R��e��݄ȓCɧI^��H�q�啙I0��&i�bLQJ���!��9$���r���@.�9�$	�iQ������-��H���)M& ��SM�T^hi�ȓ|j�م�5Q"A��!Մ{V�p��_��k��ӣ"t��4˃6�T��I��S'���82�9a�F��J��ȓ �	�C�\�P�.WyԄȓ	IZ	��=q�b(��Xx�^���2՜a�a`�ZȢUyEbP�Q�0܇ȓY^@M�C�M�^��ᢎ�L��t�ȓ7F)�U�ML�^(��L3_�N�ȓ����!��7I��  �B5,�����iO恒�U�c���V ��'�����`��9q�Q�(�v\+�	�d;�фȓ5QƄ` %�7�����'P���sl��P��ܞl����hC?E:�؄ȓI������\J���Sw�%$8��ȓ&��ز7_�ހ;B"�wѐ��ȓ^�
q��L1�-sD�6d�}��_�X�!� }t���U�r����E��,	�$N}�1��eN)�ʓf��{$��	}���(�nÔN�C�I�m���+�-�+:|@*5��ijB�#,Rx!7��5�P0Z�mؔ~q>B�ɵ<Jh�FA��M4�8�$�6_�B�	�\��XSR���=Q�xD�ǈM�RB�	�9��S*(Lf�;�Ø2FB�	���h[�'$���b���<�B�	�-�b@i4��`�p�� �B�I& 7����I�4��S0pn�C�)� d���Ü�py�q��0i��@E"O���4�w���0���7�$� "Ox��,�5.TC�Y:���b"O��x���7P� ��͖�&�li��"OP���G�/l� ��&�;e�8�!6"O2̚�e@�'�h�kB��
$�V<C"O����
�Z�Rg�-D @t"O m��/SI�MH���/��p"O���ԭ@�
�j��
�} "O�ࣅ�<cv�0;� ǟ�A�1"O�sp�Τ!�x!�F�=&i�Ő�"O��p�I�D��`���ܾXp��1"O�d8T-ʁ0f��s_-	_���A"O� ic[0+b��J���C^j�у"Oج���'dq�P��M�V�@�"O���0-WRYd�����Θ;"O���M�#
ٹ��E�.y�1"O��p�ȭ$Z�3�O�%����#"O�\R1홧�"�)G/�3iB�J�"O��P�G!\<Dn�.[^���V"O�)���_�6�RAP�ZE�"O��bvCI�t7F1,�����h_\�!�D���C�j�'��`R�Х]�!�DV�.>���JR�d � �!�1O>��s�� L����.A3u�!�	��I�U@�2\�Z���>W�!�}���A'��w��A ���&y�!�$S>L���CP�^�Z�1�BS�<3!��uo�	ӥ�K�%t�ɪ��ñ/E!��\�`~L҂��*z���HC�	S�!��L.� ��N��l$s�F��!�$�}��!�!j�7"�J̺�卑bW!�$ӸQs؈�� a3xH!�N�aG!�^>O5x`Pt�Tb�� �va��;!��)�B)r�.y稬ɢ ��@&!��/B��sHB���da`j��p	!�� �V���mR�u�����t"!�\�m�y�d�=�F�*�ˉ	�!�$݃P����mӛ�b��_Y�!�"F���0.T3D�� �̄ J�!�$S;ڭ;J	l�L���c�!�䜑�8���ĸ[ZJ4Z�o�3!����p= լ�Fp�R��-	{!�ΤKO�eۥ���]�i�VӴG`!��1��Q��&�8��+-߮xh!��(���ړG(~�p�l��i�!��R��*@�F!���K�!�$�1m����Tv2���IV�v`!�D�';H�=� �R�L��C��\!��W'(*he�t��t��z�]�X!�DȽJ����c��;F��8B�$Db!��{�Qʄ�@���� w!�䔛02�P!�m�|8
�)`g!��<�A�Ʈ��jtl��#Ȋ�f!�$�7
��zE�ג	c�%9��	�mJ!�зkf�,Z2.R`��{Ħ�o�!�ӰW��5k�, ��bӯ�!�d�8J��y��zs��#c�v�!��[y�P�7&ތ\G��U8$�!�$�����W�@�|*E␘;�!�d�V������~�<�����E�!�d-j�8D����0����I�#|!�_S�,��`�/�8e �(B'R!��U?z��u�˷�ԡ�%�2/A!�� ���5b�O�*"��Df�ɣ�"Ox����EC^���)�5G��"Oa���8w����j�90�2�"O���C�W&c�\�hF���T+�L�"O�t
Q�H����E�w�ij�"O��{
X�U���Z���
(DqQ�"On�pV��4eq�ڑ�s�"O��8�L߈|wT�x�^�_��0�"O���l*xm�0P$E�:��u"O�- �d�5z�t���W� �4��C"OR���3>C�tA�� �m�1�"O҉@��H��is��(S()ٲ"O�P�t !�U�T��<�\��!"Oԕ�5넶)fB5Je�, ��"Oqs�C04"��p3��X:\�j�"O`�B�$H�\�Z�Z!�	�VAPhx5"O��3�l��	�Lˆ-[2���	T"Opy3��oQ6 #�Z*m���@u"O��-C�*�� w����X���"OB��B��&vX��F�g�K,�y���;r,�vk�
�$���Y=�y����� �j@
lT4B��G��ybCN�!Ԥz4�����@�e���yB�C��,��  �X��tM�1�y�Í���ʆ��OD����y�+��0���PeȰ����h���y�d��w|�K�fQ�
�p[��3�yRF�~tni��*��S��Sȟ��y��Y�c
F5�t�1P� ,r+޵�y�gE=A�$�����EV �0���y��S7��2ƆǙA�2����L��yb��$����V�
6Q1d���yҬ	�l����I�:l% y�#l�-�y�I'���A���h%.�2ȟ3�y���Y7��1S�2��� �yhǑ��]�&�Kp�]s�CG5�y����1<ܒJK�<�F��@ߟ�y�B&�|��",�gB���DǦ�y�i\�!f�@��\�eS��IC=�yrΎ�\{��S�T�\��A��/��y�O�)��02��O�n��KZ��y���-J^�ȋ+NdC���y�'�4y� �OU�b1�1����yRMB3"d-�v��E�B�����y�W�C�,��m�<A�řeK
$�yb!p>zԙ��2�:�y����yb#��>��X�Q��"$����t�F>�yB�Ǔv����R��kgf������y�d'�Lȓ딿k2hp�8�B�I0_6�2dÀa�E��eX'p�C�ɜmPK�0-Fe��	�'`� ��"O�xŊO�^�pH�aF5QbaS%"O>�����#��Ȧ$[�jC�V\����(Y�0�Ӣ�z�C�	&&i&���޽#��Pk����B�	��}��t��:�ڱ۔G �y�Lw�ݙ�!��7	�Hz�FQ��y��I��i�2�>���J�̮�y��D�o+^<haĦz]�P"Z�y��-�ĩ:��'A?b�ТA��y�:2�$�#Á�Nؤ13�Щ�yҭ�O�ZdK�#F�0Є	��*0�y��C:��5�3
��ِ��U �y"b�"q�8t�����
Zâ2�y
� ~�q�mڦ)��M �!S�H��c�"O$`�CB^-&���F�QSU�y"O6-[�g�_�M�wlҶ nB��4"O��*aN!��b�͉�D4 ؓ�"O��)�#ͬ�I���*{��p�"O�Y�CQ�Y�x�v�J�zm��"O���\,DO*�+�2G]X9�V"O,�h ��U�􌋷VT�	F"O���O�y��3�L_�<U���"O����]� � �4�����"O���r@BT�T�"4␜z�"OV���f�i�
� Jƻ���'"O���T-��c�g��ƽ��"Ol�1�Tf�|X�k�:i��
3"O�rJ��*C�y��c� i��"Op��R-�,����-i��BF"O	�Qڙ���2�..��Ze"O\��J��#�ȉ`�#^�$���5"Oj��%M�w���YEb�~��D��"O�JI;+^�L;vCG}6����"O~ѣCG��P�T��N6MI�"O�Р�JD<��Q�dM�:�k�"O����ߔ7g����I&H��R"OD����C�>���hAK�\E�"O��@�ڧ��@��D0~�<S�"O��(g�N.k%t��Dž3�@LQc"O���I�nn�{C���)�"O�ͫ��B:l<Θ�5d�l�~�
�"O�l{����0��Q�c�%]�J��r"Op�����"M���t���e�V�aU"O�Ȁ)҉Z��1*T�1Uh�"OnX��$ ҵ� Bûz��=�D"O�t����:"��p.Ϙ��]{4"O"U�b�Z7}� 8�P^?W�@�qC"O���2�ة�bt���I��f"OVP)c(��D9Ѵ��>��� B"OD,aІ��ɹS�]�ٴ4C�"O3��#w�X�ӥ�&�YU"O>�3b]�:[d4p��F֒��"O�YA �	,T�>�㶆M(^�a�S"O,qI�
�D>t�ɇ@�|I��"OvIAC��4��9Ґ$�4,���r"O6�0a�^>9@���fe�Q����"O���`o�By���rDʞ#:�{S"O�8���%4�����I�t0�"O�� �C�.Dt��BS�X$ZU��"O98�@"[��CG�ӨGV�7"Oۙ�A q�"�k�O־U7p�R"O�Y��h@�Rt��D9h""�25"O�Y�.]5M���Ü0W7��F"OĄ�D�F IF��%‭7��R"Oq�P �1�8)�b+¡j
E�b"ONeɑ���Y����ͤ\J�*�"O��z�G ϰ��s ӊZ��4��"O���n�|�f�Տ�UJUZ�"O�i���E��F�af�1s+l�B�"O�9�c%U�iWұ���Ɖg�ݙB"O:�rrlF;![�����4$��"O��Qtj�n�"k��Xi��"O�8�5&��;|�*#�B�Z	p�"O���tƟ�D��L8f\2"�����"O�:�B#4,�h���d�dx%"Oz�z3b] ��H@���&еc�"O^��B�
�_��,��kNN���"O� j�4C��,d2h���J����3"O�t;T�^r��XA�Q�N�j�2R"O�QY'j
0���ġ�?3� ��""O��У�lG� �a�U�|�tUp"OTl�U�:
��9+p��/t~i;�"ObEzӤ�uWTm��)R��I�r"O��C�
]�a=k$���>�y"O���D�F�S��͋=`���"O����V1fu� �-2K�a �"O����
ĊC�s��pJ�\b'"O��Ƀ0�P�"�Mѡv�X�0"O���2b���	V��nw<�A�"O�xt��/Eh����
�Qu�y�"O��&�́l�,lh�	}��3"O�t3$�E�DPȉ �c[�ؖ�Z�"O\Q��^�0i�ɶ��P"O��R�b0i�T�j�菕!� T�"O�E��bK�V�h0��â^�y�c"O�Y� &�#}�>�9�%$tҩ0�"Ov�I#�;�~��H[T����"O����ȃ�Q���@� =�Рt"O|�����.������[K�qѷ"OF@(a-��>�	��ˉz/���"O��Dl�3� PJ��S� V��"O�����B	���jq"Qc�*��""O��R�`I(6�,}K0X�'$���"Oԝ�b�)O{ �0��,Q5r�� "O��i�A*g�H���D�=&� "O$�µkC� ��A;����:I*0"Of	��E}��7nS-|��e1�"O<� �/W#y���$-P�6rTH��"OP���1Q�F�tm3x;��5"O��%�NقQ�m]_A ���"O������_Q�@��+ě+ h�v"Ob��.��	˶Cr��
r�$�C�"O�p"s�ƪ\:�y��٧A�F�"O��r��4 0�(�r�
�̉a�"O��U!Qm��8:�ǟZkֱ3�"O|Y���ƙqk������k&i�"OXI�DDO-�����	 ^X�z"Ol����E�2T�U{�E�UP�uQc"O0��3.���ѩ�5b}��"O��yc�w��hMAG�� �oǶ�y2 �+J��(P"��@x5�5*��y���N�&T�eD�5�bi�#+�y2�2pM��s��0��	7�P4	�'˄�*U��,/�!�4b^6B�8�	�'Q�,Oa��b[/l$�	�'w�T�t8�d�x�����I	�'������	|k��ہK�zނ(X�'��]��.�~����m@���'T���)�:���0�@�c�����'��0��
�S�8��0�ZT(�0�'��M��D��0h
Y���2PךP �'�b��g��*%�mQg��3Y�$��'���!�"+�|`&��'-��	�'�P�94l�'K2<��`��)����'����á�
f,�� �^�\�b���'�	҇�N�p0�É�5Q�"�'eXa �-V�C<RI�u�E���Z
�'�Py�e��g�n�-:��P9�'���IUE)	��Eɠ�0 ��-�
�'^ �f°a�@���OVuyX�
�'���c�ȳm���b+]�q�慡
��� �!Z���-R�X �g�Ɓy�"O���/=q�(��wm0eo$ڢ"O %�BڻR�.�����T��k2"OD����_�=�H�u��w�H��C"Otʃ��$,��Ō��U�,*�"O��ټ2�>y���Yt�~4�"O ���C�<l>�1P�
!&s꽨"O�(�!��u�� ��ŇV>��"O@b(��wԒ(E�>@�f1��"O�c�$ԀF�.�
4�E ��"OƭK�)N�TD�a(�z�R�"Od��	"b2����Lܸ`���#"O��i��pFM��Ŝ;}���"O<̈w��(a��h0���v�6"O~M�T��fe6mJ�M��#�F=�"Ov=�M B�����@�V����"O����!�
������N3I���T"O�L��H�[j"��E>NlHI�"O�d	A��6�RE��P8ܜ�A"Ox=��ǟ:W��� �#�"���"OR(�ҧB�q�TebΕcm�� "O4zv�ڙNN����
LL�["OH�R���>>Yf�á!� D��"O��g)��/���1`�Q�lah�u"O����AznȵJVM�$XR���"On-�%��c��x��TI���t"O�	Z�F�AeX%���ܘc��Xu"OܭA�'[?W�]��M�cQ2�%"O�Q�V���9B�)��ɝ��}Г"O��gc�L����Ė������"O��#�-X�����9�<���"Oh�[�J;���s�مz�8pX�"Oְ�e2ְ����U���"Oč�$ ����Q������3"OD�j6IȊr��Pp�Wx,�*�"O�A����M�R(b�H�8?���"O����m�	y6Ld��AI�`�bD�"O����@�*�ţ�F�c54iq�"O�h��c��[��T(���#7"�`a"Ozx��+����M�C�]��'%:��F&�lh"6e�+{���'@^����׻��e��q��آ�':X��%��޼��j���'OT�C�ꖆ(�x�+CldqQ
�'ՠ���#��i(����˘��Eq�'��(��I����0e!�z,tX�'r��Z��l
���� v!��'��hBd�RD�n��BD�f�v!{�'�b��ǡ6���CbQ \�|���'*V�z��E:�|Yڲ��jܾ;
�'�h���˨�hX��K\j���	�'~�$3� H�*.���$Th��(	�'��ux�b�v�r��ɧ@�l���'B�	"�f�b���=C�T��'w
�Q �#"�]Q��$:�X���'�L�#у	�����J���Z�'\-s��2,M�����ss&<��'�-ї��2�D�KE�޼rH4Q�'H� �� I�aPbAadj�j��p��'���bi�#zgX�F�_�[(����'dĹ���G/Pj��<T L��'c�a��#��Y$���k��b�X,#�'Ɯ���?Y$q���S�����'�B4��c�}�q��̜�O��dx��� �ȡk׫B%T�!fB49��AAa"Or�I`f6���A�@)if�B"O���1dɤ&4�Yq �t��"O4�a��I�<��L;`nǢ�r0�"Oz�o��w4���f�6G�d�j�'D�,�QB̵m��)��ʖ�"��5"!D�� m�;����u�ӥ'�y�?D���dO�0
�88$��nr�j�D<D� (��� 5#聧*Z X�E�E�:D�����|z@%1�dmʴ�%�8D��rGD|� � ��4VU���e)+D�������5�UF�=R���-*D�����X5{2���k��r�(D�l���26Q�E1h�:�a�$D�4�.#D-�]1��ÔM="|yT &D�Ĉ`&�=y���1��s�+��1D�$��
3t2Zu����	F�����.D�D���s�Z��ffZ�GK�͡�b.D�l���z�x��7����9D��
�Δ+nsF�*�g��^��У�&#D�,��.ُv�t��ӕ'b�H�� >D��#u�R�E�\\;�IP:9z�G,;D���,ơmט|����{P�P�V�;D� 3�g��^c���3f)�@��-D��"�߳M�
�h�mӜt���Ђo0D�䣠��3v�pi�R,LP�;c�.D���L�u�n!����S$�M0�+D��2��2k�����Ʈ\�4��M)D�|	�#**I�2�H/j��E���;D�<.�g��0�2)B�R�(#S�9D�|��|"~@� �.��\QƩ9D��;��0��8�l͹6��p�bD6D���#@P}�P�^�(�P����4D�$F��	X�Q1c�!� �HCh2D���wJ D�xm�#JX�XD&/D��b.݌.��ŋ�V���-D��:�/֎8,p��h\�=W0�!��8D�H�e�Դ��0���X5,XaJ��7D��b�j� Y� a��A�<�b7D�\�S��{�ވ���ŗ^18m�#,)D�TJՆC�B_�B�.WS$� �!4D����m/�Qp�� ��<��"�1D�ȋ�B5V�X�h@�D003�-D��g&
D ��/��T�}"�>D�$�2È���#��_D2�h`<D����D��,�� �+<�ॠ$D��(�#A�G�(�����6	���[P�'D����!ȇ>_(�۠ �=6���s�$D�<I�Eٻ�z9�o�&��l��7D��Z��40c0�'mȐ[��4;��5D��Y0b	*dz�Yơ�dX)�"5D�(����o7>�I�@�:�4jb�3D�D)Ռ�Y��1 �B)�x8ǀ>D� ��M�!5�Є{��P��^� d�1D����ڐ �(��$�\�>m�p+D�,rF]eTYz�
	�h�+3�'D�(;"��w�`�DE�;>�2\�B'D�<2�M�2�z�t́�M�,@X%�?D�T*cbF�q�xxsl߷c�8�!F)D�؊�Bېx�t9%��t��S -)D���@�
�e�1��:	D�t�#2D���끅xmDa�]�^_��*rJ$D���u�h^�؛� ��E<vPq�e#D��+7�B�fT��n[(+LX�D� D�� ��ʒ�D�E�n0���A��"O�T�m\�<T��9M�'��+"O�%쎷.e���rF%�<��"O�����
�F���_����D"O��	���v?20��� h�L��w"O�����bp�1����3U�x�pE"OXM`��D*}�t��W�޽��"O��qkW�e���p�MΓw|��X`"O���qI�R5�	�x,�R�"OȼBd�#+�K���^�9�oN��y��܅7L�ɒ3F�^})
c�"�y�^0Mm,�CtJ��������I��y�NEW"%Hs��z�vq�$�Y��yRL׆E����ϳo׬�r�(п�yR��!Y ��7)Ĥm�`�U���y2' tPmRE�Bp�����ư�y�i�	~f`pT#!h���0�E���y"`�#/]�ISEo�����+�	;�y��kG����H
 ��%��yL��i����GƼ`���x bP�y�N^X&�e0�F�_����eܟ�y"8Yh���].Ը�6V+�yB��U2����K�QqF��2)�1�y2�A9�"aa�F��R���Ɛ�y"fR
������q�`��#�yR�݋}�.��h���##�6�yR�T
k�u�b�ϧ�"E�J�y��Q�=���R���w֞yK���5�yR#�5�b�0�){�p	e�E2�y�BŬr����k���U#O	�yr�5r5�yYCm��x=A����y�BF�#���c��[�w��(���y��	>~|�p�n�&<���'�_+�y�eFy�d��(V��y@���yr�Ε ;�$���/U�8�o��yR͔e�Ԫ�[3�"�څ�@4�yB�g�4�@L�,D�D1��V��yr��,u�P�{�ͦ/�������y��&W�� �Vs@z�+�N�>�y�f��
�iĿpS��T�+�y�L���ȼr�m�+^7tLӃ���yB�/qW����?[yP	�AM��y�/!>�{�X#k�ؘ;A��/�y�g¤H]@�fKx��TE�Q�>��2v���_<!bӧ4@������ԟ<�F�IA���@�ȓc�F�8v��d8��B�F�8�ȓA��$�c��Yq�A�#{Li��q�z�PE#ġv�n)gҋ3z	�ȓJ���T��~g��h�	��t��Y"�qd�5�a��bFz?n�ȓc6b�z�V�X�T$�b�e���ށ��dGs�&p��?n �����ۦA�
(���[�<ef4��4ߐp��*�qsr��C��+uV�1�ȓ]�	���/�%�U�T��G$�P$@��1���տh�0m�� ; (���ۦd���HEJκKh���<���==�<2�3Z*^ �ȓ'dd����L�EwIٹ)�4��E�BG*]1k���#A��GBX��q��:��	4��M����Ah��ȓj�RM	b�;zhd��Ӥ�EZ)�ȓZ�� ��ǅK�PS��ӈr���S�? t�ȁ#�5{@�j��
���5"O6Pj�f�>kf=H�ˎ�*���x�"O��瑟7u:͛%�ΏԢԸ�"O�� aR�]�a��J��� �"OVA���x��|��Jc���e"O�!�&�8W����ԉ�h}H�"O$<���:VF�����TN��0bQ"O4����q�T��A�Z{�)��"O��s%�F����`�']D =3"O�H��T�/��ѫf�ֱY4���D"OL�AC�L�x1��ஞ�J�F �E"O�	�1*Q�u`X�fNZ(u�V@�"O�l:�B�E���� v����"Oh4��&��y�R�X���Q &"O�!p��G���Q�5Q`��A"O���%X�[���K���r����*O(�GL�hEH�#��T'[?���'5�Ct�Y�-��Dj�O�K��'˼\��D�	�����ŋuy��J�'"h����O�$=�v4^�pY�'��\�d��&�4�F7)L
�'n5���%AA�5���ف'9�Q(�'Q�a�hγ&�ƹ��G��q��'F8D� Oˤ6�r,ܨ�`��'�*[�L�1Nh�$�@�2��5��'��%��ƘR��ʗ�
�9e���'q��C�.�
=cp��%܃G����	�'U¦�F0$���Y�����N�<9��[Ҁ� 5�Vm�f@�E-�K�<�S�X4�p[w��-��tiR'�H�<�ԍ��A�u�_��✛���k�<q�S)&��ʖ��?;�a[��j�<���% J(�D끠Ju u+p�e�<�!�Ye�!Sg2������y�+#",�ZW�ʐ0L��pP����yr��:w��|�A*�� (ּ�7, ��y"��������>�H32@��y��fT��攴[�=�1cۏ�y�d�R�RFMR5R�hPT�ߑ�y"�@�xX��@�Ɵ�8
�CJ��y'B�[�ް�&�ю^���P�yb��y3����A(.���#!�-�yr�ղ۫�V#Ed���.Ͳ ��B䉋!ml�RB(�Z��xW#�l۸C�ɴa��{�iV�RP����7�nC䉳f�Խx#(ɚ�J�oü;bC�	/(�Q��((<zf��q�B�	�
�Fp9���H�U�r�\�QpB�	�S�@YF�9�D�k([�z �C䉋���`'��F�^����vnB�I9�A{a��>��S(�9>>B�I�#��0�'ח@�&Q�햤�B䉮4bjh���|+��2oӉmv�C�	 =m~��'I�u̔!C'�!\�,B�	�V0)�N6\��n��C��!���+��7p�Vab`�OM0�C�	�*6�y�4���C���RfL͜C�	�PQ���0 ��<1eN�i_B�	:���p	����0�U<(B�bڎu�qU��,�7�F�5�C��$˶pUL͛%��}�����C�I?�ldaD*��DUڍ!R�ǳf�^C�	�-�Yڅ��z��:L[ )�B�I;i��s��*�B����r��B�)� �L��پ9����si�壠"O$h�ՄN,��D�2"Ҁ)WhY��"OrX�e���"�~	�1̏=>����c"O���+B;��-�#�<�ld�"O���hWa�P)�
җ@$5��"O���O�œ)�A�x�"OT����,�R"Vw("�P"O����Q�6���FC
)�"Ó� `N7N���U�D	P�dh��"O@U	1fU�7�I�s�B��"O:�E�:ĳ���Z����D"O:<I�"V� ��E���A�����"O2h V��e�dŨ�H;9{&!B"O�$�bE�/l�瀲f@s�"O��Rci[�f��Y�2��5eDּ�"Of=��i@/P�i�hŊa;��z�"O�4�Ë�Tqf�%I]�%ƒY�E"O����a�)	˸� ЊMhe��T"O(��m�MTP�,nM� z�"Oppi��M5`�a��L9|(=p�"O��kVc�;����98م"OT��
˗S���P�	b�"O���Bď:r�M���Tp���"O0M1e�ԝ	҂|ʃm�S�a�"O��P֍��^<�ӧ���@�6���"OT��@	����MI�+~�L}�"O�4�`A�H��lr�*�"�(�!�"O����OT?���f�'�-8�"O�P�� 4W���D��t�Fљ1"O��$��⎨a.��k�y��"O�A3�nRC[���2-
C`(M۶"O@\��ڭQ�8���߉2����"O*i���-;����4//D�!9""O�,����!'(����R��B"O&)��$�:e�rlʗ�]	C�`U�"O�xC�$�N�p舃��U� �;�"O>���� �@���g���f� X�"OjTa�'׍t� �#���%�V|a�"O����''x�����o�vA֐K0"O����ȿ~<LѪ�OV�X��e�"O h#�0�y��]<��(�"O>hkQ"
<&b����;U���#"O4a���I!/�  ��J#�J9B"O !#��3
�1��^�#.�`"O�M)cCݲW��4����%�ʶ"O��j�,��yŮЦ
���r"O䌛�됚Y9 �� ��ç"O����±�U�� �d�lS��y"��2j�0���~����6n���y� 
��$RfS)#�:8������y���y���3��ޥ)�n�D��2�y2kL+OX�]zF��!�� Xt�ƕ�y�h�2J��ds�)ԓ4�\�3�;�y�.E��q�`�Y�҆]1S%P��yҫ��J��HڂE����bd�yR����*6�@�iM3��	�'׎hI7lߕG(T2�ř�$ڸ$Q�'��C�k�iL���+h0��x�'�V������^�	co�c��!{�'��DɵX���[ic���'_�,*׫�/`�(M�"�ܝb�2)�'�U*䀜l��02b�]N*�(
�'��x@�T+�܍���U:��C	�'�x��I Kt�ty���I��0
	��� |Q{TcSj����o�;�&��"OZ����V���ï�;-l�d�"O����&��!bЩ�U,�CT��c�"Obp���V�~58B�']D�i�*O��;��E�r���4h�,ψ][
�'�N�x�#��O����l�2���'��biA��va�R��].͸�'�
�@�X7;Oj`h� �=��d8�'�����"��1�Ə�����'�T�1��4cgH;�f^�v�*L��'�D�C��_(&(�$H� irt4S�'�Xu���m��@����b�I��'�<�8g�Gɸ�у-__���h�',�5�DO�$1p:���*XV����'��	� K�ps�F�;S��D��'Sz	1�嚥���+�NM?��ɩ�'#H�`���)>�>Q:DH1e3ḧ�'���)�g�<{����%Xx�5��'P0��'!�pΤգЂQU���'-&�J3+S�QL�P��6ES�	�' Q�
�;[ �27Omc����'V8ŋP�+L��)����X�>�(�'�Th�B,Q&i��Q�AI�Q ���'#h���M�6t��ca����I��'�A��:��y��ǘ
��1�'��ȢD_9C=�)�� }� �s�'6MY���U��<�iS<x㞤��'n���d���6�Y���Z x�5��'-tP%�Ľ3���y����h F��ʓ���An޸dhN��abٲ34 �ȓ�|,)�Ք[)�p��+X.4V�)��)���t�ѽ<�ڱ�'�Pͅȓv�� tUNd!p�f� #{�4�ȓ+ꚤ2���51/J��a��,�"y�ȓ_��$�uD p|�#��'?Fu����pDոG�\A�5	��B����ȓI� <���1q���R#�[)
؆ȓ�f����Զ��yV�#+y�]�ȓ4��)���Z%O��`�_�x�x�ȓa��yw(����b�DF,�����P�sM�Y��ԩ�:��ć�*������A>PW��� �A9ͅ�2���j��)�2��1�E |c�@�ȓ_­���:<�̠���!�F0�ȓt�������л�+бf( �ȓ"4x�2bΞ�5DHxkf��,j.Ňȓ_,�U��)�o�B1Ӄ�P)���ȓK
�l�m]$NE�,�P��;9Ξ��ȓC~�:4A��Rx���H65]0��I�yA��w�|)��� ��!["O����{x�H���)�:��"Ov-���U/���H�I5b���8"Oh(B��h5��c�6��s�"O �5-^(*r�y�BY }��m��"O��qo��]��-�1��T�x� "OH�U��:��#�`M�5�<�ز"O�ի���e���x� �'��D�"OҰy�΁ X�G��8e�\��e"O�� h��}�ʱ�%�/�h�P�"Ofh�$o˷$J��1�$Θ��2�"O�
��5t���I��`��dj�"ON6�+6J�����K2�"�'L;D�ږ��!�-z����>h�ƍ:D���d$]����LڜA8(r!.D�� :ط��M���[���R�b�"OZ�� ͽ0��s��$a�	 �"O���P��'S�u@�CC;�R�"O����(b��y��dT&����u"O]I⧏�N�䍁���//���"OjM;!������%�<>��г3"O�����\�4UBX3�j�)"�����"O�LC���B��i�2*[�xa�"O��q�k�:p�rf��,��K�"OpE1����
uRp�!)��~�X�"Op"�HA:-tE���V:1�Y`�"O�(a��>�x�ؤ)�0f����"O ��˓�)ԙѷ���&Q�f"Ox�8᪏�Le� �i4IlV�	�"O�͠���j>buQ�ꆗ111��"O$���@-fG�i�� �z^J�"Oȝ�S+��z��	���q��s"O2�0B�sPi�iP�<�B"O�-Q�R4u	�q��[h�P��"Op}i��w
P9�7�9'x���"OR𸧤��xD$��G�k��@"O�t�7dQ�d��TV��9�u�q"O~�yB�K<U�A1_�P j�"O���OQ3QnYjW���j�"OrY���B�7�m��.J�&\*Y8"O2q8��X� �í�Z:���s"O,�I��$�h�l�3�r(�"O� �%��
S��C��I:o2�I$"O�P��Π+����� S��a"O��{�#�Q������A!���"O���ce�(ApH��#THq"O2P�gԶVn�Ѵ��6�Di��"O\�A-U,j����A�O��|���"O��u��\��p1&�U5��r"OXĒgM[""ڭ&���d��\�f"Ov5�DN�T��솣ӤT��"O�<���ؐH���A�MZ&��k�"On�91��:c%�tlR�c��Jr�,D��і��$�h%i�nY�#b����A,D�����s�5��Ɩ�+k���C)D�B�>��I��U�a���B�<D�P���U� I!��� z�Q��>D�����O�Yp�^�i d\�7# D�|�&	��\�d�A(,}(U�3D������&`j$��*7�9�N%D�ؑ�j�8H��x�R���r��	@%�$D�DCvk�$p�nH���<��5B.7D��ѕ���Aph]�c
T�5�i5D����^�0��Bi��Es��5D��p���LN�8������r�3D�|��c�i�ͳ��ҁqT�)�g>D���g�ڲt���J��Nb�ĕ��(!D��´hIO'~ kb�_�شc�I#D��4�ƘAk�cǏ�c~e��M,D����ܼY����rnL�NEt�+�*D��H�	3K^<L�gD�0?�0��*D��y�	W!3\,��� ��N� ă��,D�L2M�8c:��Q�i@z0�	��=D�*R��f��m�t��6[��l�:D�`����\XJQ��`A�mڤ�S,6D��ۃ�Ұ �{Gh˒"֊��C&D�t�C��b*��)A�&}i�#2D�؈��
#�ҍ1�a� �3D+.D���T�7}!z���b�h�.���-D�� ASe�>r�qòjJ�Bd�h�"O��ط�4,���h�@���05"O���ģs��EɈ���q�"O�1
��N�#
4J i�(FP�I"O�I�u�(3�%��#.��"O$d�1��1�@��$Ȓ���bE"O�aa�jV�;ƀ�!�4���"O�ĉ���+��<�����z�@�J6"Ob��3	���ճ ���8��"ODE�E�Dx��!����:�Ʉ"O�<�!��o���f�M1n����"O�����#���C[���'V�y�+�l@J6��5E����yRgۑ
5� ���>:]��b�,�y�S9U/�B�F3�J���)�+�y�)O>la��޹'x�Հ�y���	P%8��^ h}*�)7�J��yB=3m��; bܡ]� ]�i��yƁ/o:HXi$�[� Qb�
+�yrA=zrFX�3HXT�Ͳ��\&�y�,,�x|6�ϝI���c�y��:xܦlC��	8ng�41 �ѭ�y�K��Z(v�R��H�:�{'��yR�����	܉���o�3z!��w����]�m�D��l��!��"bL|��`�3�BE:���nk!�W c) r��D��i�r!�$I?)������F�nP�G	E�*�!��0;&�цY�Tlr��W�!�U�)Ш�C+�*0B���>e�!�$XqK��xb�;���*B%!�!�Xg���Iw(�s�n
�� j!򤛟3Ф:�#�g�PD��� �!��X<zF��p��C�ڈ
U�_t!�D 8޺96��?	�~�K$T�!�D�j6U#FoYOْ�����!�DG�#�\9��LSڔd׎C�	�!�$�9K���z�bȜqd!��Ϣ>�^LY��-+��Ah��K_!�P5�*xx�
"3�(9� 6<�!�D�
#�L�Fc
-���A��o�!��H$*���ߏQ������!��Sw|2QІ�ֽJƠ9�9e!�� sBzM� JI(��,��8!�$>B5EK��H�Y��0$�:!�d�<*�Pa�kT�z���:4c�.3�!��^�R�<I���1� �"WA��f�!�Y"6�n�˦g׎y�D@wO�$-�!�d�ʴ�ȡ8#�)tl�-r!��)e�|\��#�A�!8 ��!���3o�(�q�%���*ƫ�!�5,��ӧ����0�%˛�:�!��I�,4CA���vY��JD�i�!���X�h�zw ҽ?݈$[r���S�!�Đ*&�v�D�Bl��
@�U0?�!�$�x2`p  ߯U������&)K!�HX�(�07G�(2��G!�$��9F���	;b�����ߎ !�:%9d�;T�dн`�A�x�!��l�	'�L�0����daX��!�C!.T�@k��8 ��p�#�w�!��,XV]B��0�*�Y����!��BP�×��� ���Za�O�/ !�Y�<ȸ ��d��.�๋K�;f!�� �*���HB�c0jU�p��yq�"O�dc�C�.yR,�ʣ��d�BM1�"O��ru��dq�Y��hK�NBH�'"O�4��Ț~��q�t�G��mS�"Of	0��ܥ.���مH��E�L) @"Oz������LtR�ɓ\(ƩR�"Oj��wNN�4vb,�l\�}->�k2"O��j���9��`r�C�N"b�%"O*Р�!�e^0Ը��]�L
<�"O����� c.U2U&*c�f9�"OȄ*�膒|���J06�f��"OVQ��$�g���
��a�e"O���L�-wٰ�Y$�ڙv�`� #"O�X����S�`  ~\�|��"O��j�jJ.9��y� Ď��	e"O(	 ӦV��4YÏ��V��l�"OH���
�j���X� L�����yR���^���ɉ�%��1�����y���9%�p4q�lK�_H�I��S��y�Oś1|�iaw������'lG��yr #�F�;E�[�F
�`)��y�)�_�E*Ш�"Fxf�Kg���yB��8\H��rl�!l�n ɦX��y��	>_�mjVI34�&��E�؏�y�
�h��̘PM��* �"��,�y��P�@�fq9è�$j�Iu(-�yRaۨ&����֨J8$�*(����:�y�EA�U���y���ش�S��yң�TN��!b��	L:T��$�y���Ob8Y�z���{����yZi>d�Mǚ3qʁwAQ�C��C��KJj@q���m� &�C�	S�LШ�!ޅ&�x� ��'xC�I�5MF
���) ��q��p�xB�	z�ڤ��i	 !��$��q�\B�ɮx��rt"��ͰY��͉?]�8B䉲u�݊'aڐ'���4G�'t B�ɧr��H���D1w���N��'�C�əO<.=��߶er�D��p��C�In��2E�!-:�
2/O�m��B�I2N7�qA2��& :PZ�	�
ʸB䉹6����3��#8 r�,	"��C�;>q������,��G�-cL C��, �\��&�5$"̹��3��B�	�#�r�@Q-�4@����r�U��B�I7�������H��B�ɗ㪝K��^8&xt�A�v��B�	%'�2H�T�HTkNTYQ���E�B�	g�4%���d�$����C�0C� 2���c���V�zF͕��C�I*O����&�<Dr m@�MмB�I�^8P}:0m�$)��-���2ܸB�I%^��lYF�T%��]��F��B�ɚk��}��ԣ3ozXT��D�LB�ɹSXa�'��1'DTp1���B�I�d�@b��٦+�l��i�#�rB�
'W��hBAA���3��G)B䉒K輕����l��QJ	��4C䉼5hl���LX�"��"6#H7=�B䉩	hY ��!����G4�B��.&���e��&B8�Y ���@��B䉥r.>��劝�)ޑ 㞬u6�C�,kۊ�+A�Łz��a�a�:-�`B�	�H�֝cG�K1g�b	���Ҍ1	�B�)� �A�R@^-r�6�HL�Ht"O^\PōƠUB�� j)�t"O�HZ�m� .�jDBtM���I:F"O� �
��=cq�1_߬�K�"O�	�#��.��@�:��c"ODI D�8q�T��/��9��Qف"O�JA�C�(�1�� Q�v�'"O�Kc@ɤT�HL��퉵"O� � �ר��M{�ޏT��\q�"O�l;o�=,R0Ѡ'%��
V"O�0���X(A ��	UI!(�xq"O|H��[*��9P�i�ز"O�!+�!O�$µ��S��Ts"O�+�g�{"b��4�^$\��|�s"Oxy�+��K*���fD�FζY�1"O�����O+"qsq��<+��T"O�[1�ިU���b*��>6��"Ox}��Q)u�&�R���	��pW"O��[eG. ���a�#����"O6�����%X���ՠV3�2��""OR��<S�R��s�޹b��A��C(D�l���V5�dY)���.�ȸH g3D�h�7�;=�Le	b%ښ1�vs�C,D��9 �DyZ%�V�cѠ��0�)D�X+��ߒ1�|�!�!�[���)s$%D�(3� +A����b�$�h�#D�a�*��m�ps�]�S�`\▇!D��BA��~1 n.)-kO2D�p�F�^�4*r@�4��$K�ȊA`2D��xRa-S�āz`��K��lc�b=D�t�Q��7j���
�(j�HC/D�����#��Ms%��7�td���*D�4h�G��*�
�/��U�|�H�B>D��j�&�Y��U%L�_:�fO;D�\ �Nۋ�6$��CG�W&(K�%/D�$j�%��p@̐�N_>/<�g$"D�|�cF�gS��X�-�>���1�!D��H�B� ^vi@�
u�*|S=D�H(�wB�rO�JX(C��<D���� �:{��k�i� �A(��=D����M�7�)�@&��z���6D��"��B�y�wȪQ'��d!8D���4E���>�B���(R�mJ�G0D��`��7Xu���ȼE�V�铯;D�гWJ�b��|Ce�@�{10�X"l8D��KE���3d��abh�#�*=��5D�Ъ�2Uݒ٣���NQs��3D��i�V}���18tl��l&D�PQ�/L�B0��J#��89B��Dn/D�P�T��H݌xc%iS�):@��M/D��t�djHY���X�*�v 2D�p
b��%��`P+
<s��!�a.D�����(2Ly����f���+"/+D�h��J�޲J&�J�	Il!Z�J)D���t�B�l�'�G�A��^pC䉺5�2T�E/�;+�$�	ɒ�E�B�	�XЊ�c/\?�P R�8�B�	�P�9�P	]>�K��qMBB�I�9�XÃ�%���8��
[�4B�ɂ��H	KF�JN���e� ?�B�	c\Τ�L�W��y0	�9WnpB�	�P�l=��.� `F	Ir��6B�I�P��∷p6���=6�C䉭 e�ap�O�3@�t�`�^���C�)� l| o�-Ipy���Cf����"Op)�@�b-$$���]�2�8�"O�t����p�zV��4~���#�"O^�iר	�,O0�R��i�""O��(��P�C.ٙ���Lh�� "O�I2�`�T;��c#�M�A8dM��"O���Q<n��˵�Ӷ[1d�U"O~������n� ��-lը�"O��ӄj�|e�86�E�G��a �"O���A͕'@�����	�
?z� ""O��G�V�	��H�N	���"O��p���1H�"A����8=����"Oҝ`�M�H��0��,��q�"O����V�%�J�=�*1"O*8BU��2t��!�%Z�2q��"O
���f_

:h�X��P�jy��JF"O�՚W�FKH|	������,�i�"O��r4�@}��m�Pl�2�����"O<�1F�"��A���1y�]�c"Oؙ�OZ�)��pp�Ç�*A84"O\}�4�ʜ-���5e�!3�D4J�"O�hA �HZ�޼)5�W�M�\x��"O�S�H�'�8]�6��!�t؊"O��Cv�O�
uxY@ƞ<�8���"O���b�� �&���%�,^�.t�"O���t�H�F�����㕑K�XL�"O�)�*�OHh84��7~����"O�l1�ɕ��b��H�5��l�P"O��I�N�禍���W��S@"O.�����*Sw��'j	�Ia�U�B"O8T��k?'�B�`5'�x_��Ȇ"O��P��$�qr��8^:�� "O�@b����\��D�?oTj��C"OjH�/ΘN�T���ٯ��9ʄ"O��p�,6�H,I4b0�aN��y".j���0���kG��õ�y�E�<t�j���d�^<�'`���yH���4��L�k�*���y����>I��@5IH�����yR$[�'�R4Ҡ�6���� ���y���(uQ�!A!w ��s�mV��y��-E��3'h�r�N(��h��y�+ �b-Bq�2���(�nCC�<y$�>ǂ@a�2rF�q�o�I�<���4<`(q��[�c�<�%^G�<�
R�r�� Ό�,�:Ѡ�I�\�<Q<����$��Y��M"e��Y�<1�+^�wˢ0�gƌ�ʄ��Q�<�c�.?~:aA�
IU��kIO�<a�����l��ER4x�}c�%C�<��m�'�$�c� �k��K���w�<�s��v�v 2�V:����P�j�<y�(�?�,�E�c��y��\�<���z���L��_N��2OTX�<!e*Ǿt��h�Q�²f ٗ��P�<ycL��g���eȦz$1�u�f�<$��8Rt���"��[�
��d�<YT!�?����D�	5N�P��\a�<"@�$,Ҕ��rḅi'�O^�<Y����E���I$�_)�xYe��Q�<�g�L�-�\�[��L�5��@&�N�<is�L�zjx�v�RI�zt��O�_�<Qԭ��P�p&�Ƙm� ���A�<���ш"��=��&o��q���V�<� .hu�ԡ?����JJkf�r"Op�%�X�wk��Qw�*[��P;`"O<�[�g�):�����b�W���2""O���iG"7�(H��C��ޥ2�"O����I1�����<b���B"ODD0�K�%>�TlJ�D�C�<p�"O4��V%I�Sx�,#�i �	�JС�"O��*����D<D�"/^���u*S"O*���2|0Dz@k��j��,B�"OZ�s�/Z��%
� ��2�u��"Of�{7�Ǽuj�!��.C�-��$� "O��P�«B����m�'�-��"Oʰ�㓦0�٪��@�j��"O���F� n�`�R�8�P��"O^�K�΍�(�L��#��2����"Ov�aRAY�<!a�.�j%Jy2"O��C�L�5!*܌��Z,a�(��t"O�����?=��[f�G	�h�9�"O$$�����v��dA`n��x^���"O���Ɂph2 �A��.<�sw"O>yT��*MG�#@O�(hp�۱"O�Q;�B�IT֑�d�ѳ�<҆"O������oxat�S�"��Z�"O��Vʂ�gƶ�z���_��e"OT�#J̞ ��ҔM�)a^8+P"O�u2�_�@:@����+���"O�Yڅ`�`+|l���zqf$�"OL�S�)���N��+Y4m��"O�{�f���I�A��8:�H��"OH���b����Un[-8���"O�0*a�MZ���͓=H/��"O*�SE����	auO��2��iA"O�@�`H��䌔! ��@"OLQ�mΖ�<rT=�H�"O�I�'k �Qrd �A�K3ڠ̚R"O��Pă]�5����`��v���v"O���u�O�C9VuJ� П/z�c'"O<�I�mĠ�|�����y�6(�U"O��AS��Q���J�lL�)�9��"O��ri[�lqP��#{��B%"Or�F� �0���S���I��S�"OP����yp�"0
V���"O�7Łf�"�x�̘�e�Uc�%D���g�1y�@��/fM�c��$D�4S���h�QFV	ŎA1W�0D�dQ�̍nL+ӯ�>m�,���8D���7��>P(��Cu�Z�0dF�!\�yR��x_��9�$�(z��b�`�5�y���,��X�
͢q��@��	��y2
�(9@$@ʂ��=���2l���y�K�}���B�ԋ	���дf��y¢ � �:XA�&�(�����N;�y	X���y͚���y E�f!7B���p�ʧɓ*�y�]7������<Lj�X�$̡�y�m����
��"D��Aˑ���y�a�"J� �dpU���J=�y�6@&���kO:���	�yb��p�����Q��f�y��\�}�ļ[ *�\}	� �y2�K�8�N��'`T�(@@���̎�y��hT~Dx��%�vd �Z��y�U4�x4�AEU.!y���I���y��S�!�zp�B%�fh<jІ.�y
� �8��
��fbLaV��nW�*"OJ�@�-�$=٥�R'N�NY��"O�Ł"l�
s��e؄��W�,�T"O(:� Ip��
2�K8&sހ� "Ot`�P��h�e^1y`��1b"O��h]�d
5���M���Ї֎!��Đn�l���')pP�Ǩ��!�E)g�@���$ZH��s�jG=�!��#o�t� QH��g� �j�N�m�!�]���E�ȟ�6���X�ٮA�!��R�q�٣���	��@�BOZ�!���<�'`��g�~�f�� m�!򤜲jt`%"��ԅ>Ε"��ՇCn!�$���30E�*Y))��]�4!�䕍:ڴ=��.�g9�q`�B!�d�=6c���+ ��4Ìy"!��ոR�F���O�t�Vp1�%F�,!�d�-<2zX�RoƯ�hy�5��C
!��3k��ABE�}�4����b�!�E�In��G(ADA\���LXj�!�$�
�h9�e'���d���R+!�< �����,�9Z��h���l!�$Ke�,��D��QD@І'��/!��L�'�z��D�)҉s��,a!��:�Ze 6�6�� �Û$m!�d;e��0����.9j���P�!�d�62���j�T��ԦE�x�!��Nj�T���6%0x\�� Ki�!�$Јv�R��P�j��F ��U�!��0%\� �hX�/c�-�ąƵ0�!�$�!i���"eJb�ش�N�s�!�D�,X���`&�yFƹCQ%�:W�!��U<CXre3p��H.La��cL;�!��Ыn���""xdљ���!�d�-E��X)Dƕ�6�V\'a[�J�!�dج%�(�P�!��:E��OB �!��al��qFW"
|e
�� 6{�!��;bش��'�&i��d�Q��y4!��B�1K��K�g�X=@1���)*!�$E�1$��@'��X�,��!�!���]~4�0�/D�;��H��l�y�!��G�8�b13�V�H0��\�!�$��0ʚI�`���8�D,q�f�0!�O�06�y�����, ��{�J�8W�!�đ3��� LR�l�¼���ł�!�ě�w�4��V@�15,��x�F�=[�!���2��pʁBQV)L%8���.�!򤓐�13e�(1������P!�DU(%?&ܰTD_�!�0�N�G!�dߪ ��� ���3LIs0�Ӗ&!�$��$#��jHL<d|�6��+`!�D�Q�b`z�"�{ ,����ڪ�!��6x��M�ha��	�A�!��;B�l;"��F�a+��K�H!��,d��u�ՏL�4$�s�◦6,!���gyB�Y���y(�U���O�%&!�='\�LS�пZ8���D�!��('�xAb��-��)�J+<0!��:�6+�"XN@���?!򤏎!I���,�*$ �'�=�Py�kV�9�ވ(���İ�C�8�y�fZ9B���S=/)ꁦF�y�4�P�#g�,w��cf����y"�ɜ1>��t�L�qW�I@��/�y
� ���"> 4`� $�|u�v"OZ����N�"����	��4�p"OZs�.ԱP5��`� ��K���L��p�\!s��'+*�Qr���d�dh�������3�'��3D��I�t����wx���'�@���5cAD���ڴܠ���'~]
fj?�X-��U ��[�'�~h3��<4�~���>s�|=��'�|�%��B�`�_H�̢�'Y�a�0��	�Yw�O-I�(��'!���A��%zt���R����':N0`曞AB����(M��q �'�΅J׍�k��UdK=F�I�	�'�zy�����;.ʬ��ɻ<զl9
�'W�8��[-RC���a�.f6Ԍs
�'a�a��hR���YY�a�^px
�'}V�
�IĤA��*� ˖U$�z
�'�� �/P2L��r	�N5L�3�'�īu�ډ;�T��uh��jcδ�'��\�Ƣٹ��i B��Sê8��'���9d�1~�U��Z�TA~�'A�(�""���#�H�����',ը��Z�;��������B�2l��'�xAJ������dٱBY�>ھ@j	�'XT`㡠��,a�f]�5C���'H�DQ�G:]�T0��C�#� �PH>��@"�"��<�}���V�l��E`��!�$Y�  a�<�!UH�d̂*��J-c 
6sT�%��B������#^~`��M��~L�
�Eͅ>��5��.<8e���	�b�NRe��%(�`1��
̔6��ax�H�aE�6kh�0��;t�ؕ+O�y#�D�G�ҽS Dn}��H�-�9��cQ�q��!9W"դ�yr�O�Ux��Y	`v�x�ʓ�����e#���r��(KA�M�V�S������)�!Z�"q{��7@�C�IIWHqc�$Ì
$��h�<�Zi��eT�WN�dR�>��)���4��d��h�4)�`��Lit��q�ݨo��}b�]�n�ޱ�&*O�xL�œ�c�	~>Tj���@���D��m=z���v�����C�n6$��z�@Fz�f��K�H����1IR^��=x�Ox�]ZW�8{���"s
�$O�(��'��*��
ok�@����=J�I 	A�`ʦ����˵-R����ІA��F���d��4��L/i	��p�v�L��ȓ_���#`�UӐ-C'T
n� �Q@��<��hE��w�N����|��9�Ӟ��$؃�H�5\��F�L�{�%�k�� i��Z�Vj�n�E��\z!C�/ֹї�"Q�l��ͤ�p>�c�1R��P�ף�u49�eRa����\j�D�f�>��2��>�(LJ K�d���׷LK<�0E0y�@]�W�
b�<q �]��ly`�J��xI���-�:��Q�jׄ`��]�G�ڌ}�P�C`�=§�y���gd~�3R	�!�$�Ӆ���yLG�mۆ��4�p�+%��g��̠Q��7iSp[p�?U݀-^w:f��剈.��8GNE�`a�5�g��7lt�������H�cj�0��d)K%���}	��0�I�!�N�Q�f�1QKvP���'q c�N�9G�0�ۓ��)�L���{�,�x.^��Ӂ�(p-�"wA�&T�'�?8֭V|�V��2͎�$ɺ��@E&D���`C�I�0��D,O�x��0xW��/=�x�d��O��(�w�K sب��@��]��y�Ȝ<�>� G�:Aa����=�y��܁B`Ty�c;�2��G'&�) ��6����H�j@ʡ�܀ArxEy�'�V�Yu-�5),�T�\�p=�������K'%��m��0
Uk�@$��G�"3r\�	TH#�Fy�6��X|�|�"�3*2ũAMD#X�I@ ���'��<�o՘TJ�1!	�n+�<q@�� �B�8�ҁ��g�&9��}a�a�q��B�	�s�\jòdjz����-0(�z 'c& &FW��"��R�Ү��O[fDλR� �@�e��(���U��4l���ȓz��ѓ�.�uJ�	k��-��5���<k�r�7�[D�8���
݂z��������ST�5�T�k��{wh\a{Rm��|� Q��KA���� :�X����}:��׽I89��/ӎW���Ѡ�'��y�7E��'�h���lH<�p���/a榥�P��=[LL�ϙ���*f����j�@
�!8$�I�`)�C䉟raKo��<4ܕ��/E�5+������n	�s�=?E��'WT�ʆ�L�q�*	Z3�M83�
�'���$JȾv�y���~�X`#�'C��� �Ow�R��D��gАDH���k+@�9ƍ
5R0!�D��5�4�C"d��AtMc�.ٖ:!��~��4�ŹH��$m��c.!�dCl����O�B�U��n��K!�X�7V) R ̗fx)Ƀ΀�o�!�DN	X�<�sEsD.T�M�u�!򄍟3B�S �U5P�C�&G�!��'�,��i�$Q���*@�1�!��+آ�[U%T����֍�(r�!���o�Z���ꍂq���Ⓓ/�!�$I'�Q�JN�T�y���O�!���x�pڰiʤi��X��ګ�!�\�YO��ǁ��by����A`!�䌎?i�f�@apPfI��`� #"O|��+�$2v9dƒ,:�f�(�"O��W�סT�0Е�٢��@bU"O�8&�������I7		�"O��C��X�wF��A�C�@PV��"O�'H"�b%xa�I?TJpzU"O�XG잇6.`�@W&��/@���"O����h&�~�3��ڕs"�y�C"OXU{Q,�)��������H/^ �"O�|@	�}�T�A$G �Hx"O�� ��s��\ Pn�&�MA�"O�1�@l�d�
�˴��pGXmڕ"O��˴�:'͐\��m e:��µ"O�Yy�\�/�P�,� Mq2��b"OH�Jc�-7��Kzr�1�"O4A0�	��zA"r$�P�ڴre"OEjd(@&7@aɧJ�E�H=r�"O���@��i�p9R��7�Ƭɲ"Oh��Qc۟J�y���'l��K�"O�!D�ͱp�:����2dN��Y�"O&��P&̀A��Yx� K7j��a""O�u2eV�gajK�@��*\��"O�(hr,�5,B�@��U;DZ�(�"O�@�F��%g�1�I�?r$�$"O訹0,�
�Z��s��)0�9`"O�hI����j����,Y�Q�]�"OB}
D�%A�~�R�̈G�%�"O����
���6U�g��%B���)�"Olh���9Q*�ezp�ɛJ��f"O��[�&�7p0|�ȓ`�(<*R"O�8A&h&}V�m+�������"O���P�S�E6�3��2n+�  5"Oj8�tĈ>�ѻA^,vc�=��"OnxR���96Zh�-׵"�Z	�S"O���Fv�҄-��l�|H��"O2��A�f������E�`k!�C"OL8�%���0��ĨC�2'v]@"OPق�¹j�H� ��d2��1"O��ъ�PRڶe�8�A"O�5����m��o��D	�"O��!��Cr]:4�]cW敡�"O�y�e('�Tm"�脌����'�@�֩L�F��U�a�r!L���'>�`�#Y;=�(26�;M�!�'��q3m��d���I�1��3��� "�r�����:�H��0BT��"O��"���f���&ƶW��Q�"O�Tb5⃆Po�M�!��
�"�"OrhaG�ѵH(��4�ΒW�>l�t"OvȰT���E���Y��4*�N ��"O���qm�#Axd`K�lA[ͪ��A�'�l����Y}r�X�g�3��@%U��a�5����y�k΁�.��4���3Z�HA��W
��'J����K�]q
�D��N��#odL� ��4�F����y�oM< Gz��c+B�/8L���K�%���+"$�(:�剪/ޞ"|�'����UK�W��1�E�V���	�'���9Sj�&)�dDz ��/ ���F�J�1��u���!����I~��|�1FΠZ�B]ؕMR�+n���X�L}�MS-f�ߴOh��!�	kj����F-Q��̇ȓ$,�1����l��!�fGJ %��R��.=Ś�B�E�5"<G��Ӊ:޲���I`� `!ڋ�ybkQT��� ܭE����wJ� n� e��ʝ��o�l��MAu�g�IS`����2v�LQ �](^zbC�I�Y����5f��v4��x ��pv���E�<Yh����I�N���*���3��,w*`�aa�;t�,��$�[�|�R#�q�Ez��X�H�8�뷄]�<�����]��V`��Y�����TF�b(����.vø�%��H�[X�E��cJ�9֘F�D��
�|x k�N��@���y£ͽj��8P���->�ؤhK� 6���Vh�F���	L���C��L<�T��,�m��#6c��`P�GH<q�dW8�B�sW��2:t�c�>~��	�9r�(	+��G��p=����/|	���+�v8�%�C'�Bx����وr0��3����R��n,R4����@H��y�wa�P
'�4M�P,F3(�X��J>�pLF�*�V�����b�#}j� �F�H��A]�a�n�Y'/UP�<�̒�T�b)��)�8~�V��l��
�&]auN��
3dJ>� ���E��r���9��3V���3ᆹ�pf�=��4ڦ�݆me2.;d���SJ
c�8��D��G d��S�	��	��-|O2�lް����s*��CKO��45Ãd� !��W�#�����w^����P�B"!��Y�G�f�1ui�5@HF]�r��p�!��Kq���!6ڬ9�!�&i�2!�DP���0C�޸_<
Z�(��SW!��=@�bԃY�{0��a�n�!�$�%�hD��
V�Ö�"V�!�$1M��i�ɂg��<�@#(�!��ƅx���*
Ǧ�2��s�?K!�䓇H^)�&�L�,�����1j!��M�$c���@����Mх,�!�d�c�M����=��Q��	�7�!򤌱T����h	W��(7�ީ�!��S3iG�B������M�	K�I�!��Kc��Ȃ�jёt�d�Є�Z�s!��1Gpe`q*]!H�H�1ш�4!򤁑[R����",r~�!
�[�!�$F=C�q��O�au�-Z!%b�!�Ĕ2�a�g��j�!ר�2a�!��=��:�
�,z�'(3[!�ѵdԐ Y��@�M{����ޘ@�!�H7v��U`�Ŋ |���b_�M�!�d�6z�0	��	ô.@���&+�hy!򤋄�BIza	@Rt|�����'q!��G��iQ�⊔CJHiC�E}!��דF>��"��.�
!!q� ch!���N������H�[���M�oD!�X�e�h��UX�L��Ja�ܙW(!��!v�E�o�'�hP'��G!�Zq~t�B�͝f$�� �F!�� 0D���@ �^�aӄN� �Z���"OP��Ď�z���DA?vq�X7"O���̎ D�����&l��-�"O�X�2�X��z��a�!m�t��"O�S��֢U3ƕ�R�T4��;D"O�Yf�7_;L���M���5"O�T�pA9d�+RM,ޕ�"O^����1P6�:�R
0r��"OdMZ� µ!��p�s�����"ONefϏ�[l]��W�0L0C"O���!f� �V�a�H�hS"OT����+�. �RgF	m���"O���*	�/ؾ%0�ǖVn(Y�"O4�mN	@�� �g@�!{n%�c"O�̊�CO���RP��%ZP��y�"Oڰ�s
΃>�`y���
#M�U�"O�,�4l�4]�.�1��i$ޜ	�"Or5CTᑊ[�ޭH���h%Fȁ5"O��K$��3��y{�o�>.���"O��d��1<X����N׿KI"0"OHP � ��?�֡��`�98(`4%"O�����C�wz����.Ӭ~8TUpe"OjA�J��dL����ؕ$+*IB"O��F�Ɩ ��hiDm�V�4	 "O����:[�`�Fk��N����"O��jUb��;-<���*R�N<��"O(ł0����9:Š5mi�Mv"O�<��c��e��͑U�V��(x"O�q"L�?x�^1үã)a�B�"Oډ���F!+� �9�#�+S܉C��|�N+Q؍K�y���������Ǝ�a,t*��Q!�yOF(j?r�
G�B�_4�B��Co�b��N<��ǆ*ڱ��'�"�p���&��ī�K<0��uR�'�D(��F�;;��]X�N?va��I4ʮlء��n���>���H�}�@̡q,�H"��Y׃�f��#F��`^�Y*q,���$ԟS��M�*W�d�ȗ�ޫ�!��۞�$�j?'Da(�R�X��	(p�x�P�ɱN�l5ۆG �_���� ��j~�a��J6�܆ȓ}�(�2E��bMn��FN�j	�'���Qg��ɁZk�$�`�Wb�3��>T��p@��S��]�$�	�4c����I�5a��s�^�W��h�D�V�]��	�w��91�fY���K}d����'�4`�UiŨG��aS�Y�@���a���+j8ŊԂ�!�3��Z�����Mt������	�AB՚H�2C�I�dQj�UD�� ��m�m�cP�X&%�RC��8LM��u���ŋfS�>�A(p��k�B�7�j訓�Q!�d?g�L�k�	�����z�
K�+���;&N��U�~�@�KY(D���ò?�H�K���p.j��)Ǎ�lXf	_4�{���f� ���#��t',lj���$��ؓ���6��%0���%b�\R�<�p>�A)G�u�
m�f�O�De�3N�C�Lx̕3���N9�2m�)8�����x�Uo�?rH}P/�]tX���z�<i�.-,�Hu2Ac�	ɢ i��ײD�L���-�9��@��P5n9[�n$§�y ��p
b��F�*��,�QLB�y2��:����G-� -��������S^l��y��1�2��De@]w�J����B��Sa�4~����CC$z^���=%@�ؘ��HPy4�؝	�\r���K P�D��C����@Ȁ�D���Ƀl����C�W{�!�sf � ф��!c�Q�m�P�Ơ̬7䁢ӮX7��O��eJ7_���AFH"o���'������'}���Kb�whիR��y�A�׊�=#)}	W�>*����~boj�E��@�g$�C
	8Iex9���'D���b�ͺe�-j�CFb�|0�P�/�ب3V�!Q6zPHvhF0�d��"h;aQ���f5rQ��1O=x�Ⰹ%\O��K쒍�&P��K4��	�DHn�Acd��T��G�5�T�D��\8�(Xe'��0���&�jԉ'�(��d3��K�䀩=��8�ɽ4�ZY6#�����R�:[��Z�d�<ؚQJ�2�y
� �1@a͓&m���+ć�G�XP;��*E��jK�F{V�@j�41�9��Ffo������#c9bU�ׄ@�{�` �U�/D��Zv�I�)M6Ց�*�� ��7'Ȭg���RD�}������	yu��RFa�[�'J�(��eM�JȲ�!2G&j�X<�x�h %B�� a��@����N̩jn�ȥM�2{��h�ѡ^�a~�����m�"�ʽZ�PQ%	���'�b0ɳ�K>J=�dܕz�l�J?�iw ?S˖p��i�hs0)8P	5D�J�gu$ř#��u�� Co� u�h P�R8q��S��y�G�_���k��ƞyv-Y� ���y�锯Z���#�ޏ uF�+%�Τ�~����z�#�?\O�	�{�p��#�1t�،Xq"O�uA-�Uz���Ǐ8�:�c"ORY
ש�>��l��Y
�<�y�"O*a�QM#�K�N�)����"O�9I��#	�x7炱���H�"OlE1�m�%j_p=�1-�(,���#�"O�d��'�8����M�:Iq��"O�QB�߈.��yx�n0_0%�"O^���3l=�pc�M�)S;ĉ(�"O4�p���y�����F
HD@���"O���4 �4>��I9�&�4��6"O������w�Č��F�:)l�h�"O<��A0Y<m��X0%1l�b"O�ظt��j�м��ϻL���3"O�+�����d=2T�U�̌q�"O����W�	o@d���ؽn��y�u"Od�	��Ij��rǍ��KwR<@�"O� �a��R�аu��&~ح��"OniR����T�7��,pv֘�"ORu�!i�0\����(��5d:��"O��xb�אm����6���r"O���ƒ^(��pF��[�8(�q"O�L�(Q*e;�5Ѡ$�0��D�E"OH�"gi߉40>t1!�ܖy"����"O,q���Y�m����уR�u�!v"O�����WSV���$��c���"O֘jD�]Qx��XX̜(�"O��)�DP�}��T���߼s	P]�`"O���B�G�~{J�ħC�g����"OȄ#&��T(�9W�+	��|��"Ov��B��b��y�B��c"O��d��I���a��B�4ݫ�"O9S ��;�*pV>��"O�UB���C�īE&D<N�6=۠"O
�K��
b
�i!EK�
�&	�w"Ou�� ^��U��D(|��@�C�<i�B���z0�p|�J���<!#IQ-�P�(qg' J9Re�p�<�MV�����kU!T�f����X�<�$L�"'X�8���#�~��V)�|�<��j�%WA4�X�`G	��)SD�t�<i�
�xHj�h���� �Q"PM�<'M��_+ dyD��2�6��lPK�<��I�J�t�s�@B:6�ɠ!E�<�%K�rGt4#�/�EY��u�B�<Qs���7':���d�*bu��A}�<I���^��X�1`X&t�sqER�<!���U���7�!qqx�n\I�<I�Jɧ{�\L�'�Ӗ*�&� �Mr�<��gS//^�D�M4w$P ��s�<iUO��Tx�q��8�`Ы O�@�<)�aʫS����C�u�0DsԌ�I�<�AK�*��AI3��9a�[�m�<�� (8�";b(DO��=�.�P�<�  u3u-0�\1CS`ZD�\Б"O�!�J7����FO��7�f,b�"O���D�6����oU8� "O
��7'��Qrq�`,���"Oڥ�hG�B���I�-�Lc�p��"OJ=�v�X)U��aHM�rAx�I�"O+�.u����0˟�m��Q�d"O�Fͯn�@��-�~	�Q"OՑ'��*nH
�	 ��`�����"O�cGE@�9���
�%��� �"OB�
���"5`��r��Zy�c"O�h����or["� q m@�"On�U�P�t�����דz��+�"O�Qpd'3<Ӣ��	N^�.\�"O|��������r�8v�Ԣ�"O�|�&��-cH�QȀC�?�:���"O�D���G�@�*QB;_��1��"O����(A"% �b�aˀ�f��R"O���ES�&�x`!��9r�8�E"O|�i_��V�ࢪ#Q��˵"O���roړA0�t��I�9 C�0C�"O`��!ݚO+��SR�m��,y�"O��K���08����9	y"Op!���X�?z��A,,9�13e"O�%P�F�7_�E��F���g"O*����?��ɗ��><{l	H�"OpȦ���I�� ��Dy�6(�6"On���M�S�5�Go�D����#"O�d�5e�-Xɔ��c���C����"O<9�Q�k��!b7�L�k�J�K�"O��ZWmCkt��1F��p�F�u"O��[�0vP�9ӆ�E<n�"�q�"Ov��gB"��S���F�S"O�S�+�QpBAJ�O�tQ \��"O�D.�k�Ł��)7(,4�F"O�K��yش�3e/�R���1"Oc
ɼ[f�y���G�ϠX��"O,M;4�R���c��xM����"O��0�n�.*d�hPR�@g"O��:`����hE����!t��"O
L��B�H��P*�-a���"Oz
�§G_({�)J,��	"O������$��Yp!��|��J$"O�
�	�A2]�����i^E��"O��J�2?�ܤE�H�h��ـ"O4��2oĎJW�A��B�qZh�"O�T�琣A�ŀU�bŁ�"Oթd)I�(d�á�(A�v��d"O�q�Ш��o�>�X� �`�.��*OR)�5M��
Ea�o����'y���g�I�iф���f�=f���'zP[ �@�z����6!Q'o�բ�'z�8f%$?z{����>���'���Ӗ���'�
]�u��I����'���`���֬X�?}�$̹�'��R�㏂U��ݡ3��3vF^���'���'��U��@�;�8i�'�B$���*5��@�Y�G�lȢ�'��]1��K�1D8Ұ��a_�8�'s���A��j2<J�+�bXꌢ�'e�Q)v��0O��<
Z[�j���'��2�ŹZVp�uA�UY ���'����@�
;�Xa��7N�����'H�å��~�n�!��5><�]���� x-��n�W6	`	R�	�����"O	�dAB]�&��t�P�v��"O��)�KOL� h�dW�T|�R"O u�Gh�#B.j�`�bY9e�(�h�"O��@k}���VA�@���{�"O�pU˟�/�@���3Ζ@j�"O�ܸ��=��4R����XIv"O�ܓ��=&aC��M�1�"O�h�,�3� b^1��a"Od)�k��,�`��Fl̃4t���"O0�g��$�� ���S��J��?v٠�9b����&?�I�|�ԯ��ҳ�՞���B�ɞ�v��A'��J���6v��E3���� n1��'���|�5��;%���p��!�({r���zH��DҐ�t����"���k�7O&	1�o�0��%��}RI�B�<�x��Q\ﾱ���Z2��u!D�CwH�'ea��K�	x��@�C�rmqD���,�vm���>����#X�?7�H24&�;�o�9&�lAA�b�#Q��'M�݊����M�;/PLqu�֤E���A�mc��+#�$#<�'Ÿ'��=
EJ�sb!�4!�-���q�@Q���I����៨�p��<��x�2M��`������ۚ	V��'�����S>�ۓ��\�1&�;K�fY�b�?=���1���䚨��d�'&�� �H?V�>�س�F�Ts���'���keʓ=*j0C%GP ^�"�F!SN"�s�G�z\����k0��4⍱|&��7��L��'8Z��:Cā�i4)ys�b�遳�N-3E���f�7ƛF�C�������Ե�88ʶ�� GN�[Ԡ\�%PJ�=w*6��9E�P�OWF(��B�+wEެ���M;|� ���'S�Fč:	�ذ�כ���(�ӵ��;��W|��Z�Z������1��0{�����$E��a���٧ V|��:zj�EZ���)Ӡ1v��q4NOZ��Y��4��&��O�?��6��9��0seo%�$1�O�O��;���>a"T���fٛ��۴v0��P����9>��>�Ra�(�v��t(
>�1�G�əQ~"<�~��!����# cŬ�p�@��@yR�@LX��PgH
��ȝ��X1CvUir*>D���ă4�IҠW�.����
=D���B�_����2mVJ��C�>D����% �P-���Q+9�\�D0D� ��A+I}���c�ɶ��o(D�|�ūQ�M2�H��I�z:�;D�$#rN�<|�t�����%�pi��%D�|�e�۞X�1I倂 %�`�ţ(D�l���[�K�0����́C6~����(D����o��d�*g%
-x(Aҷ�'D��+�ႎcvU��"�9�Y�D�&D�l�b&�/��x����9��a*D�A�K��A�L1�H�M2��pO6D��I���S����0&��p�.D�����L�@��a���a9Xx�+D��H֪l�(�Ї��>}1�xs�4D�p�EABH<(�kgoX/g�,S�=D�P�ҭ�8`���1��Յ�~��G�9D�L)�#�L����L�  8�+ G,D�L�G�Y�|�x�)�)#Z=R���=D�D���?Y�"u*�%�8HLF�T�<D�("q�����8�%Y~�L���;D�ȫ�"X�R�6���BB5y���:T�`��NU�/�a�p�Ƹ@�2��"O,qcc�^"h t�@Fm�	+�JԺ�"O��[��߯C�	�"�,l-[`"O���a �~� ȑ,��Xr�"O8|:p
�(K����`��O�.q(�"O����雡k!��p�lP>mHtKp"OT��%`�[�`�Ë�[7��
�"O6���"��k$���c
�+nH�z "O� �*�
� [rH��f�ٛq�.1C�"OV�h��T�I� �[9k����s"O:�7Nݗfu�� N�4F�A�"O�e(5�J$,~�xv�\=_�l(�"O�Iz��V�� �ڞs>�% W"O�h%�ӢA
Ju3A�E0q<q��"O��$Q7/r��5�M�U�p��&"Od$�B
��T����A�<�����"O�p)G��2�h�p�E�;_h�;6"O�H�����G�xq,͍L ���"ODJ#�C4o��ep�_{O��8�"O"|�u�U`��!Ǜ:=Ha*�"O:Ѫ!�8Q�0�f+�0[�"OT����Ӽ��7K�H�9"O`MQ���Zd:�Ӥ]�g@>��"OXu��*�#g�"`�4�ڙ *�Xj6"O�݉f$��#fi+�AʺJHZ'"O8�E�i� �(@oZ�'�ĕ(a"O����Тf�v ;e�	���y�"O�I�0`͏��Aa�S)Lb4���"O��#�i<26�9��j��=;$"O$���B�L��q�
�L�HW"O. �)�<y3�]#!�`MI!�2D�̹��E�Ŭ�!�Ȋ^�'3D�ti:3z0c�G�p+�xd%2D��MۭN���5�ʗ|�34a2D�4�ׁ�P+P�#p��#D(d0 �5D� � ���a��+�ƐH9tFj2D� ���
Q����W�^;�E�@E1D���F�
BReN�(zh!h*D�x��Bͨo����4�J�q	���H6D�亀A�8E���qA��N��} �+8D��녌��OMD��֭�,x�)���6D�H��NȰg�~a��B<���"��2D���v��#8�{P�8HXj$C+,D�$9��G4������f�}�7�'D�xs��M�� �+;m!t�I�%D�����0�N��㓭cP)���!D����G�4;��ж��<l�V��v!D���D�
z#�a ��k����!D�஘6bph
�e�w�@$ё��;�y2ˁ$mg-��Q�����E��yb�U�Y�\�'�J9������y��?)����2��4�"�A�y��*�֔�A�X&rU`3b-ʬ�y�hj0���>T���� mݥ�y�$G� �.=���/$��I���y�2^��7逬xF��ej�I!���u����ߛd���0���W@!�� �R��2ឰ �l5J�K$p\!�S+9��U�����K#��s�EC�B!��ț�(D���!��ʃ��?!��V�E�����u`�	�ʈC>!�$S������`��%F9�Û=�!�J4���6cĔ=`��c���=�!�dY ��uyC+�&mH8�b'U�Yq!�W���uj$ˊnD(l��ƈ�E�!�Π�H��C'J�'�I��+ ��!�\����r ��?2P��Y!^ !��:;��Q�X4[�8B̗7t!�$>}��3ԀP9Y�����}"!�D��o��`GE�0�N�16��Q6!�Z1Y��  !L�1������^�!�D@�Xr
�)�/"�n��l�"B�!�� ���fM�|"f�:���>��L
�"O*��`-�?F����(΁Z� �"O�qC��~�q Eȃ&y�P2S"O�-��gќ,`�<��G�n�5cr"O�CՃ��	��D�xidY�"O��6`�<7�)�T�yX��"O���E�e�l}�Q[5V�̒""O�:"�>�邔��d-dE��"O!K@�ޙz���"d钀a2Y�"O�d��H o��P�0Ti�G"O����j΅M���W�K&.s%�`"O�@b[+���h���!]c��x�"O 5��J[3*���S��(T�t�@"O�a�#��S����t��27dQ�"O�A�v �!M	�y{�a$cI��Ѷ"O��A$��2�Bq��&G�3�x�"O��c�K^�v+�a�t$t֨�"Ob�0���F��� �=4gd�)�"O��5EN U�"��R��jF"O�k%Gٖ&�HH�eP?���G"O�|����p�*�d���`!"O����jғq��Ya�
�0؂m��"OȔx�#��� �sR��#�.��"O�dZ#�T�p?h�Ad`�S�t�*�"O�};^�a	�	`N��k��)J�"O8�S3M�u�S�BJ<
�L5""O:�Q$JJ�Cր*�bE�K����"OV�K��Lgp�@�c��z1��"O؄�!B�=B� qôcX<���R�"O"����˧JɺA@r���K\�R""O4� �Kp�Ј�^B$T{�"O�qᢍ����C{"�A�W"O@��wGlB�P7H�.t���"OR�����SU}��&W*���Ñ"O���Ei�?ZSl�Y"�R A� �ئ"O*AB��J�Q6l�'DV�'v(��"O�t��P<zfPq��"��*S"O`����(�&P�a�F��,6"O��Q��W�e���%�H/�8ze"O�,�#�W.$��c��Xk.:!"O�q��`\��c��K�a��"O"��p�uͼI�~e��a"O��yqD�TE�����%S�:�"Ox9��X�fV��$�	`DR�9�"O�@x�,�'o��XKcč%�P���"O�e����6~�g�RxXi�v"O X��2��0�􋓅�@��!"O^X�F�[��tT�k<i�����"O�H�(7a�P�$�J,S6(��"O���Hw���`ܵV�i
�"OL�2*^�e��y*E&լ���3�"O��FY88= ��עH`���u"Op��������s��,.��"O̥���&��#����T��"O�͒� PS6e@S��T�VA�'"O�ekdOǵYW�A�4·�k��4X�"O�ܻ�囃D@���R㆐z͢@)""OJ�r�G\�(��A�|��ba"O
A8�Oga�͉���.7�IG"ONIpn�t�����ڠ~gN×"Ox����v�]0P"2k�b�c`"Of�P&A&Fn3�!۷~�D S�"O���a�(Ģ��e�ڶO����a"O�d�e*E�J3 �ї�T��$u"O� v�R�R�Q�QY����}����`"O������t�2b+,e��Qsp"OT�����E�~�y�K���A�"O�D%��s�B��0�ͰlN=�Q"O�����0U���Ib�R� �T�#"O�ࣧEδlŞ�Pf�ފv�&�{F"O6`�i��v6��hG�m��M��"OFE0R�\�F�L�[�Gѳ,3|��"O0�H�M�UǑ,Q�Px�"O���ϕ$Mt4��&��3Yp1"O�����P�u�!y�ᓪ-WZ�r"Oz�JQZ�p �e
�7PVթ�"O���B% J�I�E�s7�`;�"O�e��d�:Z��b�*I�\(l9S�"Ox��$:����X9r'�X�"O.�ñ��#\L��[Fo��9�XB�"Oؕ����?u��58Rg׫�� �"O$��3����֋I+�P3�"O�Њa̖/tD�`I�DN0��4��"O�Q�ϓ_Dh	��-(���s"O�{W6�Vu fC��*Y0"O\�9��\�������B����"O��AѴS樉�0�Y�/�vTS�*Oȝq��ʱ��D�W��(>��@�'�F47��,?(,�`��	0��I�'�ꬲRĎ-U���;�KY$]��'�V�ɄLDw�x���o��Q�zd�ȓ'�X)����N	��E/_9���%�d��N����.�5�b؆ȓB���B�R�&����$H
�����$��!BgQ�*�N�7L�/uXr܇�Q��Q�*�t�H��.+^ڐ��ȓ����� �<5���ክJ�T�ȓ)��أ�C.*�@�³(��,&~���^�|��#�9�Z�H�O��&�V���Adh�� ��:�C���u����y�2��MVm����'��� 6�h�[�o�Xh@��Y�#�����Z��ql�>zab0i�x���E��4�K�	ȼć .i \�ȓa���  @�?�   u  g  �  M   =,  �7  �C  `N  !Y  �a  �m  �y  ��  -�  ��  �  *�  l�  ��  �  2�  s�  ��  ��  =�  ��  ��  �  ��  |�  �  ��  H � � { Y" �) ;0 ~6 &:  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h�>��4�O�OL�$P�)�*��1#�� x�j�'�.M{#��.��OW�r��۴o�����Y��ʗ��}]j���[1Vl���0D��镅�'/d���u֭o���j6�a����[��u�GZ��𩁮ޱ�n�������v
L2l@�]�6�8�Gx��]n8�p�e�N�1W�Ă�e�e�f�j�*<D��[��5|
��(Jp��g��B�1Ȩ õ��r+Z0P'FͮVn�0��$.�s���'�r<�s�؝j�j`��M$ĥP	�'L����-$(P �I�#��t3�yQ�8D��'��Ԣ��Y*>Π�RC�*�:��O�R ��*�bE���"Y��xg(�O<� ��C�3Ǆ� �	�I�qS�K#�S�O����b�=
����ʄp�iM!��wd��ŉ��=�q)�JF^��Ty��@s���'`�<��I�=uytEy a��]��	s}b�x2Oǖ=�4���� 3��$#��Y��T(5�<�GH�<K׌P9�-�|1o�RX��Fxb�G�=,�H�ՉMW|�A��&#@�0ؓ�Q� a~rV�%��q�IH�#ߌ=�V����$/�I�<��'��VZ?��ɰ\���*Q�
K�4�#D����>+��qw�����s��`����{"�O���) )ަ|z�ĩPB�L�h48�'[�@����@+���7LR��
�B�O��d=|ON(2 ^<
��]�S�ȟ�Dl���'��I�C�� "uH�7/�(���O�u���P؟��ވY�<mڥ��&s�X�R�(D�����-M���P�ڋe=�|r F3D�����yu���)ƚ)�,U'-}B���%�֝D�A�xx3��B �ɐb	�	>/�(���M��F�1D$6ˈ�i�$-�G�J�<)W��I�����I�1�Ȥj� �D�<� 2�:�#�^f��!���c��8d"O��P!�L=8Զ�(BI!w͆ԨQ��ݺ�HO���xE�
�A �X�̌=�"��=A�5N&H�UΜ1}�AmDE�x���	�<���Е1$�<X���#K>Ԡ�dX����<p�ԴL�f�0��#c=Fm(U�Yi8�(Gz,Ǒ�~��DO˯@��!0�I�y2��2P��$`�遘.xZC��B-�yr���
��A���)Cv�zv�	��(O�(�㉠4� Ӣ���-Z8�@'J(9��C�=)"Ĉ�dg	�"��Q�a�&ك $�O�I�{�ʀ��]g3�\@��6ci���K?���>s��9����T��kJ��2m��'�?�k���7:"�#��9��4��k=�Ia�'?�O�D�11 #V0�կ2�U{.Oƣ=E�$N1,>U1ቆ$�)ۂň��yR�?Dd6  ��l	���\��y҅J13\��
=K�4+�OS��D%<O�7�ǟ�(�憞*#��`m;�I	��.|Onc��he─<���Bd�dFle@�<��4�Zx��`��a�ܣ�"��v��Ї��@�I�U3$mYf�"p�����1B��B�I? T�*CN�cA����!I0#<��)
E��,=�Hq�,� T�$Pթ�X�<V&ۑ(��P)�P7O� ts��W�<����@�LI�2�2u��hc�i�T�<A�� 1�(����"1R)+Ũ�N}"Y��F{J~:��� Y;�)��e��V�QU�\K�<���ն%)
�1�a�A^e��H�<ѷ��y	���E��:K�k��F�'.�$;�,^L}�VhE�{5\����˄E��t�ȓY��9�R"'X>�#r.Y=*b��<1
ϓ�?�e؛K=��K㩖9W�.hu��_<��;��D��f�A�z�����m��O��	S�O܂�Ȕi��0��D	 �ښ#~x-@J>1����h��O�M�i�?'�ZG"A(�j��>���	�d3����60
 s�B�&��۰�IEy�4s�.��Ǚ�/aT�s������D+�O�A� K�(GH�Ik땅z�t����'{�	��@r2�.Dz�����EG��'#���pbj��g?�*�W"d4�m9��	��G�� G#6.8P��t1n���yNQ�VФ��$�~�|�j@�0��?�S�O�L!���[`�]�� 6��ыy��)�Ӫ(�ݹ��ރsOP���i��XOR83��M;ĉ4bHx��G�(Q����W�<a����<���g��L1:�[�RX�`Ey���/���1d�
�����֢��'ў�O8E;�N@?r|C�2\7����'{�����ж�"H�(>A�8x�'�:!hi���1"�^D�x���'�2  v��9>}�h_�H�$!
�'���90i̺j5��y6a�Dw $i
�'�10��79�tDK��IF��
�'�� �@@��2�4�S!bΰ8�\-@�'5J�ca��!������\�zΩc��D:�'<�� RSM�-x�E`�J�6S��ȓ*�^�{S@��fG����F�z,��s� ͫ�$Vy�"��U�C�1)���M�����A	 E���"B�E�GMxd��//bh�W���:A�M�1��;���ȓ[n.H�a�ڰZQ��{׎�91�!��Q��p�Q��+�;bFL�p�^`Dx2�)B�@X�c�Y"��_9Y/��0��QB�<� ���"j���<��3K3b5i�"O��@��W�(��,�=8�,�"OLi�3��U�<�Ӏ������uP��J6@%�O|��B ]dq���z�pۅ�'��	|�ĝ��pA+�&^�jtqAh�<�!��dU���.SUl�ҁ����>������≬F1"���g�:^�i#Ճ\	�yb�Әw��c!�����
����3 <mڂ'8����"|�'*6��F9��h��ֲqrJ�i
�'y�U -3O`�U���f���h�'k���ɴG/h�XF��=�� �CO�g�J��D�>�M<yw*.G1�(@���5��5�HZI�<5@�5;b�YD�8�\E"���B�<aSȄ�#N�Y �
(5R�cb�UE�<yq�ҭqJ:���ٚ<
��C/�D��p=y �Ӧ`"�+�%l�#�CH<ѱ�מ8�d:��8,E�(�f��!�������u �N�(�!�h!�6K�B-i�(��Y7dKwaW����R��H��,(�J"]Nd�ₔO(��"OF�+�H�(%ڹ��@��l�ܵ��"O�m�C.R;��wO��DnT��"O
T���G6���Ԏ��J�I�"ONq8�a^�Tgд[��}��A��"OF���OÊ�@@�+s�х�TM؞��=Q��R�ޝ8G#����y�@KT�<I���u����`��=����P�<� h z�H����,.��i���u�<U� V�y�Ҭ�!Q�v�;D��)���YH9[e��6�ƴ�Չ-D��E�M?$�.XS3.͸:�DJ�f8D�ࢲj�)��	�EH
d��@�*3D��`[�Y�\�`�H��c}��$b=D���dΑ|�b9SFf[uϠ�a�K.D��j`�A+(I��J�n}Dt���'D�imG�Vp��b+ƈ<�&`���8D�,Z&�E.���!&��<���P.$D����>SX�еG��]��zcb#D��[��I�;���ph��V`ʅ��L#D�ؒ��V u��8���5p�-1�<D�p3FD��L�ҡ�*j��b`�9D�$����y����!E�����J6D��+��[�]�@��1� 'F��1 D�Ԣ�T:��2㋟6�R$���<D��B��?��C]�q�D@Ae�:D�`��F�/TA�z��Y�{���x�B=D����f�w�\�BO\rӴ��V�9D����(�%R���A��@7 =D�Tb�$�^�x�[D8=���R��;D����R+h&b���"�S|��n&D�<���(:*v�!q�0�D���!D�����_mƥxԄ �ʵ�3D�H��G�c��]�Wf�(\YBHB3D�|r"$�8&+��P-k�޸�c,D�d�UŃ:~��� �L�]+�Ĉ$�$D�\J�L9;�+�1B�PDԉ�y"�N�{%�H�$��x���5�y�i �s$ç. �C>e�ւ�ybꗢKbެ�2i���\�!����y2�0J�"�hFk ��Y2a�/�yR��>�|�&�ܓC%�(���U��yR�J?G �W*59X��8w����y���H��(`���46z0�&@���y�@��w���Ε&_�	�i��y
� ��S��1P\HU���ޖn��%�V"On�Ic)Q�N�p����+�ruy�"O���2�?�Xa�9$�<�"O��ǩX`.�$�2�� �\���"O��ʤ���/�()z�ꖂ6�����'���'C��'s��'��'�B�'T��H�脭{/ڴ�:i��qa�'���'��'���'6��'��'�T\�r�U2xI�2�ϚA01(��'���'b�'>��'M��'(��'��}�a3l
���A?L]�8�`�'Cb�'���'k��'���'N2�'F����R�L�n	"p'�~+Nax��'M�'S�'�r�'�B�'ib�'O\����Սn0<鸆D��?���W�'���'���'�B�'f��'+��'ά!*�a��g��<i�GH�^ �����' �'a�'t��'�B�'B�'/TAi��R䭨Xk�2���Ο �Iʟ�	џ����d�I�x��򟔁�	/4�X{fƖ���A���H�����	ן���柀�Ix��񟬚5�E�{b2��FI��	�U�����\�Iϟ8��՟��ğ��	���ßD�%b������jlV�!���ʟ\�I͟���֟`������Iڟt�I͟��3HG�{5�R�V7t`��g�韸�����럄��������	럀�S�E)fw�kdΎ'm̅�����h�	�T�	ٟ ����L�I��M��?��Y,)�А��%CBf���G�-lM����������!Pa�D	2Oȴ�T��/��h��e�N�)���4���ʦ�b0N[&R�P��󮌜C��R�ş�Mc�w]4���4���)<'
�)ׁN ��)IWbT���)R\ȴ�RD	;�Pb���IHyB��H�L�����'@����ü;i>D��4�j�<	���f��5Y^^eh��&z+�	��o�To��M�'��)�ӡe�\]m��<�!��$�`=Q@��u(H����<c9��)i���$�hO��O~D����'9R�{���?�T|�=Ozʓ��ӛ�_��'�p@C�� ���AF��EGJ�����y}�d���mZ�<)�O=�U�ҁ?���g"B�(�Z�b�Ta%�"dji�G9�'n�q�;e��L�)�@q2d(;A^�x��h� X���ay��������9�p��V�#ؼX���z������4&$?��i��O�)���Ո�B85�ıf$S�O=��ͦi
�4�?�
]��M��O�ı�$\�JE�yp�K�3�pAzLB�0��P�޴7��O<�S�g�,V�A ��Z+6*ڰS��Bm~��']�6M��d�OP�$-�� 9�Ac��#ـ�i��@KA��O�mZ��M���x�O �D�OB����%C1q(�5�>Q���7�B�!<$8�S��Ҳ$����� \�ty�)�3�t ����F;��ғ����0>Q`�i	Hk��'�<9��jÚ�m�p�ڼ<�ĸ��'w�6?�	�������}�۴~��k[�hKF��I�9N_;���L��LԻ��d6?B$;��I�_����l�NG>%�:�4�M�]D�{�)��=�#�O��˿u�ۓ5RXnARa�O����O8`n�!H?��l����|��Q�o�r$a��G$16��b.�/�O�`l�)�Mϧk�ԙ��#RQ~��Q�g5�A;��R7�x�q`�5�:	�"����"5�g�|BZ��?a�	���n����#P�	ph�S�'0�7���.V���O����|�f	�.,�v�
�臘,�(	�n_j~")�>	Ҿi*7M�{�i>Y��L�b�(�L�Z�Ni�E�{��&�*�-@�Ȓ&D�<a�'B��@�l��;�`1U��!��u;��=V�䝠�(�A�B��]B)�4��|�tp �� =	ye�7z�T�a��	��ᨑD��a:��Rf�C�I?�(���?��K5�ںpLl����+��H���	�Z���WN�+��#�i�>x^J���*ǞZ\�iVb��D�|��@S�
<	�B�p	.�{ �Ƞ?P4ԑE(v@젨�g��9,p�[@�Mo��ܨ����?U��a�ȏ)܎�装ӒP[ƙ@���1�lJ�0F }�1`�*
Ɉ����J$��c� }�\p�#>@����ӷ�� �-юz���?q��?I>y���?9�/	�,Oz��%b
�o������tQ�����d�O ���Oxʓc��=h�O�2l��F�i; -��芓�T]��4�?I��?qK>A���?!�hE5�~bc� �:��F`� [�ʇ�Ͳ����Ov���O�˓)d�},�����z��n���B�$�ik���y�	v���|�	����=���֣q?��;e���n9B�9e�����ڟt�'��!Q[>e�	����GV0�H��+���x���.��(M<����?��EV+�����"*]l Ҁ�7�L�q�K(0�VU��������?����?��'����)i��\�+��h���x��Ųi��'�<x����R�(���g�5~,��`�/��m�R5��'HR�'��s�4�Iğ�����| RG�	�r(�w.��M;���������ā�oUFɪ��]= �9�%3%��nZ埠�Işt���ty��'��'��� �T-8x2��Y4�qT����O���cf%�d�O���OP��R�lT$��k/�T�v��ߦ)��,
Z�'��'���|Zc���;Th��P�\�%�e�H���O��4��O`���O\�,:إ��dY�����2%]����c�B���D�O���Oj�O���O�M� ��x!d�~�Px�`���V�P������?����?�/O"x���?=���%�x��X9���P(w�j�$�O���5��O��� t������ �"��`��Î)so���';��'n\��
tL��ħ}g
�A��dkڽ�����6��S�i���'���⟠��$q�i�	P�)Q�u�ʌ����!8�>x� .@�Λ��'�W��"f�Հ�ħ�?���Ƶ]�uȠ�. ��+$F�Ք'���'�,���'��ڟ��s�ɱ��?���u��i���w�>���=�*9[���?)��?9�'�����z��
��OE�T0{��iXR�'��S�A�����O�,8z�&�;���� sr,�ش�j�ıi�2�';��Oj>O�����䄜z pH]��q�l
H�&d�!1�"�'/�'�D_>�J��)r�'p�n�U*D"b���㦵it�'�� �%}4�O�)�Ol��ΉY1�V-����i�R��W�iR��'\�_�<�J�g~R�'����Ow ��ÂY���[p--67~6��O���A{�i>���ßX�'v ܁��g�d�9'a[;
���o��D��#�|�$$���O
��<!�m��7a�<�3%ü.d����p(�8$�x�']R�'|�	ԟp�'"k~}�fܗ��i9�$���d�O��O����O��R���6��ܰq�Ƨ?]aY[Ф�_���I؟���Xy��'`��ӟt8��G�,�����:c}�E�R/D����?y����['>1q�����ųpl�GPH �m��M����?�*O��|�����IO����`Ջ���{�-�Vx�mޟ�'`�-X�SI��۟����?ט�	Ĥ�F �*�n�Y�ڳ.�tOF��<q��BI��ug�4Vò�"�j�}rP�
�CZ>����O�D�D��OR��OP�d��Ӻ��)�
���:fH�d1A`�Ҧe�	ay�T��O�O�61�A�&{� �a�D�#���
�4W�Y���?����?a�'��?5��4}~��T
Ӷ1 20����-g�"|ʤO
<%�m�@�T�b- ̊��C�:'���' R�'-(�BW��'��	�|��\��bT=M�6��ɐ�'Y��1����n������I��<�b��$-�˓�^�}���@��M�x6����i�b�'��'!�맴~��5��D��
�{��]#J���D�!`��$�<q��?���?���]Q�5#��/+��P�]9~�f����E4>�v�'R�'z�f�~/O��d�!U����$:cz�KB���@<�LP�5O���?y��?���?�v`
C���~��U��$��1g�*5����4�?���?���?/O6����\v��99��1a!�krH��W=4q�e�'Xb�'���'�ҠC7��6��O��DZ�]�`��6�4 ��-ɂ�n���P��Ɵ`�'�f����>9��Z�eE�@����G��Φ���ş��Iן�3R���M���?����fED��ZI!�":z�H�q��V����'��͟��4ax>m��]y��M��b���	2,_B�x��e�ަ���ߟ��aE�M���?�������?�A�/0x�ЏI�)A���6)U�7��	ǟ��ˋ�����ןl�O��'/��;D�\LUiTJa;��n	p0��4�?	��?A������?���d�+��3���-��9�wJ��Ms��ݹ�?�+O&	�O��O!r��v����&��!�t��k��5>�6m�O����Ob�p�Xݦ��	�|�	ԟX�iݭ��f�>�P�T"�/3�(�۲�p����?y&��<�O"�'x�fU�W��	y7���Q��%��L��6��O~���"����ԟ������Z��X�I6)�`�{Z�֘J�Y;kƌtI�4�?��,�<)/O����O���O��DUs���*%&�u�rQUc0H|����!��ӟ��Iџ����`��?�PO�%UrG�,'.�qdH�r���?����?���?i���?��n�f�D�=�l�pfV^9"�.P�,w�6�O|���O����O^��?�k��|jeK�\�(�9�����y7���L+���'=r�'���'����

�67��O&��"O�|��#$�?z�*� $��D�2�l���d�	şX�'��	�>��$�>ђ.M�).MitJ�J�^(�Ԃ�˦y������˟$���^ �M����?1�����eN6o�21RTm�&Sg����!?4���'u�Iߟ%����ON��|nڈY�\����[���م����6m�O~��Q���o������͟����?�IW:f9��t-
�R���'m
��O��$ GJ���>�4���OL��Hs�ޤ"��l�Q��+�dD�ش4J�kb�i�r�'YR�O����'Q�'��a��K�8��ȅ�s
u��ef� e��O�O�"�	�O�y�4D
�o<,�!�-@�oǦ���矄�	>�­��4�?A��?i���?��Y�r���R�T�0�R���="�ln�I�0@t�)
��?y�OM�� R.^5
&xT�e��"�~h�4�?ɖ��V��v�'�R�'�ҫ�~R�'��	��Z�E���CuH�k�aګOd���1O4�$�O��$�O��d�|b�ナ���ޜK5,L"6�D�k\��xF�i?�'�b�'���'����O�9���i��]%I �&�}�˛P.��O ��O���O��$�Oʈ9�ۦ�!"��ȴ���D�`� �Z��M���?��?a����d�O���?��Ơ=I��+v�>&�Pр��M3��?a���?����?�0�O�V�'z�@�3o� �����Ȑ����sFL7��O����O ˓�?qA��|
��~
� �m���|n�a�'X�c�4,
�i��'-b�'t�8��a�`���O��4Q��j��������@�Ȧ��	~y��'G�`�O��T��sӼ�`AGZ�w���c�'��nf�Z���Ol,�"G���Iɟ����?)����L��-�.s'daӥ���B@��P���$�O��!�ON��<ͧ��S�%��9��)�Fmr
$�7�ϔX;��m����Iß ��&��'!���d �f��=��N��?u�\jv�z�2��լ7��R�'�?�0 �f�(��gM�_�F=��J�&�'���'_(m���<���O|�����@`��T��"�Q�Y�� ��w�
�O`�43O��͟��RË;'5F�Ce�OVYr�A��a��';w�؛K<���?1O>��t\:bd�> (���n�=)��'+Y0�''�	ƟT�I����'A�R��6cKT���
.-7|Q�C(�9'm�Oj���O��Oh���O�X���K�25P"�Ej�B�R�&p�1OH�d�Ov��<闣�<"���@���]z��Ƴm?$]��L���ʟ��I`��ʟ��I%R��Ik+����9�~�����M����O���O����<1��(i?�O�d��%آ~g`�G�6�谷�n�r��.�D�Op���'���"}�iG�">)�1+H����c��M#��?!*O�	r��Q����S�"�=�H�0[� ���M+|2JN<1��?��K'�?1N>�O���Ũ	�F�P�c���t^���4���U C�f�o�����O&�iIz~�-	�oll�I�"��C0�����E�MK���?ɠ
�<�H>�~"Į �<�K*�zr�����\Ҧk�����MC���?1��ҁ�xB�'� p3�I!M�L��J���^���|ӤI#-�OR�O>5�	�&�|�DBV�?�<�!�)S0J�X�ߴ�?A��?)�� ��'eB�'��R�MJz��&'Fpf�x�	M2:��O����.�D�ON�$�O4)�Q���4.�e�P�d:�a9���馭���C6��qK<a���?AK>��@|�l�b�٠z$ea�C�7<���'�6���'Y�	ӟ��	�`�'�
eSr�X�E�x7.ʇ>���34�+��O|�D�O�O~�d�O��1��G�j�H�
�I��C��X	G�N���<9��?9O~*�!�&��
et�+��N Etqp1�^�?	�������O�������M�r��3:~r�*(S�w�:�8"	��>����O&�d�OT��<��J�kD�O��u(fG(���B҇�X�]���j�.��7�D�O,�䔃f	���+}2nG^���9���L�q�G��M���?�/O�E:p"�o�П�S^���S��W���l��*�@�5zI<���?�k��<�H>�O5��0��II���S :$���+ٴ��䃨�,m���i�O��)R~2��c_V%#A�N�;tV9Agi��M���?������?�H>�~
W�^�.ў�����k�T����1������M���?����Úx��'��U�*�~)�ì�`[:u�Bp�ly�a�O��O>M�I�V��Q̾&�r�I�]����޴�?���?i�N�؉'r��'����)�`V3�>��$�"/՛f�|dǪ�yʟ*���O��d �O��[�O�gndtbl��m�⟬�tB�6���|R��d��Xޒ�Rt��n��Ic��� Fp��'W���V�'}��'�b�'��i>Uh�!%, ��G$Ü7sx93CCú�'xB�'0b�|R�'1�B�=~d�27d�/�|�z���`k�0��I�����Or���O��T�~t�7���b %RbH��cT*��P�W���I���$���	�� ��Ť>���J��)�vhɈ��A��H\}��'��'G�	�
	6�I|BA��5� �z�$�*�b���~b���'��'���'.��}�K��m��(��ų[�����M���?q.OJ��Dv��ោ���ms𜻷Jϛ���Ef��*�`M<y���?0/�A���	�o���2�ǋ;�0PnG�C����'[���8$f��'���?ѕ�5����̳6j䍉hתlz���۴�?q�%��b�Pl�S�'0�nt�3JD�"GB*F��h\V\m�L�~=��4�?����?A��;ى�����'u�hBd��5D����ק1+��6���f����3���@	�.W�'~��yѣ��#��e�3Y���'~��'
�Z��Ok�O������-�����E6	�(��t̓A���@����'�2�'t���3fSjv��g�7i.XK��i���D�5_H�'����ԟ`&��X4�z��F��|�$o[	n�L-�9�<A���?���򄕘hQ� k�
t�Ics�R�&�@�D�r��L��d���H���T7V��"B�y�>�q-Ol�%(q�0��T���`�	�t��/[8�M#5%J�"�J��%A��-
֢//��'�b�'���'O��ٟx�W�s>51d�#u��4��p�&�����Mk��?)���?i5Z?"'���M3���?!���*�F�GK��o�����ԋ����'���'��ޟ�"&e>a�	F?ɵ$K�A� $�)qMF]�`��ڦ��՟ ���,h��J,�M����?I���J�hV>�1葚1,�yK��:+J���'Y�	�(��hl>A��؟���M�7��%��(2 �\/��!�ʦ���ߟ����M����?���B�'�?�f�
/L�5"FD�20���i��I����MK��P��Cy�O��g�? x��&�T �4Bd��r8|]��i�����|�^���O��������O6�D�O�I`E/�.k@��&�.5�����i���Dޟ��'��맼䧧?��+[L7�质^'5񪁃�!�Z���'�"�'��:�D}�|�d�O����O����di�D�1R��'��9Oq�J��i��'���蝧�)�O����O%�`�:Kr�y�Gr����N���I-K��ȹڴ�?��?��1W�_?��G<PR�L���B�U�t�&u}��,�y�P��������`�IFt@7�!Z\]�oL�&��`�e*¾�M3���?a���?Y�^?y�'�rEńLaN����dx&�hjƉ	r���O���O\���O��d�O�9��@�æ�9E��;$&�5r�MλAf��ˠ	�*�M���?q���?Q�����O�Ӣ?��!ɲ�9�x�c&�G�BԞp�RO�b}R�'a��';��'�ypD�yӜ�d�O�h0�Hʰ1����LW,`��XR!g_���	؟��	dy"�'~!�O���'��b�jى�l q'؎D�ިx�Jh�����O��d�O��������,�I�?�Z�J�;@,�JBFE�.36�2���M{����d�O*m��2����<���ѵ+ӕHE��j�B�b�4If x�t���O�\A���Ц����0���?���˟�tǍ
=B�	�$�ަ�)�g�0��$�O �@p�O���<�'���@�]���@�h�LMt"�	a�H6��b�RlZ蟼�I��D�S�?��I��@�	�b� 2�D�)A �xE�D74�@�4G���`����|bK~���nC(qa�M>I@ �d��.CؙU�i��'���][,7-�O����O��d�O�nS@��f�ٛ>�ppYu��=����'�b�'N�uꛧ���O*��ONÂ�)L�z�
U�t����ަ��	|=`A��4�?1���?�� ~�SV?Q�͋�#ў���G[��z�B1˞�	��_���I͟��	ٟh�I��ДO�pp�Ȗ��9��|�P�(�E<9�6m�Oh���Oz���P��\����"~�e��ɪt�9���>��%ڥ�y��'A2�'R�'��'����Kz�0�a�
�21Y��s�cBY9�!��#
Ŧy�	���	��@�IXy2�'�H�Oi��)w��&)� <��c�T�K�c�l���O��D�Ot�O���+bnӪ�D�Ox�3,�ir�d��ٍU>�AEc�Ħ��	՟$�	Xy��'�$(��Oa��O� �%/��8�θ�P1kZn���i�R�'�r�'>X)�T[>M������)y�|`�Va�5q3���H��)�=��O���#jN�P��T?%"���(d<e��ɐIt�@K��~�2˓$V=:f�i�맲?���E��	n���a-F��~l���р��O��h�#=�i>O(��f�� �$��ō�(@�U�i��4 ��'�R�'���O
��'1�'kZ^��Q=�cv�\�&q"�4M�J��Th�g�S�O��5z��h��
��_xtIZ��`�z7��OZ�d�O謻�M�o�IޟT��H?�Ĝ~���!LX�C Zo�gu��<����?Q��s`�BB�\�,�B�bpaO 6�L�к�e�i|�sE�"�$�O���<����t�R�J=hf��a�E�*�tz�S���3e-�	ǟ���P�'x��X�d ��z��0AS�d�,�8GmѼk� O����OB�O����O�UpJN4o��d��+�"4=�aj "W,�1OF���O���<9v��(v�	�7��|�B-�#d�Z���(^�)l�	՟���{�I՟��	����X�Ε�Aܶg���*A�6~����'�d�3 l�:c�U��` IH��Yt
W�
Ǆ��f˓�_�)�:��$N�"ǐ�kĨQQr�<�ȓ)(X�� �9b�éO���A$� A$wZQZt@�0`�SŐX�p�7 �S+���тE;sې�!+�$\<�:f熷7��ē���/ު�cVGM�]
����D!O�`�[�,�:hi�4{�a�-��U� t�v�ʅ�Zo�Xɒ&��F,�&�*���U�,A��+Vʅ
 q:���ޟ@��5�̤�EGF?��-�W�gc�ÃJ0l$,�J��JD�]q� �q�D��'F�0�򮔌(��Ya4��S�\�xe�Ũ��q�#���`�d9u�_`46�ݳj[h���CA����91qH
���A��'0O���!����?�������|"��:�`D  �( [�������y"�DC�E{pf�	{�>��E����'�� '��|��Y��psÃώR�F]��L�a�P=I��?����*�������?q���?�Ҵ��d�O��wH��s� ���mx��U�O�`�'�G+)�i�q�Q9�퉄q��ͣT!Ėr�� q�Ė�ro��a�%[� I��D*��� �?�SE�"m}N z���b}�#�p� �ꤋ�(��4�4$���~r�U��?����hO��TgH��$BB�|s��t�M=�H����?�q��W[���&j��V<B]��F[�gؑ�����'��%�1�t�~M�C	­�ҁ�1��&"aB�x���Od�d�O����>1b|�D�O��Ӳ�Ub Z-(�\�S�e�4qGl1�c�
Ig���I�Yz�g�'x�Mx��M�P���]B�ޅ,��x��Q�7�8ݠ�#D���1D�4��-���|B$���?I��<�6�p�ڙ;
X��aJ;Q>��h��d)�$���V��Z�@�lW9%�֔��g�'�$��ۅd���Bȴq�؄)�'�B6-�Oj�U����i��'���.��a�D�*�Tyf���K[�����A�� ��ȟ��v��7J�\*b�N�ո	u�"|5��%olx1yu΀zf�r�B�e*Q�,;U�]?oL�7�N�4hX;�h˔s����''�jqcE/E��D���Ӥb!Q�@:"�O:�$ �	�O� �p���U|���+ޛ��X�A�Oz�"~Γ_al:��[,Z"���Ǡ=����I���#|��I�7���d�L2$d�W��%c�Y���IO���ۇD��'HAn���qе��y(����aP�(@%�������՟V�T>�|�I�H���R!�/��* �^�e��
6M��{�E�cȉ�5��M��S��?���^�l�0����׵T@�#@-�,K��%����?��O�O��'\��k# �3g?�� Fݐ{T )p�'c�m��mO���k�K�(Ȣ���k����1R���r��w��R#��V�D�O��@�c<��O���O���;�?���u�y���A*�R�!r���l:��3䮞7Z������CܘX��`���S�v��y��&R8u�๹��� m�i�D��O�3u(��/x�� �џ�"=qF�Ƒ|�P���$7=���#�k?��
����4Y0�'��'��	1���r4AZ�*j�����	R^C��5p��C$],W`���'\��E Ey�����<A���I�F�^58v���pf�*Or���E�:���'?"�'w�P�s�'G��'sN0rg�Uñ�ٙj� у��O0�#���=�^-���<<O�
���-�������(rY��Ua�H�Z�zׄ �c�i#w�-<O^�z��'7��AfbԠ`�<�P� PҠ)mZ͟L�'���?�����C��p�EI҃a"��!�6?���ӏX��dAf�Y,7�ޅ	gđ�%gD�	��M�������'s@�oZޟ���s�Ti�Uz�Q
�/��iѠQ�c'�	u��00e�'��'f����Cx�Ju	� ]�n�T>=RV&;@�-ڏQ脁8ʓqRd�3� � s���W8Q6d�O?��d��	���u��^�\Y���$U�O>B�'5��!RE���=���#�!<Q�:O0�*�O���b�p�k��$�Ƞ3��'j�O��c,5��8�ڂ](h�z�=OҸ#�+�ΦE�	՟��O�6��'s��'nF=r�V%=2r�y0�[!~��g8}v�����[�#�����O��L��0xt�Ak0��#S�)R6�C��衒�˙N�Ԋ1�G0Z���'� �ffĵ`LU	G�.{�}�A�РhF��'��)��4�D:c��16@���m�@�˲S=!��W�@qg��	��p��ܭ�|@���?�(�|C����)�I#贫g���ɫX���$���P��֟��I��u��'��JN�&�օ+#��j$�܀���}�8�ʁ˚;�,�14%@*Y~�a�O� �<Q0JE�l��	[��Ɵm�A� )�ٞHi�׷>(f|�!�:�����u�Ja�r����x���6��j���� `Θ3n��̵�R�'v�'��'p�	*N:��P$��$<�iJ��@�E��C�	(f축��mR����%ś��}����?��'�"�v�y�`xՃ݃��X�M��w���˥m�Op���O4�Ǣj����O���M������tT*�(2��8XŸ4H�
S����e�ܑ�@]��)�Z��+Й0�6���`�6����˲W��u{�!�#hf���Η`qr��m7�T´Y�ɱ�M{DgƧa�j��(U��򨱇�P��?!���?A���?����?qM~r��F�{C��0O��Y��hO� �ȓG&x�
6 �ty3�D�\�8�~Q��'��ɍi����4�?�����I�PC�qpPG��ID䜀eӱ2��u`��O��D�OA"��\�V# ��SgÖ~0�I�t��H�5!~��ɁnI�	��L�?�(O�x��JQL�ً�oT |�����>x��kGǉ�;�5f�	�aF�����)"ߴ�?�.�H�4�
D���P7T�hԺ$f�O��"~Γi�@�y�ޒ&~d)� �(k*�����X)q��
-dp��f\%j:��͓Y,.���R�(��G��������'Rb���e�Mk����x��#�82�~�%�ԯF� �� 	Tp1n�|R���\�Y���#���f��Qz���D�*�`�I��έS�L̴Ҩ���}jd]�q�7v�b��S�Q�SN^lڷ�'AV7m�lyJ~��'���Z�B ��m9*e�5�A�!��ރ6��B&C��幢Ϗ������OX}r��(~=���� ��E��녦5�r�'���r�C�|���'HB�'��ם�D�I,=�VY�L�wW\p��ErP|�̙.K������,|t%)�#�?�Gz%��pB)R�K��|�wfˊH?�����R:l�|y���Ut��O���3g�O�:9#&�A���Ͼ�`����On���Od�̔O��	v�\�Yd��˷�\�6*Ъ�'A�|�  C�"ߦX�A�D��=�2�S��X�p����Mk�/۲�|1�EϸN`�pD
	�?I���?���|�`��?�O�AH�LJ!��mR!jP��L�%���1��ʦ���G+;��]I1�ՂdeQ�`QuAǽ"�Z���"�Q�rM���ҒEJ
hqv�)+�Ԃ��|+¹(�"ΌP�Q�����O����5`���DបC��Х-Q<4͂�D=�	U��y
� �����;1�V]p ㆜T���"O�db�,T�w�D��Bƨ�b�s�:O���'R�ɩ=�aٯO���|�`)��a�E�Ve�����Ѣ�v
�x��?q��~�ɣ!͂P�Ve�E���I*)����Z()�:@�P�1��)iS�I�*,r�B�19��Ā��(��h��!wzHg�w���`�K� ��;L���`��Or��9��4MZ�% A╌>g�8P��;f���	ǟ����5_�� �\�"�~��ժYu���ĈS�ɝ7��	��W(w�lqb89�@��:\�*�z�O��D�|*���?����?�&�ɀtgnLH�,Y�;�� :ƦŅg�\�1�`ˌc����N *H��y.�Pc>��A�4���Q���~�����=dxS@�L3)�����"rK������O��RGӟ9����J]4=7r�-p��Rg�O��m������O��I-
������#?�N��0��#[�C�	�N`�Ӥ�?I]2�sC��S��"<����D�F��MB�i�.B�8���l3"���O��S␦m����OP�D�OF����?	��4n���o�eO��10�� b����Vk*��Ygi(�s�*:,O<�����jX�p��D�\wJ1²��+m{U�u��}*��U�:<���I�2$)j�
�l�$y;R^*>N!���'�����4��?��?�.O������%0��r��A�f�`u"O�͉7�T�y�Y�&�'
���T�c�����<���0fr��\_`.-JЏH�9�
�QEB�7WZ�6�'�Bˬ[��'���lOl|�P�Px]"�`�	C
�Z�+�NR� �L&��@��(� &�V�=�w@I�"�Bt	PG�?�@�ZV��+%Q�lہ˃(7�,ER�
ԧC����B-�hO���0�'��6�Z%@�s��&�4�� 6+|�Am�l�`P�>�Ix���cG �, ��\���C䉶��I
�H�*�rP�ĭD�%�r�I�����<Ya`;7����'��[>I��m@^�C�N�3h��c��-�\!������	�W� �X�r;�Q��N��Xv"��Ol�2W�XA�nI�%��-5�t@��$���3vE�QТ��g��Z�Aä�A�
��N.g �iF-��.�9��ɜ�W�1O�=���'�07m�]��}�a<,���c��s=�����A>�^��������,&�4ⶭ�=�Z�Jc�&g��h�'���p� dmZ��0h���Sb�Eh@H��C�8���.9�M�+էX	R��?����b��#�?���?��h�Jdq�	^ X���:��
Ȋ<p����͛S�*�^b>�d�&K��hQ���,�$D�sNR�>�d�(��"jXɂLƍ�$�Xe%��xR�鑉	��`X�q�	�c���������*���'�����U�+r���+Ò_#Rౘ'0"�'?�M�f�)�l�g�	Sl�0��dR^�����'��9����y@b5��OV�ճR�'Q�
�x������'R��'�R��~���il,�2ȑ��ʕⓅ�$9�<����'����#���6ٓ�L�UF{���2-X��{ӨX�H��ؒ�#lqR(�b�%�b��&��.����hO���JU�.��W�Ā/>	���O|㲡�O<!lډ�M�gy��'C��X�]8�$>ܢXg!�`,BC�I�sNՠ�)�� Ҝpc�T��v���h�ħ<q��Z�=�Ƨ-83�Eb�lY� *�Z���p�'��'�q�O�?��=#���.
���ğ�H!:�#S�C�g�̀4�'OEW�'���0f�F���
�dx�Y[��װA�`��Uj�rHiӓu0a�	�h��:D�����A��1�S/�����	iy��'��O��Y6��C��,5���+��%vVC�I;� �d�o��Y��9��I�����<1�$��<��	�ؕO��P�s��:��YE��� ���O�?���'dbiZ�@��Q�RM���-� �O�-@ y���XE
�x�O2£<�gR	4A �H��͈h6�tAH|zǀ����+W;5�dѐ,�t�'ƔLs��?���tȝ�gjrAY��=E
�(a1kG��y��'r�}B�N�!�Ni�'�H�;�	r "�6�0>QҗxrA^����	��:���'#Ӏ�y��H�:��7��O���|�uF �?����?y4�-��3�]��]�!.O{�9Ђ�G2
К<h�͕�.���Y>�%?�;��̩M;^^X��@�!��sm����cȿpud �1,��%�z�|�*K�r�`Vn��_��ac� 	2��T/�՟ �ݴ,;��'�?�$λcS�P@E�A/tof b�N�.V��OJ���OF��Uo79c@ӑ+A%%�t��$�I��M;����j`�Ӕ)g���,�1S�^�ж�,<��I��Sk�GjM�I���Iɟ��^w��'a2L@�d�&T�\4k�ގ	���P!C�2#��KFIH;OW2y��)O����ɿ*����J�1Z��ʁB��-�@�H�n4z���6(M̐{�f�?�GzZC�$��ևQ��T��C�=i����y�����OX�O��d�Oh˓������/+��������h݆�S�? 8i���)�LAs�
�I�0�3mLi�'����'�	8��a�ڴJ_�uR���d��9��dO��Ld����?9���?� D��?q����4��8bZ�!�'�<�:����&L���Z�f��T�P����Q(F�c�L8��Y�o��|�7�2�D�����xbSB*|6����DI� P$�O��oڛc�&͑��Gp�8!p�����4�?�(O8�d0�)�� �vB�)�#İ�sdJC�<yB���"B��eK	qܽ�GA�<9�-��̕'Jn`H�{�y�����O�����n9kv�1�DH?-�R��^�m�b�')BN�$J��i���f��S�4b���0�n�$Ea�$I�Ղ�(OƉfd�7�.t��2�S�/� Ԋ�/^�����ŧmt�<��Fܟ��۴.�O����_�(�q�ԿA�Z=�3�W�R��s�����3�fz���;�<qwg/�O� &��҅WG����GM�����rl�,0���M���?�/���bqf�OX�$�O�!I��Ҋm�����đ�h/�|҃��#s䭠��J�X:��1�d����'���?ф�<(2��0TaU��^Y`�	M?�x�!�SS�=Q��0���'C�(*��P3�u�1L�=O=�1#4d��R�?���O��J�%׌\��W�dX��*.�C䉡e�ؐ`�	�7JJ
��ޖC�"<!��)
�	 ut��qFC1:�>pk3���?�W�@�+AkN��?a��?���8��.�O�N^*�Y8���:Ph��P E��<%��dx a��K8i���"ߟў��#��� )��JД;����б�?����+B�����GG)K���3ړ$Z�"kV�+X�9K�&
O ���Y�R �Ɏ�M�x2�'&bV�|z� �:��9
�"D�-82<�a�'D��y���
9�Z!4�6�yU �#�HO�ʧ��d�Y�j�d��oD��ӳH�t�s6M����$�O�D�OX�����O����O���� ،��E���E�I�P.)�S%G+&��]'&�R��x�
�+��8��됃+�^X��bݻV��"��h��;�Rqzڴ����!& 'L3<�O����'-�
A�s�t�i���#�Ő�rO��$�O�O���Fx�ֆ�[h,82�*�堂3O��=A���Фj�p؈G��7��=��h�
�
���˦y���l ڴS �y��iW��'T�w�Bx�A�\8F R$��.ʶg�0�� �0z��'�2j�4?�<�ˣ�Qc�|����sl]��$� ��=��j�{�'�9�_\��� "2�RW��2y3N����5#� �<)	 ۟0q�4��O���Nշ>%P%��/X��ȩ��'	�O?�I�;`|=��@�}>����G������p�ɗ*>8��7��  0Q��H�c޴��?�����<��M�p���0�P�a}�]0cK�r�<٢�3�e E뉛mV�;��c�<Qc��.�8h�`�	��^�<i��֮��*�W�Hň��Qo�<aB�E�)���K]�j9�Tc�<��/ζK���{�.\�;':�eb�<1'�S��y�' ��,��!"Dc�<�RG�򄛇o]�'c4�VnJ_�<�F�4nB\����=k/b�RkVq�<y�jK#*Qx����*DR��j�k�<�R̗�&���j#�-1Bh1�6�Yk�<�b'H;.�,�:��ǝj��t��!�e�<�!㎧hTR����L�}��GBF^�<�Ђ	ЬlV(��<�M0�.�q�<!%�(*P��Ţ��@���k�R�<A�*� S	��IC� *tƱkQ
PV�<�eL�:Y2A�;Y\a�l�P�<�JX92��(r��ĺ4�ވ `/OX�<a5a� 57�̓.^�y���p��]R�<I2dY�k��K��]�����x�<9�h��P�،�7�ŢV�r�Z�<Yĕ�9�����K�tl����/�<A���P3vג?B���y�<I'�eĀف��=/����]M�<��+W/~ ������"��)�MJ�<iĨə^q$���L���i�Z_�<�F'K�rvz!
�O7>T��VhN^�<ѡ�! �4Qj�-�q����hT]8���@��V�S�? Nm��bEv�V�kn&i�PB��Ė/�VE`�eE�fa�`�R� Y�)2��(�Ѩ��I�$�+�!^�)l�L�'rH�S�S\��|�I�i�Mc��"4���
�A��
�BZ�n�@%Iün���B-�O��[�����HL�Mn��`�M�4��'���b�[��,�gjYr ��F�'+��Gɚ�J��8x�H� X�Ȭ�'�*���	5�axb�P�{ �! �����`�tB�?4`LY��B��9H%����A΄5��O��s��Ld����@�H���pig;�B�i�'-"���ӅUМO"<��B����ؗ��8��PS�#ҳ8�1O�QQ0#ӱ<�4)����=):H���i�v�r{��q&��<�B�2�hwd�[�Ą
Bm4eP�ӧ�,Odp#���=ɘ�jSHD�7
�y"�ך@zvї�X�2�T�:#�_�c�z��o�0}I��hW@T�w��{N<1s�]X����C��k�t QpN�sg��'W��.Oj����_>rg ��jq��K��F�X�U�C�#�R$Qs
7
=yj$)�'�(�x� T0��O�nФ*f!�O#�d�!$S,�.~9�a��1,9�=�CY��-��ō�v������"5}��BND���	(����/n�� �72��rBGP	��=��B��Y���;�"'ғT1��%C��[��Ɗ"r U./�~���J�
r!|��e#]7�88��,FD~R�V�.�RprR!I�HTHQE&���O$�S'��+�J�B��օ7L��'�剫�f�B4	&�Ջ$��R'��q�xbd��k�P	ǉ	 R���Z4��8Ʀ)���0� 	�Pꔉ��/�,Рi�!���%�A8዗K�h@�b@	U�yW6".b���W2@� eΌ���>�O@��*E#^���%gӿ j}��D ��OR5�1�ϑ�6�i��')��⎔�
���^&�y�W(�5"ў&�j�)O�LW��'m�h��{�$Y�B�6�y�e^�v#���'Hl��ۜdmF���G2�%���$.j_���!c[,4�њr
g��|r*'h���mϏX���@�� ���I$���)4#L+Ƭ"9R�E��aI��" ðj�J���Q���Dvz���b��te3��I<u�^�Jش�TM��Ƒ�,����D�bV~��p!�4;93����ɥtS�T��W�
�����4|
��Ь��'VHqz�n*->�e���Y�BPP���p<��m Xf�'��2�	�BD-	Ȕwq(I	�?a�AՐ4��l97aQ0��4�� 6�ͦ�M�;o8v!I�/=���'��=|�v��<�#��<!v">���$e,�2�ܾtD� ц̩6���+�&т��D04�ʝ(r�]��MSfOb��I��%}BL�o� �*�`+,L�@�����-Dtc���{^: RQ �(ؘE�&�'S���g噯i2p�*T�VopD`$�XX���B(妅H���H�E@���O
�9��РS^�}l�77���y����CJ8�����yq��Ͻg���ѢWV�]�����'J����oFv�Q�l���i2��Hp�#��䝲%S�9r!�X��5޴U\��f	�g��1iu�X�X)�ş�{b 
��3��ky�ODJ=��<O�N��
ݬE�ˮ\@y*g�K���' <���\���T�b��H�'��`��Q�^�j)�	f[4�kA���$�ȈL��p��j��Jq�ՠq�X�����E	ZV�F A-Z'��(��O��~���2Z4 ם�y�`ſ���Ĥ�:-Q�*%{�Fݹ�'�Z��- �1�P�˟�[u��T �
'�ǛyGj$�jА�j�Oj%��O~��	D���9V�'�n�a7�X1ֈU�R�(qO�6��Q[�˘7�O�`��K�Z��:��wKd)��jуv��!iq��E7��P�i����V�p8XpN�Ae�b��6����A��D��#d'ROW��À�گuc��2���n̓5��0����"T�pmLh��3?)T��1x��;&"�7�a�F������#�rlBu��,<  �?���|�O\0c�fT3`n�Y<ոb,	q�1�`VCf�9��C�kF�G|�w�.�� �$������6�p������a�k\x4c�.7�zH��O(X��_�f�RDyӇ�?���Ӵ���E<��	ԄK�h�����k�O�ݯh�p �M���2�&��x�>�(D�W*Cx�">�����f�Z�����V�n:��e߮1�^�� ��ğ��b����~�"�%0f&�S��Fԩ�y2'��p�ni�&9=�<��g�R*�ب)�yb�B
V	ة+P�F��ѷ�yܓd�j�;#A��Yꊩs�@#;\��I��[y��'��PIb6O�I�k��"��|�����T�H�Qc6��pLH����tuP��&&��pÌ�X�'��6Ovts�M�C���`E���'�}3*���.N�aS�L���\�R	]���G|�`(��=J�j]+�h@t%���$�OJ�=)�V}�R����Qx������Ěc}`D��"Ľ��OX9�gO�1�Zw�w�L�s5�P�H9�����dR�a�Y��F{�OV��(E<6L�q1��?�f��$���f�0�H�F
6�1O0�J�V*v'����c�	jikB���KjpP�V����{s��Jj�'-r��)��Q��%)`q�Ԫ��wgn���>O佑�b�%$H`3!gfY����D�;9�f\�E�S�qb��=��y��h�2 'I�'b��z����M�eD�C�%+�LܵO���f�A�'ژY �h��tF�i��I�Y������%"	�hKcL+�	q�'D� I���;3C����D�IDz,��	�t1��qÓ��M �c��������>\�}�S��<��l+�� ��=�#j̴��	`��Ѣ�� �9�7t1��C�N_nT�����w�� ��*\���v�=��'p�q��,�,��<2���c��R���k��'?N��Д��C:ʐ�5Ι	�y�(њ$��U��a,m�v�H���
�KvFN5����2d��*����:����⬀4CP��d��\�LQ��!ٯh�
I1 -�8������z�\�#�rZ�k���;Y��f��p>A�O���GI�;Kq|�;�	�G�������?����I>gNe�����ov�A�'+	�p�fj�4o5�A��M`l�E{|D�2р|���Z�|\��;��҄p{l;���N����xr䇧c�$����64��U�f���'9��	��X�"M�m���(���r����,���2�+̼ _��+֌�P����![
�yBfܤ'e m�Ą�B~\R��J��LxV�^�LI)��7lO�`P��W�f�f���Η.R�<sC�	q�~Dn�V����J�'��äF1��[�i-2�v,Ɖ��E^�F��X�'4�ɱ�^�O@��!AL���2`�H�����Y�����$ %;�\�
4M�zd�݌X|����V>BZ$-�,N?O_x��'y�I�x�'?��,O�<م��	S���ҩQ:l�J����\'�� �s�`�b"�>!�:4H�E0��'_p�M��+����}���<1��{zt�۞'�AqΚ%�D��#O�\:�c�<)Z�D�;���3C�é3�f̑��>tn��Ӈ;��m~r2O�ԣ��W2, }�Bg�4&Ҷ4@d�K?����m�Ma&e[#��ա���p�Ȕ��%f��1E�S'k����M�lȪqb� <t����O��S��u�DT���x�&�3Om���ЈvN% �O�'�X(������d Y��Z`f}z0�uFky� ��'���9]���[�'����Bb?���� QB�3��4���M8>��S7����Gg�lC��x�.?%�ި���HW��ٖ@�A`��ac��$
 ��t��-� 5 nL?6&��B&��O��O�dg]�0:(\���ַ_^��B鐒	~��
���k�h|���U-�	�`oMN��ѫv�8�dO'a������x9j���ߨ��u�ē�^���mBWE��� S��<���U6�2ќ>y�O��m(a���r��d��{?A%��gMlei��
&�����h�lx�dk��*f<����`�RxAS&c�)SKK�7{�Xc�@�0p8�Ąɟ�r�����A
��Y�Q�4�%�M��Ѓ�l��p����4���maA1fCK�F���b�!A1:p�'cv4�i�=f�|r�ۦPV��B���N����gn�~���d�W�:q�7��2l�8ū���c&r���:�-���Cܟ��5n�17i�p�Or��i�I��˟9F��� pXQ�5:$�����/7���##��3;?4Y� ��#~ �p�-�-r�8�)O�����tw������/ I{��O�d��N��DlBqm�hqpQ�g�'���ڀ��" Q�ᠶ�İl�T���U�#!6i"e�@�z�����E
��	��ě%�*�`���i!c�~�|o���"�#��r��Ț[b�O0z᪉�u7�q���^٤ �u�io�50��(Br�b �կZ��3��Z�wh���Ugٜ]`Z���c	�Tx�ؿ}�y�K$�f�@���l!���7���E�TdF�J����z�f�`7�\�,�
�)T�C}�O��e�􁟙mv*�#�_j1�(���(F����
��ce��z���Q3Mͦ(h (���� v����u��Tl��R��S�c`��'t�����o�P�Ѷ�H�1�tE� �y�Z`p�/,O��T	$or��0���?}ZV����1��M��54���A?���Y/M�����e� P�y�b㙯x<�Ԑ �ʽz�F	�'7@Y��K)j���ʤC��K���K<��A�>Et4�k�y+A� ��ӥ�ˑJ�v�c�ߩ�����E�3d�.��� �
]h��wJz�8A���)Q�ԍ�Y�'�@��Q���k��u�!I�!(�R��a��Z�
@�9�<��I8eaH�S��NW;��ePOX�N�>I���4ht��$�/�O�I�ƌ͚�J(K�.��q��C�4M�X�H"���$���?B$�>QH�a����$�%O���1��? 4e�B@ϔ�a{b	��,���	H�Li���{���`���=Du�T�D��O����Wv�|�BV�O>k���qx�c���$� U�@�O��QD�Y��%�7ꚡB�>�a�� �O*F�N�r�dT@�$ϘF� ��f����л�-��RH*�DN/<�S�MTɟ�yU%��B��U����uXD���%$���u;�gS�:�:d�B���w�����AI�c�6t��SnD{�gP�zYt8�k+}�Ƨ~�$i� m�����͇<z�0� e���ТB*�O���G�2!�$��TL�8��B�,��x8�)�O:�)?�<���t-���X��� R�X���'�\�D����X�]�
��90��M�Gl���R"*�b����-Ob���c�#9X�x�JD!jm $���O#wD!G���e >y�0�W�^&�:��1u�a ���t��'x�x'n� k�u��D�8� B�Oވ� ��]�L�`�	�ߠ֨O�ܣ���E)���ќ$����Z<^AX�j�̋DHB��p<��j�l����!.�#����&Z�:+ց�"<�O9H#)^"���J��/��(�m��tR��!�'r�)�5�L@�ۃ-;<�q�!A�w�}�%�'�h�2IH4@��(��h��a����5C�(�FzB� j���Th0��b劁���WkU�iX�a�X�n�"�ى1a|r�1^HN������� y��cQ'����fF�P�XH�
�Ds�X�k�f��M��eax���*r���[7h���hKG��O`�*���dFp�f�97Q*��՞����I�5�5NC�YҨ���@������S[RHG���)�8�c>��9�-��4�HؘV��&���!�$>�|�;?R��U���Xdl�է����N���`� ��҄K��&Xj\A�0�Mo��\@�'��S�&]�4��i�'�UipdG2J&������H
�=f	��hT2Nd�5��g��|5���PX�tj��M�v0���G._��$G>@Ɔ��
ϔM�$��AhO(!2Q��&+W F���ߴi$��E`_H���<"*�]S5��D(����a��yb�ے�d�j�%R�Z�!��פ�y��F�b%�F'�%�:��oҬ�y���:���F�X&F��5�b�T<�y�-�>�$���+r�Ԡ�d���y"k7cx�+�lez��	�y�&N�4/��1#��t�>0:F��'�y�	N c�,i��)��R��1�N�ybB�kXnm��IG�*���3��*�y�cW�{�,{IW�v)B耐�yB!�:+����E#2T��!Ɯ�y��3�J=C�N�-_�z"el��yb�L
F h��.�#VW^:c-B�y�.C��(�K�4\d��s�R
�y2M�z�\��i@1?a��pO�
�yBFR)�[�,�5b&��o\�y§�#T¢�;�	 \�J��b��"�y��fZ�a&Ĝ�A��¢���y��8e |(IƬ̾9���3rJ��y�
��I�^%n�B���pd	e�!�d�3xHm�jL�=���6{HC�I�rGЭ d	Q�~�f�����3fNC�Ɏ]�Q�g�}�2YspaΥ=O�C䉘%����'^�o��Z�.�xU�C�1)��"a��#��Ѐ/T?�C�I�5���q�r�|XR�FD6i>B�	�r̮ȸ���?B�0K1�EwC�I���m��@�'P�(���(E�R
0B�� !�4��T���i�c�.n�C䉽 zL3c�ۇt��H�Ø*@˲C�wÚݹ@�SQ� °.�VF�C�	�7�,�@���A-�P���>$]�C��+Y>�����ѼS2��G͛�� B�	�\� [��7�<UӖ녜#t"B�I?\�q)3�A�P�<MS��ևx��C�I>D]d� T�i��403��Nf�C�
��+�I�UHY=]��C�I.��x�2�\Ҥk��(�C�I��8�h`iД5ȷf*xt�C�	+����F�J�����A@B�I�l#����\&XhHtX�h�6 �bB�	�'�2|Q����$Ġ��LV�B�	�;���`)�� ���D}B�I�9�p�IY>Jad��Z�P]B�I.������O$�3�eب{�B�I�z�m���D
�P��TP�.C�	�r�X�R��)��q�R)�EOC�I�l@> AB�6!��I��U�8��B�	1}�B%�h�P��HͧTX�C�	�ON}PQ&+K���`���-��C�ɤ_�B�{�i_������
ӼB�I�l�|�%Ƈ�r͖=�d!��B䉹8BH�0�EB<���*%+�<N&C�I4(�XH�����ڂc�T�BB�I7&?ґX��0��i� ��68�C�)�  1"�B[ O� h�MyT��"O���0�Z]R'	ќ\^�	�E"O�D+�FT�L��+�HȖN_fP
�"O(����=U�|9�0G�md�p�B"O���g^*��r%�Bv��W"O�-�W�?+ֆ��3+*=�|陖"OʩKV����3���?N~jX�S"O�1�GƓD ��S׎��`S�U�a"Od�r�����p�$W�L��q"ORM��H�>�"Uc�%ʬ�hT8r"O��7�5��q ʴkL���"O�xH4�.]E�j����4]R�"O\�T��U|F��,�`E�5R�`���	FRͦ��U���` �L_�Ps�$�S�Omd�g�ؔ(�DXڕ�� °��'J�\b��[/=�a�BGP�x�05��O�����Uڲ�k��ץe�@�rd�a~�T���gU�&O��yq.�/!T�y�F)D����c�2�E;0�, T�l��4D��S��(=���t�]�0b	 !" D�s�Q�:x��2��^ V�;Ө<��p<!�Z�"�R� e�-#��ĩ�P^؟���zM�giA7���r�G
~# (�ȓ��|8���Z�A^�Yu ��ȓ5�v�:�/��;���Yb�	�7tT�ȓ���u%�u�$�wg�$��0��k�����N��n�q�lP�SM�!�ȓ|������d]Qe��L�еAqG8D�|��e��Sl)��$\:h��7j6|Oc�\Sg�J:j_�8�瀙�}f"EҤ 8D����CJeu�eȄ��3avg8D�\2�!�.F��@��U�Q�հ��4D���"�����#�B�k��n3��A�����n6Pa�,ϡEI )br�ηQ�FC�	�9)a�@B_�OE�pxG��U���I_؟D��k_�i�d�$��*�����=��ˈ��Er��O"�������N1�"O4��G�8$N�Kd
�(r���8&"O���g6*R�x���11���S�"O�UP��'�dX�R�	�1"O�X��v�\"���	"b@�"O,� C�8yj(ؤ��rYʧ"O
5i���<5vV%B�ɡ|"����i�ў"~nځEJ�#r/��e�Lw-B]g�B䉞;Pt�{�E��mhFy:g�LvB��=̂�i��A�"�:��ý �2B�	.0��H�6	sH���]%D� ��$*�$�N���	RE\$>c�q�U�N�!�� ]���gO��7k�-���	�5�!��<
�&�@�AAz$�렬P�&�!�D?%���ë(_y#���*�!�Ğ1�J�ؖ�XF�xɧ�N�;�!�D��?�
�#�� ~�Xagǳl!�$�o��8H��Mg&�E�2�ޯ	��DK*�TT�ӥ�>zI��ZE��
��O|"�R��9|Z�����0.L�	X HB���hO�w����c]/"��Ya�:9df��ȓ+D���%�g�A��ۊq?�ԇȓ}�����ڇ~�����N�aOP�'�@���D%�ɺ(|�Qsq
� "�� W�� 8�C��!t|�jr/��a��wJζ VC�	��5�vEG2"������T�C�ɳ]JĥE���	zX��	.D�B�I�u������(lW&�*����Tbz"?Y��� 8�R(�9/:�\�		8a,(�`"O�]aF�M�w�JL�uHH�Y�S�"Oj�x3/Hl�)��ge0��Q�"O���C��Fȁ��&�6h����"OZ}�q�0�̊�C��G��Ғ"O��[c�F:s��C#K��L�"O�E�a���Z�>���[60�49�Z�('�(zçF�<u���*�и!㥓�N.2��ȓ[�4�TF�q�a¬U?\*t!o�M�'��>�I	��K�" <�x#�;B䉃'�p�2�Vyx���ܩ'���'�ў��>�0��>%�օ `��z� ��KQ�<AA�+;�5��^�
6ݺ�+�N�<�g�����IBa4���r@�ZL�<��4"�\�HpB �w{Rp!VJ�<��
����Xr��%�r)��^�<QB
U�1<ZI�AψCˢ�C��П��Qߖ	٥��I���M5kt��ȓO��T�a�E=r�J�;�f)l�������Y�-�8*�ʂ#|{��=����c�aK�
O����t̊<��hJ�a��*5<��Q���6<��؇�<9@�f��"cR����Q4>�r�ȓ)�j<;D�� b-�N�U<n0���?���e�X{惞�A-)�ҀW�<)��N>\�|�����'�<�v��w�<�tb�
8�kF��8Rs�����q�<i3eS0�Ac!Ϳ,l�m���p�<�TN�n���Mк8�-���i�<��&ߵ��c���=���c䌕Y�'��xRc��7'$��э��r~��ʔ�ӳ�y�܁?��Y�.Jq����0F��yM
����QT�Hhg$��y�"�+PR�b�nH�F���F���yR�E�OBT!H��R�seFDfKF��y�×�E��ڥ�޽&|�����y���Y�U�>@�JȐuH��y�����A�Tj�r���H�y�D���ݫ�-Ya�z�PPb� �y�g��[�,<�U��FDX�'A��p<ɋ��0h.01��B֎aޤ���Z9!�$4Z�|"
���P���Ȯ�qOl�=%?][sV
gҶ�{DK�R9+�H+D���� D����tR���.D���ǁ��t/l�#5c�#AQ.�ӣn?�O2�{P����wZ�ke
��\���3rɤN��x��8�5���&5���ȓv�R�[�'J��BI�?��,���pu��Z�_���@�ucN���}��p
G�Z����g]�CPR��ȓ'x���gϖ�f��AdP	?$�`Dx�'�� bɐM��� g�R^�]��'�N	EM�\�
Q(֤:{T,`�'?�D�t��#%T�Yە��.���+�'X<a�Eݼ�KPM�|�\}*�'d�K҃�DFl
o�Fc8�'x���* ��a0�M�-�Ա�'7�;�e1O�dA �L$+�!�'��)�Q
��&�!�u�ւNč��'���	U%��}������P@����'�@dbT�Ix�L��S�@�K��	�'�����F�^(��+u�`C�'5�0A �2��Y�H�f�)�'�D�$AR�=���� 5��|�	��� ʌY��ĉ,L����	^B�C�"O~ ��NUc�,@��F� B"O����$,ˢ��"�\�X^6%3��'>ў"~�Q�
*S)��H�Ϸl%0i�����yҎO�%Q.�����T�S�O�y�Α#�b�k�fE={�l�!�HI��y"��p���Ƶ(<f]�%��y��K���Ate-"@!���*�yҪ 2P<f�x�j��Fʸ@�G%�y�엥x?�u����	���1W���y2" o�h(�	�V��ɺ����y����/�@���,��H]���r#��yb	6O�\B3���;M@���	�ybCܝw�hh��/�k�+ޱ�y�݈(���)�͗���A��Ǆ�y��Ja���;�)�;����kB��yb�F�S ���b
/c%���덊�y��^Oj1�B�Vdn��'�y�/Q"d���n��e	�j�\���'�#���d5�ӯ]��|��'_��Qs��	�m�� ]!eCD��'�!���$Y������]��ik�'֬��F�$�\�(��S!f1��'"hyS�&�Lu�5�ː�H&t�p�'��eU��KB���GZA��:�'U|��n�g�ʐ2�$ԚK�'�e;���3/�@��ć����'+X�36I���<:��9vjd�
�'Bm�D�=cE�<���t����'�T2��`�M;� �jlRi��'��&��	�kĦrk- �'�h��d&��k�!�"��s��͢�'nTA@%��+^��Q ɏ�r��x��'>�:�_�-�a�(s�Z<�
�'��ᢆXlI^��KB.=���R
�'�P3CD{�F�Q���4�	�'kbR��kC����?@�X�		�'�xS�۬0nH0�h 59O����'�� DW1��yc��f4Hs�'�<�����E��p����e:����'ׂ�Ȅ	�!p�)Ua~f���'IJ����:��-3TGFӀ�p�';):v��|bH��A�6O(LI	�'"L*�����,_�wM�8��'�8�M-(������hp�q3�'U�l���	�t(J�mҝWR�y�'����G�w�ZU�p�֍�H�y�'��,m_3��z ƍ4�Y��'�h�A��C%5��"�Ɨ.1�mh�'�jM暭��؛��Y�!%����'���!F����k�O� ��%�
�'���!am�GN�����!�*�'��P%`|���ba�L"��X��'��	��iX�D����ˠ_��"�'PtbP)�+Op���L��P%f��'ۮ|��琑:�ҩB���1ؘ|!�'���)ЬRp��ǂ"	�%S	�'� ��ʴ���	E|�s�'�$1�c$�79�&�C���}1B�c�'4޴c�ĺo� �"��t��4)�'��a��G��MUP|1��eG��!�'�X1���S�(��I���bƒ�!�'7*L��$S����$.M�$�j
�'�By��狗A��񥣝6Y�6*��� (�i�/I��l���9i=���G"O�S$UԦ�����n��P��"O�8��Щk�" Cs���K�)+2"O:�2V��`�%���h��1�r"O��@���o6��C��L[��ȕ"O�E{!�V#a6�*���8QE�D��"O�bd@Bi��H	���$6Z���"OXŀ�'�,�z9;�`�:����&"O<���(u�f��U�F���! "O�ã��-G�L�c�Ɏ	��q�"O
�F+�s���3�S�2nJm*1"OH�'9v�<M�u�ʀL�С�"O��d��w��]b�T�0���"O��`@W�o�Z׫ղ����C"O&�r7'��)<���ʖ:Cz�	�"O`�x�Fy��Q:�d��O�r�a�"O�Yk%�_"#��퓑�:�L%��"O�5�ak*,��#	�6�
���"O����*�t|�=P�c|���V"O�1)$� he ���~���"Ot�� �dѾly�!V�9t���r"O��zSiA/+X�x��ʖsX��B"ON�����F�	zao�%V�p"OZak�B^Z~�Mk���&�ZA6"O�X��B��5��e�T-K�ݨ}�"O � 7�J#V��|�gl82���$"O|�F-�M������ri"OT,3��� F��ؐ!�ɇ�N���"O�|(��ǝK՚9 ��U�]�vw"O�-�B�^����J�`�A���"Ot�gJ�43X���lŲ+�<1B"O܈C���@N�;�
5oJ����"O�((�c�>_:����*&V4�p�"O�(�t�ϒx�L�ceyH\� �"O����M1�Ph�o���ؑQ"Ota����Sl�A�o�X���"O$�2'eE�	/F��1M W��1HV"O���Ë�d�:�mI�=/��	�"Ot����&e���K�,�W8B���"O�a�!��$(pZ1)M�42�	"O|s &��B��H'������"O��:f.ӡ?�*�"�Ⱥ�nѠ"O^�6��}[�x�A`�aՀ(�P"O|R�͚�^v��6�
�3��,c"O�H�r�O�2l����]Ŋ$�$"O����-�wft��aP�SL��С"O`�Tm����Ļ85������@�<iQ&�1e}*]iG�%���FU�<�����������*Vd��q1b�O�<�chW9��;�T&C��Q ��H�<q�HmB6�ف$�7
���hP�<��^>���YA1_�H�� �W�<9ph��othiӑG���� FL�R�<���Gr#vx��?�@0� X�<a�g�7Z%v�1D��L����,�U�<a󉆅@d�g#���f�Q�<9��P�&lʔg�#�.�X�fEQ�<�n�4\)���;enN�:�LUI�<yr�Ǻ%#��1.5W%L�RQ�Gn�<��H$>����@�w����g�<��h��M���%�z����
e�<Q�I��y��1�-f�peN�d�<�Q��"c�m�wHF�/����]�<�v�F���)Vi!	٤)CnY�<� �A;P�8iF�E�$�R-�9"O�9Z��v��4
��T�MV�i"O�@P�$\�O(F�!w��!S0@!Y"O:�3&�W&)v�W�-iE���"O.��b�U�v)���AT�r*�59�"O>Ȑ�`З)�@A%�E&I4��"O�qt+��F :���n�l:<b`"O�M�J�u}��"�,��0�p�[�"ON�� ��` .]+A�C3S�Nh�"O��i�k�Ld�I�O	�p��]q�"O�	IN79�xIw��:~u* S'"O�9:�j� y�����1znp�"Oa�՛+Axs�'[�AY^�E"O^��Â�3"��<9Vm]�=�l�h�<�GΌ;e�܄���"�$`
��W�<�&��<WQD B�˒J�~-�BmL^�<��O��2�F�7ў(`u�-D�)Vh7.��Hi&J�,��#)D��e�ʞT�$��fSN�̠`(D�D:�+ ���}�$�Rw����#�&D��k1N0|�	3	�AM�u0Rk$D��B��!p�ҭcj۳��Y�"D�lB���k`@5�2�ڂ.{�Q���"D�@s A0}�j@ja!s3�1�B�?D�L�&�K�y�5�b��U�)!�!�DU����!��$Q,�/�!��{c���AI�+62�"���;�!�� ra�,�6RM���
�-�!��D���G�'n.��`���JK!�Ĝ�f��J4i@�	3��ۧK��I�!��-L�$����6~t)�Uj24�!��֨e�eHMpc,#�XW�!��
�c���G�U53Nd|1���=�!�D�4�Ѱ�P��`!A@Zh�!�d��{� ��^)|���[��
0j�!��A�E*����Q�P�9��S>�!�$U5w"2�IcN?<$���TRX!�$V.!�x��D�[o`�Uʞ[3!�˥'eX�Z�Ɯw�D���	@T�!���S~�q@c�.�L�� ��*�!��
���IZ5�C�p�ݘ"��b�!��
p<`l肀�	c4���h���!�d߶*���J���q/��Qcf.o�!�D��N�t���O�]��dJ�5�!�$��Zu�s.Ј5�d�`�/��!��K�:��u��dV4hٔdp�
�%{!�Z@��t�v"Դs��H	a��/p!��QEM�`��l��=�E�1�!�$@+n�|Lj��(r����@�L�s�!�.s"�2e��aP���b	!�d߰=vt}1����hy#%��	�!��ߟ�N�X"��J�r���-�8�!����"IF�/%�Qm"<!�䏌:'<-��4�48!�L�;!�d�!�	˓��1GfF)i��өK0!�$Q�!�L�q���`@]'{%!�9>�n��qρ�R�B��eN�<mE!�䀽~6��d�LV�V�
�!�!��@c�\{���C�v�y!��!�"!aZ�Ia\�X��Ӯ��!���!~�~ha���F��B��	9M�!�$X9��)�F�� ~�I;�o\+fr!��BJz`��bP>iΌ��M
d!�K%�XV,�<^�1s&�\�[P!�� ���sEۗ,'��˶�Q�'���"O�q�p��w��Y3cR�^a�R#"O0����B���@*%�T�d�,a&"O��K7R�.-��)7�z��0"O�F��gK"d�DΙ�C����5"O�(+�+�>\=��	ЌN&%�*}0"OPm8��E������+Ƨs�<+�"O��Z6��/3��xA��p�V���"ODt#��K�.���A��Ʈ��`�"O���b�� g�Xj@ˈ�i�PH��"O�Y��
�0jz�rH�����*"Oʝ��LI|�
�� �",�� ��"O��qĘ<8:P�[QM.*rT�a"On݃G�K1]GH	LΑl���`"O6�r0��m�@����B�"Oh`��DQ��};���a{R ��"O\��(��_�$� e��F�AD"O�᫱/�8<�5�(�"O�i�TmE��@Yd�kf��w"O\zǐ$|Z�£S}s�0z�"Oj �\�c�Upv^/t^x�e"O%zV$:&m�E.B���E"Oq�c'=NW��p��Ӥ �"O,��gJ��J�4"A�I����V Zj�<��cU�J�Y�fK��vD�EIb�<i�F��� Q�&��[��b�̎R�<�C�(���\�\k�A��L�<��	0�XIQ��g���`���@�<���_1G�.t8� Q�l���a��y�<Y �#x���XA� $�]H�%�s�<15�H06Q� ��炓*}�]⇌ x�<Q���4#ԂV)Eg��U��)�s�<y',ؑ7*��@&D��dD�Km�<ᡯ��U���c@E��m�YRn�d�<9b�ٜ)��8JD	�*`��Y�$Cj�<���V*i�ycg��?���2�Kd�<"�Z�kIR���D�7�n	ôOI�<q��A��$�HU��-^M�,�a�Qi�<��Fσj�x��
�-�� ��`V]�<��d�,E��a���)N&�\ B<T�4�E%	FD�������a��q���?D��rV�Ȍ-Vδ���@;'Zй8B&*D����K ��h�K���i�U�vf=D���V"H�|(|�;uHP�X�n=�U;D���r���/#�(���A`0vɉ��=D� ��G�6T����e�AE�@u24&:D���K��l؂��;�� 7D����(X�P���� ظA��d
F�6D���gH�la ��S���j�ry9� D��c���~Wr�i�_�	!H�RdJ#D���@n��`Q��G8ɪtG D���N��Z�0�b���3�v��?D�0���L�8 ��냦U)਀J5�'D�� ul�)_�&�@D)�uZ��`A%D�T�r���fxSbT�=9�E�L!D�� � D�1��lctoӍM�r��"D��"dC�L���6�\��2+"D�$sr�ܓVJ( 8���0Y*�E:D�d	r���K!��ZP)ʉŬ�s3G7D��X2&�Oe����[�@s�Ea!�3D��B�>�>Y�př&vd�q��j7D��P�B�i9&$�T@�L6��K�F4D�����в���1���$X�<����<D�(��$T�AU�%�1 ˩oL�XR�:D�� ��W��[���:�nx�"O���զ�Od*����<��ˇ"OH�8�疬D��Av��2��͡V"O<�
6�Q+pt�۱m�-����"Oܠ��V�����+C�h���)5"O�Q�q�O
WX	��*2T A"O�}dЉa�
�Uc��(JD���"O�q�ة2?Б���H( J� ��"O�!�v, o�ʸ��:uF-�a"O2�3����������|���"O�d`dA��hh y��H"_����"O̴�c�T �C�^��"O
���\6G�\sJٛX
y��"O���7%�%b,e[�'�OH��"O�P1��Ρ5R�c��2���'"Or,2�嘊ZpMs���c�20�5"O�1kqC<GI�4z��1̕2�R�<!C�ތpS�ā����n=qա�i�<���x�h�" K�-m�9���c�<����~�*���-��,�R؈#I^�<�#L�u��|����e��,2�R�<��A�duV����V!u���9C�R�<Q�l��YF�}��Y���O�<)�LA�
�2T`V)�Tl���a >����[�
�S#jߖU N��r�����B$$��e�<n����ȓBHA�LQ0y�1��
O�|�݅��O��R�p�t(�aG�C䉑����P�,^Dm����C䉚K�pţ�dܾA>5�d�}��C�I0W��t�aJQ�Q�ݺf�~�C�I�gF���AH�%T�d
b&B%�nC�	��V`����5r]�8z�*�H�B��P|�0�c�"�*��F[
}0�C� @�M��'��+XI[�e��X�C�	�p��\�!�4J�dP��JW/�!��ѡB�D�s�o[�gaD����'�!�D�aƎ%H�gڐ������]�5�!��"<bf9�G��/#��XӰ�r�%"O���Z>�0=�h]�Fݚ"OZ��ǥKr�R2�D�'<��G"O�](�o�D��ֽH8 `�V"O���rΒ�"�P� ���	�ą� "O�,�����Zm�ȂDo��w.� &"O�R"V.6���NG���	i"O�ah�fE.Ь�Q�@7����r"O�8�S�B��;c��Qq���"Oq@�)�:8�ѱ�d��=�Ԭ�"O>�X�B��9����	1��e�"O6	#i,c�]a��/q��=�"O�lCQa�1
xZ�4AJ���)�P"O4�!�G�6�����"�*�&8�`"O�Q�;CMܵ��@T2a�d�1�"O��)�L�=��c5���0��Y�B"O<*�)Ib���	pI��! "O����&��}!��%W��A�"O̤�S�9-���v�1@xl�h�"O^l+7l�. L�k��ʝ*C��ð"Ol���:t���0T3��C"OrQ���
�,pE�I�j"]IU"OrY�G���{J �˜�
dZ�"O"-"���v4�)s P�a�Ix"O�%��|�.�j���h4��"O���v"�7@��X�B�P'�� ��"O� d�06j׫> ,��V�ʎ��Ċ@"OV�jOL.e/�	zFmܢK�`��"O��Ĭ�8^�u�b����`��"O~� n�j
ړ$F0�ƴ��"O��c�g����Q*��.�P�"OX%���Е	�p�b6����es"OZQ�B�܀#/b�+r�r�
�c@%D�Ё����ڤ*�����`�G8D�����1���+�bF���G*!D��k���<�C��<*���:�b,D��[�bӳA����BL�64ZyF�<D�D2U�^W�M��J�!�>�)R�9D��s�3J~��х�5)	k�<D����ح^�Y����!|4�, ��?D�$��:w78Չ�lLP~`@�>D����J^'��[�g_�>kF���8D��q!ń^`���m(f <l1d6D�b���c3�M��d����4D���P@C�|�.�{�E[�v���I�4D��I7h$�F�ٓ`�Y-ԉ:"�2D���u!οP�r�8'!�6S�}�1G2D�Ȱ ��%d�lyJV�h ��5H.D����
 ��:H�R0��b/D�@"�6��=1o�8a�J�:U�'D�h��ؚNSP`�poPJ�JC�*D����ѳnGR,�tɞ&��m��&D�����աcܬ�a*R�!*�b�$D���J�o��-tX�� M�^�DB�I2O����QL�3��Dx��ʼH(B�	�R�|���?33�,��i	7t�B�I+mS`���ʤ'r@;�!�\�C�	��	�c
�-f�\����˔7*zB��l�l9S���r��Ƞ��$<�JB�	:Q2�"�$E��Ę�B�9)bC�I�t�p�p7ϛ{#���`-�0;��B�	#VLYx��N��2�bmίA��B�I�2��|�u@J7W���;W&���B�-dN�j�"�>N�zY�ƥ#O��C�IE��׮�2%���q�Ě�-��C��88FU�Dʴ'#��a�1C2C�I�Tl9bj_&8�����5E�fC�}O��9!N��b
]Z��N��jB�I�Yؔ�f�0 j5F��uHB�	+Z�D�5aHd�u(��m�jB�I�gd�����"���z�a�XlC�ɉ?^d�W2d�|!�́�znC��pƔp����0g\ݓ�j��J��B�;&��+[.�@���O����B�I�G���Q��M���!�
B�	�8-l�k����IЪ����@ �B��(���Q�r�]�6�S�)_�C�	�q���;p�h�A�!BN<A��B�I�>�p$��K+dאY�D	���B�I����UA�,I��z��͂~�B�i���7�t����T� %�ax��&D�9�#�dX���"Ӣ)�.a� $!D�d��1.o|́$�P�d��ɺ"`=D� SP(S*�L�06Ǝz���;c�5D���d���P�PD�vfͣ�����-?D����������p$��H��M�:D�L�E��p���e��/�b����7D����f��z����ߘ*��T�f
7D�|�1		�C<����x��&7D�x[��!>��a Ĝ�G�h��¬5D�� (��f��.i�鐖kU (4�B"O�({C��-Y�`]	��$u/�س"OX�g	!�\��A�B$/Z��%"O�,�+�#f4�i��ӊv�����"OJa�Q��Q����G.ʃ(��A"Of�܄6\����ߤR�B�	�"O��a�7t�(��50E�A��"O(G�6�(��J�l��f"O�@;po[1���$͞L��D "O	H�N� E<�3A��U �"OD�9E���A ᙷu���0g"O�%�V��.�F�!��?��"OȜ"��͔>y���R�@�q�Q;�"O`* �D�T̚vh$Ef1��"Ob}3��V�,����!)B��M!�"O�	���=!�8]�"#��H�"Ox��Rg�����⇘G�l��"O��&��i׾���0j���"O��b���\�����Ę`\6�;"O ���/]-:���=NU�P"OH�OƲ9n�R���L,b<k"O�(���-���u��+?���a"Otuk�䃺J� ��T��6��"O���F�v�@V��\��r"O�xEAU����F�&���z�"O�]�Qa�9
���`G�6lR�X�"O����c�R�1so��Q�8"O��0�#�'
A��w� 3�Ԣ�"O<`���y*�6�+
�XT�'"OL�Ycٶk�^�!�-Bx H��"O2�A�GZ'"�|�0h����� �"O�͙M7E�c�	s.@��j,D���.B="�@�!#K�"��+D����I����5Mʠ%�LE�a.,D��Z���W��d�p킅~=��0�*D��B��^���:�$�OYHH1M#D�T�I�u(����S6 L+�!D�!0ł[Zd0Scٙ�	�E?D��;�GV+��]���V9NTЍH��<D�h�QF2C΀�[#h�/T�ع�5K(D�\��'���H���_�ohLq*
�'�4X;c�~V�,8�b�>uf#
�'n���54h���3��	�'�@H�s V�w=�A��[�0���b�'�����Pq�����;.��K�'�ri���U�k��$�S.#��'�f�B�*-�TI���,%V,��	�'LPD�F�#w�x�@��N'��	�'�($KS�~ ��4@����'��C,�Qf���CE��P)��'7�0����!`")�s�L&�����'(.���F�2	�$qd���ve��Q�'�j�y��i��`�C�Q7q�,���'�$	�ǌ;?H��"�I/�<J�'�P�1�� =���Jn޳	�
�b�'�̄��қ>��u/RJj*�#�'B�h
���%{Ќ50���C�Xl��'Ld%ie�Ja*]��f�8�����'���P���2C��� [h"m��'ˆЊV�A�3��@���ԥN�����'A@!ku���ݳS�ԧq ���'�N)S��E}�$�p��	h����'�� �4�JD:C A)E�@A6�+D�H��%�c��q� B�UY��;�*D�� �U��!�	^�� �/�`��B"O�%��C�X,dA2儋��0h�4*O��J�k����鱂W �\tX�'}���A�v��I�� �4��tH�'6�lq"�^�H�䬞&0Ȱ\q�'��b(B�z��P�PYl`x�'����%Yd=@-�j��]=R�	�'2����A�k��YecA�O�����'܀Qrw���jw($ӳ��&B��D�	�'j��9�e� p`��k	�5!�p	�'���#o]$7)y�R���-����'�
�) +�(9��ª]�A9
�'`��π`���0���]&:UI	�'�乵ғ 	�eA1	ʩ\ԤHx�'�h�[g�B,?��q+��Z�z(H�'Q�Z��\;1X�C�$��	�'ƨLh��_��1�F�	�F@2�',�\��WRjE��+j$�<��'�A@D��Dl�qa�O4i#e��'��q�f�'i������d����'i�ݱ��Rv)Z,��3�ai�'�V�KbE�#���#0N l		�'贀���H/0�3i(-�@���'D��0)µb̔�!�]�J�EJ�'�P1�e��{��qR�P0H�#�'��Iz��ͽQ��\�m�)0�,y	�'R4�1BTg��Y���"u�=��'���K�`@�~ؤ�����@'d	�'v,j6�J�**�����C`�=�
�'��� ��N8-��c��Cnn���'�9P��:U���A8�����'DvI�d�dBY�D|G�d�	�'I� I�S�2�A�K7F��$�
�'+~�{�ʂb�pyf/��q�Z��	�'��8T!Q�*Q��:6��=h�$�	�'�L�r%c�w�ȅ�`�G�a����'i�pR�U�v�\	��W��3�'���1D
Wtu#�F[9U&��
�'��Я� ?�<;r�$H�ق
�'S�]���4�qA!�W�=�x�
�'��f�Yi��·eS�dr�B�'c��H	�(4�#ݍ���D�<��?W�x*��q6�4J*YH�<�q�N�Q*���ǃK�^��d��/�B�<)�<p:t
�A�b<d#��@�<�Ċ�8�`4��@ף�����s�<1�Μr,4Š!��#)�h�<�CP�Qg�h�%F�.��T��"�x�<)��[���%NI�D��h�L u�<)��0Q>䀸p-�]K,�`CEo�<I�k�z�y����0ӆKl�<1���V�\*�ϐ�R0q�
j�<��n�y�N�$!Z	9�x� �g�<����D<�����EDTe�1�\Z�<9֦��K��њ���wb65�gEn�<%�#@,����d�U�<�E)���T�Г����!D�]F�<����7i�M(0��-��={w�[g�<�ӋSog��FJD�r��)K�N�l�<�W��2�>�s���p+�1#�}�<�R�9|��c0$
Kk�L�cʝa�<�ACN�(4`�� g�̹��#�Z�<	FDA�c��q��D�+l�-�0�~�<���B� �\p�c��:K����B�<� HL���ϔ.}��`���݈�"O�\�1�м��diǞ���! "OV��#b]�9����|��Y�"Ov���Q�gw���tN�*Eht�8S"O�eJ���T�~D���Vs��0�"OR0��$^�U��Ȁg���Bv���F"O�B�RYFUس��7��l��"Od�3T'�0@$������YQ��"O�)YA*��b�Yp���&e�"OPa�@k��lǚ��p��8Ö��r"O���ƞ:�$}��#��p�pqAS"O6,��I� �Ɲ�W˸>�ɐ�"O.�"�
��m�l�M�88j�cw"O��3@O�.�a(E�E�⨙+�"O���N5U2�s	G�a>�U�"O |y�mU�z�-�"F�3�Ό�"O��6��u�8�1�L!}n�x�"O�͸X����)E?q�}����*jZ!�d��i�/2<�HQ��j�.'-!��&��)q¯�oF��7�]|�!򤑚(=�qj��O Dl	[O[�N�!�� (���+��[ $kahO�h!��¢@�b�����ա��~[!��\�;����F����PufŅ)�!���_�����Љ#�v�+��Z�!�Nm�|;rf�8.!"فQ�� �!�Ą�&� Q�U��+"$\c�H�:r�!�q��p�񬝁�T���4�!�4	9���0��u�fQ&��%�!���c�I)��#�~��(�'D!�dZ���58�<~����,$9!�G.n(s�,�	z>*9r�D��f�!���1�4��0�N�	䀓�D<�!�B�	���"[�)���QMF(R!���:pǨ
`y�G�Pf�!�@0��`�l��34��î1!�wBY�Tm�V��e�SG@+!�DD�P!<��Mѥ'|Ԕ11lc!�d+Mێ�(P��I`�0�؊�!��d ذ��7�:��j�&z�!�$0%gN��0l��~=����N�6�!����$�K��$I���Dh16!�$�Fag(��`c�����N�m�!���'�.����߄�p<X�B͙.�!�Ė�� Xa���ِd�fT!�YR za��$�("�j�Q3f]	F!�$L�2��M�#��k݆�R�KJ�*�!��՛t`HѸ!�ȱ)ʄ��^�w!򤔏S�C'�Q	;����
�!�Ď#�٨�@�4���$	G0ge!�D,6�<�ࠬ�\�ݣv�ћ8E!���#*CVP�g�U4A p�V�B�o&!�d�c:����o�8m�"Y�4��3%!��������<G�|e���K�f�!���
0 I��D�G��}� �.O�!�@?�,r�`x۠���*�(�!�$2|*Q��pi�����E�y�!�R3TQh���!�	}�L�p���1.�!�$�$e�xkׁ�
J��-ۥ�!�Ҁ����.�'l���	�m���!��M�!	d+e�׆!�� &��a!���p�i!���*@���jK�-!��<����*B+D[T������r!��8l���§S+]Sh!�$;s!�� �CaC9%,���N�|bмY$"OԠj�.��H٠���%�v"O�8@L�\�L�����7
4��"OD�:$n�7:�H����'=i��٦"O�D�3 ;Ȧ� �Ǜ�a|�d�"O��bT��uZ&���Ίe����"Of���,D�e$����2d���"Od���+ZO�H�E e�}"�"O�I�m�0.{�0��L�E�HZ�<�a	��J6ؑ8��L#h���.BW�<�eJ����q�/BY��p��Q�<9�B�"k����l��hW�^P�<��,��D�[G,E�dj���kBx�<M�l�˗ �k	;F�t�<Aq��8+h*�#�.8�Z*�X�<Iq��W�д��(��LB��O�<�rA��S���BB�f3t��U OQ�<���0 ?�0WG06H�Ԋ�D�N�<�g�W�N�~H�G�xƍ�w��b�<��mʒ�&���H%Ƚ`N`�<I�0'�l`�mku���_�<A��R]D�BV���^�Z�+Z�<�!$�]p���T�Y(<�R#�V�<�R�3V�|�R��E{�rTP��R�<aP�v'�]Qsf�*�r<H�i�M�<����D�p(
��!;��SU�L�<A7���M	2E������HUkL�<Yt����dH��,���D�<�$Y�`lV�B��f[|l��A�<�w�]�R�\a`G?.(����<qr�H*\~��B�-8{8�;pjCS�<�)�3n���}�z�r�y�<A䂖�aO��6FP�is�@+�~�<� �i��ݻ��хr� Xñ+�{�<a���+�� !5b	���`��K�<��ҭAr�R(��s�^�0C�K~�<�sG��3	�< �(ͶL5lip��O�<1�"ć��<:���"|�SEo�I�<�t�4TtZ����{����B�L�<I$ `U\�A�
U5ȥ�JG�<A���$VV� @�iU*��݋2LZ}�<q���5@�r��#v�x�ۢ��z�<I��3Ѝ�)�����LR�<��2���A��&,�
��r�F�<Q���4��P�aP�1t�y4i�f�<�3O#m�|a�"��0I��)AM�<9䡖�&53��P$t���я�J�<��L�4m;��5aQ���/�<�K��3�+�f�UN�8��ˊv�<�U�A�{RԊb�2�mi�Ch�<q2���hV�d�b��73���zTH	e�<��JVnjm���f���z�JVb�<��6f��a[ N��c���JbeCC�<ٷbA#�Rt��l�-�*����_E�<��:7ۨ-�&X+tB��@�<���$R0N�٥ �$T��-�7fHT�<q��͔I�k�cD!�
l�PDV�<a��p(����<}HE0r@Gw�<	����7K����GB�#���"o�z�<I��A9sFl!q*��b��գ k�<�Q��8^�~m� ��v7^��`�k�<)@�?:����ƺ:޺`2�'�}�<ɱNH��`��T6%tE
�b�p�<��Z�:�zaj��xYB���I�f�<� )���^�#�P�``A�aa
	��"O�(��+��r��iB�mE���"O����3@�]�c�w����"O&jB�CS��"ơʣq��:�"Oു�X�b�B���R�,'8$P�"O��U��v٢j�C��Nt`8P�"OQ�1�H��=qD"��.jt��"O��REe�~-@JV�)j`,#�"O�\�U씩��	��?|���u"O1��ӡ.�}RG�K'oWԊ�"O��1d��'hs�%B�G�DJ:�7"O��"g��Y�2 #4�_9.4��zW"O$)J$�ѕK����qDT!~�R"O0p:���2��Q*���,		�'���KAÕ�:�� '���h�
�'�Z%�qB0m���q�BΜnJ�!	�'令+�O٪Cw�%pSIq����'�8ܢ&O�,5x� �Zl� ma	�'�:�I!��{˴ݸ7�x\$���')�dPUƻC�i��˄h�~���'���
1ۜU��jS3Z;|U�
�'K
��&_�0�R,��M�WjR���'�`
�R�6PPEN[5:�:�'�XC���+�rx�a�C��5��'�u�"�#N�l����#8�nY��'E��C੍|n X����]	d0:�'��yRhX�6�X�!4�Q%^���[�'��ݘ���+tA�Bm�,S�!�'|�wn��}�VU!�*W~��1��'Vm���Q?~��1N��wrXL��'�&(���m8Ѐ�n1B%@�R�'�rIp�NS/	l�i��VF��YY�'����L�
�:܂��5;#�a�'Y��脫��y�,����I�-�̹�'��5�M����[E���Q6��'R삒-�nF��BV(�C"EB�'�M2�/�(��q�-N�K���
�'�0)�\��#r����	�'�h0�F�_LsX�����!�'�8zR���M�d �N��|�TI�'���J	�Y�PE��$	!I�,��'�P���?r+�M�k�5ZĢ�'Ů��6���I��Ӓ�=+�'<*�f�� *�U�Oح.���S�'��'h�p$k5ʜ�%~���'��KgC@+t�����J��L`�'�θj��c��$p����\�	�'ܠy`��W,[��I�#ώ\�#�'���w�Do+r����#M�B4�'�h%�G��8=f��t ɏ9F4��'���¦C��E]�9aJ/;h�]Z�'uJQ4k�632=1瞿8��$��'��T�r*�1�d���Aа�~��'�N�z�"_�gU���x�����'̔�b����Ve��劀e��B�'BD�P"���_��H]-_���''P�H%��U$�����R�m���Z�'���tV��T�6�Z�j���	�'��B�]�J�Y�_����'�^13B�h��@E�_�ER1�'��(��A�$HईC�ϊm��Y�',���C:a�-C���(a$��	�'�"=)���^�x��B��V��X��')zh�*��R��� �ML�A<nr��� ��C  ͒�� �%E� ��{f"O`D���.�aS�K�{��T�"O��+r�V11��f�C,FHd�"Or�3Q�D=|�� ���/*���5"O�P���7��=�䠜?0t쁡"OH<�`��QK�بdo��{���V"O��G(�ƒ�z�/d��q�"O���@�B�9W�YҠ��,M��1"O��BO� �R�ę1���y⍁_,��ҕ�_�|�#�)�y�]J�b��&IŎv�}���Ŗ�y�X��v�h��M)k�� �5����y2B��R̸Z��ؽ]���o�y�"ӨV,,債i�[���`"�6�y"%�\�v�!���$}%�P�t,�yR/=w�AZU�: �&a����,�yRB�~�H�#�D#}�Z%Z�眬�yRL'z���֡�A��U0F	�<�yB���S�4�ɇ�ߚ�8�"�K�0�y�ݢ+��i0���t�L	��y���4&�\��2j��S\���yR��$).l+��1�:�2E�V/�!�d�܅ѻ<0$�Y�A֜x�Vͻ "O|�X F$���Pᜐ�\"Ox��%�[�R#��#ł�A��J��y�n�!���GA�-o�<�f��yb͉��m�0�W�_{v�2�@���y"W�SC��jrAQ�X�^ ;�X4�yB�5I�g���x�>��AΖ�y��2J�BtIG�B� ��QC��y�Ȍq��I��d*�fL��y��5o���d���(�H� ��݉�yR�N
:����\ 0���V)��yr��>���놪-u\-�c���yrH�8���&��:+G�Đ����yM]��v��Vg�� �P��3(��y�
<a��l����&DzM�f��y��X6���Q5R��*ѕ�yB(x^��:�EW�X�� �F��y���6��u�֨JT4A�K �y2'_F%r�w��
G���ɓ��y�-O�r013��,�P�� hM��y�)щ���B� ñ ����%��y��K�$R����[>h��D���y���a���G*��X���y"�Dv� ��4@�-�9��ڦ�y�˕�4,nE	B*�4!�51`hH.�y�����x�Q@���d,����y��Zq���y�Mġn�P=�G��%�yb��8w6-���̎m���36-ڼ�y��M��4�d���e��y���D4�y��_ 0��Q�oF+�,Idc��y��:<p���0�Y���PSº�y�m�:�X�3���)T�Pű��֙�yүԉ[}6�	�E�N��p[��Ƨ�y�$�.,�@�p#��.(�Th���y�G��~��{��� <(Z�C�#�yB��~����[�	���R��6�y�ɓ0s�>tkD`��|P!���O �y���������t�^�hBe��y
�!9&)���<B��h�����yr���<��J�%�Ei�J�
�y"c
84xD�*F��Z�c��yRnţLF��b�67�e��.S��y
� ���إ��p �$R�%�5"O*]
�B����B�RE}��"O�4�wjW4W��R��A�֐�	�"O�a($kU�q).u�V���q��"O��
�OM
q�,-���A:/�B]�"O�q�2��"Q�	��d��p� "O�q 2n�6h�R]�hR���$"O�<��DϽ"�t8�f��	ά�*�"O�5Q�k�	��IL1h�A�"O�\Y&���R�e �*�"�"O�5�q��-S���7D������r"O��a7&��LFn��]8IH�D�G�<���Z�l�)v.��w���p` ��<��o,�%��)�zH�G"Rz�<i��$au0x�i��4��@�<���&g�Pj�睃U��%�{�<��G�4�P�P�f�y���B�<A�l��6��8C�W;Ns��[7L�|�<����5� L�� صNg��@i�u�<yg��+,
`ʠ��-y=��n�s�<���qc���08A�=�&Bm�<aAk�x��A���VZ�`��[k�<��4$9�\S�D�)kf-Ywg��<��/�!P����c���2�T�3��w�<�̟��� �cR'e�X���}�<�s�G�(�T/͢@3���S��|�<au�K�eQ��a)�d�rX���B�<�T�E�v�)Ӆ\�TAe�ׇ�Y�<y�MNH(�F	�?@B2��`�SX�<����;vXz	���I�R� ātcU�<�S���|�����8^+��9�JS�<Y���*G�����nB3;.y��P�<q�m��,w\dP�M:v ^�QfPE�<AKY�%C����I��eJ��~�<ia.A?��Ss�H�_LĬꔍ_C�<�W��%P����b��3/J�0�J�B�<��*[����R�k���@�ΚJ�<��ǂ F�Py�������l�<�5��;��d1��"����B�Q�<���+|��C%��+t�yY��L�<��	'&�u���Y��ac�<�1gL���}PC	�K$��Sa�]�<y�����-�	b�q�a�<�%K�s���w��1F9�U�bI�F�<i!b�< >��.^�KF����K�H�<��B �8Ab�Ƅ�j"�`�z�<�6nٲZH�T��.5yd9���b�<&�!,N���]-a�0i�]_�<9�eW�{�"�ih*T��+A^�<�U	�CS��l^%G�Q���E�<����T�K!���!x`Հ���X�<Ǆυ2�Lh�奛,�0{��QQ�<9rIv�b��ьͳ2�b4�׮�X�<	5ě"6���J���D6j� #k_T�<���e��ey���!G�ؘ���!m�1��h�;�<x�u��m���ȓZ����
���2`�4�ȓ	�^u0�hS�dS8,
6 ñk�Q��n�L��37��9�H�5�����P�40��7P�]`fB/�Ԙ��X?����KW�}����5��/v��i��$1L��[3f��Ǫ�,	T���ȓ#���5	U��B(��F�/O��5��Gu��yU������FEũh����S�? (yRu	]������R�)��軦"OFDÔ`���@�"�B�"����B"O�ñ��KP�I2u� ˘M�`"O��0'B�{�������8�I�A"OYK���W�0�qV���Dɂ2"O���F�y �� �ؽ&�䴺�*O�m4��Vאe��"&��!�'�����-y%���2��+��P�'flAPW�<LC��C��O�Ϯ�z�'Wb���\�T�����;V#�YK�')~� u�5%��h
S�F�lA	�'�,�h7��5r>�XS�͝Ax�-b�'{��v0?� "fd����
�'�P�Aa�2S�ƌ���.����
�'�����S�naʽPƒ	ܤ�[�'�� R��ҧ� �˴���|��}
�'�Lh�� і�2�C�#�&pN�+	�'�D�#��O09��4hT0����'�:4��EݛDњ�����n�r�Z�'8�%&
�%�*q��N-l�~��'�\B6�2N�*I[�f]"�	Q
�'�e*�HZ/E��Q��]
2��
�'�8L��W�2�@Xc�@)>�A��'
�]  �׳Y��}�1+_7 0�@	�'SFuS���$��5	�&�}�֕�	�'?RԺS���<��A0E��+�\ �'��5 W�#9t���3 P�UNlDx�'�̵ ��F�j�$���X.Gw
$h�'�&a��ؔ)T��5CO?B��1�'Fb8Bѣ�*[n�[`#^�2�([������rq�@���kO��p��$�!���;���G��d3�i����\b!�DċP��8���+5ֱڗA�mM!�d\�'����g�Rv��\�TcَU���'�S�OzB�p�%қ�xv
�&j^����hO�"2��e��BEeɅq1"���xr�'R����
M���ʱ	^*ݸ)O��GzJ|B�OLza�7n`����ׁ�����"O�!���ݔ|�8�s��42{&��x��$?ړG��K"�ȥ���nK�-I(�*�'�����J�mH��G 4:6b�'7^=��)�u��bj10Z�T:�'U��@��J�F�~m�� ��(;�8z�'I^�R��מ;E��sDώ%5xP��'U�		�Q)>���;T�	&�~��'{RiI�-�+D�IBR�Pt�
���'F�00��SV�P����'Xvt�@�'���� �Ƞ|�2�zg,@/b����
�'�u��b&<�*B R�id��
�'`�ms5]Yj����-�ͣ�"O�d�A�8Z7���"!% 	5�'�9Fy"��!����+9X�����ź�y��O>{�"b��OW0�͹�k�ݘ'	�-�	t�S��OP$��Z����Y���]yqO����u��T`Q�S�����%Μ<��&�Oҡ�&��;2�dqn��|QȐ"O��j7�h #�D	+r<C�"O@����.ߨeˣ'�M�VȰ�
Da�����jȽ~0F���ȍ�]y$����ٳ�yr�'�j0��䌻O[�x�$v",3�O��$�_��Xu ��*J$�l��VEl����+�$��Nd�I`N@�&��I���^Y�F{ʟ�Ig�ƶV������[����"O\�5�ڭ<�J��@;*k���S��L������ $J���-a�N�#A>�(�c�"O�`;F��x�i�O����i��'$.؄��$��}�EB.8*����
������/�?m���!�/r��DB#�l�!�ٛ!� =8jFt*��%O�HL�P���?)2a
��)~hEJ"I�n�dL�m'D��;3�H�6�N��V��_j�y�cD��hO?�dT�S�&d&���&� �:���,\�!���/_b����Z!�>dȒ���b'VQ؟�2�a� V.�q%Ӱ&�\��=|O|c���v�� RT! ��Q�HL@����'D�\��J�k��� ό;*�k$D�X��̉�u󔭘RN�(A����&LO���!EF�'u�6��@$��k�F��q����{"�t�0Q���$w�Y�A���y"I�]��CbIZ�!�N��̝��Ms
�''v�b��R�8�� K�)Sd�杣�yB!�K�~c�p&��J��܋`�A�6���y�fB:,O$⟌ӵ$>J8��DP��"˗R��'����Ϙ'���0JϘ+*^�����%&)ϓ�O�T�&L�袐��h_w*4�w7O^��$4J�9p,Z4SwJ��ƛ�o|r�|��{�Պ'q:`�t�%�x0�r��-�y��"#~�ęt`�b�*9�Be�+��=�y��ɍ��0{B�S*Y{�-A�ɐ=�y"kZ2]��c�R%1��s���~��>���~JFQ�D��*OC�9!q
]@�'��O���q�t�.*�2+��(�x���6��0<��ƚ?@hY���3�f����e�<�ծ��x��s�{u��F�L�<y@Y���p�A�,@��5V)_t��&���"�ǔP���+a��<#)$����4�O��oJ$2�H�r+.��P�P�\����ȓK��d��$C$=�޵�gkܻp�fd�ȓS��M�3��-��P覎LO��1���s��`�hI�)4����L&@��"
O�0ط�]g
���"�Y�)�v��d��a{��䍷2�9�dv�4Ȳ@����'�qOP�'��@u���F�B�8 �V��/Wz���ȓU'�૦���ڰAũ��eF.,�'}�D.�)�'?64�PP�E?��4A � 5� ���)��<"�ԘR� �'G�#�����kd���t~J|�>�1J��}�Q���[���+Q�_S��T̓v��Ī%Iƾ�v�8w��3%�<P�ȓ_0�u���E�a����B�*x���G{���O��Z��Y"j��A�({�v	�"O)�۴�|�yӏSU`:� "ON�3���6
�"i8�.�)F�B�"O -8�
��D�~D��@��pٞ$��"O�q�c':2�H��H�rT���"O��:$J�����I2���qX��"O�ͺw�G~)�1"c,
Jښ���"O�`�EŐ����0cj�Vlؐ"ON��
�~*��T*�6�̠�t"O�p�-;R�uuD?
���ѡ;O(�=E�Ĭ}6�xS�ˁ'������yr��I
q����aS�����1�O��+��(��,�Cc̰cTt��"O�y9cdG�aX��z�'DIY%"OLsڀO�P�c�`�<�(jS"O�5b���*�x��_8R��"Oaس�G
4bYy��<1�\0�5"O>I�%��>'I�pP�k��49�"Od���I%e=�J5�OP�64r�D0|O� �8ȖB	�y@@�	���zd�vO��ٰ~��2V"�q{��Vm�z�!�$ˡ?�#�E[w( �	��$�!��T�#Oti�5&9$w��1T�J6%�!�$I'b�0!�=���h4�قs!��N�}��u�%3��@%c<]a�ԅēe0��"�:B[�)���
�P�j��ȓ@��]bR#�^|ej���*3���ȓ 9L�pňX�4H<��f�ک��n�R?!���O~�S�D��i5,��ĨD3Y�~�0q��L�Dؚ�'��}8��б�w!��J�-�	�'�X�#�&��T��Xd�
=lT ��$s��ϓ��OK��0�$~8��Ӌ]�>.��ѳdl��B��Hn)kG��~&8��&�1]r1O2�'@��O	q���#po�����B���4BȰˤ�,D�<��_ �P6��7�܀ұE&�	I���S�9�T��/�8H.ܰ ���<HB�I�c���P�-_ܜ�1%�'c�B䉙!�ȠRA�;$��h��St��Ɍ��F�a��N�qR�Xr@E�~�ӕM6�yR�JA� ����!�6�R� G��M�)O�јM��g�v���5�Ʈ|��@!�&x��Ć�)��ݺ�%�mA�D�MĤP���Fx2�'�V�xql�"T~ʱ��S/R���'X�
6���i�t�A&.�sK�i�5O>�)5"�;S�e�r�D�y@"Oa�G��(4���p���*;̈�"O��や�_�, ؁
�I�*�"O<��`g]�$��*��¡(R��"O�ԁ�c9Hxm���N0y����"OB=µ��P�{U/B�r���"O\d���+V��g�^!#̞���"ORP�d�ʉn�D0 2�x�����"O\E�W<9�Js��@D˘\�C"O���EW�y+���t�X���1�P"O%xB�\9S��IQ0���IZT��6"Ol���ʼ, �X:W��C܀ �"ON R�l{� Q3f3��0�*Oα)U��y"ѓ;���	�'�2%�Sc
lR��1�Ћ;��+	�'W��FJ�A���k��]#/`�!*	�'R(��@\ZE+�P\�"���'}rL�q�^�|N��kV�+�͡
�'<�ա��:*�x����3W�P	�'t:uj#�>�p�B�ꖝy����'��@{'��@ȼ�ʕ�[wܸ��'������|$	�	?m��P�'qh����J�.�J�F�{��e�	�'j(�!�
Ȁbu6�g��oBx	�'`��������:}6�a���'�D�:�FR54���3R0�<*�'
J=��JћߨmP���"��
�'g�D��D�0�(๵c�]�܁�'����B��*Jf�!�ˎ�M\�P�'��"a#\�}�8��#��1�\�'�2�
� � i�t���A@�-R0�'p�|8��؎Fǒ���ꋚ#����'�a)�/Ʃk� j�g$ou����'c�P�3�R, �����Y�5t��'�^)�����Bc�Q;歆?w�$,��'� b�*��!��L+�k�
�$��'H��9ceQ�<��ITO
�d���'"R�+�n�T�-��'ٚeۚ50�'~�B��F�b�Ri��N�/SWJ-R�''v�SV�T?�
�J�E�"q��:��� ���퀒P��p�Ǆ����!�"O2�r���^�|���&�{^��"O4��P ��l�r�Q6��,Hfzpy�"Ov�5�։~��Vl�#!�ҹ�"O�\s�)_��$:�k�6}��"O�!��4j0.Y��
۲v
V0��"O�e���1:*�|��*��|�yp
�'�j!�� �	�^� �*�a�����'�V��D�ύ{ެK�ޱ_�� ��'� Y�Pi�"'�3@�9O��ܸ�'��e[���i�$���  ���	�'#N����.��QC``�HH�	�'��t: m��+
�(�P킺���'�\�D�zU(����<�����'6T��WjP��L�``m�2*G:z�'�|KCА�B��a��t��ȓPR���!A�L����cw�U�ȓ^�a��F֣IE��"�(ՒC-��ȓoP��˶-�KzԂ� O�tZC�	'�
d@�
/o��=hb�C�6"PB䉏����VD�&r�ui�]d�B�r��zb;(tl���ܞkhB�g�9��	�g�q�cW��^B䉋Q!Y��K�H��7҂0�~C�ɯ$�~a���4&7Rl � �q�0C�Ɍ^b�M�Q�sG��S� �	>�C�	�~#>��f�ց+$��QMD�r��B�I�:6zx�W�W�W�d�(>�B�	� I���Aȼ.���A�2f:N#=�Q�ѐ%�ʢ}�b�/�'Ȱ"$�R�<�
־f�$m����r@*Fj
:�d�Cv�ҷi�ɧ�����ar����؟5ބ�Jԃ��y�,��~�4�[�$%L��i͔��yb��V��]b���]�������T�+���z���T�$�O�+d�/��KE�ɶ��r�ìn��� Q�-x!��W/v�J��1��%�ƵJ�។2k���"&��X�p����=X�47OE�D!�d��I�@*�B�I*~!����9���	D���q��
��>��D��>E��'��𩒒5���D��'�,���'�����(�y}��R���N4H�'����G�. bх�!oZ*x�u��2"0 �F�]���D	#>��D�6,|@��(O����@
�?)�U"�"Ou9aNͰ=����2��p�$�I<��,�ܛ`zQ>�r#'.+�N�8��+[�����)D��b��R�j1V� �k�#KH�a�s��-$q�F�ŋ��S��?a!�Ûy1� �'EI2h��=r�� ��m��[�g�8[I�!��| �����<��e$Ъ��d��{�h@Ò*jӬy+r�"*��Ƞ1�W�j]X��S���5P��1D�H�nTc3ia!�DJ��� �I�?C��q��2,N�(jѪA���� 6����)�g}"�H�w�Z����J�v>$  m��y�n���v��r��/i��%�ȇd�L°�W�-C���&�T��lX�

�%H�i����s�D�C 9\O](��]�P?�8(�� �_��z��V�U�]k���L�Hm�U�ڭ�xr��!} ii�E�:kj��#�ɀ׸'���iD��*y��{1�J�(ռ��|Z�F�$b�e�W��!6t�u���<a�A�+���d��9�J\�@�	���S�bNmC�x��D��HG�,O@����A�{�F�"�g�)1���"O��s,@M�A���^~��0��9����ǘ%z*�E��axr`O2*�=X2��z�DMK�ĉ�ݰ=�cZ�h�,a� g!��"wᜂM6X�B./�Z����H,s!��!d4X#gA���}1�N�KS�|���n�<x���?G�P�p!@'�h!�$�YU!��#$����%�� ��s�䀒1D��/h���>��3� z�����kd��B���  �'"O�@�&�&Bs�0R�j��"OP���/t�NĲDO'#�fE�d"O�`�`	�8��d���Ѹ�&]��"O�m�.�"P.	����#O�fc,D��k�i^(Z��i�a ��g22U�BN+D�� eb�!��`2��u�`�5�S%N1Ј􉝹z�|u�&�
h�V�RR�Q�u����ܽZ#�QA�A�8G|v����8�RAhB��$>�K�Ǘy�S�OHj��%@������95�$r
Ó.���D���A����T�W��TZAH5�h3?a�*�$����$#gÈU����H�(\��g�3wq�	{�.E� m�P��S��T�r~�-R6� G�^�Zf�ѲA�\��R��1x!��V�" I�/�)Z�z�di���O�2��H��)a
؆#�qO�?g���c�o� rֱ���I��B�>b��q��ʌ�oO�x�f�7�@�r����$��Ƹ'c#}��лB�():�M�Ы��r�'��	���r��xJ|Be :
~)��G� �8���i�m��O(,��ĘDt�<p�H��P*�n�+��	 0��l�ӻt��S�4�R�v��S=��ը��V�0��\�l�	m�L�3�)ލK:�~r@�o�v�{��R0|KH<��j6�\��эy�gBrE��e�5Q�`@�w*���3�_�;HބБ��U�j�Z��Xl@0CG�H�"����R9$���3�.sS�@A�`N�<�`��=�`�'��!���}��'�Dy(�
�P���fb�n�a����U7x����� ��Y ��[�`X�<C4�s�,�O*TʅL<W���s4OV�t���?�c��Hv�捱��� �Lp-��*"剟A#�	Tt�i>	a)�6K��ĝ?p����bK<W���cw�+{7d<;���/)��sx��8��fs<@ە�	����1�ɜ=r�=Q0O�l��D<4"��+�PY��OчB��L���{f��B"O��q3	�1��[!g�=v��|�R�Y5���I�;|�����`��>�(��aê܆$P�[���V�B�� Z�$�����?�����ٱ��<��B���2`�]�~&��a��qN�U��B%S���a��=$��X���=��I@��٘��UjD�1*Y�ÊF�}*^�b��9���d�u��D^���<a�Ɇ���	���<���7~$� +�.}�n���WS�<Id*����U����������f�w�ɃHt��C��-n��?e2����Z�R�5rS��o�!��W�`���_�SRN����Q���a��|��ƏS���h[�`b��H	p$���.v�.O"!ȱDIfn��e�?#<1���<��jp��Mst���!��ck��S�*><OvŐ�a]6bh�̓��P:3�{)�qqB(zЧ��Y:�#�@0�O���ׇ�y38Xc�
�L��%:�	�"c�̊��{70H{�M���/r�4 2`/"����W$Q�B䉽�,m��C7v}�$P;RwX#=���>��ps�"�A[v()s
�"3�ȓ&v�H�q� oz���BG�������M���u�D��0�T�7Z	����Ts1AH6��	'�A=D	�X�ȓJ�L��bn��&��Aq��9;����I�<Y&�8 U&%b`�S,
E#ӡP_�<)D��_]@�3SEApz�,CWH^Y�<�0�L�!S���Fۑ	�ȭ�5�Z�<y�� 0W�ث�M��J։�W�<I��n��$�Q�и֦��AL�<YM��*�D�4@G�k��黣�IV}��� 8hX���7���ѡ��.Z� �YQ����ć�d�Ԅ�D�@����G�eZj1�uY�;�<�D"O��gc��XQs��*,����Q��53 �qn�03"|r�n��<A	$OB�2� D�!��F�<�����5'���G@����D�Z�N�b Ï=��$B���$�;j ��	:���� C�ĸ�ȓ/znP�+Q�vТJ� �",2�hlZ�kp9*Q[�EN0H��'�Z(����gT��S�N�3�� [�2�ܨ+��+.��IR�l+� �dJ�a�1Y����D�\VD�%MfH<�ЍT�t�~�(��ݗ��Yь�ϟ<j7�M?�$H�b�j\����O�`Î��HQ�C%�A٤C�. %�5�N"(/!�$N+�I�2�R�}�$��4m�B0��*^0�җ!ʂk�d@ۡf+	�A�r�� ���h�n�
#Rt,�ҩL'-.E�ĆF4V�|Z����^r�D��'�)�cg��I����.S%T^�KR.0>x�@�ĉ�a�<7�� rL�5�G��j�2a�a���K���0;m�u��m��R�lZ�Q�`���3=�	�l��$5����)��#(V8Q��P;O�4�����'(�8�.4M�dO:N�8���A�+�4�r5�IkT�����Id��rp���?>��E^)F�̓d�����m_����ĊH`��"�ƞ�<2�����۰��E���{����(��T����M��] ������W�:���J�;/
��TL,WS��(%,B*;ϴ����N�@���IU�.�����>'��tLE,VW�.ՄW�����J�T�7o_���2m[�͓J��y�h?{w�!0Nth`�0�xݛw����XԪp�ƺ�F��\����d@��> �1O����&\��%���(��s�߰=��`�$yvL��k.^j���3IBRS̀(Cn�&[>Lt�g�J>�0T@���	0�\�%�E4|z���C�	uP���+�@zҍ	c$D
��⟌�"��(X��&8���[��Ɋ,(m�N� �L�sT R����x��F�B A�:C*��I�]+�<T�
��V`A#��8z�n��Ղ�Cs�8�1�ii�m(7OV�2��O�Cr�(�Q���6�>��fޕHTD\�Ch`q��-�YF�(��"D�|��A3��ٸ&�]g¬�dN�6)NU1��؍kS�aXvl
�A���S2��͐f�G:�'�`ܠԣU�M���i�뀽=Vjy����P���c����C˦Ւ��ց_�ƴ����-=<�d.��t��o�bX^�AU�ϨO��Eo��Cm\�V�@+Vk�Qg"O,!f!�_��PU`�V���P"O���$
�R7\hAo�%^z�"O��qj��[l�L��'�td�"O��'!�#:)c��Z�5���@�"O@� �Kʤ�l�a7D�6�0�"O�5{"nL�G8��AdK�E�`�"OR�pp�ҩ3����f��+����"O�-�D�D A*J<��H�|�Q`"OU���E�=M�(8����#B"O�I�saQ�w5tM�e��c�����"Op�f)HVnݫ%���x�4�$"O9(���Y�uQ�mo �8�"OZ=�k�L�{B��|i��z!"O敢D*Z�9v�i%O�:M���"O�,{@Z�j4y!�.�]�-I�"O��SaI��C�>��f����L��"O2�1��ߵ(@��� /W���i�"O�	�!$�u�28r�ⓖT��1"O�M�BeR�d���P�%�����"Olݸ�ʯ=~��5�M25���"O�0�@�7yE�sA��0+U"O��Z$jߚLաT2k���e"OT	�fi�05r�բ!������"O
��D� �{���=��'N@Q��o�5�M��ə6#�:�S�'��xQ*�q֪��"C׼����
�'q�h*W��
qlF9��L(Jߌ��	�'���q$���.���1��Z�܌S�'��U�0� 	=�<�Ge�^�P�'���$�	�sk���1#S"R��
�'��Jo!����2�������'i��2d�Ơ�Ĩ�QAð@��'��Q�&�;'6(H�FpӒ�3�'Mj]`1# � �r5��F�*se&0��' P����S�""ܹ!�G�|�h�'Vj�S� ��r�~�A�e<FRZ}q�'��y����
èQ����'7�V|�'R�j`���{'&̐��<��D��'HPJt�Y6|�&YВB�2H�q��'�r�I�_���r���B�  �'Kڈ	K�$v�Ăq�H�ߐ�B��� d����2HgP��G�`�)c�"O�!����0�cƿ��Pa�"O��J�M�&��� ��B�zǄ,˴"O�Б�� }����ՀS��i��"O�=���IVx1�a�2�DȨ2"O��ё�*Y7�<3-]�]��}��"OP���F�p:���`��9R"OX"�Ң;�I���	-pu�V"O"� ��
zuJ80���x�"O��'�Hk�>**l�颤�,d�!���2}��cf$��0h��F˝?�!�$R�[8�8�ʓ�ؓP�T�'!�$�#"���p�	�`$L1�J?g)!�$t�V����Z(q*�"�5!�,A��1�۽|�,	�`OY��!�w<��!�G�j��hJc�!�D,X��OF��%�	�1�!�$�]��� C7(t��_�!���h4}0U/�-��Z3�:f!�įm����/;R�ʵ X�i�!�d�!tDJ`Z`�<>�0���X�B�!��M��p�@�}���D�Z�>�!�d�E�Pp�U�;^څ�'����!�DL���ڵ��iW���@��\�!�ĺ$Y\��QF�4>��&NǤTj!��#��rv�[�)%QI��W�O�!�$��CW��t�L+ 9��3箖��!�$Δr�\�2%�19�a�q��(!�dD_r�Q1��d(�mIW���Q
!�d[%&]�� A� `�"$i��'�!��� �phI4�ܑ#6�"e�@�!�>WZ����ބc+�l�2D[Y�!�DP��I᧛�U԰�$�vz���������Ɂ|�
���=��$cQ�V�HD!���B��|K� T5Bǎex�dY�S� �8�H�6&DQ'�"~�	�S .�[q�PݨHI�`�'>C�	�4����D�\��x`�
 7�� O����j̶W�z�>F,+BH	�2w���R+D��0>��d��_+�e9C�;`T)p����'�P`9�E6U��(�ȓC=�Hy�#B+@Sܠ���p�J�Dx2Κ�b����D�O�r���"<��;$�a&��X�'����eX���擂Kޑ��A	}��� �OK��s���qM��7aji���?��x��)D��x�˒8X��`r��Ŵ?���j�.f����+
%asLPӳ�'|L�Sd�ǐj��h��+E!�)��_-V(�`P'="�)���|���	U�D�")�}R�(�h�<9�K�1���A�R5>8�Dfl�'��8��\�UfpG�k�,X#�U��v���Kド>�y�n�=Y�n�2$呗c
�p� �D�г5HF,AP�O?��ڀl�H )�%`ܰU˓d��~��#j�����.�p��E�%N�����%h��$�1m^<S
ߓ~HX��ߨf�L���FЊJhXF|¯�)���3��I�'�H��$/h��=��č'�4m�ȓ4T6��4�˅8���)�GsL�a�	Kְ@�c�Z�a�t������L9�Œ%mZ���EI	/:U��b�,D�Xs����ƈ� ��H�G�<!�\&� ���]�0<Q\��UQ��@O�1�QCax�8�!"��%�D�R�<L^��f��.p��Ic፡I�"͇���X�c�"x�W�\�p!F{�HA=��`b�ɟD1�z{�"�&����'���"O�E�4	F×�-��{�g���?YÀ�3zux�r�Aݽ���S��Dݲ��W���N wD ��ȓ1_2�I������� 3��'�~t0&��J
PԘ&�'g�s��x��+���qJ�Az�qH�YB��� ��'	S�A���	:�Ѩ��y�!�Λ�.���Ò��`���K�ci��i�ᜤz��iH��)Ыe�ڜA�E�B�<MCp�t[!���p<���2���
�lB�G.4��֖�\�@G3���0iȧE͇`�}����qVB�ɷ`�HJТW�}�)�-ɂH$D��b��Ѿ� �ʧꀻ6ܵ�d	7D�<��G��D������܇f��	��f2D�dBB�� � f��N2����1D�Rc�C+k���7K�*r9B�[��;D�4��&������+�qB١��6D��X殆
h̉�Ӥ��2�Ғ�*�(cw#�0q �I���I�7�(�"3'I,Y�ON�J��˻X(��80�S��\��v�'^��j�Ā@��'��u�_�:�(Y��G�<v8��
�'��X���8̾��4욓vn�I/O�8��1hH�Q�M��|J ���a�Hӓn^�D�\��C.�q�<�,	�@��T�%Ƀ�u5������2]���f\[Um����gܓI����樉�n�2d�s�+KN�P���%K����@�дd��ɛ�ʝ6��(��Qcv�'/�E�ρ�h/0�w΋��<Xۍ�DD�(���˞8�ħ8,�d�,��Sl���aY�\�\Ԇȓc[����E�C��;F�Y�b��m�'/݋bo�bj�ݧOQ>�H!���3mX�V;d�X]K����P~ )��' Ҭ�El^`� �5�ׯA�`�D`-}"�B�[���eX>�@��-	�j!�'7��cUHM<g���K�$հ(���r��75��[u�Y
r͘l��� �;�J�/�� X�"ܳ�yBK�� ������H@��	*�*,�$.I�ఝ�GC�!�axB!�sL�l��|��UeT����u8u�P��7zҰtpu�>�Da	j����'�ll�7 Y�	���Q�&/ȬcJ���⌢L+qOq�����������[	���A%c[���!���>92�-�`���5�`Pq!�eX�l��:fh��R�x[!*_79ɸŏ¹�Y��a*D���T�@ 8�;���,C�u3T!(��eS�p��H����H@g��/�d�;����$�&"Ot��	��#4l���^�l�&�A�Ƴ;���'��Q��c'�3�d٫e�L����6)N$=9v�@}$!�$�P^Z�8�X- ��� mZ��3E%�U���
�-|L���&DͰ��ՇL�^����ɡO��I����$�剅�n�3���Te�]��ꈛT<�C�I�7�<�EP%<C��9g�%7�O���.čLd���� ,Cb� ��eUSZRݱ��ڵ@�!��"���s�G�%g)��#E�ԸLld�0B�|R��9Ni��+2V��6㍏/������E�@�>�����8S�X�f@RM�aG�K���hq!ڍ2w����M(i �؀uaHb�����)tJ!��>0`��\;�ܴ+���?A!�����u��ký�\�X7m4j7!�D@��P��2l���`�C 9���\�
dH�L����Ї�y�
T'�A����k����w���y����V�� ��Z*��æ���y�G|xMз�B�RU�=(���1�y�R
����;V�n=�&��3�y�Щs���Q��ۇG"re�F��y"D�A�^�Re��;R%9����yb$ݱ-ؾ,����'*�(��ɮ�y� ��m����2F	;
��S��6�y�e��#tł�댤;F͡��F��ybK�Ei�-�匀2��8+�8�y�n[�H�f�X托�r����mą�y"᎞k��:���𚁲���y�EDDJ8���e
��#C. �y�j�I��`�U���M�b/�y
� ^H�EӻU�VzDj�	:e�թ�"O����
&R��� Ɨ�P]���5"O
ȋ��[Y;��d�#S��c�"O-z��W�X�DUX�C;���"O�WD�~L��'C�F�(DeL�<Q� ���x٢��
Fe�$�e�<�@T�r�,Hu*\:j
$�k�<9e��,\F荋3"�&d�ӗ��S(��EĞxyR߲s2J�$�'��#"�I��;3��x�P3v��� VEݾD �ȓpq�l�gɌMtp��Daɹ>�ȸ)G���}6���D'��M���ӎ�|�G��Oqx���Oe��E��vA�E!ط0 e��'�pl�{C�x,:���1���+&���2t�۴^���3R���>�&�Z2���A�UӅ˹ �V0��H2�6&���B����#b�ĿS\J��?�7JK+gX��s.�O<�;Ǆ��z����W�E�:f�ّ�E��e3��"F��:k_@T ��\Wx�J�ld��Ȑ�g�p���IX17$���@5��S��'��	#�B�ix� H��b�h������?�ͻ"Ǵ�6�Ѡp^��F�P�%�d)����%CN����9S��5owT�9����Ӄ�����9�Q6hxL��*��pА�I�5�M���2�F��$[u�<�d��K����;`��d��*k2�ѣf�%�Ms֤��Gj��1I��omȴ���bHZ�ڰ$���5�M�
p@p�El�'��R�Fсv�g)�7(��iS�"e�9i �9�����q#�ӶjZ���`��Y`��A".ȴ|K�l� U-5^EJrh�!�T��'Oʭ8a�E�j��"���̆�2�\1V\�h�Oࡌ�*@I��c�i�
�qb@�:�w��H�@k@�l�V�l\�c�m��'y��4�^�ɸ�*#�2�Č�Ӈk�@d�n��A�ـm`F��'	�R`�M�	��$�O�7��!wE���* �m�tH�@�'Q���C�<�'kƃB�@Ƃŝ;[�beί�f8xD� e-Xة���.R���3��88��◄$+r�`C�a�مȓr����NS�)nIQ�@B8t�����zg� ���EPo�a1$�2�)�ȓ7����c�����%Yp��!��a�ȓT���C��e�< `�z!�I�m�<�`�P39�6PS`��A���e�<���Q��ٹ���q�B�����`�<ٔR�n8D  ��a]����Cj�<��N�!h1"O1n���`�KGd�<9d� �q���e��-E������I�<� �X���+Ԯ@
��mZG�<	7��7�Тց!�h ��+U�<���D+o	�聳�=nb�dC�C�V�<�G�G���\!�H=�bv�R�<����."����-��tÑ%EE�<B��3'�9�H�o!��`�C�<���� ��H�S%X�tjH�*%,�b�<iN��G�PyLV�5��e�*\�<a���<��1����B\�=��n�[�<�.̹Q?5�aU(ZD����A�W�<�p�J�K�t���+�~PZgGM�<A���(.��l{ �$h뀼�RaTJ�<�̄�2y�u{�� )xT���֌�A�<'*��fsƽ�צE�j���ct�<Y􆛼'� ��d5 LZ�h!D�Z�<	��~�t��,H͞��5�B|�<IR��^2̓�#� ����cD{�<�lD�arF�т �)1ъ)�qg�t�<qC���@\�%+P�7:�s�Eo�<1)� dQ���q�D�R#R�o�<9FDA�\�N��jW ��$S�o�<���PF�
�c@ 9mCr�YN�<�0'�7,�$cua߉.i�$V!_I�<	�FȈ9X������"e��uh�B�<)��D)*���
C"N�r����~�<��f�pҀM���_B:T�!�@�<9ԍ I��T+�DѶ]"Z9at/�@�<Qd���N�.8�ˎ8Q�D|y�+T�� h�Qv��J���qG�w�V��q"O�U��
�D�8Ɯ��B-�2"O4�X7�P�p��82T�̙V˨�j2"O��p�4	��l��
� � g"O
X�cAT]2&t�2��!.��H�@"O���OR�G9�0	򅆺.R���u"O�R0.O�$��Հ�#�Uo�U��"O���WN�V/ݚ��ͦK\*��8Oj��P.>G�P�4ES?9������&}�I��<�O��02�{�V� �rp��*ȕ'>}�'� ���1O��(çw�h(�o�*7wи�Ԅѷva�=a��{���l������8Q��8\~&�,ba�)�Ӂy�����|����Ik��P�B�<E��S.��@��cS(Q��UA��W�M�ua���~"�T��s�4(��-�h�e(K�z��� b� ��	Vy
çO�f����^�J�W�A^	l��"��9}��+�0|���Ђu�n�(a�,(��Wh��Y��Ķ�dIQ�U<B���'���>�;%Ԉc�@����81?Cr�'8h)Fy���(��-[����K��}�A5c���2�(O?���*īd�`1��.*H�Q�O�:�Q��	$�'	���VMн-e�E��#V'!�*�Ex2:�S���Z�P�v=��EPp}:���N����'|8"=�|���Kpd����� ��ېlIT~��!?QJ�"|³��n��4�'(N3L���I�$Z�<��	s}�>E�T�Ap��A
�Z�t��sF����$�(����p|�GɱEX��G��Q��!�d;p�sA�+~���	�2L�)�����$[�c�j���-W��R�	�YH�Q1������S�O�>A���?�Թ`-Xrz� �S�. *��m=��O�n���Yr�,��^}�遧�F�!pY��OX%��Oj�E���[���1���
Obݢ�f���D�Y���U�O�
�yg�ˮ|��H� �x
�O�(�'o�\ l%��"i�e�5"3b&�EiS�5fV`�P}�4+v6��]kvA��a�%_s�O�(P��H��y��&�I�p��B5Y�6�A��ݬa�<�؁DH'X�a��%Vw3�S��V�<(�bB�rY`�x'#��EZ�����0k;^�
�� R�|�j�N/,y!�Ğg��H�/�C-�}s�bG!򤁩(�9�7���ZJ`h��n֭�s
��<xj����(��$�H:V��[���gZ�k
��ȓ'��A�&ᚲ#�,�2��ɘ8bh=�ȓ:˨e�d�S�H���<�e��.�����SBDA��CF4B����ȓb�:�RlI*�ڕ��D�ĆȓiN��q~��L�1r)�-p��r�<���B�s��]K���ENexaKq�<�Q���N��)'��U�[H�<�A��8#�l�z�R
N�P�P�<�'��d�j���OHL�6d� ƞN�<�P��7/���a��
1 F�H�<��D�{�>YǏѕx�� ��E�<� E��%�O��H9FBܬ0��C�� z"�:�B[�'���#�^~�C�ɗ:��1��٦=�>]y���`}�C�	�,_����Z�w�Dt"�O7��C�	�{��B�E�47&� G��	��B�I*l� �	�Ş� @�a1���~B�I2�B5cf�S�Y �=c�`(y�PB�:G?��3D����1HEaK�kbC�ɼ[.��ѷ�۝L��P�>bU.C�eќ��7�� �(a��<�C�	����t�Lr(Q��k�w��B�#'Hb�Vo]�p��&]B�I�<ԙ��Ņw��1r͈�e�BB��"	,����ߙ?j�%�Uo�� �^C䉐:|����.w�A���%JXC�)� ����V-����g��H���u"Odhӓݿ��Ġ�R�N +%"O� Q3��ki���b�����"OZI��@�[�\�+�OC�r 0�K�"O�9!���J; �P����(�u:"On�:M� ���ւՖ, h`і"O<��V��%+��:c�Zq� ���"O��G�C�"�a��ۯsozhz�"O��c �>�j䲰�ƦF�͈7"OV�J�$~�x��/�~�T���"Op;�'�au&qz!�O7m�\-��"O�lq񎆉D����3���l %"OD��F/V�5J5��� BW"O*q���]�윩q��"O�`#`e�>ʴe��`�3��M�"OV݈@퇛Z�2A��oO8|��!��"O�$��$�~:�ɡ�(H�.l��"O�C��X
iT�d�oD8�A��"O@�'G�l�*��"�Q4�.��p"O�j�N׊"�͂�n����4�"O��$���^5�g��y�J�V"O��%������~�����"O^	xp��h���Ö.W�t�Q"O�1jA��b��b�� T|��X�"O�L��@�<N����J�'
p�M�"O�ђc�H����#p
K�\`�(�R"O̔�*�/V�
!���N)pg�Ī�"O捘e�]2��hҷP��]��Zz�<�Ø;|�$Z�*X
Q�ޱ��eJw�<�N�5c h@�FQ�Y[�Hu�<I���e�|�@0%�8q��� ��f�<a�bF>iWMR6��H{��d�<q��N��0��P:��0�Yc�<A��Zc��)���*؊��U��`�<����Wq��C&��<^���e�[�<ɰH�R�X���/+1��FN�<�ClK#.��l[?�v��WD	G�<��V�fh;�mZ;��m:w$�z�<Ѵ&SP+P�B!�
�!ʧ��p�<iL��U������0>5dȞH�<i�l�4q�&�Rc�0!�\|:BgDF�<�rC�*��e
G퓁��ȉf�D�<q��� `#@iA&(���E�<IŤ̗h��ebů�C���{V@�<i��� � 2F��~��I���z�<	7ǟ|����!Xs)�� ��AZ�<��ΪI+��H �G �9�c�]�<�SGL�'	��2� ^�T�
�j6��S�<1��ѱHȪ,Å��7��H����N�<�Mތ%-^�C��؛*u��˔
OG�<y�#���FJn
.<s��A�<i6�Q�m)��Ї*Ɩ]���'�h�<�n o���s��[���=2 d�<��}x�!V�B)���1�[�<�dFǍ5@�I�X�$]�1h�l�<Y�g�'* �+q���>��5I���C�<�ӍυK���u��I`����Dj�<	1#	{DTI�х��C<�Qz��h�<�'O�;	%&�s�G�H��A�g�<��5���ޮh[r�3���M�<��"o�RPb�*[�{��K���T�<icDF��*p 3h1A�\ +t��k�<�JG�*G�8����0o�9%�Z^�<٣!� uo25#�F�*nD)�tf P�<� tp�s)W 1lp<�	��o_����"O�I��@�}zuꃂ�r^f�a"O�ق5$�,
@pi1v`^1H\\U"O(`8d&>JSڤB0�ݵ5g�TXR"O�u�ダi����P/�,^�\ds�"O����3/b\�b�g9'��@"O�l���غQ�>!#��@>��в"O:�;'.�$=�
y�S�-��ǩ�yb�Q�uR �d�1#�f�#Fn֚�y�%�X���@�5!۾�����y�-�M��zD$�H��aBf���yB�޹>ւ�b�_>�\U�V��y/�C��1�
3;B�i$�\��y�}�X��p/'��I�Ӫ��y�Z�tȺq�+�*~�̩�	��y��;(��Hk� �9tQΕ3��L1�y�F��TT�$�߹<�Y�W Ĵ�y���w��Q�H�+8�6N 2q!�R=SJ��@�GuD]�a��9�!��<&J� :�-�T�p$b���{�!��E��D���Y�݂��)�:�!� �I�Lh��=,�T(���S�!���lhs'R�(�
XCuG���!�d�i����V�f����&Y
(�!�I�-�$�3�f��X�T�r��[	�!�˼p.���d�q����~�!�D�6	uѣ�`��
1)�{q!�d�E�hE,�c[� ����nA!�Σw��8dF��UK���F��z�!�ݬH����.IA2d���Y�'x!�D�30�� �=VU¤CQ=/!�$��RQ~���V�H���q�O��!��˄w�ب��Č	V�=��m(�!�$ޘ#�0���'�Yr,�5�Q2�!��_�ϸ3���9J�J}���\�,�!�$��=�5i��s��s���!�d�@��mB$�	 kd=;íHn�!��t��Ixd��OLL����C�J�!��#z��bQgƒfx�8֪�=t!�D٘aC��`�m0!�_�7f!�$�<T��dy#�ݠE"ؤ �U�EK!�,�V�Y%n�0.{��ۢ�ŜO�!�DڸY��Q#�� n@�ꀉ&!�$�? h�R���D��85�ӕTg!���;~nV� H�`��9���QD*!�DR�(�D�� 4H� \�6,�
!�ą�y	�}�F�Dj��@"�m�!�D�(P�X����@�s"lE`�!�dҩ����B�%9�
��B��j�!��V�
�h��%���A���!�\��y�V:=�<,*�RZ!���C���c+��C�� �d��!��5#>�چ��[��y��̝�?�!��N AR������	R�����$j�!�dA5gS&�S1�	�ءb�F'P�!��R�x�bUDƈj��̃� R�!�d\cGބ��kR�t	ݚ�!򄏵3:n���L �)�E+n�!�φ
[*@;�#�%�hQc��7�!�F�OHF�j��!C
��𤊐�A�!�Z7v�����CE��i��.�!�T/a�ZakN��KJ��!i9P�!�D3N�٪���^��#�04}!�DջEXVYA���D���fͅ!�� TAIӡ���\	���˧Df��I!"O�a��a@7�}pS�߹ngH��5"O�g��)M���
qHEPf��$"O�D�Tg6e��,��"VW^�0�'�ez��T3�ՇV0O� 
�'�ޔ{��O�#��:�Ї TI�	�'	� �0�� TaɈg.��:E`�'�ȱf�(G-�-@P��0���'R��	��'�R�A�M�t�P��'6lh��͌x���0�_:x�6`"�'���#A.&�r����	����'7�P�R&L�_ �K�#N }B"���'ф�9i�
�l����xH4z�'k4�b0�ۜ����ҙhm��
�'z�Z��Q��tZ`$Z��x��'"�T�#H�]6ȥ�פ�;)aFE�'ހ�JU�D�ҨXw��kx	��'p���߼-+�|#�G�/L��(��o�@�V��2v�ŲQ	����G�	���� 0D�ucůK�\��]D"M�B鉀-��p�(ҖE�ȓ
]Zaj??|8X@4��'c�($�ȓ)�.�r��ƃ~������֣d��̈́�*��Eل%��apX�����yV�͇�\H���1k��Q��)�)��HԼ���1!�h��wg	vG��ȓ��l�PM��~���f�,t+Nɇ�1������O�v���ƈ1M�f�ȓ�=��,��]��d����5j��ȓrRTd���X�r��C �00IBt�ȓDr�	Ջݎ-L�˒�c}�����+O 4�qq%G�]'E�ȓ%��\Q��.��]��/ǈP�lI�ȓ=��dQ#JB�yWm��#�ZЄ�a���rA ��l�����`��ȓ�H�
1�I�YR!��j�.�`��_!pq0��D�E$����bD�^�@|�ȓ#�:�� @�?�   ;  =  �  f   �+  �7  C  �M  .V  �b  �m  !t  �z  �  '�  i�  ��  �  /�  o�  ��  ��  6�  y�  ��  ��  ?�  ��  ��  B�  w�  p � g ( c1 A8 �> �D �F  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P���Gz2�~BW�I68�A��b���l�G�r�<�#%��B�n�p��w������f�'�axR�W�T�d�A��:.�~Pq����yҭ܌k����b"�]3�	Х#D���ę�=(�aEQ${}:���K�6$�!�0K9 ��΃/ \�hӷK��Ց����	�2�����qRa��+�%^�OVi̓����Og(�X��ĻhΘ�٤kʝ@�'_��B�1)�ѱ�脙o�s�4��'߂1�'��Io~rƞ�9�h�J��	INP�F�Ț�y�6JP@dȠ�Y�QC�CC�/�~2�DN8����?s��mC�͍~8t�*�%K2���#��G�ư�c)��6P��H�e��7m#�S��M�c�M2q�xl�#n��l���G�|ܓ�hO�O�N��ܐG��	��58�X@����xr�~��z7�(�A�����=�0`)�䝦v�ZH10���.pRF�WD!�$�2yh��a �<lxE�7dB�
qO$�d/�)��ٽ+.���K�^gθ�Ec4Gw�{B�8�$;- ሧ˕�d_ ؘ���!��Q�L�y!�ʄ*U�=e@V%:u��	%s��M~��� |<�t��  �Z5���m�"O H�%*z��j$l��R����P�x�Jt����
Y�i!P�����?#�T9(��-�Ov4`�i ~�R��Z:4�*\�KEI�\��'O2�3��S &�̙����:a>a�	�'��$��G`� p�e��eH�q�	�' �$�.���;5���]��s	�'��t�����<F�AC
�S�RDh�'ј�btG5[��M0&�O�|���ј'xو��Mx�X�k��5�\5R
�'���h�&��2��D�+qF��6�Df��?�'c�-�]ɞ���yxT@���,D�����ּ�U���V1*��E��<)��I˷�yŸ�V�5����V�#�IY	.ޒyr���e 	�ȓg6��3�ޤe�� W�?�̑�=9��������;[N���*ޑ�i�iX��y��";\:aKs)��\���#�(��d)�D0O<(0���1 ������9<P�{6�'�	��H��"��#��RsR�n�q���8��r6U�dyx�����K�nx��GzrF:?���̲Oa&�9 H^�%+Z�� �K �y�-T#�j��F�2(vh�S�l] �~b��oZb��ħ$?^d� k��7r � �$B�^��'D�x"�'Û��'�
%�ţS!qb����@u2���<���<�|�g�>)&��M�Y��W�Mv%�e�W�'��V��'>�z�#�d��h"�#�S^*�{!(���Ʃ�q��@�Y�r��)y���	 UQ�'��O���& J8%�2|����x,H���'m�˶�׿l���A!.��ށ��4��D1��?}�(�'f\j##
��Z�1�֊�x��'�>d���=3��a��`s�{b�g�f��>%?�*�nK�d�I��Ϝq�6�S�6�O�ʓH��u  ���q	%�4Q�%E��Kr]��35��#k�/|B�I&]�L��$醣-�p(�@-ɻ5޺��u����0��p�� B"�1_��(x'�'4��p�)�{�Hq#���_?ܤ����b� H�'��%I��+�����UC����Dš���>��q�E�[��u�-c�ȼ�"O��q�-�- pZy0sZK�|��e"O�B`Z2]ԭ���9Q+&�Q���,�S�.Ūу����p����V<d TC�I�#",�`�ݖ3��%Y¨�30z#<�G�'���i6�_�^6ҝʕn0�<!��'R��',�F���c�$ɍ6�Q�/5ʓ�hO�IŬjQ�$c���Z4#��j�џt��e�Oa��c@&ύ+�"� ��M�ܸ����hO?1��X�"D�DJ�'TY����l�<�Uc�0"��`� �"><t�t�^f�<���|�9X�E�,������_�<��-)����@��w�b�5̘[�<�Š���,�(�<rלYs��YX�Lp��dRn��ŀEkϼgx`�k���-Y!��12>�7nޖ1"��zta�4�'aa|�%K���`&ǁ�w�`���4�y�H�Ne�)�`A����pG��y��ǉ!p@�v�؍��[7a���'"=%>���Nԙ!�ZE����Mcd��D�:D��B΄�a@䀙���Jb����(O��}��g|���Ԧ�������Q�?�p��u�ޜ���]/u��eq�	�}i&)�	a<	���7>��?˴�TG�_�<�ծDTF���F�\�Y��[�<� ^T ��6$j�"��?m�(xp"O<��t��!A� 	��@c©�T����3S��q��*��!A�i�/7"�B�I�u�,#vC�A2Q�C�TB䉧	Pq���?"|��"A�j��C�I;_a6���J��{��x���]?eְc��F{J|��N�M���B$�˗N��MF' ~�<y��b���b@폓,q�q��W�'r�q��I�fP�hʑꆗ>��3�̡n�B�ɐ`�����dՇY��l�1������y�\��$
=�!F ��Eh��W�Կ�a{���Z��1@$���dV�A�TOBr�!��6Q�<�q"݄�v4)��K�!�d_;�p�������3�,F-�!��%w�dh� (Ƽ9��ԃPkЬ^���hO�ʽy&A�'��\P��M%�.�f"O�#��\ʢ�G8/��d9e�iF��N8�4� ƙ&n�l��D����,�1,�O ��ʹ p��+DT̐',ʗY���1�O��Ms�'�z|*�!Ps~(3u�XG�Q���$(���2��Oo�05k�P�ցYc��+\��j
�'�.y���ń�t����qT^\l�t�I;\2�)��2�ǝ?x���*6Fi�Ԫ D�@���ܜ9��\�����TK���e>}�'Q�{��2\��}1��$wH��b���D؜W�Ac�aN�M]�ȚDcR��PyPx��ʃ�V���a,_���Of�~$��"T���̖,FR�)�w�<y�l8������('�1��͇v�<����h$�4�*=��1sGYt�<i�K�# ����m?v
��nq�<FFΔz4���c���a�	An�<��%�'u�a�!L�&	��1r�j�<�A���a��B��OV@z��pc[e�<�1�-FQf�y��Ac��ѐ#�e�<S��yv�Z��]�z� s	F�<I#E�(Ey�`ݝ#�^U`�W�<��!s��L8�v=
�+A.�K�<�Ũ]��\m#���"��a�TFPS�<pD3��3��G����I�<)��D![�ZH�4�D�Т�Ν~�<�����M�$C-�	�xru�x�<Q��,�  eB�U;� fw�<��Z'*�8ڀ�H (�n��wDY�<	���L��L��(N�o��л��P�<��&�M� ���@�{��	�"`D�<�d �t�pa!�U�>K�QS&�~�<� I�M=X�(���@EΡy�o t�<�"��6x�͈�ɛ�k})-�i�<��d�$;��d��(��eR,1#bb�<�+���=P��/Z�R�H��K\�<�@	T%e.��I+@�IP�, A�<A�P2W�\�KƎ_����T�<y*˲�}r���}��$��I�U�<Q�
P�e5��Yb,׎6���I�/\T�<ѣ#-V9Д�G�p��`���	x�<����;]y������4n>�xg�s�<�ˁB
`�ӢjA�B��a��]Y�<av�*J@zQ��\(�x���UV�<)$�j��*16i�0D�R�<�4��m�l��7����h L�J�<i�l�,m�p�i��H6�ĭڲ�OJ�<��94l�(@�?�P�Z�E�<�ɂH`�1�۔)$"Y��[E�<� xEA㌉%tB����߼}�g"OBi���F7T��	��5�ʨ��"O"��L/iwx̺��A�ب"�"O.��/Ԗ1SJ�!E钻;�Lp�e"O���H�$h-������"q�<D���'���'o��'|�'���'���'�l ��W�}Z܈� >��{��'�B�'��'3"�'Gb�'���'�x�#�m˟o���$�I"H۾�c��'��'Y�'r�'b�'�B�'�^!��g�K�Ɖb��#������'R�'K�'S�'�r�'�b�'D�M�+A���X���/��p�'���'CB�'%��'���'���'��M˲�5�.͓�%�*3�6e���'��'�'�B�'���'���'*�Hv`��b� ������$(��'�"�'���'4��'3"�'[��'����	X;��j�$�=�xMx��'6R�'��'�R�'ir�'�b�'���B3Eߴ��	ѪD: ��ҁ�'T��'T��'R�'��'���'��B�'Z$EӶ�B�"t�Q*��'~R�'*2�'%r�'(R�'�r�'�^���r-����l5�њ0�'Ab�'�'�B�'���'?��'Ob����C2r]8�9ⅈmD�g�'�'Eb�'��'K��'	��'���,@X�A��cƼ,VDڤ�'�R�'A2�'�R�'�RHf�,�d�O�h� Oܮ9r:��L�,�Ո��VyB�'��)�3?� �iMV\� B�Sa�y �>,]��g����A��1�?��<饲i*�k��͍Cn�mh6�M�/&�����b�^�$E�%툽	A��xs	�j�C�~���ٓC5`u��L��RD,��f�v��?�(O�}�FoG#q:�y�m�W[�1��e��J��& 0��'���Plz�A�D'ws�	q�葚�z]@Bc�M���iW��>�|�M�Ih��.=�1�d�"ј1�O�+eKn%͓[f^��l�&�Z��4�����S��!;GNܨ@WR�#W	�FI�ļ<AI>�i�Fq��y�rE]y'�UA� �R-C�a���?i�X�\rߴW��V=O�h�Nx��*S Ji*���85�9�'��ԠAAYi'd�*����U!h�+�'�m�U�Ȍa[�Ā���Y�X��%^�h�'���9Oܕi&�%)rb�����(� 9O��lZ�CQX�m(���4��I��z��I���i�]�7O�$oڀ�M���NL�6AP]~�ϋ�K�(
0��4?�ֱ�&�
b�X��I%qX��H��i>͔'��Oш �Ӂş�^,�cf=kD���OP�m����c���z�&�m[���a[�%lTk�'�m'�	�M[Զi��$�ퟬ��-j�=H�̐~��G$�RX�7N���>"�x�r���M��1v�>����T�҅�Q:�MXCʷ@5��՟�'��IU�&�M��M�<gi��>JQ�&�yc���b��<I�i�"�|��y"Cl�l�lZ��LJ���/CE�ubs*�?{����Z#�\M:T�}�\�'!�"L���[.@����@�xwm��[�_���(�[5a�cЏ[�<����<E�d���[2,)I+�$qT�aA/��ݘ'7-X�-��I!�M�����٧)��R�]�S�k!l�����IP}�$x��=l�� �3oQ0����������D�waR���n� d��i�T��"!�:e(�&
�=��F{�O[�	Ɵر�c 8'E�e�7(�&1.2-Q��r��'�<�4#���<Q*�Ի@2��@*$���0@i�4�����dW�=#�4�yb����O
��j�79p��FB�H��Ia��� Q��-��Q���$⟲1⑧��|�0�U�<��p���� �!6Oz|�Q�~8�
 �#�"�2&Ţ���G��
$V�S��7�����JP2�˃D=r�.\�Ī\4j��F�3bq�xk�F<Y�\h�DAU.qr�s1��b���'�~\�Cز0x�yK���%�L��	�=`�ssMؓ9�x��l�9>������99˼M9c��	��,Bp�$U�a2�KՉ���8 ��7f��x(&m������#�4v�Ç���t�^��aM��%j<c���(J�V����˕'�a:��	-(w�q[cA\C��鲡�( 1X��L�#m�%+L<y��?Y������O����|j4`j��Z��\����Q�hQ �#���O���O��$Ѱ}@���56.�8[K�A�6(�h;<%�o���d�O��d�Ot��?!��Q�ܰ�O��%��'A0~��Q�RI��yĨ�C�O����O��D�<�4��?^Y�O� ���oU��t����v��HƠc�r�$�Ot˓�?��� �x�~�V��8&'Y9�h_,|�ح��������I��'+�R�<���O~����D
'D�?$L��Y4*�e���҄�i���(����H#|��禩��G�._%�es�-0G4�Ekw���SNv2��i�v�'�?��'��I�k6�5�F��2����V��% L7��O���?7�H�S�����^ߴXQLP;cPf��`�K5�>,n�tX�Qqߴ�?���?��'^퉧�ǂ�J4�카f�6���V�W�7M������?Q���<�BtxcG��+J�&��NR>E
��ѱi�R�'�⩟�<O���O���9L�yD�}ܞ��)ÆW�TI�')��'EڹY�yB�'w"�''�`��ˑ�	w��"e��V����ct�x�d�.f���$��ȟ���gy��Q8j�l��$������L�:�B�'�Z��y��'���'��I�d4dy�C�f�;��pj�)󤗽�ē�?)��?	+O����O��� e��A���lPcܡ{�� ��%h��?���?A(OB��plS�|·��(��	czĪ�Jz}��'�|�X�Hh��>� D��g昘k #Da��4!	�M}r�'R�'!�	�vz$�H|2 d���;4M��d��0#"�7J���'��\����ӟ��w#>�2ARh�؆�h�B�Si�~��7��O��$�<�bV#]��O�r��5�@	(,�S3.C�B�]R�)R�����$�C>���dlX��UD,i:Z�1a��)��nZky2EQ�4�&6��l��'G�t"?��m޴HT�w/�{#@����M��ɗ'����O��h�sӢ� i�n��eْ>��<�&�i~�{`G~�����O��D�<�'��ӊ@�0<IGh8s��\u�)yD0d��4<��T
/ON��O���D�O���� �5����fM�<��؋1	���������I�J8!L<�'�?Q��<6����Οb�Z���Ε�v�dEQ��	����2���0�����c'��h/��ۅ��<��-X�N��M��rD�@���x�O��'
�Ɏh�
|�H�@�虲+�f6�A��4�?��C`��?���$�OV����<j)�T�D�C��J�(��N��?)��?���'�mxq�\�],�+��%����� $2X �Oj���O ��?qW«���&��"�WPW@"cc �<�M{��?a����'m��'�E��4n��qUj��F�j�J�J�y����'�2�'��	���CD�m��O�}b�Bw�������A��ļi ��$�<aBO�c�	B��E��! ���#u��V�J6��O��?�� V�����O��������Ur�r ���A�;n
�C�P���䊭T��#T��P�4"��H�c��WmR��?9DcU��?����?���b)O�.�VZ���G��vZ�Jv/W(��Vyb��O�O���[�`0Ѣ��p,vEݴU+�����?���?y�'��4� �č�-m&�8 D�$����eJ�|�lm�'��ڊ��)�OF�sMS�����Gq@�Bt	����IcyB_<L��i>Q�I����uM&�K֏]-8��F��'��� �	�ħ�?���~�ˮPI.�Z�o�ghܢ�`W��M�����p�+O(�D�O��D-�	�/4� �lJ�T���@��Rqt�i���÷�{~��'��]���	&^�Ȇ�f�A�������R
�Ny��'f��'+�O���U�C{�d�1ωP�"=�R��n��x�WG�eL�	����by�'�Ԑ��֟��at��[��Q�JI�k�A�i�B�'+r�D�O�����+����K'*zr
G͐�L6@h�#K�����O��<���^��$�)�H��"�*͸���,ԒZ�V�~�n��p�?���TX����{�ɭCF(� �G�n���A'Pjv7��Ovʓ�?��������O���䟬P�A�١��h���4��5��t��?1u���x�M�<�O�\�B�#j��׏�j�D䐔ɥ>i��V�i����?����?������"�XFF�
c�\�U�M�
8:-¶[���C8N�;&�.�)��Y�F|����8&�a���`�7ZS9���O���O��	�<�'�?)5"ԝ]�2���G�q�<��IU ���v�
��y����O�;��ܛ@�^ ����4AD�b0B7��OL���O�Q��,�<ͧ�?����~��&D�A2�7��P�P��@b�D;���'�?Q��~�$��Q�x�#��J�SM��KC�Q��M���]זm�.O����O��8lE�Ad�D���䉒 k��tN=�u �K~��'��X���I�k���N�7x�Y'�P�p���Quy"�'y�'��O ��N�Kq��%�	��p�$-|���ϸA��	͟0�IPyb�'Et���۟p�J#��l�A�f`�1L^=Cúi���'�"���O���E�Ҕ#^��`��Px�9�K�&xw虃!����D�Ot�D�<��yv��,���D_�V�h
d���NL��j���P榹�	}���?�EI�,��E%�|�7iF�i5<��p�ȩj��x���fӐ�$�<i�e8��,��d�O��i�!:��1��U,'�Z�^�$�>��.!nT���S�D��-�z�ɴ͆�c��Y��Q��d�O���-�O���O������ӺST,��=z�Csa�>k<�bB\}B�'A���n@�O⠽���2N���%&K*u{|���4Z�D���?��?����4�X�$x���ʷ��(��X�.��#��3�4�:�8���o�S�O��)_�bC�)��lZ���԰���m�6m�O����O��E�<ͧ�?I���~"#A`�hff�,|�K����c͜c����oV.�ħ�?����~�b�ƀPƚ	�h�`�����F?�ʓ�?����?Q�{��@29/z����xt<q�kK���Č�}��= T�����ޟ�'�R��>~0x�W�[w� I�H%C/�D��V�d���8��_���?�c-B_I��c	G�N����$d�-[�`�bkSO~r�'��P�p�	; �r����@Y�� (\��e�c��mZ�0��ٟ��?1��wLZ]�sH�������m����(p��0lh����?y����d�O8T3�ν|��m���Qg��k����$�e�{#�i_r���OJE�r Q-���� �cF���Pt�DcѸЈ<
��i��W���>}��5�O�2�'��č�a_2�+
��}��eQ0.�>Yx:c���	�8��2@/�~b'A1,�1C�g�����~}b�'5��
4�'�P����dyZwlL�S�F�5�l���bBqLz�J�O���`tu�%����!�εr$h��-#fX����z���$Q�b�'�2�'q��\����@8���ъ!�_Z�\aQ��M+����<E���'�b�8/�3{V��)[�,���`}�H�D�O|��<��|����?q�'JޙSG��.�6�Z��8��,�P"�	�d��� O|z��?�'28���X|�x.y�.̊ׯ]��I���<�'�r�'���ě	+�f�Y��B#�D��)Fl���(�"���%?���?�-O��D�����x\��Ғ��-����)�<Y���?i����'�"�"���P����}�|�r/o��#(�?>���'�B�'a�U��������D
�/Wp�݀`k�[�*=8p�D7����Or��#���Op�[3,f����+Y�!wc�
���Cʇ:}�n������l��_y��J�c@7��O���2@h�x�B�4iƩZ7��00�@Xl�Ο�������';��S��d�'!��X���I�R���h�zfk�nl�v�'u�'�m�57M�OR���O�靣'���¡�/1�v�c2�ޡd��Em�ߟ��'��
����|��Ms E06�U�f��'Ҡ����ͦ��⟔X���#�M���?�����'�?�L�h�a1D�C�!�ĥ+�g5�����0�����	ty�O��U���A!�j8�8��N�F�o��6�Z�4�?a���?��'����?��Zt����Țf�~y�aC�v�A�iy����'�RS��Ss���<z�ċ�<-��GK>x�>q0kV�M;��?���	ql�J5�i���'�"�'�Zw���d�
4��IRWD�m���y۴�?���6t��G�E�<�O��4�'X��oC��cf$��!�P�U:(O�6m�Oj��������I��	՟<ٮ�����b
( N@��xa��e�*1�y
����?����?����'+z �醇W9&$jU��J,�x�g�R�{���'��'�Rc�~�(O$�$X 0�D���K�V��]8Ü4'k�u0B=O����O��d�O~���O��DZ�edxlڃ����q�*IG�A0�T�7��y��4�?	���?i���?Y-O����!��U�}�|���D",F��yt��/H;.tm�ϟt����������	��nI*�m�џx��>T[�� b��Q�L_+��#�4�?1��?�/Oj���	`j�I�O��	(?>8[SkA�m͒h�U(��g�t6��O���O��V�q�ql��	㟈�ӂ��1��aۿ`XD ۄ��4 ���޴�?(O��D�3+��I�O���|n�6*`��s��L0_e�yKc�\A�B6-�O���-f�o������џ��S�?��ɧ,����F�ީ�^4� o���#�OL��ײ x���3��3S\i�ӎ�1� �A�l�]ڛ,у*��7m�O��$�O�������Ov��I%�-�b�3�I�0x��n�)2��	ݟ���������'����}���*%��F���j�B���O���7tZ0Tm�d�	ԟ��	�]�bplm�'!�G:���N[�6M.���/=��?���ퟤ�I[4���Ŏ]*���IG�m�(\�4�?i�b�㛆�'��',ra�~��'w:�@�c̉z�������f��Q�O� �P>O����O:���O����|�p?�<p;V՚Wк��k'?3�c6�i���'���'�&�'����O��z�CCj2TA���3/*t�z �U�D�O���OL��O6�'3r��p�ij���spf\H2��5HU��-k���D�Od�d�O����<���f����1ST �M�u)�LX��b�t����O(���O ��OyTaSC"x���O :V��}L�-a��l�a�C@��%�I����Ly��'�JH�O;��'7J����^�J�s�@W�E�L��q�
�02�'��'�Ir��w�����O.����B��Cn�1�l�vD�.l�b�uD�Цi�	ey�'��<�O�ɧ��4��T�G y�2�����9nZ۟��	%m�H-��4�?)��?������I���ap��PEp��(�- ���X���ɝ;.^l�?�g�ɾ}G����_��fAv��6M�)=zz�oϟx�I�x�S�?��	��P�ɟl$�ɡ��4̊n���q�%E}W�fe��4��|�O�O��$G�mХ�@%CS�A����526m�O�d�O>YB�Ʀ�����H��ߟ��i�@��6@!��O�@E�2+b�p�O��a4O�S��������@UA�6A�]Y�Ê�9w�xQ���(�Ms���~e��i_B�'G"�'����~���NpIiw��7�f�3�߬�Mc7ݑ�x�ϓ�?���:���?���?91�@3p��$���3F�$kDÓ�	�@�i���'��'(����O4�����mE�e8�`_�r�`'���x��<���?9���?���~]��(кi��x G�R�_����c���`�J��s�d���O���O����<��:� �'e��$KW��_��P9���.n�5p��i�r�'�B�'/��'��i��FaӺ���O�U���;JN���l��6�%�Ǧ���͟��Fyb�'�,��4\���~�PS4�wn�� E�v��)l���L��͟L�I�:y�!޴�?����?��'\�� P.&" SDc�]�h��i2[���I4��l�i>7���Q$��C�FǐW*���/Icʛ&Z�X�"����M�\?����?i��O��R��/:��y��P�4�:0��ik��'����'��'q�� xLzM� �|�##��*:�кӻiVZ�aS�v�P���O��D�:��>YM@�I����&hN�~��{�F˛f��3^���|"�	�O9JW�"#
���?��p!�Eئ��	��$�I�?SZQK<q��?!�'�������i���X0���ڴ��1K�\�S���'#�'���;�F�0�=82탍\�"Q)'F}�����'9HVp�>i���d�Ok�*)͒X��.PFE���^�e��ɐu7��Ilyr�'k"�'�剛XۚeqQ(|���Z�JU�&�l�3eJX����?������?���p8p͚��X�mR(+��A�`L�Ѱ�+��<�(O����OB�d�<����?���-�X�Jҫ��%���n߿B��ҟ��I|�ҟ��	9&x��	�R�$4CE�-AT�1r�T;m}"ˬO`���Ot�ĸ<W�<2m�O�Pi	�I�_k �۱E�j�N=ɰGc���d/�D�O��Q+2_�$3}��Y�{`��07k�"?��R��Z��M����?Q,OnhK�}���S�{߂p� �"�J(Z���v8�M<Y���?Ʉ⁽�?�L>�OTʽ3U��1 lp򠗌"��b�4��X.E�m�2����O���NQ~B�ҝM�����XوVoI7�)o�ݟD��:�!�?�~R�A8Ag�� I2�=(����Q�p �.�M����?9���xR�'	©"��tD Ԙ�ʋ,I�AzT�pӀG��OZ�O>	�I%8����&�$5���R  �6o�5�۴�?���?��I]�zr�'#��'���\G/�\��LR�tmLZ7gC����|R��!�������O����%��x1h�Q�YI��$?h,�oZܟ<KvB�����?q������sOΚ&޵�CM�3 ����s}��.i�2Q���ߟ$��Dy⋏<^"����">�f��G�W ;�pٸcK"��Oȣ=)�w��Ð�8V�����;H�6d�f�X'�?�,OJ��O<��<���5��9c�tt�V�	u���(�n����HE{2�'A�Q(�'4�`��4��0�ΰr�t{D&q�l���O�d�O����O��r�c�|��Z�ʝJ/� !����\\�P�i(�|��')�"	$=��l�M<A�ٱsUN���C��kA��	%�Dܦ���ϟ�'����F��~J��?��'v�<�P��
�s����d�	CR���iK�Ozܚ��)�	�?�ؼEB�����~|q�pc?�67��O��d/.�d�O��d�O.���O��ƢH�e�K4WXr�¡��|�$���i���' �"e��=����O��q۵ ��p�D�@"��T�E�ݴ�y���?y(O����<)(O$�����hi�hUk�4��r�O�Ʀq{�P�S�O�n�%U�M�ƫ��mJ;�S�b�6m�Oz���O@���W�	۟ ��A?i��V�Uh"�auf�!Afd�Z�bb�H�7<�Iџ��IƟ���@�o� �i�=^DI;"���M��>k:�#��x��'B�|Zc8��A���s3%Aa���Oj|����O�$�O�ʓ�v�zE��w�]���أ	v�R��+�':��'G�';�Wbfm�fg� p���k�C��Ptn5J��5�	��Iڟ�'���UFy>����Г#���a��%v<J@�>���?iH>�-O�<(�U�����	7"�!1��(ޒ��!O�>a���?Q�����G�e)�&>�!��*&=6E����=+�$uP���MS�����p<��1DYl�5Cٸc3�u��NK¦9�	ϟ,�'$��{��8��O`���Z�둩Ѫ/��a�ĹO ���M�)On���O��d��O���i���零b!�aDP�@,�޴�����6lZ���)�O��i�@~2N=kȤahwa���||��JV5�M����?����4�6�<Qdc�2:x�@�V�ڕi��]�Ə��=����� �*q
^.v�:\h�4;��=qsFťu�� ����U��2&�^�<���g<$㷈��\�ɻ��
`}V�X�G@5p���� g��]L����kOl��6���d�){�tU`('&	 ��Q҃%�<X�(����Dv�P�k"3Lz�#�!VDa酄̮��Ic�fӱB�VL�U��P^��Q$�X��R&��k�5#�I�FLa���.�?A��?��Y��O��D`>YqvgW3!�ֵ�2j[.'�@M8�U*��Nч9�h9s�(��԰<Q��>tM�L�h��hU"�K��V	JԌ(�Ԧ��Ҵ1U��'D@ay�M�q��S⎁=T@�)& H��2�x�Ȧ��ڴ�?q-O\�2��$0��[�"4������� Sm>B�ɗ�T⡈:_�@j���M�>b�0����˟<�'��5�3f�~��L�́�]�'S�T9� �g�@ ��?�Ђ��?����g�>A��)d�D�Qj0��&�*�48�+E�i@���C,^�H,����i׌|DyB�D^,P� *�=Ί�X3�F/4��Rg�qS�B�.�B���epxEyr���?��i���kszh��g8X��d1���,����<�����<A�%�
yv�k@���s�́g<�T�i1�����	`2` ���@T���'��ɷH�Z�O����|�BdȔ�?�w`]�?����`�E�El��va�.�?��� ��7���Xq��Kd��8�1
(���'9�����:	����viH�}�4L�OJ�(r_�@����p��w_l�S$a!���Iݞ��~4�<`Pk�B
F�C�d�1U{j�'��0��?q����O� TuÆ� ��aY���u�i�"O�ҹ3~Л�iH76YlA'1��|z��9Y�e��F]�>�.���5x�NU��4�?����?�TM
2=lC���?9��?�;X�fTUf�t��08"���|��!&�'g>�p�Ɏ�����7P��X8[�`@�j� s��	`#��xR!��)�x���H��Q�g�I�/e�`�
�V�ly1��R��D~B��?ͧ�hO|�8�"U�s"��3V�F����PA�<	E�ۜ#�\����r�<ؒ�h~28��|"����ā�)a����0J���a� ��b�#TXp^���O�d�O��;�?�����n	"x�����AZ�N�+-�hM�ӄ�8�:�c�\��q�	Ó(��k�>�l{�g��[��[T��fU�2�/W�1��e�a���6�תq9��s�H�N�qAƗ'�>�d�O6�=��"=>������;Xh��&��yrJW����u�Z�8e,Bq$]�ǘ'��7��O~��>0��_?Y�I�8��p��F7[�PG�v�|�	ß��w��ğL���|D�ZK	��aD	��1>D��*��-� <�1��7lfZ�Q��ܞQ�������n"l�BШ��<;�#�Nd���p@�52H%p ��=;�,(��C��O��	@�'G2S��i�F�#2M"��w�*n��D���&�	j����֌Bm�H���\GG�('�7�+ٴ'L<�6�ǁqJ=c��asRi�����d\r1��mşl��u��MB�kI�k鸽�3�G�aE�����9���'c�0���!0J���O��{�fuJ @�~�*�t�� mĤA#��PF$�@��Ü>as�Dl����p �{����J���O����ɀ�v�
�:�#ӭĊ@�M�ju��O<�d)�I'�i�:h��0�F�: ���A_��1O��D<<O8�����C�9�I�^��#�'(#=f��>>T����<�D}�v�M�j����'
�'2HT0T�?{�"�'~"�'�7b��;��ᪧJB�_e9��/=$M�y (�5H��PkfAV+7�:`B#��:�D_ jt���A2�T����(�*���Él~�-��-K�M�4A�!�	<�D΀v�����H]�}�� %�H�v�� l�����P(QE�O@�$���=:^���&ͽkc�M:%��2P�!�$ʍ'��,H�� �hUX=�F-/��I��HO�lZ�4�'�e��-Ѿ����b�̥ft�ja��g��-0�'!R�'�Bqݽ�	˟��'Vz���K�!��r����Oa �@K[���z`�0A��TjWR�F�r$�M2�F��}`�ϵuX�`�UF�A(�rbJ\57It�j��F�j ���R�Ҳ��r��+ʓ4)���2�X"(,U���c	&�����Ę�4\�v��W�|'���2��@ezQh��V����2, A�Ǩ��8��Q<�]�<a�i��P�\j��8�M���?�e� �j^��IbAI6N�� *�ځ�?)��vsJP���?i�OfP4��.sԪ�Q�׉bC� �u�Ʊ� �{cJV�Kâp"�ޘo	�"?1�&C�G���\b3cUOY8C֊�P�Ri����Fæp����2V|���Op���O�$��.
"+Eb���UN`F�3u�<9��������"�a��]b䢁��+RT�%O!mZ>5����M�L�����Ǐ'�����}yLۗ+���OO"W>�1���B!̓�����K�t��I	�(�	7�\(*$-E�]�4�K�)'��9��G$@���Od��!�%� ԶbaW2"�x�I� 0�%	�,D���%�l��EG��uM�DӢ�?Mb����ծ���Y[�U�~*�G:�	؟lE�d�'"H�#��2`s�I��,%k����OJm���T��Px�FT�>T&��'X�#=�WeV!|����bE��!� �~M���'5��'�| �Q%7D���'���'���pt���}@������>.���k!#�jB(���Y�rp�s�Fe�g�	�mYx��Vㄼa�H���L�RT`�ڷaZ6oY�p���_�8)4 :�3�$ͧo�5PL��q4�p�n¡p�ran��M[��<(��#�S�gy�'��Qc�K:���"� ���ONi���̷sY>��AA+Y�������{��D�4f�d�<I`�4i�Aۚ7�XLAU�LI����?���?�����ݟ(�'gfbH
�e=?��isp��	d�І'8BX�U��n�/6�pMA�&S��O�� eJ͐B��|"�Lc�� �'+�6 �����F��] E���B�Fh�A����(O��	6@�����BI��sn�<	���'"��'����<�?�2��v����Rb��e�R���k�<y��>}{`EXd�ƒ=�+�K^̓J�F�'8�		rjB$Rߴ�?i��v[�j��#Y�p4��U�g��U����?1�	�?�����Iθ�������Q�nU�ųi�.���K^:$"��a���ȝ�ǓX���WbC�5h�|Rd�B 8��=�7n�!S�,�CO�襸5��M��E|$J�?a����k���W�Q 24���Wmy����O�$(�)�g�? ����W�BO<���O�,V����Olګ,�b ��@:ƚ4�׌�fO��	|yB�	���7�O���|B1��?I�aL hq�a�VZf!�w��?���)�����f�"J�ޤ�i�(��3U>՗O���q��*v�D:E�1X�>P�I�H�'Q$r����peM9b�C�IR�~�
M:U�?e��z���B�r�HI?}�o�(�?������\ڝ ��h%�dT!$��`�<����<�D�A�D~0 e!m��09A��hO��y�'b@Ey&��8۞Ձ��62wR���&tӮ���Ox�D��F�,A�!��O��D�Ot�4�D���=9�v�򁪟�	߄<҇�Ȗ�iM7&�8Q��닢J�b>�lڊq���ɬ3�6Z��̪L+w��'�q��i���>vd=[pLЂ9�fM�'�\1W�it���<�h�U�O-��-���C82��UH�J�Ʀ)�۴�?� ��5�?�}�'@2�ˢ�(�᭙  �����`�S��!ќ��eE���5���O�<Gz��O�Z����ED.Td:@�!��,0s� 1u���ߢ�� ǟp�I۟��	���)�O��_"nyG�S�� ��4Azlj$i�/H |�N��%��n#O�ś�
����"�P���V�6�1Ce��Jlm�i'"��L��<n���EɵZ78�Ol����6 �dX�&AF��Qq���dyra�
)l�蟘�';�����|����[�,�7C%�a||�`��?&�)�GG����QR���'ZL7��O�OИ&>���`�D��0ҊD�nB@��-0D�0��d��{��T�0�'���v0D�Ȳ���=�1Q4@�9�^�+V�3D�T�rj_	4tةa�ŗ�p�P}��1D������6���U;h05��0D�ء�-�2I��$hP�F�V~�� 3D�,�ҩ�&n�@;�z9���SF<D���kG��1��"C�$t~髧<D�L9W�ў	���#PF�l>��{�/D����iR�-d��1c^�[b�S�+D�٣[���d�t�ڰjR4��1 'D��)���'U�A�@�:�x� �$D���`ВwҞ��*J����ƈ=D��3��$O�m8�o�(X�a")&D�x6'�SrXt���B)>6�q��-$D�����V:>�
��6�S�r>��!N>D�,H�a�t��i��KA�lE1�?D�0ٷl���X����	OI.�JB�2D�p�c.0J`�)'
�=ZWT�y��/D��rP��|� 9a��םSk�x��1D��1f&O���h#�"�:c����.D�d"Qǅ�d�L1�(A9-)�1r�7D�X)�&�..�nI&�ߴ3#��&5D�(�_��������$m��8�5�%D��0�Z1��m��P5~�F."D����.אG��H�F��~Q���>D�L�!�AX�|���Xu��`b;D��؀k�lU�d�-��d��f-D��2q N ;
�#�m�( �j�4j+D�DR�#ʹFܸ�u��"x�Hȣ�*D� ���"��49��Ǣ6�:�R��(D��As'Q�}�8#��?j�4��P(&D�X�Ԉ�!W�l�!.Gx�41%D�th"
�$����'Aw
<:��!D��K3ñF�q��,F�0I�w�5D���H]24��a� �*�y #Y;
�$CW# 9��E��{$+�?�=�2E�@����c��"fRu��"Ys�3����UI�@��*̳nsDL9"��D�TQ0$(F�+N<�2OԴc<0��I-xȠ|�shE�yB���"N/6"<Q��զp�@�v���z��($'��ӥ0z*0�I�k���5�d!��ö(	�ɰg��k���Xeo��<m��ȟ�H�fX�R̮vh���3��[dcR�S�d
�.*�"��D*�X�<���U{<�Q��,=��B#�-qL�Z���U=(��+��l�RQͧ�Zѫ�(=�9�'��J�AI E�^�C��)k��[
�&oXI�,ϰ�T��g�<Y� ��-
�|�Aɣ�^�9���A�~X������|j�Ԛ/O��?� zQ��o�(yJ��8�Ae"���I�X!���kΪz����&�[�E�O���`�ͬ:�&EF❬��A@� �LV�	�72��	)�3�I�Sq�A�O HcR%��/of$:i �Z��%��.D�k����"iVb�O8��I��M��^(��d��&��J�k�d��8��'�LJ2�W<���j����e�jժq�фd�|��b��v8�i�G�^��~�2,^�^=󄝓1.ճ�����A+>��8��'��a�?�5��D*6��\�c�/CLP����1K�� �`��`�b(,5�X�#/�E[�S��'��8h�B?-WNRs���T��"<Q�H����s���>ڮ�(��H��iZ�G�Q�7F�)y�9+�h@f���y !>��ɠvLd�'5'D��TB~��B
�I�EK }�2���.�*[�.��4��4d ��'�/l����O����=& D��t�W>g�H0���+��aH�	gz�q�ő$}~�p���-g>4�2��"Fz K��^���p�KS.j� `�����OPiBw���$$�="aW�O�&����4az�#Ň>�zQɝw5@�eԓF��/S�f��XpM��	p!NFyB��n#��2�O���Ag�E�\ICm��-^5h�.�)��0���!�FP2=���=��(TDM�\�OT�ܑ�c�����)0T�xt��eh���R��^�Q Rš�E��I��2�N�
�� ��HT��x'E��3�~�㠡P�L��������3�D�:G��y�d\j|T���'g�IR$Bh�8
ʆ�ذ'K�cAR�)U$�}"�!Apb��rE��@���J	��/�nߤ(J	 �O	����|�"]�$�VMrލkwb	����LLx��#�O�bfʊ��֔C��\+���'-���P�CQ%ܕ�@�8i��`�O�(妜5) `�O�jq�'�4�У�#?�m�5��Y{��a��d�9{�H�%O�-�v8��c��򩗾%�>l�P�'��� ǡ�~Xx][r�ӆN,qԢ.2�ꃍǕ��O.!
��B�$��Q� �K��9�G��`�>��c
JX0A��#�3<t�S2[(p�	��л���UҲ̦��9� � 
8�|J��Im���������*��]�HѰC��oV��^bFp�wC�H��AP�3��ɋ��D��@�F��ws��e*C�PtvEi��f��B�0>�a�ևQ�f����	�$�v��'Y�Z�¹IP���������m�*H����I�:5t�q�X� ��ׅ?���KK�-p� �բ-� 3Z�C�	�O����.��`�0�`Ѐ�@��9&-6�	��p�չ� �s}��^�@=r��5F������HO� 
RKٖS,(l+էP.4�6���a�`5�L{A�Ӕ��@a�X��Dɶ�(m)ѯ@N?�X�M[q��:f4����k�\E�����UG@誧iV�o�X����"h�u�S�fv1���D)8)����#��]���A��d��ylH�7Ra+F̏�C(�A��X>�0>Ae "N�@@��Ьbz6`''��ȱ����h���',.�mڥW�d#�^390����'d�\�u]��4��	�i�^���f/y��u3]2��AT�	�q�!ڂ�:-����C�M��!?��#TF��B�G HJB��$Ʉ3>5R� ��
4�z��,L9�W+E-p�<R��gB���t�	w�(�"�aL�;�l�	���3㇒
bm^�F{b3�*���#0"����d/7��rU�i�peB,Ʋr�|"�4mN��DcI���C���V�nAq�'<�ě��8 :���v�΢|"E�O�*�R�r4�I�c752�;��%��"�s�F|r�փ��4s�w��8�P��r\^�dG�{��T�U먟����i~dX�'jHؘ���3G�^�C�W�a���oH]l���}r��R��rC.�yϰ\:���)1@����ŷB�rp��'��*Ը�� �D,SL\k�'��U'�4������¥]%8�b �f��&XE��s�*= ���P3eF'��l�Ql^w+��Ć�,u�fu1O��17"Dd�����5޴z1��]�I���� �M��}�Ofh��%P"(:��V�9ؠ�6��ْ=N�)���hrL�p�*+Z�,��<O�����c)���'P�3?�"�ȰyƔ`���$}�
�V#�@�e�(a�<�2��W�Z�%ړV��A�m�!P<�� ��{X1�WF��0�0�kp���	���ٜ�MKC��<���!"��HP�O���M��]K ȕ1p*�
�l8It	��d�!!����#`Te#n�&0�I-0����g.؃NJIz`mĢ�6�B�ʙ;}�X`���C�V
�t�c&ȣA��deԂDn&� G�H/Q�4aJ�� �dh�Ő�DP��E�d=�<C��B5��y	���)�4/Y�D�Ex��@7B��r�b� �M떁	��l=��fNMP aO�.��Ɍ��.(@-tcT=��Ѳ�M�q�$�o6n@��'��uȚC�Rѹ���;�Dq儙5*���G�Ǖf#P��D�ƈX�Ve�i�'&���u��(B��8S����_�>�ȲƓ�q�:aBNL��?��䃍l�<�	$ ���{���D.��2ƒ�u�*7ݟ:Y���d�XQphҮ}#.T���O�`&��g��]������y�?O�09�(@8�P�k�J�8 �D�@ ^*G�����2��C�F�<��n�?�i�B��|�DN
Q��D�;:,pC "$x�l0��� /OTc��� s�@���&�~����uG�֟9�QDW!9Ex(zCeY�\�z7¢4���h��-�	�N�{� -H'�-�I� ��x�/ԆlwKQI����ɯ~BL���@�P����U��݄���I���uJ4�|m�����}�LD�s�Y0 �> A���h����T�}'ў�z�K��֘���B ��/
i���c��q���'�(�#�kB�q� :��A#L)�ȉĈS8�M�����B�㔏qxn�z��L!�>��& @`�'V
 L�[k�݀��y⓮�� ��j��'T��l�V�G;|�@����M�Bq0\�+-l��	����G��'4����� ��M#�ٷ�Ž��2�e�*V��)�0�ڲ9J���D�3��4�������m�Ӻ����eT�����#�Ba�Ď�,�6�2F3��8�LB
HȰZ��
C�!a0�$�:t�6<p�D���6� ��d�#W푞�ӉUp��()Ā����-A>\��*H�89Z@��Sn�^�P`�T
+�����I�VЀd񐈋����Rd�R
��F[�0Q&�� (�֦e��/	�$��4��-��	ꔓ�.m��	[�=��0��{��4⠨X�:������䃗\�H�cF�Sdv��kH?�	�[2�@�@�y�(-!��
�h���c
�\���ǌ�0&� � �t�D����Xw:�b�����١��1��8����j��\���=J}0��g�#����B�O��䂕4/�Q���"����D*��!�,^D��l�!N���^�7����A���]�T ��m��gjj�*�(xļT��4�Z���DOZ�x��F 0�b���E͙Em
�ѫ�#�z$0Ŋ#m�( 8�a]<l�6@!��	!ټ�b��3����
ߓ'�n\���	ކ|Q#���V� Ix���5HA����e�'�)e��C�}Ô��=MV�]���Y�]��%�ϑ���i��˪aqL�
�O:4.h0���Z�̀�É�31��3�"y6j-��:8��2��Q�C�i,����@ā�xr�Z�a��Px�wj]�6�t�ȧŌ�%�d-HÓk�����Um�<,C!cQ-���8�L
�R��:w�×F���r��X�w�$�j��ػWO�]+����4:�@�+��y�B/D)����uk$՛!_�stB�Pe��AQ�R�NB�Y��E�''�EpFN�8-=�郕��T-D]��a�%l�Ix�	\kx�0���+�&x�2���wp�ч�I�޸H�Ù�C"ZTQaE�!G��佟Ѧ�2,c"-x੅�E'��aL�#%��0ҟy��% w�%`N�#$��d $��;�0=1��2�2��4H�. �GpN����/HSĽ���9[��q�\
�?�0MԻ!9ؽ�'x'���3�u'�Ͱ\l^��Bԫ�~!�q�He�>l�Rm�9c\b�l�Ve�#�\�x$��['��S���O哔?�x�jp!ɞ9�^l��ϐ�-�Z��_�"_̘��ݦ}>���Ua��)�-ЬYl�OV�`��1+&�V�V�C�< 
!g�-�Ј�jҎ)unT9���P����u��L�q��ސ���O� �2��K)d���0c�I!h��yj'B#=��@2�[/sF�{��H6NzM��W*'ތ��a�O��?����)!z�s��@�?�~d���@f�Oǲp(��0z��D�$҈D`s#�u����I2)�"����J�5�}��@C<Bh���+Ҷ�Q�§)N��B"�<
8"A�%eî;���S��Ӧ�jX�0ɑ�brM§�,T�����$P`l�<����`m$.�<*��@Q�����'G�n̓#͍=d��"��2~f]%�\�A��-w��yb�.b�z�(��<����V�À[v8��%N��x��N��Mt�S���)N< �eAC�*rl�=��i	6�C�	'[N*͂�����=	�䟤���x�~�E�ϳ ��H��H ����YX���E��p`܉�����'�P��Ipn�}YS�۳*���"Ī̾*�T�8�D�"�(��4*z쩦EŬS�H%*�ț�|���C��w��)ʧTh������F�6N8+�h�<�2FkijE����I��i���O����U4iKu��Wfe�%B�q�h����'J zaNA���g�E<�a��T�p�,�wL��A���[�K6iHd
���">G���_�Ot�'X��t٤�C�^r ��B4^��Ɂq�Z�j<��!�0�Oͻ7(Йr�h�s�;7��`�'�+��� ���u�9IV�E���;�ɳ���`zt@r�L�w��Հ��'�:!;c�ǛXj��D��*|cHZ	|��U�>´���& ���4��,A^��'(\�[���H�>!Aq�R&qܴ���O0x����&�0y���2T�(�}%h���ԋ"�a��y��'#l��	�����d�^����xN|�>i�jX�0� �ȥn(`��Aҵv,���	-��ć'	W>7]?up�"�լ��φg3�z�&H'7�B�Mk����Ig���VR� ���h`�C�hDRu._)� $���i�����x��S7
���:�A�='���UM��$?"��ę)uFTQa$ٯ�yb�\85D��1b�Mg0Q��K��dר�4��@%D�o�X!��	�(H��DA�KF����Ũ�8j!�d�0%C�P�A��!|j��s�9K!�d�)+���a�߅anp����wJ!���|���J�(p�,��C�b0!�DC��~���J�n~z�i`�W'!��ݢS���`�Y�7"�(!�$�7{Z�p���G99IVd 2#�6	!�d@5(��D��&ؗ @4pЂ�¡�!��\�z 	�v�T`?�AJ2!�N�!�$� ���,J�A��9����C�!�Ć1W5�A#n�6,�ʸC���S�!��ͨǸ0�D�.d�UjEH99�!�DB%��5ʣ�VSR\:G �$q�!�K�F�0��$	�$:eJ!n��!�� d�  �L:3��́�Ѓ)<~1��"O�Y�3A�ĥJQ�֖b�	�"OFm��K�0�U*�υ�J��;�"Ofӂ��;���ɧ�X>y6��"O�Q�r��u�H����O�P꺘K�"O�X��^98�����J���PW"O���B.�Фb2Hޞ#����"O�@$U�jF�5J��Ȼ� �"O�u��K�b-Qa�l�=?ٔ}�d"O$����%+��[�+#�n!��"OLu�qm��x��H���*����"Oe���1c�Г���ZVe� "O����8F"��G��<\�F"Ol��m�+2' 8���^:�QRR"O`��)�
0�ъ�g���	�u"O��7��O���@��"h �"O��S�\�;��h�w���yFu@"O.0:�eQ�@�l3"0,�;�"OL���"ȥ����I�y\A��"O<D�4�_����!#l:h��"OL���%{�JX���n	Z=i�"O�i�fB�#�>�pᝆ_\��"O�H� �ˡF3�@���u�m�c"O�0�t�63�����e"\X�"O���i�%CTjTTe�|V�%a$"O:$���=qz���C^�4@<B"O�H�F��9e6� �b	>0&�h&"OT��&�O�+1��"�aV(��B�"O���f]773V���)\��20@w"O���@p��5QhЅz�r;#"O�Pdߒ#,�\HTf7C��"O��`�I�m�ȴ��x��+�"O`��S�c�\�W�кC���� "O��2�i�:R�9��-6yN�"O�4;f�1��m �Nրe�Ba"O �����o�~�
�D��=B�"O �C�O� 
ިi7V�H��ѩe"OP0#���s$��+qsP8��"Or9�m�;[�pRQK�_����"O��"��3tC��2��HZR2���"O��i�N!잤"�-Q-G�Yb"OH��&'�+f��A�9<"�"u"O���q$��[�r��$+\ake"On�� )��mFf��'oݍ'��@"O�'��mq��
Q뀉@�Pq`"OH%5mm�����2II��	�"O���É0S8*A��g A��"O��2�	FqAJ��gя%Xl*5"O���#��yd����Jlp���"O���GǕa�<��"�k��v"O���c���8 ��+W�3fv���"O隔�޽Ine!ƩG�%��"O����+Y+`���B!�K],s"OTQ�Э���Tjϒ�x\e��"O�8C�#��x�pU_t>��6*O�}�Ң�1.�̹���,2�"�'���*�j�[����L7S0i	�'��R5��);�xq列�C�� @�'��j�iǐL��U#�:,zT���'��b�۶de|��dbU�Yy����'��m���i�t"��Q6x���'�0�����n��q�m�F�l��';N�x!Oc��l�5"|& L�ȓ/��ɲ�E�✼#P!�|-~q��S�?  0�a-�|e�qR�(�!�-
�"O^�⌞�:��@ �2|�:l�`"O�m)�oW&ea�p�ّ>����"O&�*U�3U3,��ݡO�D=��"OB��V��6b�Yk�a�x��ز0"OvI1PE	�2��)��o��(���u"O-��狓��I01Y;h��'"O�x��d�L�-��.�<8�E(p"O�0�bņ낌��-C�v)6P�R�'Tў"~b�f�I^�m�6C�xf��#����yb�K$kY*;|d����ǲ�y�����@�/�"9���+�O��y��=o�p;A"ߙ0�n��-��y�K��4��i�|������y�
�N�Yy�*�vR��0���)�y��=5�	�fD�v���#+פ�y��E�?��U���\F6����y"�"hyN=q%ʅ#]�$	��E5��'!ў�Og0-p��B2���%!tӌ!��'��)�ס#̜�tdI�s�8�a�'�z�97D�?��{�l�C�xI	�'��B�����#T�=7��h�'d����%Ef�4���4ӈ��
�'}��3�T=Tr>���\[�f��'�����By4���#\'}��PC
�'��c�'�^��yf��i��[�'� ��E�	����	S��I�'Ǩ�y$F�_dL���cW�P�~H

����""e��2��4�D�K��P�!���2\,TA5��dq��3�ɤ!�D*�b�X�,ּr}���H�:L!�z� ���(	�e��R�脉JE!�d�+Y~�jR�ӓ.@���Ǯ.(!�dޫC����_4�A�N�CSў���I�b ��c{6NL;��/ `B��*b�Mh�c�i�z4	1$D�}zC䉋I���A�����QV	�6�RC䉂f�n���@ߗ�,PK�/N�}OnB�	�pt��#��{_*Рu�L�S�B�	�_������`�FJ���B�m�J�[�`"`^��T��%c�B�?bITtir#$UlE� G���������O�����&�P�;�
'_�F@Ia"O`iC�MX�fxl����ˁjt���IB���i�a������ �F�?"!��'��HxQ���:��4���6$!�؃U�:�3�+�>S�0� ���5M&��pG�ă:0�nAiV�5n�<9����y���E��̘�a�`phA�vi�<�y��G:`�(WᙠEl䵱�_��ymܰR�TIð$�EYL���A6�y�0`�`��ϓ8Cw�-�4F��yr.�qF���$E9�������O�Dzʟ(���MB9V��u%�f�(s@"O�� �CV�(�69Z��1|W��@D�'O�O��D��O&TBAg�l
ix�K�5b�����'���q�? ~���ʕ,�����H+D���NS�_�9���P�k� %D� �ˎyW��6�O�B�A��8D�p��,RX�ӥ����.i07�7D�p�([�\C(�JP�>W��Bg�5D��෍ @ ȣ�$�:[�b3D�h����=IFtq��ʲ1
�a�1D����'�Bd��df�;)M8샒l/D�� �|�E�0Wؘ�E��p�ms�"OqR �$g���m!5�BՙD"OT�У�??V��(r�]cw���"O�`�u�;Tb�`���bn̺��	M>�p�J�f��eA��-j$��؁�&D���rbtsj!�CL
�����B#D�l�nMC�0K$던Ԯ,z�+"D��bC�� �<�#�'��GH�B�<٣�x��bBb�WB<�w�A�<y���MnVmIB��*0^R5���|�<�d$˦f�h�`׋u� ��a�^�<����'=������J/��J6�\�<��dU�6�n�+ů�'*�$љ�gW�<���%TC��	�٤!���Ae��]�< ��g�=*GH�eZ�wn�]�<�W���B^ts��L#H�ȉTN�T�<�� ��6��Y;G��_�� �p��N�<��D:z״D7i͗V�	$Fd�<� �8�a�d@���|!�l�ᦍ�T~z��µ[��҄*�W��ą�-�"�{DR�&y3�۝/�p���
K����F�E.%٠cV�Ȇ�Q�|�AViۜX���Qa����ȓsR\�8�ޑ+lB!�֤T�,���ȓu0�!�	9$�:�p5�Y"	K: �ȓJe�(�^	TV�P�M�%q�r��ȓ"�ƙ�3I��A���6��
)��І�V#���Ə�"�Z��UxU�Ć�o�Z��JE6Xcv`QXwB��ȓS�b��jH�K��5M̆EU����?p%��N(.R9C��i�e�צ��Q�"��홶{f$����*�8��ȓu���AF���)���;��ȓ\�8��,�+M6�=�cA]� �T��t�2u�+tN�H*�霠#R8H�ȓ"� ��@�Ԁ7������2��m���LP�Ʀ�.wl���z�A�����aʚ�hHc��6X
����.�2�
�IB��%͓,p���ȓP?L�q�T/��)P+9��D5O�dБi�1>Đw��3)�h=�&"OH�r�ĚO�2�"�A�,��P�"OX1 �/yw�x2 �(|4"O��Q7���0˒z=�!�"O�<�夙]5��BF���#(��q�"O���ca��:A. :F�	V{�I#a"O��P�� ��.=��+w"Oj��
��v(p��
S�?�h\�a"O@�"�
Ӟm<HǨ�Ϭ�@"O�<z���!��d8�)�5 h2"O�)4�O�Y,���(H.%��Q��"OБr��<r�.��VH���4 �"OD2�%�e�@����N�@�"OD�����y��0�!�[��#`"O&���a�k�!�ōj��8��"O��w�;4�� r[t�jQA"O2au�" Q��I"
��8��C"O�b`��_�5�ӯ#��s"O��e�\�8�	���N�r<��"O���G �m� l	�la�зk [�<�q�A�9�0�Q�t�)(Ǩ�L�<��+N0~�^�0�ί��]³��_�<����D���Bm/gR��3D �v�<��c��T���q�AB�	�,SF��\�<� ��Z2���%�ҡpU�hPv"O�-���$cx�J�U&8���"O`�yD�H�l�Z�
 ��"d���"O�\��D��"~��D�w(�ܛ�"OdMP6�6M�(�:���(	��أ"O�!Ub����������ٲ�"O���#.��6�c#��;]߾�a"O8�Y�\?
�L|Q%ߘ���D"O��K�K��� i���$��8�"O4xcE(V!E�� I�o��Ȅ�"O����B��D�л�͛�W�*�#"O�1��BE�~���o��X� e"OF	S� gIVxK�)�]W�P�"O�8��!�4Y�ch�3UA��r�"O"��Z�LKbT�æ�"G*��&"O ��É�!I�X��f�����%"O�<:���%q��hC��D�(��"O� ;���e�d����Q/~wT��"Oz����\�������#���)"O�)r��12AiXg#�8k�"OT�cŋ<��Ժ�%S18���hs"Ob�@��V TD��0")
}@=�1"O�h�AJ!*EF��!��2kk֤c2"O�D�`��6vBl0T�_��x��"OT�� hր��\���	�=k`�zb"O�ac���m�B`+�.Th�j"O�R� Ӏ4B�{󀘅3_(�W"O~�)G��:�T䩃O��)8b�;G"O�9�w�[�<�6͈UNÖ&�@5"Od�:D-ВD��LN�Tk����"Ol�Q!��7;�<�2�+��}= �b�"Ob0� `t|�QV%��y!��"Oh������Y>pP��04�G"O��ҖJ��e8*X���$3�ʘR�"O��rj9v�Z\��!�o�,�y�"O�,�1gF�T��]��n<��"O��A��`�xĢ'�N�Nݴl�""Ot���۝_� ��C�?J�8�6"O��Q6B�UL|�E�h`@(�"O��zR폌,��MD�W
c�Uh"O�q����6as/��Ng�a"O2PbP��@�șDA�(�]�0"O��c�:JE���Ʀ��=�E��"O��y2J����H����-"O؍*e	
$���veN�(�B!cs"O�
�f�8�0%*�d
*K��ɨ�"O8��o��7��Z$�['#�X��"O� �!��{5���D�/<z\-!"O�\�Db��H	:���i�"O]p�A�����'ɳp��u�"O�lb�Mґ[�N ;r��X����"O�}��X"D�KֆW8F�MZ�"O�ЋC��a����^o�Ѐ�t"O��,��F\�
Ƣ�l�l�93"O0��]��MYF+� C�� y�"ONl�q/�y���;�@�0}�^���"O�R�/��q��E�G�#��34"O�P�T�w��]r.��,�d�a"O�X��Q�ޑзM��B�J`b1"Oh�pa�r^��2���o����A"O �cDƲYuk
A�p��"O�hSa 4%ٴ�i�
�0<2� �D"O�iXV� l�n�rc�<(rE�'"O@قRE�2+��!1�E���p"O� ����S5$p	k5K0>����"OR�)�a�x���ac Y�|�>�a"Oj٪VC��cj(t���
�$$*�"O6LbgX9"B9X��_�B�x�"Ol,�@'ʿg�l)�r��W����"O�|�'�� 	���sC߬@�z]��"O�;S���|ʴu�!���P�#"Ol<÷Ηi�rH�QиR�!k""OpDJ�� �i|~e�aMM��$"�"O�h+��*VJc��^��("O�S����&됌�3jÍFA��"O>���&[L{`��fD�j�fر�'��D��SrL=q�M�r�%�ȓ&#h����2_\`�g�xe��O�� ��O�`�pȴL�
p�ȓ )�A��� �k���y�Ƥ�ȓ-V�AS�J�n��Y�
���ن�"��i�|���DAW����� �6�8�n'�\��g�<o��|��;���1��@/"9��� ��%"���ȓvs&���Hn`:��虰_����ȓux�Hv�F(�r�;�H%4����ȓt�D���gīH��o���8H��l�5ق�P��f<��R�H!��r�BYJ���0I�C�˻V�n(�ȓs4��7�χ*�����KCP��_�(T�$.��\�\�r�	!	^|�ȓX��Q�B��b4�H���%�=�ȓ=d|�P��ű~�&�(bꈻ]�65�ȓ
�$�S&�&@��!� J�cK4����8�sŕk�8<2�E+X�h0��ER ۢ�X�Q.����D�TZ ��ȓ�rTKN�h�����(=��ņ�7���TF/hݲ���%K�~����|9�L���;����$��]�ȓ\Z$�ç��j^�S�dփ�",�ȓQ)�����B��C�I@6x��P����e�R�`Ț��R;8'B�ȓ&:�q�*�"��{�!X��ȓ9\�/T�t���K��զT��Ɇȓ[�P���R4p�>#���.i�2��ȓ�>dQQ�O��X���W3��u�i��W�!k!`�&>��ȓHh�����R_����(&�6y��a)�\����(U�H3b�g/R��I�J���"��ձ��Ilܮ���q��@	ԓn�X!ρ��@��ȓJO�q��B�riCR.ke���K���DL�����x��XI�n���i���X#�޴�*Y����Ό�ȓL�v�Y/�)��"��a�ȓe��SJe��������-������t��j0��9qf9�ȓ2�T s�M�X�pyzw��y@ԅ�z��4"S	�
M>a"��UYx��ȓ|��x����47������a��M��5���g
S8KSII��N�St��ȓ[�� j"O
�J/<$"y�����,�����)N=���	^�ȓ7qԬ8E���0��R�%��"�Ȇȓ6M�u�b��u�\}ZT��V<L�ȓx�����O�>B�À+��$��w���Ϩ�9aʣ � �ȓ]jmS�a,T�x�	",����S�? H �$�^�Fq�&5=�baZ�"O.a	q͜��P8zEI�D|t�c�"O|�g��E����B;_o*�8d"O��;C�%,d.�����`�o�<�GBW&�d��udнH͞��&� V�<)�+!$}���ař:�D���
I�<�Ģ��P�ХO�44
�2��F�<Q��K4��0 ��(S�\�Br��k�<��ƛ��Z���Hˋy�*�Z��|�<��PV���5
�-ʗ���C�
a7���ߤ
�����k�fC�I�@��)C�M^<<�cDёJ*C��B�к"��mV<DI�cTJ
�B�	1t� D[��$� С'�" �@B�I=e$E &��
&�"҂	A�B��1)4P���+��A�ҶF�`C�I�P@�ء�Q8�4k�Ѓ,B�ɝt�.X�2F#ZF*��6�N�)��C�ɋ#��iB%��A�
<k��
�s�B�I�GK�(3U"�%�����hJ"U��B�	"�Q�X�$c 50`�F�B䉟)�P���K�iT����U��C�aP��س,& �#�4g�B��q�t���$�]\�i<�B�ɱt�, ���	����J&�Y4�jC�	/?��̫Bi�dI@E�aY"~m>C�I	.`;1N>� }� �DjB��,���O�"q�Px'��t�4B�	�.�2��<J��T�2*Y�`�*B�	�N�k�#�� �2���ָE�2B�i*�E��NH���O��W061�	�',5�g�U.s��3�-PA�t��'���8W�D8$sí��$�٩�'��t�5�W5,H&5���	nX��'ȸ��ş<����a��9D$0�'4zi10(�)B3������j�f�x�'���d�+Rx6�h��16����'vy�F
jJ��3p��+l��Y�'~Z����َ(밵�`�N1�
�'�8���#�.n�H,Z�L�� n�2�'��\��LS "�K��.9b�<Q	�'��Iږ�O9Ơ�� C�:6��xb�'��L����tf×2��y��"O�)�� í( Px��Y8'��4@�"O���3*\+];V�h��V*{�t���"O�E;���z��2c��
��`�"OԤ��,W
w��b�"ңp��+%"O"I�7��JO�tz�@��b��	�"O�4Q-�W=8��F�ĺ0F4h��"O���wΜ�7���3��WE�9��"OҌ��j?Z�����F�	شy*�"O�Q;�' ��q�cf(43L�� "Ob���T�xb��J�w��|P "OR�⥋�/(~�R��U�5�Q"O~DgJ�*3�p��y��)�"O�����;y�	�Dφ>���c�"OX|[�Q�H�F�� ��늠�u"O�(1�ꕑ_�`%�w��^�d���"O`T)��ǋ�`ى�
�0m���P"O88!"	����`�萹*w��5"OB(��+=u��a	 �(6"O0͘��	�Gu6I� h݀T�6��"O�H��JN Y?�q	��Na]<�:"OֹX�D9 ��)q%B.�v�$"O� f|;҈�z��5b$��m��\!"O�$x��
1!��}�ТXf��P�"O2�c�l��&,V}�w�+��a�"Ov�RcKU�n��R�cG�T�x�"O� �,o�� EO��X��"O���w
R��+@Z,C~��0"Or��娉D���$N4Fq��� "OČ��	��nx������i�Ґ1�"Oơ���@�sSJU`eE�W�1�"O�|��\s����J9����"Op��՘!�2�U��!��c"O$��g��)C��2$� �}	X-��"O20�⅒b/�{�k��$E��"OROȿa~\y7kR�,���H�"O�D!A�M�Y����E�N�|�8i�"O 	��%8krT��h�� �#6"O6�:�(�7	��D٠�7��X#"O����h��H�@���2�<��3"O2:AF� ��KdX	n��"U"O c f�i~|p�6�@��%+"O��փ�:�|��d,ܗ���W"Oj�8�'�Z�&lH�!��F"O�}��Eb������!*9�"O`��Ht�b�x��	hW�D�y+�4�REF�ԌH��d��y�K˄j[� �'G��)�8����y�ڀ��U�T>�$9@�HZ��yҠ���= J,*��ڑ�L��yR-��C�h[ύ�r̸@PVn��y��P ���z�n	�=��Db�d��Py���t>�+b/q��8*���c�<�"��<Ő��!Ϭf������\t�<�6A��{���BBMT�|��!�aX�<q��Pq��S��i�B%�G-KU�<�ӷqD���������hR�<��h�BLY�G��x8�b%�N�<Q#nP�ݪ,�e�	*&Q`�`�v�<�$I�M��M��Jc$�sRNq�<)0�]�\�",H1�ir�I*D��� # \P���:oz��#�$5D�<��b�:`�T郍�U��`)p>D�L���">=h��GÎZ�pt#'D��� �;����u$(f���h$D� ���(�1����O�D�"��!D��b�+��u��b�		�N�>8�?D�h��ąuqܝ[S=N�	�>D�h�B�U�<�Zc��n=� �N?D�X�d]�)B�11Tjz��"�(D��ڲ��&F�=��$^�Lx�1��K$D�ТŠ��q�����ğ���	�'$D� !qB��z�![t�sV�9a �/D���&I�F��e�-Z�����-D��D �.KDZ�b,�,/`��'H+D�(뀮��X�2b_2@���%(D������|:��]<t�P�%D����H�$aC5��_Ėa 1�#D�"%ǌT�t�`1T�l��{��?D�PbH�8�0��W� ���ᦈ<D����ax�k��#b�H� 5D�`Y�d�6�4�1V��2�N`��*'D���1�K�|�%��%n�F(a"D����x��[灂�	O��>D��AJ�uDy`$ߠL�p��H>D�l��#L /��uX�)���j'D�� p�3	Z�, u˧�!h��:�"O*\�u��}l��r��Y�D��"O�0ӓ�.��r�.{k@aQ&"O@��ΗxLz�k���(J|N\�"O�d"d ӌ��԰���=��IA�"OP�ZEm׌�:�Bf������7"O�ʔ�>I���2�φ�;�,I*�"ORH����>�j�2�Ԝ=M�2"O!���*T�Ѓ`F"0�ݫ"O\�B��ڡpD:�꠮ȪG�e�"O���PO������/`��M��"ONx��?h�f����<D����q"Ohl!gCE}֌�3��E�fha�"OL�� F�ʥ�1L;rr�x;w"O��`k�0)Ԝ51�Kތwi�B�"OB���<��:VJ�hV���p"O�lA0?�A��M *i:�"OzM1�bA�pG�II�',=ȡ�Q"ON苆��50�;`d�00����"O\А�h�!^I����"�?FH��"O�y�Q*{�2���?�A�u"O~��E��G�(-y�g�0[�"�"O���C�YeH��u�߹I���"OPh��T"ȉ�R"�J�h4I4"Od��|-�C��&n���"Oƀ���A9Cu�	�c���"OxHiA��H/.�iSh�[I���"Ov5���4�P����#:N����"OQÐa	E�xgAE�j� ف"O�͘Ӯ�/Dp��9�!Q�h�\y(�"O�:�W�_ ����UW�H�"ORU����i�<ZҪ؄4���CU"O�eB�0[0y�%i�j�&(�"O��R$i��n)�'h�]pZ�Q�"OԽ"1�6g��	���I?dS< 1�"O|�R����р��q����"O�ErrL�'���BP��$�H�q"OJ@dD#v��i���N.4�r�A�"OI�vj9A�<cf�WSFx)��"O,����L�HL��s-R�"�8"Ob�c��-8� 7
�����89l!�P�Ń��S<O.h�j3B�[g!��;-���cP?�,b@e�"f!�Z;}�T@�}ݪ�ȝY!��8���k@��� l�⁏��!��� O�uh�ǒ�6z�a�R���c�!�T�\��X �]�Kq"��&��/�!�D�#[
	�A ���q`\�!��Kw����ɈH?��!����!���@��aQ7�eSG��g�!�dP�CeP؆��-YP 8���~�!��h7x-[�	L:0�H�aO�H�!�/[�2dzd�M�X�b�>�!�䇃Q������l:��ŃR�M�!�d��^ά(�ˎ1� +�す^K!�d�!'-��9u_�2�9A�M�|9!��i����=p��!��׉'#!��

�4B���^(ơQ��x9�'C�h!"
�./�|�0��_L���'��H����\4#Q�Q�n��p��'^�����.(��D�St��j�'���q���s��U��HT���k	�'��� 6�׭j�Qp5�*���3�'�R������},��%&M4>�� ��� �hkD��?�4$+",	�]*-�d"O���G�*t���� �nO��{d"O��.�
�*���֔~�Z=X%"O��2�C�3��T鲡��{�*I��"O�I��J]�X���T`��ܥ"O�MW�ɿ2̰\�3旧�PAv"O`p�B��=��ӥEM�%�:u"Oش	eV�o����r���⸛"ON�7����u�c�
s�Rh�c"O�@�IP~�8�6Aǫ�p ��"O�y9�F�7\�Z�X�'��a��"O4��1�Ř/�0�Q��/DL\�@"O<Y1�g�����0�Ǒh!��"O��;�j�"n���B�bA�LDja"O����%������C$+.�y�"O��f������b��Z�!1�"Ot��"��X����ŁL�#��Z�"O�<��Yx�H��F?[�&���"O (y&	Z1|u© K������2"O��#"O�%�a$g�>5����t"Oh�  ͘k�R$�s#G+m�A��"ÓQ6a>Ss���J��pJ�"O�Y�#g�V�Lh�c�A�Rdz"O�ɑ�, �B���j�퇓%Ҡ<��"O�YS�+��1���8q��]����f"O�u:$"?^�lX��!&r΄�u"O� �fdN#A���	2F�"OΡi�I[� ��`/���6m��"OQ���8Θ�*1�Ǘ�^��`"O���5M�D��� 1�ֺHe����"Oؐ�@I��+�zs��4l�����"O�Q�ś�RS��Fhͪ�P"O�a��TF.l�1�N��x  �"O���Or��L�g��`�4H�4"O��ず���C�ݥ~�����"O��8s@L�n����efc�Ie`0D���→1R�4��ajN�k�&d3�1D�(��j��-8\-g����`Ew#0D�����J
J��4:�n�#4ɪ'/D���Xy�A[+-��ɻF�.D���uKI;0�̘��/2�l "2D+D�sb�%r��{�'�>�F�q�d3D���1B�q�0C委"k6�D2D��ЦҙT����CFM)l�R���#;D���R�_ �� a���[��\���7D��@ �C�p-�tb&Ky���$�"D�|�#����*�J�ɶSɨ�x'n!D�Ȫ֦�4a�Hػd�'*�6�P�$D���l�8S�qӳ�G��Uh6O"D��r�B�'c&��g��x`|i�t D�(C6o��2��Z�C�j��1�0D���TC�2a�)AЮu�T82n]�<�6�G<xI@�Ħ*[@����X�<qG�^�>����%�!C�R�*1�]V�<	 �^54��n��@�,�Df$D�4��x�T="%FQ9G�e�a"D���i��9N9����<01ܕ
W
3D�Trv�[�Iu�k1h�=b>����0D�(!���n���jՅ�<��6�*D�k�ɉ"DQ���v!�d��t�"�*D�T�cƋ P^��H�)�!@��lCu!'D�T1�nY�f�����"�&d�3'"T�7�߸Y((d��
!j-B3"OtEw��8X��ȳ��( 	J�"O� �� kٵmU�=��"�
,�Z\1"O*�#�
�R0�a��c��B��1�r"Ovyc�[��	��ʤZ���*O�`P'眍]�|��q �C<�|�
�'K����lx}�Y�@X�@�d"�'����w�F�+�f��C@j�J���'/����$��ň�'g0�x��'�@���A�QM.xq�R9`���'�p�g/��K�s�-S'CEx��'N��U.��8��ah�6PZ�j�'gn�;w�-%K*4�@�ӌ6˂1[�'6�1�#Ɗ�;�����*�`��(��'M�2凍!I8T1 �_W�!��'�n��@���8 M8�G�{	�Y�'��ʘ��N�ʣED�.�!Q
�'�^�)D�̈M9�Mi���+�L51
�'v��
��@�/���Gl�hp�	�'�ʔ��a�%��L�&��
V�	�'w�43�)��3���qf���cvd,#�'���i���tP�TF�aK�I��'�6�`�l�6 T��C���[��Z	�'.}���'=2��gc�"ZK攚	�'�h g�V��h&HBb���'fh��ܔ�褚�@��2e>��'��`��P���*�Y4[�B��'���x��
p46(8���l0��'�����YjPz+U�Q]rt		�'Ȕi�$ρ�_V����"�X��И�'������r�����}M��'<<�䣀���[ �@�p@�8!�'��zCj��:ǞuK��m�^���'� ���ʹ)�	ADH�k�d��'t�WF�|s�t9N||���b=D��;�):,@��-=J��>D��)�ǥ��]�f��fT�9a�<D�84C�r$��COʾa=��j��.D�$R��������MS�nb�
�))D�X ���d����a�E �1D����"I�+��h�$��Sֶ�±0D��!6'�B��mL�M�<ȢS�,D����ߍ0�����h��E=D��I4�D���l�ҤJ"�  O<D���cF�R����[*��#��!򄞏A�"X2!G�^Mt�󐧁"w!��H�K��ı��̃�&�'p�!�N.�����j:7qR��2Ł+�!�ڞ P�m�vH�
{����&ٴ(u!��Ҩa�z� ��`�F���R==q!�M�iB
�U d٪ū��؄ �!�$���j�?,�,�Ӵ�2�!�d�j���sŢ�:�n�+e�G!�d�Swh,��"�>��bC�J�L�!�E�$����o��&dL��D��,	!��"_��9����\��#%�[9x !�ï��q)�Rs^�J�$[�!��^�~4�OǣRT�����<B�!���:{g��[ҁ��gNR�Bc��'%�!�$ Ls�T@�`�;K 19� ��!�D�؈=�0�7�N9�&��QL!�DŴMF��*���|e�u�LT3!��w���7�T
�tKI[��!�d�%��%���F����(��!�D�>Fd��j�yR���d�L�W}!�$y�E�%�_HX���&�j�!�� �%�/��Vs(�rq͇v��m�R"OH�8�̉<e��5��*-�:�9�"ODia�l��s8��z6� �%�jv"O�E{�-�	���8׉��H�	��"OYB�"$PB�A;�iU<X��K�"Oly�2� 98E�iP5(��dv��f"O6���*:	�M"��@[T���"O���ֆݷ/!�1H�Ǎ Xފ=��"O���g�mkބ�ԇY��X"O^y���Ɵ��<rQ����Qy2"O�	ꅼ7�T�+� ��4��H�"O^���cE,5�r�P�K�Δ1G"O��h�Y� �:IIvZ�<��&"O$��B˕[`�0,����@#�!�Q�g���IR50�,P`����E�!��T��@��u�X�!'l΃I!��:����'�)X�,0�6ʃ�y!�DS�QI�l@ �2��#l�!�DOO����^���ڔ��N�!�䉳J��ћ�U'm�h�,B΂"O�B�=(t�)� 6�����"O����
��?g� �/�?(z0��G"O��
�"�8vi��SI�JTް 4"O0���ƙ66?ƭ���D=��"�"O�Lz�^������&=����"O�����\JQ(a ���+`�Dɂ"O�e���ںK֢)��@Yu�� 5"O,�"H8PZ�|��ɞ�!��"O�����W�1��Μ�]w�RS"OĐ*2@H���9I -�ol��Ju"O.@�A��b��W��=J�����"O ib�H��
n�)�	Ξ�+�"O�1@��¼m�<"K�͔�3"O^X�Wh��O�n�q`	��k��ո�"Oh9��I�p���r��j`z��"O��H�%(�.=2V�QT�ؙ�s"O2��� �a�<x��v��qS�"O
�I�G7&��!�SA����*P"O𥁄*��*��fe�+rh�x�t"O^]�ĕ1� h��C=@abE��"OfI�&�aq�x�t�]4L��i�"O���@
�zЈ�C�xAI#G"O@���3�h��c�O"$�b""O�1�a�t T$ �@�#���"O~����%�b� ���s$<#"O.԰b��F4��XB/�$�Tȡ6"O�D����(K�"�{��B�<pLpY"Ox|� �	B�I�a�G6 b�m;�"O"�	u.�+&L$x@0&B�zc�0�D"O�� *UI��� ī	��|s�"O�$�t�KU0�p��F%u�@���"O��pc�� ���N�u�p��T"O�A"Շ�$�n�� ���k�����"O i�B,ݺ"h�02$nO����"O\a�WG�B%�(!���:�B��(n!�$�Ɛ�2�ʌ}�@�!��\%FC!���Pt�a.\��� �-��=!�DϦ{,��5���W�r�w�2!�DU�O�Yr�l׭sQ�����R#!�$�!ԝ;Ä(<��LYiV�z!��B�~�n�9��ɉk- �@F�!�d�I��A�mS�< ���%%�!�d�&\HFA!4o���)�n-�!�D�E�Љa@^�\>��lL��!�� �\�ԩW	�v�;����9jx�Yd"O<L�$d �p�q�_^θy�"OҩgM8R�jh)� ��Q_@���"O��EjE#�:�Sr �[ u*"O���P�ū^JB���X�U��Z�"OL(�s< ��$	��y"r%Rv"O.��L��K�^�i�GMJp���"O�m	�)�FP��s Z�L��2"O�FȮ#?�mB�N��= "OL�b5m��V�"q$�ͤj���u*OF�{b�0)�����D�F�ĳ�'��y����?�`�z�Jȸ?��A�'�BT��<^n�� ]89�<��'���#��	
�,��g��;?\��'��8��Fƽ=�`$r7��-sL���'IF}
d�|�T�U�t� ��3�y�J��_ h��,� m��qC�nʤ�yNB(@C&�#h���6ά�y�MuT��b�$g��(#l%�y"���*q�<g�S\W�Y��JP��y�%�7�.0 Tm�5(��I����y`Ǭ
�%��'ҧ&�l8���y"�]�\��r��� ��Hۖ�y�
Ǽ`���wϔ4�xH��,���yr��l�5c���0uW40���yBBR�؆-��ũ^L`�$"�y���P]��B~r����-٫�y�ƫrH4y�B̳{t��� /�y��H({aΘ�cj"�"�O���y�'[�\��Ad�
Z��{��\�y"�N�M����]�R xĒb���yRB3'�xԸ��D�`��G=�y�OI�+]rؚuh7f� ����!�y�BK$$���s�_��!b���yB�Вw
1s1.B&#ҞSA����yb�Y:y�E\K�9�狅��yRI�?L����ܼM�r��g/�5�yBf�J�a���9Au>�+��ւ�y�T�T"v\��K��gs�]b���y��#}(V��A��];����^��y"�'b�n9s�B��{B!�ƍ�y���;��p�׎Ɂ��=X�/ҳ�y��+N�h��'H�/w��G���ybN��T���I%�$ �ԃ��ޜ�y�K�|B�������%�0`X
�y��!���Kԡ "&� %��$�yRȬY��MV/�:<X�e���y��5��]:v��||e�&@!�y�f�m� 0���ݏlVH���k��y��ڪg���W(T�V,K�	��y��&4��X�$NDd��S��yR�������cI��J� N��yG�+2��2wȁ�B����	J3�yb'0<�T�RV�];7y4��oK��y��M|�<�0� <�^�Z�_��y" ��0<��S�3�¡R����y��+9;I�Gᑇ'�%��<�y*�5n4;6�K+"���gJ��y�j�*?u���g��d��G�ؑ�y�OM�^�2KVʐ�T[��
ǃ���y��R�!�8=8��`w\%i����y��	����ӂLߡ#��;Va��y�-��gp0��Ј�������y2���;�(PΉ�yP&�㦪^��y
� �ٰ�m�
J��}��j�ԙ"�"O�8�G(MEVHimZ�8��e"O���@V�:��}���ڳ\Ǌ=(C"O4E�S ?]aRY��Oj�^��"O�0���̒A�f$���8�T��"OD���

0(�f�Sa� ���@�"O49+���p��0��-����"O�`��DD�}:��9Ɓ��A����"O�D�CH
)pL��K��]'�`Ȑ�"O~�85�p\ڰ���=�D�`B"O�!X�
Gua"� �O[�m�hЈ�"O�����t�=����J�V�D"O~��ǯ/H2|��f�.\ІE�@"Ojm��GM-E �CM�+5�X �D"O�UX�B�'3<Ѫg�U�7��1�"O�	����0C��VW�#��K�"Oҩ�r�Q$X�<�� ����uB�"Ol��1�^�G8T�R���~�L��"O�0������`P�x�Yj!"O�cO��ֲ]9m9,ʖ9�"OL!�2q2��e�Z�Bh��"O<� �c�t�
��"��{�&}�""O(��&�	,��U
G-͔Q��4�#"O2:gk�3	<�5�3�½���{v"O���疻���Ie%4�`- �"O@���-\�/���ɷ���=Q����"O����+�F��S�M�L���"O��vAD�,(IQ4��?=2�a2"OjAR��t�IxG�Od��g"O���Pn��FdЈH��)�B)@�'"��J�%%C� ��[3hb�\C�'���ZTa��Z�`S�
[����'w48�W�߁3�ʁ�R�ۦE�Y�'��q�#�m�N:դ,TR�lh�'|��1�Ȍ�&��3��K�65��'�f����L&
�H��*
4mվ��
�'��3�޼{!�yj��\�cr���'�bp	��Y�Bu�#� ����'��m��c��i܈X�&"	't�
�'��#DE�7��+A`�{'I9
�'��Up���"��]�s��x�"�B	�'�0���;� ���.@jR4l)�'���3�̀k�*BB�Y�_pL٫�'Y��W	8 !��@?h�4��
�'��`Q��Ӫ�~ ǈ�`�����'�D\j�f(.AT��G�Kr6��'~���"3j���f�"�L���'���R��:X�ZX����C}��
�'ü����N�
�е��I�;<�ѡ	�'~ h��֭D:޹`t�2��8{	�'J���,^�^3���(�2����'��y�a�U6��I�,�%)jx��'���Pu#�/y䉑�-N(?�"�'=\�e�>8Ϧ��c�ќ$���'M�|s1/C42��(CKo���x�'D����i�`�P��5̰�c�'V����Ezq���9}8�A�'���ԉ &j����O5&���'�La��oQ�C�U�W���cH`�p�'��ZEb�&'P�(�� �r��8(�'�p�a��ٝ0�X+�%m� ��'Ib<�p�G:go&��t��Lؙ��'~vh���3\����g�G;��	�'�p#���a��#d�ߧ?N��8��� ��(��N�W�hQ��dɼ`� t�D"O�՚���O0|b�c�#%�i��"O�B���:X�,dCcV�e-�LӰ"Oʠ�[����@AR�d�q�"O���U M�dO^( 2�ǅ�@(��"O"a����8|y�U��W��20"O�Ѩc��(�����{ڊH�u"Oн��7r�"h�q��$PF)A "OҨ*%����'�H�["k�"O"MsiD=��E�_(n��"O����]�X����w@��q*�Pg"O2mc��T�����n�p����"O�h�v+ZZX�T��N���Z�"O�1!dF\uMx(�N���Ε�u"O�ubu��( �\RFL\�[�ȺA"O���6(��sz%	!�,X>1��"O�I%��:�L���I��:JhIY�"O�1��'V�M�si�'�J���"OH����V)� �H̊��Md�<y��M�H�=�p ª-�R��x�<��
�4�֐�?h�"=��O�v�<	dh�$��Yð.=G�*9q#�z�<��DC�nwb!��F��:��Y9��r�<9(6M3����FÏ+����V��h�<�Wٍ]R\�qf�N��t�S�Z�<�Ү�"v{��S�F[�(�yjA
^r�<�s/��h��R ��B�*1�$@x�<!�O.�"-xU��tɢt�<qb#3@.E��SP(4����v�<s��$ל<�P���6X�����I�<��ꕹQn|Q��P�N� iJ���F�<�R#�?���jƂU�f&%�����<ɀ�ς4s�U��aҪp�����bFy�<���\�E�BH�1�Q�J�fE��.�P�<a��*��A�E�Q*"��5*N�<If����z���'���yra�@�<!!�\�L
p�"D��in9կ*D�<�ƦN��� ��i�Y��jc�3D�̒6eY�n� ���6k~�p��0D�P��$�(1 ���%�W�N�ñ�,D��(�K��oCJ��PɏY�j��V�*D��ڵ+ۚ-��$}�Py�<D�4��C%e�X K��]�` �ا+9D��5�	�F�.�kT��&��(��:D����(ղK3���Dꕚ{��Zs9D�8C�A��\
��" TU�hŘ�m6D���@��vh���\�:�<��O:D��8�dΉ)���5x��#��5D��[S�]$*��M��璏=�z$+qn8D�t:�'�&\�,�$�F�˔�!AO:D��BET�Ga�!����f�y�	8D���nԱ'��=�"l;=��1�(1D��0ơϩi�.L1�$AZ�AcO/D�l
���(j�@Q!d¬6�z,�2�/D�0 6H[�t�
���C_%"5BL�`a#D��ѷC0�ցjg� S�Ly�� D������j�~�Yb�

@d~���!D�H�tMi=�LɆ�&o~RIp+D���&���:��e�c�!* �a�L+D��$&�;t�> �qj�C��cff,D���D�2*r�䪁��V.��W�+D�0�w��>?���:�
�@�3L6D���q@K?]�������i� "L4D��xĆ�Tf�$���ĉwqX�a6D�� 
��h7n�
�@���x�"O�����U�Z����)�:C"��&"O�ԃf�E�q���b��M�@��"O�M!e�T�Qy)ҋ��u�8);�"O�1�w�Q]�$Xf-��u�lp��"O�KV�W�*�|P��Uf�����"O* ��m�4+jڄIGFM��љ�"O qIqƙ�\�ʔ�BoH�(���x5"O(����|NbP!��[�Ww��0�"O4)�ŴפY�-Vd�Ҕ"OJhwo�PސL���� |_�\�3"O<Y�6L�4o��i��(,2Qv�U"O8�Hp�ȶbW�dK�gcPƥ��"O��I���)_�D�:�یtU,}Cg"O�`���3j��m��.l�X��"O2$AqD!X�ƙcC$�Pg��2�"O�� 	�u.J�Z�C�%a��"O��� ��,�G�1NQ��y�"O�A�C�7�n9` Ֆ=<�
F"O�|#�J$"�-�D.��4
dX"Ob��b�Ӣ	-:�@�,-И2%"OnГP�I.'��If��<S���u"O 5��MN�N��|Y��T�G�|�r"OV��ЫX�BN�!Tʩ@� �R�"O�:bc���`��'e�Ĉq"O�Т�	,K#��E���"U�M�"OBa�ъK:�J�cT`!�Đ��S�N˔46\�r&�Q�'W!�BA����O=�^��&O�nu!�d�7
�x3�����#���wg!�$�rהl��C�G��mqe/O!h�!��@�> ��*Uai�)ULO�]	!�$]<W%����d��)W��Q�+_�|�!�DR�pr2dj&��Q�4���+�!����T���TUܲ`bP�T�!�$KD��<���P0lQ��D�iI!��P�^�2��w�M:
�	si�5u>!�F�Pp&؀VFُv����2�C�	�!���\&��W��d��ڡ ���!�d
�^�|� �^6hn����Rq	!�d�M**��.Z�h���q�m%/�!�d��Dl):@��2S�xy�J��~�!�ø(�
�(�A;K�HD��oO�2�!�$�(�l �a�D�s�jPK�/�6�!�"��TPbGݕp��93Q�Q>�!�D��ḷP�]��Z��"
V$c{!�D@�I�%��*�B+���	 �"O�0�� �\u��6G$Z���[�"O�j��Y���4(؂ f4�"OI)���f+���vaD�!�2�
�"O�ͪ�×@�vPR�V�QmP-jS"O���9:�6US��^�t���A#"O�E��.Z�P��F��a�1!"O.�x�+H�8�`�
�}r�S�"O�$�D׸3T9p"���#"OZЫ$��b0�!��@�nǢ��@"O�X��Q6O��8Kq��6�J���"O@�j�w���;s*J��0��"O�y�o\3xY���+t�� �V"O��z��σ{��W�ڳ��|�"O8���V$V_�4�ʖ�"���"O�Y��>%���B&^��X0d"OP�$C�\�0�)w�J�1C0"O�!	�k�U>I���%�Aq"O� ��"����R���H��k��86"OV1���D��q���e��ڑ"OT}� DT�_`��ŗ"�H�c�"O�<�C.)�0I�CJ�G�,	4"O�p���� ��8 ���)�����"O>�`�V
%���Q�"$���H3"OD@`5��%�ɗ82�BT��"O}H"!��ow��RCB	�3�d!�"O�HS���о4�c��1�,��"O6� �l�u�%x�O�|�*�r*Ol ��dK{�ؘ%��?]b�tj�'�����	�=�����WY� x)�'B�*a^G<��y$ʋ�K�lHp�'��)�qN#N��@@����B(��'��c ���(ӄF\+Gv�Lk
�'5V, ��4[�4a���Y6!� �	�'м��vi�	��y��C�9��Dc	�'p`���Dgn���G�R�3��	�'�@5���!�4���+%68��'Cna�3
�\� E�DK���/!D�t��Ɇ�t�hI��ˇ~b��!g D�IAj����`����) Rap��"D��h� Ә:�xPض��?�$��3�+D��Is�E%���N�"I� EY3/D�A`�hp�ZT��Z� a�8D��B����ekc��6#<��<D�����t�8�i����i��:D�ب�䑛����K�r���6D���'7[o�M�����j?z1��4D��;�kV:k��t��"L�`�	��1D�P�w��N,�,���ä=K��L.D���$��E���BI�=��%�Q�9D�4W ׵O�`$R�'��Z�"D�Dp��7b��}R�"G3~1B6 B��h06mؑ��@3FࡖaH
  B䉦1�v���>Zl�1	Ǣ9��C�ɼ`R�!�Q�T�E�����~�B�ɢ@�*L;���`m��p	[E��B�I5b=�8�'Ł�ּ�P��N<C�	��։S��A
�)#go#�	�ȓ �Ҵ��Y�kR�M1.N�!�ȓz�����$�?[�ٺ��A�_Y����5Q~-s�E��R����eʬf�a��p�|���NKƸ
�(�3Fb����l=���0��C��\��!�5J�B1�ȓF+|1+�V#o2|�E�^5�P@�ȓt�ҥ!��SGcd���ύ+O`�|��!��D8�GB%�᳡N_�AW�E�ȓ=�,˱E��,ph����X�(�v���>��5�,A6>����wgͽR�>���~ɐm���9%�L�Ҥ.b�Y*G"O�@&��A�Pq���4�F<�p"OZ1ď[.F5��;�����j\��"O
�@� �/e�j0�+���(�"O4�c�o)r�� K�&\��T�a�"O&8�d#ކ���9H�BM@�"Of�Y2�4XOr}�§J^?nI��"O���ď��'xD�8Q��2:��"O����=�(A�R�%�)I�"O���ǉչ�|�QOK�_�8�"O��kv)ݚ
*���# 7�|�v"Oh�+�Ċ�,-�er�N:m���"On5��M�$���/nӜH+c"O^���A(iT�Z�-Fch���"O� �����U5DPV����HW�)T"O^=#Ʈ@�p���BF$�2�"On�
�$rL��	^-��;!"O"uY'g��|������S%P�a"O�3��L����N�!!�[a"O��A���A�:AI�lp	� ���yRJ�+N�@�yp���0��	���	�yr�J�\l�6��]��iB4�V��y��@5j�"Qr`�I�!�l%� g��yb���&��0�KXAP�B�@
�yb��ZI��aF��Q�"%�Y;�y/�	/���Ak�}�8;�N&�yR�YV��D��J��+���	�y�gy�fA߮���Y����8P��'X�E¥Q'
X��t��[�*4���=<O
i��M%m���!u)��Hh�&"ORK�Z����pi��-gf�Y�"O �ƀ
�� �U�hU���"O\��ҁјO�@L�0�ap��D"O�p(dR�z���2ʵ8q���Q"O0Ԙ��ǁ�,3��g��x�w"O���4�+qM�����,�$�q��'J�ܤO���#
�U���B��er�"Ot9J����6����͝�
�@��5�Ӫ�Px�<U����5��4�q�ָ�y��؝FT���π?�* r�J�y� ΃�V���OΩ���ڰ�y�EH�{�~hW�N�xO�dH�MV��y$T�:�h�0x�N}+r�I7-ў"}��'a8�
�Κ�s���2��}ؙ
��~"��f\J�iT��,Ji�`!�W��y��!f����k�B^�T�����Oʣ=�O#.�P��8k}Lۀ�H6��]��O�$=�I_�?q��r���t0�p6�'qF�4Γ�hO?=���]�w�|9��N�>aUV9O4D�0�]���ӣ�Y�p�D���&��c�I@�O����c�(9�) 7��*C�ZȀ���I����`a��5 �����N�bƜC䉷k�V\Rv�ȈK��Y1r��Z�C�	:\�x�waF&h��BR�Ƌ<^,C�	(�6��E킻�����`��B�	7u6"u�&��������1&�C䉬2>�ĳEIQ�?��X����	J��j����Ol-��	X�6,)�'>0>���'��D-o|���/9~���@B�|�!򄎅u�L9r��]����f�S!��E�3I��$�W���y�q�דL��6�O���$Z�Cy���!�+��th�FH���}�����ް7ULѣ���7H�h��N%D�Z�`	6���`V�Y�~���k�i}�,�O���&�z>)���[I�0�B2��=h��AJ8D�,�eK�\|�Ԃ0�V� x<����2�hO?�DD�h}tX�w�ޛx,9��O!���&AYR�c�����ӌ��x��D}���>y��$�1Gڴ�㍁!p����rܑ�dç���z�j_H���S�E#.W@D�ȓ1�=[�e��Z�X�2h��1�>��)��QC�W8	D �fY3M� x�1k*D��)@npʚ�1㖲,�扨Fh��l��	����1R�VX �Rt ^=O��C�I�^�40�� �9'b�i�$�>	H��I[<�3A[�t$:dk\����c���O�<���?0EV�:"銧֦�3�BYM�<	��]�AN(��(�"J�\��k�I��hO���'e
� �H�M�+���z����y���r��3�Oh��'!�@;u��$Csh�e
��$s����&��I�g���q-@] ,���%���=���Ĵ?�c EN&Q5�((5�C�{Y�,�ƛ3���_}�4O�`���O$L�	�)|�` �c�j����hO?�!Mb�$�3LF�UQ�TE��[}��)�'0-4	�
X-W4���@~{���']�x�����+*�*ujrm#�IP�DU!��D�9W�q���'A��@`GѰNe!��6h,(8��J�9�T�i�F�CY�hF{J?��R� a<1� �P�Z`U�d"O,�r�(W?X��	�A!v�@l�!"O�1��*B�5f��2U��$J��"O���@�2 H4k����4N���|2�)�S�9��˅��ZTK�u��D3 "O���"�C���4���%��"���n8�|�@U\�x���n�~7Z�R�M2D��r�d�9+͈lꄦ�3SR%CZ�@�'7R�O�3��zn�%��}cd��c˝_�!���8JvV�3TɁ�Jp!"��3!�IX*<���O�l��H�0-+-t�O�6M>,O�p�T�2"�ҕ*���:aÀp�|2�'�P�b'��P�NI�q�"m7������D�/�\A��j8&��9'�4day��	�����Qzx�n�l�� �"Ox�	��Re_nm�wCJ,2a��"O|���.&�-�1!��=�.��q"Oܹ8qA���a{3�/I�$�D����F�I{�v��A�@�B�VM�����F8((=���&(�һJ���C�M7Ky���ȓv��mPt�^�z�C�M��<s8�ȓw�43w�WWB 9SC��:��'�TG{��$]19i�$��K�����f+�#L��z����}�� U0X�֜I���i��� �"O�����`oi��퍬���"O�:�E�?��Ea�,Tj����"O@�q�����"�QG�A�"OJ|kgj@4�("AG�H8����O���
/ "E!�)Ec�d�bb�c7�	Fy�'�(�F��#&B�!RH��3(%[�';��
�Q3���;�l�-��	��'z�raK�/D�4�A��y���O(���O>�O�>� ��L5�D�%b�/Q���֪%D�\��$����$�f�%�%�#D����IΝ+E��*��U�z]q4�"LO�㟔�Qv4�ܛR��z��թ D�L{㮐��2�����M�U�G�2D������0|<4��MY�u�ri�PC��hO?��%̒h(򠏢}���p%��`Z�	ğ0��ٟ�Ҋ��'���j-�x���'Ϋ#9�Ps���y��� ظQJ�ݩhl�����B��0>�I>I��W%L76uhfb�+`�658�C�V<���R�d0�˲w�ScMO�[����.O8�����	����v�*2��l`��Y 3��C�I�5�0���
��tF��l� 	�
B�	p~�u�4N%z@�3$�j4 b��D{J|*r&�t����E
��<f��2�g�z�<��I#=��B�G
H�leڠ��]�<����I��8{q
X�ޭrg��Q�<�5L�,ޡ��l�V��E�@(��xLѣ
h�JT��0;�x!,̛�y"ɒ>4�Z��4��v6��RAc\��y� Ҷ@�Z|ˑg!qn��1��ʘ'<ў��~�I�&�t���a�:�Hq���y
� |��0�
���bȨ�P��',�Oh�g�Ehb�@G���&�H��"Ob �!��K����h�]M,���"Ot|A���CY(uB&_<dL�t���Io�O��D25@"1Hs�^!PZ����$,O�К�A� ��pGd��-���SC�Oj)Dz���F� IЅ���E@�x���.X2!�@(2�q�L	!��M�ċB.�'{Q�h�?�VjU�0!�q�M'D-r����H�<UL��9� !sf��R��+���z�<��όjR�T�	�@QCF�v�<�n��d�ܻ�CM j2�BW��g�<#�ƜD>�;�*G9��#�Za�<��.đr��$�2霞<@ Y�6e�Y�<�C��,g�&��Z��1Y�<Ǭ�3[����)	�^���*n�<!Qd</�� ��F0�S%�m�<�S�P*]F8JF�(c�ҕJDJZf�<1F��'b�� MP�SӰ�k��l�<! ��$^�,����3L�#4��f�<��k�A�@����Ń���ڦ�~�<9��=���.�C���J�s�<�σ:/�@��7
�pp�*���d�<�Fa0v��)�3f�$la��X�<�7�6�6uAE�� ��i�7ʕY�<�7g�
3ݪ؇�X.Y�`�����I�<�u�
�B�f���*�����MC�<	��K��lʄ�yb,��A�<A"偷��y:�@��~�򅙄��|�<9	�P��$���["-l�p���{�<!�g�z`��b!�>�6-�s*Sy�<AE�S�"�\̣��1i��+`B\�<���A-v����P�Z�PU˅��n�<�S)L/��P���{V�p�weSF�<��
��1�}+�F�g��	��@�<y�/��vD�2`84��2��^@�<��	��'fF��eC0.�����m�F�<���M���ͻ�
ٮ?i���JW[�<y��SH&Y��n�-m8�ե	[�<A��C�Z]�������	��[q�<9���h= b&߉-�6�Y�/C�<�`���k�nA�g��Ǿ���NC�<��o�?vw�X�wM�%.�p�a�%IW�<a"��F\���%y����Q�<�5A'��8��C�'fȳh�q�<�� ��N�ɋ�M�"L�	Q�V�<�5l��6�����K�4���a�J��ԃ����}����.f�2e��Ā�������g����("D�(�F�9lT 4���q���!��/D��P�аi���a�jY��+D�`!�m��
���!�w��Aa�&D��3 �c��=Ct
�6@�e�S
$D��sp�>WЌh���������#D�,��F3V��R'"�j@>�-D��2"��@��Z��;I��,���!D��aa�R�w0<�S��I�|�!g?D�:jP���nB-P�:�J`�ޡFS�C䉎pBP�QN�*8!F\�Я�iC��`񼴓u�P�3@m�V��/s��B�I'QΕ:�`��UlLi�TB �z_jB�I�V��7��F���j�ċ6�B��2{���Ӡ��,E9	ZGC$"PB�ɧ=��CgЎ;���P�k^�&B䉥/�,\���.5��X��W0B�)� L�B/�} � 
������"Odx�����{�+��u���Yb"O4u�5��y�L(��e�y�T�H�"O|J �%S��3bI�I�r!*�"O�x�R��������:������?F�t�Ó>o�}K���٠oP;|��I�?m�q�s0���%k�����0��&8D����'.�Ԉ� �+t6f��&�=������T��a�=}z�O�|2-A�\���ЌШ�>LK�'�<���9\0+n�d�� ��%���2���#(<;f��/ha���p�|�T%�)`:�ׄߋ�y����r��.ª	��a1�Q	=�p�:�'P]�T��Z�Z���$��@�f��}%J4�/�"Q<K�W��+�#�Oԝ"��_GLm[�!Y~�C-��F	�y�0�U4q�`��aӪ�"�H�n ���<�}j�ߕv޹)��atX�ŧ�|�'�Z��O�2ɖ�)��̏J���]Y^��b��a�>�[V�����EE	-r��B�h4��x�B��VՒ�F�VҀ�c���yB�:``Q%�̺>�����i:�����*��q*׋/�L����\w�����e�v���	�`|�8��U�)�$��
��!3�'ӟ\���új c������Q�W�u"�U�6�i�F��e;H6��c)��}&���
���a1�?G�L��).�q�g�\.��ԭ�t�j���b_�{>��Eb�;E�T�h��)	/��I��K&z2LJGkΑI;�-AR�Ĉ�ޒ$�#(
lP �SPӸ^{�X�����c4ж�8u�;�I{�fK&N<`��MJ�P�ք �Cصa�L�����|���G혅��JA}G�� �:R:��i��Y	]���פЊ���Ï���Z?u `mݩ~� Ze��k� Y!!��>�x Ǭ��Ql8Y�&�Ӗ8���M@s�ax҉N�~����))DxP	޽R���4��*+�씊bD�s���KKЈL�p���hN+-KjtBW)޽Q������
�@��ƮA�
V��+a#�/4)����D�; @A�O~�֬ �
�?V�:�� ��!Vz�$��ԵEk:!1!B��X9*�G�
Z}+Tf���6�̔�Qy�0���5Dh<-!(BJ��F��,J2ꁑ`"�D����I��c��X���ɚ;�b�˅�G>6TH�!��:���S��,�&E�f�;f��iӄ"�!:��RHh��7O.�=�#ޓ.� M�Fo��d��}�L��&��KDyӤ��`y@���k�8=�t�2E^���v{@0�v�IJe(����lu(g�� m�"	� �uD� a㉔�N�#�C1{�d�˒0�R�jA ���Q��g���s�>L۔�RI�X�q����u�c91���$Y���e)�y�(�#���5��ɦ99�m�@��+����B�".GRȲ���?`�����.�k.n5��Dį-�j�C�N��(������x�u�tg[){}|#ƍ��'�ѷLQ7Hz������d�
���{�A�4��xuTsf��$����՜Ol�b���-�(��e�Q~R�J�S�a���ʽ&�ޡ�s�	�n_�xpE��^����(|aEI������뗔|WB����Y����{P	�I�~A��%U/□�)<���Ȅ�y[TѤO��� o�͠�ΐ7����/��	��e8�L��[�U#1N\/����po����å��v�ӕ&� ���lQ�M�����d�!g��}Q2o�
Z����-O�	b���$�
J�c�?�:��ƪ<4F�P1$(A!$=@�cjj���;��C�R��<�<��^w��i�%��`q��C��P�"�Lb�������D�"?��m�8{T��N��,(b� 8��q (Z�f(�xK�M�2���3��Q��E@&�δ4�xxQC/��9��I`��ۇc.�dC-G4���C	^.0$�`�9)E�q�$dQ�hФO����Ƞ (�񘡅F$lYG��;k�� ��Tr`���߱N�����z�(+�jV�9�t�_�:���
0&&��v�^3J����+��'�0�!䎄0j�y�clǏh ���C�@�N0��X8�dܘS�8� �	���5`�]��G�k:��sN�FtX���c�A,"t�ê��	$z8�6'�);r=�B��?�^В˓2Q����d
P�2Y�#o��V@�`LL(E��iՍ�4:��	�J���Ĩ�k�@����Rt���.IVX��<�z]0��rw(͂��'�~U
 ��su,��	���4
�잀$��e����}j���H ��!��O����Ȏ(Èj!�#��M�D!\�~m���BlH��RqA�؛����`��j1`�˕�d������'n�E�7K� T���o�PEV����5J��Cŉ]�^a�C"I�`N�1C�=v<B��eH�?&�:�D�7L��S�C�K̓A���t�>B��L�s��I�~a�ON�� Z�2��Ѫ���{��i�w��[yR+ҢVE�1@֠�8�(�PЍ }0���3)�e	�]˃ϓ �<�G�Xx��ڄ�B�g�UKD���a���H$4��Q7G�y��q�\��4��c�YS��ɤ�	W��N-(܋�b�BbHC��i�����N�	+t��D�L��,ç�ٷ2�]a5�\�x0J���ϱ~��e�p��Sʵ؇���K���w*X�<�}1U ��y2L�є�33��@�Qi�wOz����NS\ȇ�I�vLp���X�HXH�sSn�$m�h�"'c�JA$(��"U�g�Z���j�(v7j$��D�)"V�{�/8m�j�
�ǀLN>�r�=f�P��V�ƫY�p���~K�9��+ظc���<����9`��<ȅ� �<<x�㗤ܒk���S����\�V�;#�>�Q��(;����Ǒ#��R�Ҿ�t��1#.:{E`�I�!�.�C�*��1��O�`�%�W
�0���!��hjʽ���η_�nU����+MB��f\	>"�P��V	�6��!Ţmaҙ���c���(c��`x�Ǿ1�&Y�tG�B�Z��)Ά�t�3��RNvayB��,k�R ځ�oj&�:*y����F���(��FR�!j������M;d�P$��TJ%$îV�ͣ�C�}���3\���u��L������ē�����!�W1 8EG(�¼� ��2Bc�MA� H�E��^�[�/�(&?���$�˂E"L`����v������MO��Bń�Z�C׿ƈ�`�-�)Qx�|���U�Q(M�,0{hSE
T^�'�\U0U�ӶVN��!����?��tl�ed�
Db��t���JG�ޥJv�A�D-��1p)��>��x1T�ܨan
�b�]_}��
$l��7�
1�bK.;?��!@A)C�,�j3�i�Rx���&0p�(�SlDz���X|f�A�A�W��(���6_)�E�㝋<��Ae�z�H�5�X�2̙���YT?I� �,�4A�nĞT���թ~[�t�`$�����8��##�T��E	4Mv��@��ɦ�z$W�V��6��(l2&�V������G'`�p	�	��
�&W�j>��H$b\?U�Љ5��t���#�h�FĒC��N(h��҆DO�@*�cЀ,�j�����"8GI�tJ��(�tɺ@�#3>U8T��% 9��![�0�I��=��ύ1#��[��˳���2 A���s�!��S� �)+�O�4-��s��˳���s����u�0;���`dR����F�t��WN�12R�<q�&�:
�|�c_wOҡ;���+H���'��)җh�G�:xCnP%'����4�W1���#��R�3�QB�jM�O�j9��[:G�<=��&����tI׳���cD/K�"<\x�S #-Jlx���3��$�c�;�Ba⅄C��1�'8Pt�C��J���2v����,�>̎�stn��X���x1��P�ҍ�s�	<C�d�5-��2�B�J܋=Ɇ�[�G[���x��@�Z�α!�
��L�� �˵d��*@:�y��H2Ťl��n��&�L7�40�lK5�u׃�*�(	,*s|�s�φI��Z%��$����gV�A�v0X���)Tְ�
�hI캃��P<	\4�Bڟ��/ƶ+��}(�b_
�f��$o҇�tD��)c*����+�.K�6A��6)��YxV�	�|�����dd����C �a{���n�j��҃Q�Xd��7E]fT���F�A,5���5�b#·F6�� �T����\C��9c@�5_s��A�/�[T,1���[5Xq�eG��d�%��XK��#�T�\{��	!���YU�D����y!�"�6z^@\��M�y�w��(H���5�~���<�u'B� l����FI
�p� ��}�ꦏ 4On��˰
�W�W�j������pH[@j "��QQ�-��k��lI��ճ �뮌;,�e:GȑvTeX�C@������O8�S���
�Pf��"�sTH�9�"4���de��9qK[S��,@@�7�x(�����Y��ȀGrqs� �"�ٱP�ۚ�u��� ^���~�2�M l�rIe��=G>=a�JP5/4���ΗT�N����Q�]�bc��o�bmX�+Կ8O*)i��P4-1� �1��l��yWm� PBj���lZ6&��v!q�r-:u�VϟlG��fN~��v�
3 �p�i�g� <��Ir���nG�8s"�'{�	�#�\%B�r��S�"�b�)1':��u$�	mB�I�0���ލ	� �-M�Yp��'a�-����z�"P�لv��I�sm��k@b�I����W�ƑA��JF��%x�.IP��0S����,i4�s��@E�1Q�ܽ 
�E��0'�HQ��${�ܙR���v���(HadB,mp��带�#d}�sE�B�QS�نx�pRᖴ<UP�*�������ѨH/^�ҁv!	Ej&�P�� ��Ԣ*:bH�h�f���!�!HɬX�����	��		9)�<���NyP��.B����1�� Gl>Ix�� ���T��$�@����Dmh��K,F�������q|�
6��%b�� �� �xyv`0W���eH�Rfx�'�����̍oO�� G�(at�0����'�����d��Ev�b��w�tUy2��hG���$Ʋ/ll�P'�ה#�k�g�PL�/ǖ�%I�� n�fIΓi�ztьQ�PPH��/6�đRW`���'a�Dd�AE �"irM�e��'^�N [�X&V[&�U����(�����҆�^,�I��녑�$����j�5cɊ^�  :B�z�y�f?�$�x�)0��\>���U�B�1�*,�G �c� 6IZ
R��K���g���g�������&�0a�I!s��BI�R��<;![�p��\S!�ߤI���
�"˿y�<f��09�Q�t��-f!�̛���a�,�S���L���J���>|�R���>	�m��HA�H��Ȱ+\zC�D�� �a�t����x��ɱ'�>�F���f��K~n�f,��E�J�u��]����@F$$A���,WJ��H�L�t� ���c ��z��
r��u�.�BA.�NM>,#�m���J4ЙR&�,NE���l�#�
,u�P�y���y���p7)N���K-_^JPӐj�3h���X����@�EŶ�P��I� ����+�/[U^H��
T�l���`��cWJ����b���wA��O,��p*�Kͺ�r�'�;(�2=K¯C��E���yr�l;�	ʂ��``S�� $����'�4��ȑlN�4� !�Jzx�Xs�	ˀ��|Pm҂ ���mژ#�.`;1�� rwf�{Um��R�)m�7��-b�'�Rܦ�5a%�4Lk���sqt�#��=Q��b--Kq|@���"?@)� ��<x���'�@t
��ctC�=��#�O{LT�Iz����1�<	�����Ǡ�<ZY����U����j#~���e�j�R5x�����1��'�c���=��=���'I�p�@1<!�_��nZg�'� �c U��D���S	I9�	�l�:d����(�,��$c͓g�r��&]�>O.Q�")�
I6�(Y���u��OܪX�t�[�.7��qvh�9W� 	Aׇ���hOHT�FM�1�!r����KJ��9��E�kٶ��aE7s)�@!�W;��.�\9�f!D�p/�dq'C֍>Ŧ��m�lRp3��Ns:t���,��+�F��a�T&�����)
�2��14牊o��	�� A�e��1� �Y<��vJك(�<
u�$�J6��a������u��<r�M�fnΐQ�o�j�JT��!q�0�*�F̙e����3��+Yp-#Faj��2r���p9���b���f�E���ڭ&-N�S�*]z5{�ᝇk��ZR�v=�u�GQ^$����-.���Õ~kjp���D mY�ErL�P���H3b��1���=��ӕg	<H�2��FZfa�ը Z�Zt���ӳb��	�&�9��E牽H�0ם^�:M���D�8��ɲ�ҩB� �>�)S5�X��I�8�>�r�h�Z�6��Cj��R�u"5���G38q�Am�?��pMP�T���#�CR����C�ʖS�����0�Fh�PWl��S#�ZT"�k�#�$���:R�O<غR�ݢ6�<Y/�n�����¬)��-�Q������΍`��(���!+R�xsI�B��s�TO�h#�"2�ny�LN3a{�� �dL���'��K�M~�H� Aɷ�n����A;W��`��H�Q̖���i�:.���t��f�9QZ�lC��)r��Kp�".i�����4Qat�b7�A�FayE��h�Du[%G&k�DءsɅ�Wݺ<����6Vrrm�F�D�9�R�:Um
MPQ�'V$l�Z�ك)�,WТ�w$�7TpTq;�
�i��	���Gz�tu1b�'�b�';���e8Q՚)�2曽R(\��J��F\2�b�Aʾ/n��;U℣]�d9*���e���暿V.V�M?M��M��� �\��H�<O\)�#Ș��\((�ɂ��P��H�89BF���Y3
�Xʧ*��x�����1�D30��������H�K_�K��,33NQ���GB��(O<�a���/��,�GD�+�$��@�'*��Z1HI�xIZ���J�8�O���JE!�'5rIhC���4��(d�Q�S;d�$�6�� cC��1�v"������5�:�j&G��H9��+W�	�?I�bx6p�4C:s/�������0� ��GC'N4��ϻ����TFV�PR֜Z��G�gaTP���31/��Hv/ԕ1-��7�L}�
5�
]36�zxq��݀|Z�8����1��)K���4'�%�g�A�陏�?qDʜ�3*v`�����`�Y(�D|�Ȕ�u`DȐ�%�-:&��S>���N�:�ni�1��]�,ݙc�L�^d�Ѓ#��$�������<l��]�:�ў�p��_ ��ݓł��z�J"o���$-^-lдH��U�x��OfƄ8�+T}�V�3o���l���d�Ra&�Z@�<5�)�z-
��d�4x����5�3e����g(K�l�E���O�!��?@\�l�Ԩ�=MO����I�`��E�7�y��Tz^̓K_;DHj��t�հ?i��(1�`
�c���]
���`�Ľ#��Χ>�Jq�^'5���Y�I�p=�t"��*��OvRʒ"�8ƆH���J�"2��ONh0��М&�K|���D�N3EbR�Ԯ$���Y����D��$cѤ'@�
�IϚSA�E�g�'Y�+�mX0qv` ���P� M���`Jߏ
�qO�(A������x>���W0��է�%,0������]R�r�qF�9�LP�|�|4-Wu�a��8"1O�e� �Å9 ��i�(Z<z6��`����.�$
͸)���(�Da6l :)�!�խ(X9r�/�8m����x������QSM�BȆ��çP�����Q@�rq!2ʎV�p��:H`�AJPD�@"0s���� �<!cA	J��5d���}��=sEPD�d+-u�H���V���?��ĽrT�!Ă����I-I��$��@�+��r��'�dh��eI4F�8�ib.]�/LD�M>ars�h�
y���$�/�̠�� P��˶���I��~rN�$@�
((Ve�';JF����4.�x��f$�x�<�V�[�b��h�Q�˒�h[�s�`B�I���S��<��CңN�`B�	���\@��]�Wb\�D�� cB�ɸwj�s�FTȈ[��3@��C�I�b*f#R:=��P�"��pȤC�	�-���)0(Ml��81�1z��C�I5��Q1��b�P���XB��{E(�r'��Z�U(7d�)�:B�I�T��eږ$M�(�$�y��\��B��	a+�u��fCI�2]���[%4��B�I��
�2���McT�k�d�S��B䉧B�Θ�*&Y(i�3.J?Pa��A�'r�1��u�H@bâ�,%�~���' l 9�w�����5Y�qB	�'��$2��OzT��w��pVE�ʓ���p�N��[�NW�F����ȓY��cqg�8>��[Gϻ
����$X@�x&�&EYPx�&'��#�>P���Z�#��;B�d���ǆ*@N��ȓ3�@���e��R�4�
T*�?e�v��ȓeZ��'��r��
�Ӵ#P΍���ȁ@	�z��Mx�* 6j��̆��(�B���_�ţVZ�lsb!�ȓ]Ǣ��,W�ﲄ#�d^w�D5�� 6���E�
w�Ģ �BX.�ȓ$�
eiBAϩ)���:���zu@�ȓ��X�Պ���t��*�E�<I�GQ7�y:-�[.�7ǔI�<��*eg�(X���i���s��@�<���;G/�Xh2��q�scTC�<a��AS@T��@���\ʗoz�<�|V����	�  2TDT{�<�4O�!� @�`Θ��Asg�w�<��/N s�>�,X0p��Y�-�{�<I�,�?͈�fB�=Z]��0� �i�<�iEA�L5`�.١(���y��Uk�<� <�ာ�Hμ�U�CKi�e��"O8p��<�$S������x�"Ot�S�-@!N�LA�E��m��eF"O8i+W�� kU�`#6	�6=y��"O0Mj0FS/F#�d��/��(A�"O>�aڴ�L�`G�2 q��,D��v@G$��dy�,�'>c�?D���pD0t ā��Q�-��"�F!D���L �Jߊ=+Pm	�Q��tS�5�(Q>����'-��0��L����υ�(�\����O/�	�`�C �8ը4n�.�r 2���m�8�3�Oj���N1$L��U��3D iX��	�Dt�5!0BǬ(�$���¥sp�'P ��K!%J�!A�"O �*�	w���d��0�
�K�ON�{vGX�0R�y���0|*��pLR4X2��/�,���s�<��IVla!�^�9��`i�#�2}|��(�����J�Y��OQ������26��D
��4��o��p�!��
KZ���҅'(� �ڳ{��[�Ț�6m�%����oJ�w��6mR�L�H)F���c���S�',|d� \�ˆ!�j��z�2G|�参/� �� X�@}L��B_>5���:~�@1�l�H!��N2x@��'A
A?djAu����'YVI+cnS)����Lڠ���'�0��Qꚪ:t�a�$�Jk[?��f�G#oC
Ahѱ|�%q�B�;7p �FD�53�	�!R؞d��)G�ԙA
�$oZ�UQ��t\�	���A2�VY��g�ĐH�ے5(��bH���Yr���< r�������.dA"�.�O�,9 ��XK�ez�)@]�0�F�N~�F�%"����Em*A�Ԡ��i�q"��_��~bh�!N�0�×3�٣6��Bܓt��Y�JAA��@@�ʅ�Ƹq�M�����G���0�͇�C;vL��ݗG t��p��#Ǥh?�]1�!0�d��
��A��<M$�C�K�m�&���)�4 ��̊CC9!�r��f��ē�f��B���ѩa�=3!������7}t�a��ݺ�[�b��G d�w W��0<��˼?�T�딄�@����������(��MO��$���:���: o��=�Z���ۍG� ��ʛ�����hP�DY~�9��܃l���i.�	� �FҦL
q
�}�SgM�2�"�+�kP�zY���)<�Q��`P�v���1H��,�R�#^	 �wAX�pA�M��;�YѠ �;w���!H��k�x�R��V�pA�+˱)3���OT���W�g[vD	Mԏ"]$2��(fMq����D��F�2����؋Ԅ6O�ch	+0J�����M�c��9��3���1o�
ސ�OF������Z8ᖃ��Hr'!�;}���.j3���@a�%vV���oX��T$��#ظ|
����z�bYS�<tyZ��B��l� ��G��1�:�7��+ٮ�V��;��On49�)�$)�@�H�NT镎���Y�2*��C,d�Ī�Y��Q�@�'(�P�R��CׅB�B�����ۓAXP�IEG�h�X${W�ǲR,��>	��՘P~��F�İsbv ;�b�-���Q
{Q�[$o��F����A3TY���E��E��ܸ@X,,!FjK#��$2�H�"��-Y4e��d�J��HO%R��Ȃ�f�� �O�uML <(��Q�`��<@�$j^\�� ��Bؙ&����
\9fHҰ��	�h��Ѧ��h\�Е#Ƨ	�� �P�G:d����aEY0vP���O��p��I�8�0��c��m�$�x�������^�Mz�iA��*N""$�` �f��Y��A�ħ��!�j����&9j�T� �@���!ߩtb̄�Ʃ ���ISA�TP8���1w��y���4�,ե �HҒ�`�gۜ�ƬIc��UV4�����ĉ�'�?mps䛦h�Z(z�+>�u{�)o�aF~�Ѣ"H}��욁D�"Xi�-ӴT]lH1reYG�@=[D ĩ<^����$U�QPNU0CX���3-^ltA���B�L)c�`+:S�!��%��'�p�$��-���b4���6�`�I�h���F�e,�P�#Z�o�dQ���Z�p( q�b=��&�M4E
��ѱ��/.{� 2$��`t����Ȫ"��"FHr� A�6@����ȋ-+p��O���D\d��Yu&��/0*���iN��PFn_Tb�����#s�!��\�`��5�ƚ�,6,$�!���nC�x�@
�S�����ȫdF^Q3���	���Y ȫik��Zv�'H�(�O�yCP�n+rl�篝�9��� ޶��0�b��|�ȥ�S���<qp��m-rd��+?���K��C5rf0�p�U-@�J��Ԡ><Od8�@͕�A�N����eK0��?'�:a��c��c]j��U�X it��#"-R�=5�4
�%�>^Ռ	�vg�= �.I�3cL"a[d��5-Xkq�Q`���<(��A�@B��]��G7�I!HªL���O����G&iZ�E�Y�0���� F�C��?v��G���S�n91��3&�3� ��rW����J�P�=�'e�UjJ����Xq0�U�P�LiH�4���ܪT�<T� M2OgR�� Aӓ��$�6� ��-�=d9��±�Ɠ���A�: �J�{cY,�x�`����<�E�LZ��@�B/��)�-��f�(_nҰ�uI��/���"OP�d����͚^��T�r��-��qƙ(_b���eg9"$��3�H"A�0р-[tT���Ɋs��ӡP-1d8��bF[�a���Y�7�"3&/m�ej��*+��!s��.6j$��'c�����02��@KE�umh�`�˂� 384�
ϓuon�[h)�qሗeq��J�@K1�8�RDLn�n�q�c�p�4��O�/M� ���85I�`������Mk�`�i��Qt� �Q-�x���%&��;���#I�`�9��ʣiM��a/Qw��h��bF5Ys>�A����`i�0$��F�`	� l������V
I\D��"ɘQ P[�;f}��d%@�z%���|
� n��)T�z�N���fĤ5.�X'��RU�7-D)=nFHB� �P~x�Y1	U�y�H��f��06���޺4�@;�S ̼���[C'ID[8��N2 ��3�/��4uay��)4�*�ǃ
jR����O�?5���#N�{3�,�F��k�f�#Co��McP/F�#٢@�c�_/}i�=�FM�t<\��!Li�hdYs�Q�4rҼ�I<����Mh�O�ٻ�ō�E�����&~�9��ʖ�	����k4�`PB��j�j9� ]�W�~I�&�L��?��
�z� �ɖ�j7��pBMC�̖L榑k'�Z�o�ZtB@4e�n�?�f.�9ia�[	
K���h�F���n� J�V�(B+�DT�8���K�R��m�&����EMi�N��nT�O�L�p�[�L����i�z�K�㇒HA
� A��-$ѣfK�><z,m�B(�����'�z���%���Ao8Dxʷ�n�H%Em(ca�u�7��('������R�$�j�ݕz�6��b�O���f��25��s�ITc��H��HD� �-Ph�t�O�S8���$�Q�A���"�i����J��MS�P.��\��H��9Z��"o޿ ���١"�)�`�b.T/p�����O�AQd��w�j��$�?ڧ} t� ����`i��ΝoV�;T#�ƞ$P�F�t���ᶥ@�A2�������h89WmO�kQ�+\w?&KRLK��ʨ��F!{<���G˜eϠ����`�҃�
|C��	�O�Τ;�i�y:�����eϤ�`��;<����>sh�DRG��_	@��sC�u���#W�&q����d��2�ܺ�؉�	|�<0Q�G��#��R<1׬a�c*\&n�~E2d�νW�<�;cڇ;��u����&E��;O��2Ҫe�C�\�l�lar��B�­ȶ	1*w�E�q�ۏw5�1j�\n݀4��g�6��Pg�����H�vmF�o1����葨r^�83�d�)�6�9!E$P`L8W%L1VA&�Ѳ���X\:� GvY�,���*�8�a!�事�ܕ7�Di��CW�H�Ԅ���kx�21��'H<v�Ɉ?2p� V�_�]���I�ސ��ajzםk�*혥��|�R�+�+^�L�`��bC�a!QI�S�h��¥���-FDY�뎔-Y(�ds�E�b�_ !��\6C6����H�%Q�`�ΕIS�� M  qɤ��_
a6̝0H&5�@җN��!Ѡ�V�)h]�q:����e�	K���EQ��\=����J�J��'@�.����Lg?I��>.iX`CΜ#bxEp"�_'F� �bF4c��J��� ��az�	P�(eFX�Ν!f~UXB)_%B�1�"�D4wU���M�a&x)�!��Q�JMcwŝ�`��h"悖 ZV�:E촟 ��s��B`�([�������}#��ab�>Bk�(��O�R$���Vb�![r��4d�����
0�Rd{Sċ�~�ҰI��<�@$�qm����KԞ}���2�cF7q�$��I��@��0��;� �I���e�ϼ[ov5����:TA�t��_����M�FL.�Z�$��z;��w.B�h��h8D�(tJ�͢��~�2�f�m�5�P�]�?��l� e�S$[X�r�,��$��� V
S�0Y���D.r�x�0�I@d�0*�%_L�'l��!��� T�Q����$J�T�|̻­���D� �,O���(�k�.�Ĭ(��'�>�(x� 5��%1Kyl���'\�jZ��7IR�X[�-�I8(y��y��D={����]�Oq|��2�]e@����\��R(�p�h�2�L!�y�ɭ �� Z-G�%��4ʀ�gy(�4��kS��b�*Da���D��1�;v�@13F�,{���䉳�Ҍ�	��7kT��2'MO�$�a퍹r�R(A3�.~��qq�G�#i�@X��X�A������H7qt0 ��>IW�ɐf��8�L�$",k���pR�8�@F��N���N3,��Cb���64��X�)���ˏ5,�(Rp�C��*�E.X�
#��p�B�O>8������ ���{qz@�6LR�S��������}���F�l�2mh� A�~������~{j\�f�P��g
Y�|p(��̶#�Tb���SP�w��@;�HkB�#B�:(�!�'6tx ���O4=�f�����J��N�u\И�1�SiB�9M�(��TG�L*� ��D���:Pl��sWļ�Ʈ�q�V�
�j9��G�j� �(A�Z�<�@+"u$���Ќ���O ����Q��a���� #��@�d8:`Z)�A
Y'L���R �#Ef������]����'[j���9>jL�
ؤJ���B�XM�r�2F��*"4p�r�B�d�v���'��:f�f�T��e�~�b2�G(2&�&(֮J�d��#J\,���Bf|��p�+;�����CW�0�@��V�
�����^4�a\��:�O�~`�'��1`����+�NB����N�'{��(k6J����T�$�X�nD����3d�����KI�����|����J�c��Hˇ(��>(�	uIȟ*��!���}���h���	�@����;b�vhx�#A ���)I�}$�sfO�36Pipi��D�ѩ'!S�d�lD(3���K�:ކY���C`�ZshҤ����73��r��d�Y��<Ҕ	�x9�T�5��)����X<��Z6^z�!�� �ءW-Ţ ��u�U��q!�ܦ��'g��0��#X����4�]�]�.(��V���Q�!��C�"uke�ƺ4�vqP�͟،�`���Y v9B'T&Dh�E+���Y�e@ƒ&~V�I�@�&X�ք��3�<�ʏ!0�~��a8�%��I!��06̥��O�p*�g�<)[���({�U`����	�)�vM:��A8W��u� �>SZ^QU"�'���B�68u8����Ѧ�h��߱V+D��VNf��b���=���
�gh�;@*�7^V8���	�q���:���3%�08���@��dz��O�9����.Mb����J�cD��ܲ{o���t�.L���{BP1,��SW.����!h�~g �v�Nxh���)	�xŀ�F 2�u1f�[v�pjBCƣ\;�QXwd ���+��0�$&�W����ՙm�V�(����4I2�نLԄ;>�aS]�����"���ɑ�> �����T�-ې̀a���3��
T0\1�Mh=a`ӇǾ�u��
P8L���1����#44��:��B�Ou��#��3Z��{����g�@�Fe̽&<:�5�ILZ������C�����S�ܨ����l�j[^�niuX?���� �"x��6j�	��1j���?Q,k"���h���H����"ѳ��?I!bQ�BFQ��#��cI� c���'꽠$�*J�!W`�0�䅐�NL!"%/�4��)���>bt���M]M~�؉��36�<��f�;X��=�4�%^%[@㉃9ov��U�My�ة�b԰2�8����@����W`s�S}�^,1��	:q:��:�a45 0m���T�K�C��fci��!����k�I�Q��$Z6��~z��q��>#�n�@��fda���tf�3�̜�PwQ@%ٕmO������'�6��R�	/o|ޘ���$Klڤ��C:+����g�H���x��3c$U�v�!��-O���7��80A����F��j���x����Dؓ5�n� ���8��y�FKU��-iS��Uȃ��k��a����O=�\�s*2"g�� ��jE�ȝ��p!Р[`�B"G�(R����� �?	 ��d�P���{%䔋`P��c��1<��|ж���TEN�FEI�2� ���L�j���3��U	d^��k�, 2<��L��N?VAJ=Ӡi^;rI����0��l�B�,O�4��ǲ#&�]��96��� Ső<�j=xb�DL��@�0d�Ԝ�c�ׁ#QP�x��̛ �� f���S5��IֆAwXt[&/Z����#(	��(O�8x���LX3��������X>U��
�2���`5�Ù���kFM�Ω c�N�Pn&�)A�[>dAZ��q)ĜGyB.֛K��	��� ������?��h�nTTbЍ��eB$�ya�~R$��ˌ` ݮ3������U�@��p�[�#�.8Д��9/��BJTiX��T��C��uڔ�K�7!fpc���C \u��'L���+��5CiJ�j�F�]�D�˸0)xD�u����_�R���!ADH���2�O�Yc�H�¸��Q�� �5K?J�Y��͸}pђ�@J0Y����#d�	�ؔ����/��Oе���p1�hK4@`ZP�ɣ�� X��#>�6���n�T(آl
�8||�,��s�#�Ml�ux��P�h��Q��o0%?�<�D�߅b���&��'.���	��hO<ԓ� �����;'��42�O�xh����L�Y�&����I�!Y&�X�u�����G��(x��
@68a�P�Y�gf�!d��6��}�J@��h�1t��8+���i��a�\�']�U�κ��CU@	X��,B�ݗEF�k�ˊ�a�9J�@�$�92�^,�&P`؟���q�4lp�\�^�f-���C_�j�S��C'��ѥ*�z#$H�eK��D�>xP�G]�'�?�f@Ĵ0�X�#khѨ�s�	�^�'�Ƹ{u#L,4�A'>]I�a��u���%��:e����˗gpS��ZW�VK�~D��3�I����s�J��i���I5q�Tt�O���v��긧���8f.�Tʕϝ,IX@�Hޟ-������?P��RD@�6�����	c��P�"�2	���fNC1��>!�j�&!��`�l�0�r�tPTK�jyeɱ���3G[!�$�y/0�a�O��`�&�!���oM�Č�|�D	_�C��tc
�'��B��H�g/&��J�#4�d���c����5�Kw��pe�F�g�Q(f��<�v��pd�����}b�ē2v4K�&��Y��=�Ʃ�-��?�@�3�y	r-@6vѹ�(�7����uR;�O��6���[���X���0@�0�'Nl��rBYr�Mj4  -��Pl�Q{aH�K��1�ȓI�����ב�@�X3�Es��H���6��v�X�h$�� q�݅�$�(%� ��g�1�q�KkWؽ��:p��XE�^�O�A��H�"	�Ʌ�+��l8�"R�R���z�GM&D�I��	~]��K�u���vbա5��ȓt"����jY��j��S�Eu����ȓ�L�0-�Z\jY��D�=���ȓ �<�㠈">ζ�U�վnԄ�;�H`�giM!5��� 81x�0��h�H��1��F@��7b@:=�؄�E�@F�)8i��4 ��|���ȓ&a���]�d�2��v��nЇȓ!�\�W�V�^�^0�˟2��l��yhD�f�T�KU�L9�M�*(%2Y�ȓP�ܵX�'�
����NI�]����ȓ	pI����-.m���������&*\�����,?������*4t��ȓZ�����b>"L���[T�Ą�f�Tm�%NC�#�i���a�.<��Fib��#�U�^��0Q���1� ��!֔B�Nؑ(��aұ�B L<�ȓ48��0~�\���E�'�(9�ȓ@]��ݜZ��K4�8$u�D��.��b���=t���
���������n��I8bGx����5�qC6o��[9��S�O* ل-�>��m�f%D<Z4�1��BMٰ$��6nW�)���*��F2/�e
�lZSKx Q�H��|q�3�S�O��L{�o\)QT,:��Q9���'�X扱���h�jE��� �Z���lC�&�҉�b��!�(���%�)�'B�d�CA0C�l����V�p<q+�h����'<u�}�`�8��	�@;|��D��Fe��b�{�"�,67���(;�(�ħ��I��nI����C�Cх�zX�ɔ�a�ͼd=YI�"}
b-�.1������˻d�H���@�a�5f�4xq��>E�� Px�r���*�dK��Z�X�b1*ŷ)�ڬ��!�S�O�|�87#ʍM5�wQ�͸Ȣ�s2���~��dY�3�[q�±m bRM���HOV��i�"7�����*����D-YU��O�!GzJ?��αY�V&��3qp��d.���s�$�����x�S��*�E$H<(z�V䗂7&��'@�-�''����-a~�{� �P�h���.u��7}�KWJ}��i+^����s�"��B�+R�'�xA�'S��񅊫�����d���T���/NYz�!�0I���<�1�Q��0|�`k�,&����)���Х%�A�ɩ���ص0�����sgO����Uǉ�?+�I�GY��o�(:O���<E�d�%t����Έ.A2��Î��M��^�t%�"jkP/A�&d�Fj
J���SUy��x��*��<cS엶vBd�;
T����'��ɉRa�S�O�
��D�
.�6�����*,)`�*O��L<IG���jT:�>�ɭIM��Z�W�Y0���	�~ޢB�	�=��!�J�,%U��; JG��dB�	���Wa�J��� F��B��q��D�	T\[^�
���?i)�B�ɋ8&t9���/r{.��͐��vB�I(y�"0`J>NK
ȶd�6�FB�	�N������L��)��lN2.:B�Ic�Չ�KS-~�e����.��C�	�b�4��l�d��dR�MD�(� C�	,=q�t )[�$̚$��*D�R`B��}��4���J�6�ܑu�( :B�I)lb�)G��8���@�(�^f�C��cvP�	A�3 ����͙�f��C���q�ҘST����W d]�C�	�<��re� J`��ԯ�I�B�I�O�6-J�A�o�@�1�h�r8vB�.WV"�hG͊�3��8���k�:B�ɨU�)1C�
��K3L�(�C�ɷH��q.�9�1�v']���C�I�'�Z��C�L�JZ|q�R��C�	�D�FE��E�4`$ͺ0y\C�I�.%�dլ"4���d��] C�I>hF����H����,C�	�r��E`��V�L�Hq)^�&C�	���9��j�����T��}�0C�	�!=Dx�%g�8s�-�g�6&�B�ɷ6}½�2�W�[�b�ke�؁?1�B䉒;[�1�$D/}�-��S-ÊB䉊|�	Q���rR��i��^1�bB�ɰo�)zb.�@�zc�̝0�rC��*7�z��P%̋cV���ܩ�pC��-?�������C@a�@��'�ZC�5!86��o�#%49V�J	T�&C��<YS�m ��˵��Pת˺O�B�IRY�����F���J��H�)H:B�	%H�����/�Z�����FB��=�h��1���p��g�G�n�8B�	�p�Ћf�)J�B1cwm�5Y� B�	�R����ʕ�zQ@�Q́�G�C�I42`;+�5\�ب�CM�z׬C䉭@%�PPD5|>� ����$r��C�I>���t'�z�pp#�
,tXC䉢�a	�"��2�cA(/w*C�	����d�ؚf� 23����B�	�e\�S���^,ܕ;f��vB�# 	�J�	&,Oν��i�XB�I�R�H4�2��s����b���6�RB�I"Fr���D�'~2М�,B.T��C��y��5��g����c����C�)� $�@�ECQ��Q3� 3fC��6"O��Ƞˇ�	�,xꌒ0AP�@"O�p�G�>Dţ�	�+.z��T"O�H)��P$����@	�(q#"O0��3�W�`cnݣ�M�vx���C"O�����|rm�T�A��0��"O!"�WҖ��Ӫ��	yb�ʁ"OE ��H�v5�#	��x_ Z�"O.�I�Ѣz�:8Z�n�� L�(�1"O���d�ܠ|�Ը$Β���`�"OR�B�K��m�3��A��`U"O&�����)1�l� c�
�Y�b�w"O�A�AK�P��H�n��Q��"O�����'Z��R	��fI��"O��p�
Lf�(��$��:7�8h�"O8L�!�` P���
y7�Mxd"O���9R~|4Ad匑:Ui�"O�t���D�/R00���6l�%�"O��1(�'}S~a(C�Z�heE"OF�B�)�'����ь�~D|�I"O�P�p�2��C�7[3��"O���#b�H#ΰ���(���"O�x�Ӊ�#�>y	�.�X'0�@�"O�:#�_�2��X��Q	���Y�"Oh!� I$����v�݈2=w"OpH	�KG�[~���ƟXښ���"O>!����>!�2YrץE f<m#�"O^8�doʑ)q �"�D¨>���"O(���	�6����4a�rܦ��"O��K7����\	��O�E��� "O~�j��мz��%���,D����"O��i� � Y�y �� |:�G"O�hX�C�Dr$� �$$���V"O�;CK�w1�͡��ǵ�&}�@"O���'Ȫ����T�I)H��\i�"O��Ql��:�B\3�h_�}�B��$"OT4�#�4n�R-�w��^7^:�"O�	
P�ߨ{�|9��
`ح��"O8�B�G�?B_r�Z2FYW3n(��"O�HC��N���JAE�u,���"O�xA��4{OLj���aӁ3�!�'�85;�LکE�����:�!���{wx��Fn�=4�N� g!��O8�p�C%��s�V�(��!�$�)+��� �"�Tiѣ�<�!�$\+ ?�QH2�ًM���9��ߙ�!�DH,J!@�6{�ޝ�S@�x�!���L��Ui�Y�5ب4YS�]!��2��0�Ֆ0���o�x�!�ػ��`"f��v�i��	O��!��9��}x'iR%zJ��M�&nN!�D־'6�;�
�%�H$��l½�!򤆇}��ăCb�)��,"�K[�!���0%FA��*]	��ۥKI7-�!�K�g�aRW�>p���C@M[4!�d�,DS�U�C-ڑ>I0����;1!�#.�H]2��I�6h�@d �N !��Ϭ�L�#H��?�Z���L�d�!�����	AD�K��@��tI�'W�`���~��z���t*MB
�'�ƴ��ǝ�,i�-�!�M	
�V�z�'����q� #08\�	�G��QX�5"�'��5c�oT 2f<S�*�?N���':.���ė6KW$�+1 "I2� ���� ����7qZ,ǀJR����f"O���U���)��
�#6UT8"O ���fq҂=z�k]�\jr�"OV Q��y��æ��0jKr0AE"O�� �,I�\������0E�I�"O0����=T*:�)��݉:LU�@"O�])�O\����ж�@�a ܕ@"OJ��&�ۮZ(%yU������"Or�)��Y�#�X�u�¹{��9"Oz�Q�6f��À��G݄X:�"O~���h��![��S-gl� �"O0HQͭ'�n�(V$ڋZ�\9�"O^yac��s{@�@�H��f-H=�"Ol�sdďe�����(���"O�}p���+;�`G��6��Q�C"O x�ӆ�Kl����L��J��$�"O�<wi�L���~��Q"O�`��U�l�L�3tig��ɀ�"OD0�MGK�,Xr�70� ��"O���e��u��P����zU"OP��d��>٢��Ԣ�mo��j�"O�85Ce�Hm�Ǩ��)T�)��"OdH�3��[�}2��=BX�iu"O����� T�\�I��\I/^��"O@���;�fm	Х̽r><�ȗ"Oj��ȶ�d�g�S̄rG"OC�
P�N��ț��ˤ%�(zD"O4�k�͎41vI㰮_�<�t"O\l��m �v*=!e�ѽ_0h)�"O>H��G["@{6�hQ�S�UX�X��"O0m9��ۂ'�D�y���ZL���P"O��k6��.Hpad�O4(��H�"O�	 K ��� �,E�z��@"Ox��f�OP���`Зn�8y�"O�P���=:�p�rQ��(��I)a"O0�"1��(�\�3�
�e4��`"O|����- ;,șԧoy!�$�/V��I�D!J�����A�.m!�D�WkP;��`r�堧f�F!�U,NH����O�T�t`�"e�~�!���J� ��FN#�~������!��^/P� !F�m�\��a"&BT!���

 ��ć�Q�D�f���=I!�$�-�<��֮�2�$�'��)6T!�$؛a��hB�6LK n��$�!��
RA.�
ą
�T�V��An�W�!�H<����é��!��Ș/4I�!�7l�ZKHFB'ʔ��ޚN�!�X�^kl����(m$r��ڵi�!�$χF`,MaV��c��,!���d|!�@_Ҁ0d�L�g�*���o�2ih!��68L��� S�"xD)�R茹1!�䝻XQ���	�����Ȣ�� I!��^�-�(m��R"@>��b�m�Q`!��,g5��
CCj2��a�m��tS!��.����%D��LT�9!�%8jE��0���B�q�!�D(G�&���NZ,4)Rb�X�_�!�D��x��¡�M7(����B8Qu!�҂1��kS�<Cw܈p+zEi�ȓs��9�)�R�q`F@�>���E,��KF�}Ôhc���>t@E��'����%b��u����b�1]��k�'��qh~T|�jҊK�.� ̨��� zu�"Ǻ��ء$��0KE���"O\P%d¼}��蚳B蕹"O�|aeo�231�8dGL�a��a@�"Oڐ�H�4f�C!\�#��5�y¨�&:��E�l�	h!"Y�cD
�y�H��X�V)a���\e�D�c�R3�y���`ܬ���_�Q>$V��y���(c��(@�L�O��YcrBŅ�yRH*~L�5�� Q�A�����Ǌ�yR��>�D��B09��u�B��y�k#1*�A�d
*'$�rʷ�y�酓!Ȳ�s ������O��y�KխrH�zf�O�i��E�E=�y���
^�EIẅ,s���0��Y��y�E/	�X]�p�ͦ N�����yB�̂�i����Mz����y��=G%�(JP)Q�4E �kkA �Py2NB�O��H���W*J����%��l�<��ʓ�Oi\���ۣW�t���a�<)��6LY�B%ILH}(e�EU�<�ń: 0  ��   E  �  Z     �,  �7  LB  �K  -W  �_  �e  2l  ~r  �x    H�  ��  ˑ  �  Q�  ��  ت  �  `�  ��  ��  ��  "�  ��  ��  �  ��  �  �	 � �  �#  İ���	����Zv)C�'ll\�0BL[H<yVCQ��F��e�P(������C�<��	��e��A��+O��$���X@�<�v�C��p�TJ��izsf�a�<�&	�P����w�&H�ؐ���e�<�0i�������^z��B�V�<��(��Fz,Q��!\:�\U�N�R�<yӅ�I~��3��,}��٣�JVy�<a㇊)nt��;G�ʏ���b��Kv�<i�B�r�8��L	�W6�}�=T��zf���R]��0/�6őf?D�haV���  ʔ ݿ���1D��[�
(m����@!\	{�� 7�.D��`ƭ�}`|��a˚t���Q3)-D�[2�ߌ=�v!����ɳ� 8D�t���O�u|D�Z��Y�P�1c��7D�LÐmֱlGfPb��U̮L,�0C�I�[mH=�W�٠d��C�l�&9�dC�IMM^� a!1�>�Ie�?`'�B�	5Jy�]��tn`���JF}��B�	�v�6��V�+#*t�c2H�`��B�ɦr9\�{��*v�h��⡍��vC�I�v��ɐ�ƙ$�P(˅��=EItC�I��9��ǟ l�����&2lC�IO��P��(����'�lZ@C�I�aS����k��p,rI�3%�`B䉅%���Gk�S�X�z'.�#�C䉙U���@
��K�V�j6.����B�I6\�qi��-d@��4�\�Y�B�|�d���a϶l	Ҭ����_��C䉈-�I�����NL�,�ب�E�8D�l�C�*&�n�h��Ώh�YS�j!D�h�$�$!��0*$�b�p��� D��3�X(q~T�אFbv��K!D�ȩrMY>n��ڵ��$V�$�P�5D�l;'N��d�MJ�6[EHS�%D�����£j|)��f�}�� �L?D�,q�
ۨP>&@���S�b��K� !$�,ö�ǵzB` ֬B�R�%ˣE��y҂��K���( Ǡ^���y�����yb�[�Wr	���[�N%�H�FK��y��֊s,f܀ GäA��$�+�y��)�i:���L���T�tgV�C���F2��mB1��/ce�,����v�*B�I�[�D�5 �c��X��8<��C�I�;Pus�KG6K:�<ȡ�G�n��C䉸{�����	sǸ|������'����O1���$�T�0o�;y-���`C\4]���U 6���'4�Ӌ� � �o�&cq�=ٰ��=>�7��O8c�XF��'��Z@E�>��*E��j�^L��'������LW�����X����&�1��x�B��E��L3�j�+F�|�(`
���ո'ǉ'G���|���jP�4|PH8-�C䉯nO
�s����eh̳�(����MCO<��O��j�HX�>����&��8?"�ї�'_Q���N��f�p���x�H�4L-D��{$�]%�u�mŨ!�Ti��,D�رf�&(��ˠ��g
Bq
��*D��&㜤4m��Z���1.O�2Fm*�O��R�Oa�y+S�ɗw6�(���@E� *
�'_8��c��pe,Q���L�����1O���@}}rN8�?�q+��Q6��?EH���˜Pnʽ��	�a7�'���77��O�_�ܩ�M�N�^I'��E{����
/mx���bϡp�L|2BOR�����'f�#}� ��YZ7��PFm� g/f�"O*8ӄ5�(J���7/���|��'i"���O�����%��3�=��'�����+~k�	b�(����'`��22���Ym�r��:=�a��'��e�T$�Y�L����|s�@��'-$�9�k�3fy�)�bcL�*��q��'t6���]�Ԁ�	� z��C
�'�j�;�T�:�s'c�B� XI<ь��I��!9����(��+@.�A"!�č({��5�'�6C?������WqO�����m�b��j0}[�C�e���R�z���)��'D��=BQ`��M��C�Q|�S֐�\�I��W��C�	�k�� g,ݎO�y2ǀ!^�C�ɠyk�
eț�K��[���>��'4ў�?Q�晒0X����/�.�T(SP�6D���SD�&J�L=
��,4�ve⒎.D�H*f נc֮U��ƪ��a"�o+D��8��	Bn��%�2�P̘��O�<9�>@����F(@*�
��<�� ��(��9�ݗ0�����fC�<�$�Ϡ}f��u�	="8����x�<��ZnI�` pd< vѰWe�p�<�A%�j�ڐ�t �;=8�����u�<�7L�g_VB��E:�,�hN�h�<���)?���"֦I3;X�]HF	�[�<�V�ة2���:�\,TMF(&�l�<y#���"ِU�Ҫ)X\aC�)Dd�< ��p<j�$���	
d�<YF\�,M4�N�<8E���daE�<Qq��o��a��m�He{���<���O0��Tf��'���C~�<Њ��f���%�C|؞c�`z�<9քi,�iu�*q&=`5Xw�<)��P%[�ŹsO�+�8��v�<A5m����I��2`�8DpjOIX���O��s嘫H)f #���+	����"O�9jB��"C��S��S�ej'��*�0|�ţ�0���!DI5\�Ir��t�<mF=(�4Չ�`�pt�A˖�EE{���i�v4H��'DHĤau*ڵ~����'����Sˑ�Z,D��$��xT�%��O����@3C �)�>��<��.\��!�d����v�ŏ5	�DM�$�!�Y@np#'j�=��ȳ@��@�!�d��(0Ɖ�u68a�C��T�!�d�4Q���S*W�ܠ�i!�!�d��iT�	)�%�l��1�r�;�!�d�=�h�p���g�4�"G���!�]#7[r�IG`W&	����r S�az���B�Q
��G+�[����ϗ"y�!�$�?^$�k#��7��)C�N��1O�=�|�k���}�B�R<e�E�x�<�dV�>p̓t�Ї;X�"�����'��𙟠���W��\3�܅0��I�L!D���F�7N�H}��o��
i,x���#D��˳b��0��`��	Xy֔�	 <O�7�#��'8�(��vk /�}��i�4o�C�+Q{��7��$)�����'Q���IR}��O ��>�#a�H7'���	�jڌP�A��%D�ؚ��$�j�ۖ�K	8M� `�@$D��'�w^�|��MՂ4W� 8�F7D��
���~�f��,�j�p��ʿ�|�
�S�? �d�TA�5Jey��.Q*8���w~Ҽi̛��x�'�� �X�K�#:�"p�p�@��yҨQ?���C�*�"�A%ƏE���'�ў�>Aؐ��j��Q�ӆ���Hc�+�O��ɥ�)��Hʪ5�ک
��6an�B�I�!���5#�Dwz��U��ji��|k�xGx��	�z��i´��(y<V�A�'^'�!��?�P�5q�ޘ�4&��	�a{�X�;!,��s��Z�d8c e����7O�`���PM�����O,U@q�"ON9�`�A	\�J2�B�t�汉��'��f�|�d�� p(1g�	��Y��e��sNb�=E���aP��I��t��c돣B+F�G}"��uG��� +[]WVʒ��?�~q�'{a�!�+�F���ߨ'�R�f����y/J�j&�$z�N΂�u(�GM��yO�=}�����Q��H��V��'��{R��0�����P 2��i��ŗ�y�e�%�`�s�H�0�H��4NR��yrW�����<%��/-���A�.��m�Y2��V�'�qO�맴M��3�B�8!�@�R������ .�ȓ���P�K�Y�J�3�P�z��0�>!�����GÔU�d݋ �ؒXI��%��y�(�.�XQ��lP�e ��v�Y��y�jC�-6ސjp�/]jh�f*?�y2�I�:{.�)0�]!L� Y����yrMV�F���a�DU5*  ���4�y)Q�(�p��է_Q��XQ��Y��yBk�r�;��]3O�p#����y������5j��768�K����yr�
�A�Lj��Ǩd�����E!�y"�u��T�%��F>Hi�H2�y"O3&LDj�!���a��yR��?��J�핽={�BT��y�+�@���с�E�wf`�1���y�霓3�b��V	LB6�HX����y�+d��C���=%�n��!V��y�&G�MI�t,S/$�$иF���y�+;$�X��ek~5:I�1�y����E5\T��]3`�`uy��	��y�&SnAu�RZ)d�����yB�3��R�ؿ#�&	 ��р�y"m 7r+b�h%��5e�<Y��-�yb'��2�(1�Q$���B'�y2'���>1Ci�=*^�2�ն�yrc_�&r��ֈE�6�n �D��y��$6=�hE�ʵ(Ek`}B�m=jѵ��4gց F	�$O�:B�I���P@ʖi^Xp�y�FC�	;Ǭpу�����UMǣ6��C�IF�|����I(4a(��f�jB�ɜ5S.�����?6x��A'N`�0B�	�5o���K@�3��!�6�4m�BC�	I�z(	jU;خ����L�d�6C�I7����G�2��xÂ5"�B�2������$0��!��e�#R�B�	23΀�h�#�-��gF/:fJC�	+ɪ����K� 	%١���X�6C�o(��g��}R����\8E~C�I3}c�ı��^��֜2Ůĳ/K�B�ɳo��"��-zך�*q�G�N��B�	� �dHz��&],~H8�aG�M�^B�?KN��hҮ�u#Z� D+�=u�B�	7H��l�I�0N4T V.�m�B�)� V��P#B�)��àQ ���q"O��)4,ٯr>Bi1�o��<�D"O�����O�^��"�O�K���U"O�aat�_�X��y�ݸz���*O�-1gg�2/������T�\xp2�'p2�'b��'�"�'2��'���'L�E�񮈄3�Y���I\�lD�'�B�'<r�'b�'r�'��'���K_6$p4���� <x��j��'�2�'��'��'��'��'�d�(d�Yc`y��Έ0T��S�'�"�'���'�'8��'�'����-XQf�-��)�('#$mZ��'��'���'"�'YB�'��'���@c�� ʝ���S�Rl����'2�'F��'{b�'[��'2��'��ɉ��*%GB���i��'���'��'���'���'d��'��ᵦߪW6��R�e��	��'t��'��'	�' 2�'�B�'z(t@b(G�q]�]����+��'y�'�B�'���'���'b�'w�$j�f�H�V�"��T/��Z��'w�'�R�'�"�'���'2�'y�p��L$��b�Tv�  ��'���'�2�'���'��'��'��E��Iʆ�: �/[&�����'���'�R�'["�'�r�'�b�'��rbb[<xXd҃�;D���)��'YR�'���'��'�T6�J��m�I�l�E�^�>�p�Ǝy�&��G$[~B�'��'9B�2�y��'��7m;p�Nܙ����G��gÏe�N��:O.�n-�E$���ܴ�?���Y^�f�N�W�Ԋ�*0՚��Α;)r�'hL��a�i���O����D_�-�2Q������J�\p� ��c�ȑAE�[��?)O*�}*u��#N� 8�wO	=$��h�Wǃ�L���J^$Ƙ'��jxlz޹!匹kg��jF}�F &,���M3a�i���>�|"���M#�'�p�	��0v-{d�bL��'۬���$V�kF:ĉ@�i>���+W�I�aC޼4�晣����RҞ��tyr�|�.aӆ������ �Q�f׀�
kR�_������O��m��M��'|��+>����'����c��' �n�";`=KF��~F"��|�����u���O8�bRn_\Ġ��
r���S��<y)O���s�t#� �8bhL�f)�����p��s��	ڴ1��'^7�.�i>�`�Sa4�h�
u��p�;ݴ{��v�'� \�6�i��I
���If� B^���eU*$X��1�(J��l<[���D.�iӑ��z��0JĴk�0,�c�=��-�����ܸC,N��p��h4��0n�(����Ą�(y��ɔ�K�-��U�J��p=�EǱh=����(�8v�u���R�eUb,�6�̫v��(#�^ A����9x�lʶ��,^���P�W�ym̃�Ő�*��Z$�.��u�6�96$�i
A�ϵs-�����]�`�r��Ý������!�$��ի��7*��b�)D-I0%��:O�b��J]�ꮔ1c\=_��#��q��՟��i>=�O��BV��1I�PY+%�L����ֶi�2�'A�U*��4� �'�<�T�I�I���(����!x�����a��ǟ|���?ݘL<��-�� �%�P�M��m��F�jf@�Z��iU�Ep�����0��M� ��ɂ�H� NQ�8a��~]6��Of���O�A��/f�i>������	0��ZQ*��w"ن¸����d�O4��y�1O���O�D-{i��!��ͱ"���Dʉ=s�lZ��h۠J܃���|����?y*O��iw/ؑ7�>8�f�Ih�CF���I�{:�c�(��ܟT�ImyRc��2nT�� Nm�h<@�$�r��Zc(%��O(���Oʓ�?��=-���O�
[�"`[$Â7}�xg�T��?����?�-O4SEA�|`�:�s�Ɉ>�@�"�b]G}2�'"�'����4�	�u�B�MӼ���*n���9�m�-X�*`�'���'BQ�$�3���'-��1�gk�5��T�֣*8pb�i�b�'��I���	���c?y@�o���Nɲ��ETu9X`�`Ӯ�d�O6˓L��� ���'-�\c`�4bwf[=2f���GZ8�.���4��$�O�� VG>��s�p	P�	]"2�����"S&W�3w�i�剐yv.%���2��������]�'��u��Og����0���+c�p���O���j�<ͧ�?��g≥�2�+ۼ~�J��BȅC�`6�'(�ho�������l������|���œ%0f�T�D�L�,Qa��-LK�f�?���ʟh�I�?c�L��"@px���0H�BEϒp�ȸ��4�?y���?�ף�#Y�����'Dr�͹c��a�b�V�E�*�
� �'
�D��?��[fM�<����?I�K��쑅��~e�UZקҽ�FY��i��	��M�6�O�d�O��d�_�t�OZM*W�Ո:��<�F8Y�ҙAuW��$"k���I�p�Iǟ�Im���	=fT X{���+[��A56p,�jb����O��$�OxM�O��	ğ��U�&� ���Q��&�è|���|y�OD'q�2�'��'���a�D�2a�	�9����TN����F20
�7��O��d�OL�d�O��?�vo��|r���3�2-�5�K	���5��78śF�'�"�'��'e�ië+��7��O����<}|�A� ��}Paki��Bi�o�͟D�I�Ж'6b��1����'q���/�lE�˅f�� i�$?@�V�'���'�"��h]j7��O�$�O����� Z�Yp��y"���0M�9#��enZ��,�'�IX�����|��M� bd��F?���*)��f�^�Q1�ir�'P��+W p�����O~�����I�O�a9%�[�Q�М��@�x'l�AS��Q}��'�|({r�'%��'����O��'��Ta댺g�6\����2�Ҙo��F>|�Jߴ�?9���?�������?A��!Uz�:��̤!n,�"��1ZH{�i�\)�&�'Z�P��P�ş��� ��]��i#U�&�����ؙ�Mk��?���� ���iB�'"�'�Zw�b�ǣ�|ߤ|2w��3>��޴�?Q*O��{�?O���x�	�·�݇+v,{'�K�q0ٸ㉇6�M���C7 E)�i7��'b�'����~�G2�bhyŇݰ^L��3�c���d��N��<����?!���?)��2�J�$z,�gk� .us�욂����'R�'/���~�/O\���H,2s��p!�M�R�	6#tТ噟��Iݟ����ЖO``yj!�v�J,��	SVQ�Kg�I�g�91TJIꦹ��ҟ�����,�Idy��'lM��O�:Dk�I��
�D�^� ���T�>����'�R�'6§�~��O��N����'tBI�3+�����Nb�i����/\7��O��D�O���?1B��|���~R
��x��c�Q<�m��j�<�M���?!��?a�C�Q���'o�'����@N��� �U5|���*ށ#Ȁ6M�O�ʓ�?)�Ȃ�|����?�� �|nڪs�9w��>�v��P��h6M�O���5��æ��I����?-�ɟ��^�/��x�� )Vv��A#"R-����OzI[�O�Oz���O����?���O�F���j֕G<R������4]L��*��i�"�'b�O]���'R�'�(%�q��.Ҥ��D��lP@�)��Ӓ�d�O��$�<ͧ��'�?aRW�cNv�)?�I�A-�9>
���'���'r,HG(a�����OB�d�O�t>Ixg��'&�:ax�h G#�dj��}�|�:���Q2o[�<�O��d�'�r� 6b���1U��%M�����'��_�7�ͦ�P�R�M����?���?i�U?���5�$!�H�z��&Uz��'�X��'���'���'K2X>��0�V,{(��cWpהA"��O�(�pe��4�?���?��d[�_y�'�|�	%��rδ8�⛣I��H��.U��y��'(��'���'���'�b��f@uӆq��˄ W5����EVPM�aAK�A�I��L��ݟl��Ky"�'��P���5f�� d�0��c-ŴIh�Ae!���M��7�RXS��?��Z?鑲��M;���?Y�L��Gܨ !!Iv��M�bhE J����'1��'�����THR�n>����@�
���8,�A��:qKN l�Z��r��O����O��W�Ri�l��|���������I0���R46���O62Y2��ߴ�?!)O��d�:��	�O^��|nZ�J�ѱ"��<!�:�փ�>36��O���PcϚ�mϟX��֟ �S�?��	E�ڵ�FL �e�i�����l��O��D
����4��i��STϏ�TB',(2v�Ii�J~ӖM�ACæ��Iߟ����?����� �	�8� V"H|jU�F�¡̈�%��$�M�R Q5�?	����4�(��P�$�?���N_��l�D�1X�z-l����۟�Su�S�MK��?!���?��Ӻ[eQ� �L��tn[�>�4%I��%�	iyB���yʟ��d�O��DQ�l�z �f�!5��S��U�Q#6�oZ͟`��o���M{���?����?u_?I��bM�k K� �Z,�����>�X�'��k�'X����ßd�Iӟ�t@U)a��	���	�R�5#_	7�Hu	޴�?���?!��&��[yR�'�` ���e�^�i�: 3->�I��?����?���?Y-�T�Q�KXϦy �}?�y�����Dn��4c���M����?Q��?Y����d�O��zr=�kl߲`?:�1h�9L����^54���9>�.9�I����	�d�0$�&�M���?Y�W+~z����Ǟ$w�9K�o�,����'��'v�	矰Ò�f>��'c
+"�=
�^�ra�R�
��s�Tr�'7��'�,��Luӌ���O����`�bm�3l��KD��t ��+����i�	Nyr�'F�`��O>ɧ�ܴR��� gc�:E&���W��n������!�ݑ�4�?Q��?Q���*�>���hC�KC@�&g�~ ȺX�X�I.c(��	쟀���d�~�ᯕ0kA�ɻ1��˒%�g���@�I��Mc���?�������?����?�$,QMB�����˰5<pc�[�6�� D0YxR�'a"i������D�O��$��D�� Xda3�7Oiz���a����O���D"��0�' �	џ,�h8����Հ8[���d	6�qm�֟��'��xӜ��I�Ox��?e:�&�g���*eR�zr�Di��i����	-kRA�'s�	���'rZck>tȁ�2>���Y��˕,��!Z�O��y13O�ʓ�?���?����?�@�ޞ3�T�V�V� ��5d)I ����i���'�2�'�6���D�O�D��L#V����2:�TC���K5�D�<����?A���?I��tXiP�ig��!�4[t����q��ňvz���D�O����O��Ģ<A��W��}Χ	q\����ȑc�p� 'A*��x�R���I�����\��:
�X �ش�?���o\R�0�茌^f� ����<D1��i'��'�bX����k�N��������厄/n�9��
?b��Pl�ȟ8��\y��6�J������:���ײ<��c5����.z��}�I۟X��6���Ip�~��%�R���R� �2�a��⦹�'�����Fl�\,�O/2�O����KEZ]��k⢐�`��8n�����I�zP��	U�)�"5©��R�x���%�JV�6���Z�o�p�I՟@�S��ē�?�nJH�i�vƁ�O(�@k�(�Lc�6�ː�yҙ|�O���'l��'��� �H�f�X���U.*����i���'��![.�O8�$�O|���(7�A!g�;v�v,8�E�7fP7-&��XrΠ&>������~��܁��B!K��� �P�up�ݴ�?�ǃ�9%�'v�'Zɧ5v�L�-"�E#	T0�*,B��V���ĉ&4��ı<����?)����P�z/�	c��@?�Q����@p��ן��	E�ן��I���P�A
	�Z%��Ԏ,���K��G՟��'>�'{�R���WG[���eGgNM�c�6�j��ɬ����O���7���O���B]�d��5������5 �6y��
�Yb
h�'�2�'pBP�,���<�ħ{���' -}�p���=M �P�i��|r�'�2Ɲ�y��>����u�v��`eݳ%�afcL���	䟨�'3�`1��?�i�O����$x�8���:b'�yx��#^P��'�"�'�b��<�OR��32�1���ȃl��(
r�6m�<�R�&��v
�~�������|�"L�!R]�6�P0\Kr�i��dӆ��O���L�O^�O���)@&-�*h�JH�A��Nhp�i�H*�z����O�����Y'���3i�D��2��>�na�����0%�R۴R�4)����S�O�Hː\�"��S6Sв��#��';`�6��O�d�O\)Q��Z�I��<�	b?��K�Txz�{�C,B�4�j�m�ݦy'���D���'�?����?��e�KY�M�%J����j�h�yZ�V�'����P5���O���:���f�! �VC��q��.oh�	�]�젶��̟h�'R�'�U�`!��Ll����8D��QƏ�p��D�H<���?	L>��?yeL�8t9��P�jpv��$遑lv���K>���?i����D�rHb�ͧWs�-cu/��w���7HI?�|��'~�'Z�'�'��b��'�0���9�@�4���I&��>���?�����dNE	ȅ%>����0I�
ei��Q�8�b���M���䓪?�s���Γ��ɋ4q��K��*'��a�"�'��6�O����<��ؙL��O*b�Oa�]�q��4�P��]6=wRh��&��O����5���5�T?�j��U�����%gv8[��y�V�d�O�P�,�ǦQ�	�@���?�SşTi�@S�i�����Ϝ-z�d8�������Oґ��O�O�	#��b3i���e��'s�l�ʷJĮ�M��˄!S���'��'����O�r�'�rOڕ*[��u��R�Q ��^�BH6�X2I�L�D�O<��|2M~��>x8���$i�4Ha���00�G�iv��'��D�?A�7��OX���OP���O�I�'R���ś#%ʊ$iEk
K����'��m��):A�2�t��l��RR!�BF��a�d���}n� �d.L����\{za)�'�wC�H����o��z��]�4�he��ڶG@h���҈zI,�r`)�zߌ�Kt盾i��\VG�&�*�
6O�Rc��;�)΂na|=2�,�V�<���ᖤ]�
�y��W�K?��3ꁵS�\�A͕�QMe5��6]�X��зlA`�ѭ(�
���Ι�xgq0 	Z��J���\t`Ũ�E�!����$�t\���Iȟ���,����	�|2�ꋃ(��H�'� D.x����:��9��ʐ������v�n��ޯ,���Ǘ(	m�"�B:j��@�<U��)sΨ�&�ǓR�T�I��M�Y�ԫf���|(�a:�	K�x{��+'�=�����I�8���y����	2R��Ф�l��C��#�M&Ϳ(H�wM'e^��s���<�*O\!GR}2�'��ӣC��E�	� ��/ѣ4C�p��!U�Q��ɟ|��bAIUΩc��U�/�� ��O�~�TX>5J�.J?7�����O3^T��%}�T(	`(bC�t�����F��Oz�i`bI��]>h��K�I��ТK�`��i�O*�)ڧ�?�∝F��q�^�T�X�e�]�<���/n�@�MR(02��V�����F�6~�ꄆ�G���4F�Z~�l����Iҟl�sj�6{�L�	۟���ҟ�]�2�0���U�D1DTYta���<\`�C�js��scH�mxN"�^�g�(mN�)1���? `���"]�F5�%�"�Z��P!�n��ӥoT�Yc�e�*�fف5���y'oE9��)����ܨ	�"+$�B���IH�O�2ړu��"$(EB��N�51<!�ȓ)�HH �O0z�&gI��VD���?Y �i>��ILyB5&��	�"el2T2�EW��s�䀍'���'qr�'��]�H�I�|�u��Gw�a�� �a?�M��e��bd���߭l�Lx�֤M=^�P��	,<�8,br�R�wdzi끮 �E{*���n�9w�-y6B�-,�
HP��$��O���#O�f�lM0���3N�fM@��ܚZ��Mv�b�nZe�����	є�<0"R��3c1/B��"O|�b�c�����G�3�nѨt�������uy�--�`�'�?�5o�v�J�����J��8�	��?��
R��!���?�O��%��cEu��B�/ˎw��Ș�!�zA��wj�0�d�
c+FI8�D�1O�:@�$ 6(%�Йw���0�W)|�H������W�x@��?�����K?"����S@I�|����� ��,1O���䈩&��a�Q �}�&��҆4!�W֦� <u��Yd�j�G�歀���O�ʓ4d�৲i���'*��7@"M�	;|�y��&v�"*S�Z7H����ߟ �^��v�Eܤ,\v}�"���|����'l�a��@n�:Es��_��������S�
��]8��k�O����IH��P��ݶ[6EK�( ���Onqn�şh��|���\�V�&N`Th�3C	�l�*��#MğX��ş��Iwx��;g+��D�B8#�I�@���,O2�Ez���Re�����?�ѣf���:��?��=~�y�����?���?Q����	M��*��F�:c��4��B�Q���\10��l	ش2�Z�Ӧ�k�g��(n/^x#@gA�k����s�Y�N��0s���.4��(��iYI�#-b��QuW>���N�w ���0�&,[�b�'&��.m^��"uӚ(oZΟ�U�_ԟ�>��?QD��u'F��P'�9f��������x2��Kc�����Yk���V"��yR�'��#=	�@�,�?�*O���g���R���,��+k�:2�@�b$�ū���O����O(����C��?��O�LYIa��n�@8 �O� p(-��	#:���
@�8�ЙI�D=,O�@�a�C5~��P�r�X ��̂ ǀ&3�<|��N�<�̓r�E���qW!S�\�ve�wAi�]���@ՏBk,���$�j�;� �O<�l�-�M#�
.�1{5y"ro��8��h�f���)��Y�W����C.J�X0TׂA"1OhoZ�'|���}�f�d�O~A@��R%Z}r2�˄FS��	B��O�$ºN��$�O瓗HI�#���|2.HB�Za�DlZ$i[�)��!+�j֠+�]� ���r�^���ɑ)�!+�(M���#F�N�i._V��#�A�_�Z�'oY&��u��H!��p&�h�g�O�OT�� ��"|�4���r�*I# "O�X���Q)�y!u�
�؋��x�+eӈ̲�,ћ0���sd��>��(¬(�d̾(��l�ӟ8��O��K��`Nr�2X��i�f�Z7�����I���'� ɒ���N����(�*X��T>m�O�Tibş�Xb���WF'`ܠH��K1�Q���X����]BD�}�w+�3%(�2�`v�IJm�f��+0��C:���S�_����2&�*;=̱�Bg�f!�D� C*<�Bo�>3�\P5�Ђ3�ax.+ғ*A�ٷ�S�A#�Z��+��U:�i�R�'N��5x	~rs�'���'��w�D��L�o�lXB`�<j���� ��5��AkA:�) �1��A2���y�$�.&t��p�(*�4"d�ܧ  nm*���w����R䋻Km�qz��Ý�����`���B��`�8H2�
йseL1a��iM^�W�Ι�i>�r��TD �*ǽCk�(���2@Y�؄ȓi6���g���@�{%D08D�'�f"=Q��i��V��@���1`�����8>�@%�SA��ڱ!%Ɍ͟���ٟ��	��u��'�r0����J��Ld֑+�H�9d�x��$���M�*����3����Ě�N6~�B���F��)zv��?ھ�Kg��@�Riz��6|O�}D�$�
yE��
3qJөֈAB�p��m̟l�'�R�dI(�����5"F8;5���UE!��ԍ*�
l��.�� �0�3B
	�XT1O�Hp�'*剒g늡���:�ċ�	�u�M�T-TH8�h@�( ��d�Oh���O�Da>9
�`˪Z ��9��:IȄ�0�N8Bۈ=��;&��'�*"���[/�PP��瘸>����!T��<��~2>Գ�c1�̄*�i������J��$������O�ġ<y�+� �1��:��ʔ�c���IVx��	%�  Nt�Թ�_�(�N��W7�hO�צ�!'A	�'}�����A($l)PQ��؟0�'Y��U@�>1������9����^�T�"�"�4P(��-߻|��D�OEb��]�:�K@T�h�Ho�^��	�|´
�(#a���P�	�,���*��[����8  UZ���qP��`����!O�Iܮ,�����p
�U��V�qQ��^��i���d���i2ܴ�?Q����q�-���ës� ��D X���'��'	8yz�^	��0$ ��?G��p�i>�X���K�PW6�DJ1dpZeh���W�܀mZƟ�I���
�6δ\���4�I���]�[v��@PLC ̌�D�ө.x�(f�@�?�thD�"SK�UK�eX�'d,�r�V٫�8��p�'�W�x�� �n-M����N�f�[�`K]ܧP��Ld�P�$"�i�0`I��R7W��)�iIN6��O�(��m�Oq��I�T����w�rlc�/�$#�zE�l�Xh<!a��i�V���u]��Ih~"�$�?��xY���R�mZ9yDꚍ9�U��,=!�S-8ɨ���4�ޭ���-6!�d͓vr%b�I�5}̄y���"7(!�Ē4v/HA�F�n�&}c"!E%p"!�D�"t ze�V�vec� �~	!��Se�1�tO�2	
���t�!�� B)�c,�����:��X8�"O��Ф��<0���
��Dj�(��R"OB���ĳNa�!9�/&ܔ��"O�a�%]�۾�a�͟%��`kT"O*�3e��=/T0����$�b�"O\t��lB�F�x4{�,�06��)U"O<��B�O�(*�w���j���2e"O�;��OtЌ�됀��<Q�"O p� ]<�0�/��;�Zt��"O��;"��*��9�-�3Ol���"O2p�,�rt.}�u�"Od�b"O�"㡕2@�PV�ۀn�")B"O$�;�Q�N` ���dD��"O\ ��)	� �\� �^p�)Z3"O��>[�:$)D�>����#7D�T9�#*N�0��G��8C���j3D���׍�j1&�@7U�YC���� 7D�d)�� /epT�u@�"x�ܠ2�7D�4k�EW!S�2�-!qu�T�4"1D�0�e�c��;ר�cv�(�T�#D����fA�c�L�q��`�P�0O.D��Ş9iv���O�|Z\�� D��K��H2GK����O�QN��7�+D�L�c�&b����P�q����+D����v~���u���!ȕہb)D�{�g&���A��Td��")2D���C���j�~ɠR@�+ܵ�#0� <�J�����6�D-t�j%�0�Rې�9�"OP�4Cj��d�E��@WL��L,��oZ�l2(,C�O?7�£{��%�D�-�����k�,ў�p��d�ɏ���H~H�U��0b�bUq�A\6��dX�bo�I���Ob���� * f�c�ɛ�e`\%b��M��f�2��	Ħ�1����"��i�	 s3�����3T�5k
-r�E7O #A�<O`����,iv�z��J�p����}��8a����	�ez�I�[��11���8��I@��"��ӊm}n�ϓ	��� ��ê)�~�AG�~�l�hÀ	c���R#e�\��4��6}�N����T;F����o'��'@ ���3���HR6eRv)�D ��(l�"HȢD�e��	B���u��>�'P��*E(��otX	��j��U��RI8�N��P��Q��/,O��1���&A$P�A��U�"��A�>C�I��)�']`�s�H,P�Tm�$e����'���d��5�T�r��W�֨>�ĝ�#�A�}�t�ɜ
5��d~�[?s.��G�|��
��\��{�aZ�`�5a��K49�B���$D-�y�iJ� ��4c��[y~�	�
~���'Ƥ~���ř?�OT! �o��aW�6^|���з�F�O�̠���`��:ń�(bHq�g�,j���N���X����6#��OH�P%��4g��dT+=�؅K@Z�K�ڑ�Z�\l83���9l�$�%�mHi�ӓ�hP��\�kMpb`��-�P�k��b̓)�@�+���`�'	�fgI/�i��h�T(��ɡo]��0>A�D\.=kj��,��C^��H2B��P��@I2�hz�D��'� Ә'�7�  q��0RV�\�{ �T�aK�8x +W-9@��!v�	(\
|Ex��[�oC��s�HF���Y����1����8�B���8W��Y5�I�yp؈t d�b]��Zy+�1�5�|2�5�qO|�hӉ��~}��s3�n�d%�ȇ�v���ӏ�wCXA��FF�1ɧu��|�� ��d[0���p5ˀM�9~&p��_�Es��eG�LX����Bꈰ��-�ؑshΠ!�J�%�~���'�Z�ا��C<!h,�s)ņy�$ ��#(amЧ8��qy�Ǖ'�21i�@^�.K�<j�t��r.O�O���"9Ѻ-����3��saN!C�ȡ`O���r������O�	�N%;�&���>�f9��if(`�e[ ��#��lŞ5;�OT-��O.a)��s��JsJ��?�ǐx2�+\���äݾ~\�k���=��D ?fm��1�bO�G&�8���͉���'/�u��(
�Yli��::��5��*Mx��͆�0����a,,O&噀��oj�	°(U;@�B� VhB�I8����.�@��`>���Dx���\U+(�:��𺅊��0?AA���-�+� Z�<�f��" X����Fԟ���[�S�Ti0lY���B+������&��rd�A�޿%!xi���4�vɦ�R�+,Bt�-�C>'DqnZ�p���j$A\���w��2��%mڱ&�x���}����O=�O� Z9�g�xL]���-50N�h�]���g�Z=.Hl���O���D�DK�M�W�)j�`�C=S�*-��$
�8������ֱK<�1���ay��s9�M�a��H>$�h\ ��d���M�O�6���\R&�)jc�i�b�����`� �JڂY�XA3�'3^��nZ4�(0Y�͏4D����L�Di�=O��JGlΝn��O��K��q��L%fk`�!ū�2���"���m�Z�*D�#�r�֑��B	"�x��p�?�ɡjY��]sF5��) + ���';�h��C �(�9�I�+^�"�҉-QP���͜�<�h��O�u���
�Q̈���ë�?Y�Ϙ'Y���'1�&�8� _�-���ƶ-����l��3��t�f��1	�{2-�y�.��e�	�P�J���,�M�4gÅR�1O��ͧ29�&�x������욇^�r��E�Mq����I2A����!��U��\+P��?���g#L-cOz-kF)��y ^19���1�ߢ���|z�cI
I���l�?wE�I9tFV�h��F�r*�?�P�Q�!n���v���f�v�J?��dj�넥�q\�yQō[�2��ʓ.��P+cI�Jy9eI�l:`Gx"����*ӸS��xa`��R���G�;!2�9�I��SvM|��W�f7-U8V�l���k٬KwE�-[���as�޾<̸p�:����4t�"��hJ(ӎ��R���#�Na�!�<n��6���yr���e�A!؄&��M�������	�B��^������u����$�080:#���e�<�!��N�?�fi!�m�/Y'~Ъb�S��Sc�6�V��w��
84 �'�vH#�e��~Ѩ�OH�A�'B�O�@���,ǎ=v�ギUS�]x��i��H�>�#ד\�r՚��,
���+WV؍�Qj3?BkFŲ�z�V+��R�`A� tݹpa�ͨ��'�xD���ۘsP�}yu��,j�b�r�Wz9��;-˷W����'W���'T��*p�iQhA�.�e��p�%�7a>���2O)R�S��.W�R}
ۓY�L����8{t���2S�d�чq�B�l�~�K�ꈊ�+(����I�,x�0n�:l�n�ǔ�c���Ƀa@X�0��:D��B%�]�(�`B�˃ݘ'��`$��@!�M�h8aF�ۣC��A��ϝ_�M!n�b�pL(�K���O~�0� �YȊ,�5�@%x^��w�6�Ic���I>PJE^����'|����|�&��n�)�<�q�.��_�9�BSQ掭`�ϕ/�~���Pb�0sd�=.|��V��hOp(��]L��qǡX/9��x�C��p,��l�<7�����K<s[��s�X�(t�!9�l����1�-�:x7a}Zc�@Y;w"�`y��-U
5��j��y�ʙ�h]�F�α?�f)+!oK�g�>t��ɽ#���PRJζ(O�|�Vh�+������I_/���Ç(%)�����	�
o�U��ؚ1�|�P��]�8�o��y,�����k!!�T7vkK<�M�N(n�2���,msX�1��w��[ �R�Fh��j@J  ��IB4@��G�@҂�e�@�,��|&�Բ�, ��F��!Wf0B�JO�qt�(.�Zpۓ�ty�Rd!PB���@�
�P[ ){A��i���"נ�؎ʟG��w�h9S5� M�~��&
F���=�p�G�*"`�)F��47���Z��Pц�
/����OZ@�O^�3sY>�ha���vL�U�O� ��Î���Dz�fS�11e/&�I�C#��*��'O�|����ƦŦO\-3G(��q��`�d�~����328��JAB��:����-b����	��  AA��}��tI��_�\�h��	� P���ڳ"Y�d�S�ܴ�y��iL6�ȑ��0?��Q��N�<h*�l��\)���]�X�X��$
�I*{e]~�*��`���˔\��Dg�=��IP��ߵY����Bp�����7���B&�<|O.|1��K$�̴[��C*��kգ_�e��A��[�8�����^��?Y�'����@�?��է��ԡ%>a��(Cm�U�#H�45�d)FB<��Y����� * �kS�� yR��'��4�}u�T�ǅe� �)���#�@�S1 ex]X��ω��'��HAp��;vC�Q*2�S�� SA�4D7��a3��b���2�*}��	��o@6�ظb�Þ�RØASE��!ze�5���p=���!���)7靿*.4aCjN��O�Ts5��X�X�Z���@�:I#f_�!�V8[�N'�=�5�*'K����o`MS7,�L��m�(X-;-T�Pu�5C�}��6��$��s0��޺[���V���O'�,�蔳̆5���W�<����G�g�NY[��	'-�i�¡��i���B�E h����Do�0p޴�?	 �F����F�0FN�H:h�\��`�8hf�1�f ��)סZ�v��S�I�c@?r��g�/x�f�'���<Y-�#4X����K�3�I���EQ�<@G�E\�E9���T��%R(_�CfI�5�xa�&T!1�"��!HQ�$\�|�>��H��\AB�H�4TP��� Ū,��2��f������l4�(p���j���a�˛��V?E��O���N�D����#�,-i"��(u"�$bF��1a�� W$\��	d��1��){T��&�ʐ_:6�e[��d�٪���H$��q���+MV���&VQ����q��m�������Is`!�	l����h�����#K�Na�c쟿D]�P�ߣC��S���b�� `�镎�N�d�A��d�6)��	V�iX �iX����H
�q�tl��N� 8r�Q��O�Ra��PSBքxiTA����]w�6b�֝��6�YW���A����䛬8�1�`�9�O�4���Ő�I��%��%�$�X1rCr-m�pa�|�}Zw��7͏4�<�*R�̰�|�;*־ES!@�E�}9��Y%F�f�F\�@��@��E#Ę���/Q���X>#����y���A�O��16i
�K0Y��]�i�����?u�=c�F���*���M�4"' �!0�P i(O4�1Ԁ��<��x6��0�I�?�9�'Lt�3���l�F���(�M�����LC1z���f�?:�{2�&C�^��%�R�@�\<��
�5;�Ap�Or��Ħ�[�'�اu7��]z�OJ�l������% I��с(�O %S�/V'b^�����<�~i2�EHs؀4��Dް<�`웰|f� k�mߩZ<V�����	s�T���Q�E�I�_�(Q������)F��U���A�}K副<AT��*P���FH r|�H&k���@d���0
\.��D�8][�OJ�0JàN������	�p��i�Fh��P=��:4+�<N4�
��d[&.T�M(5��)Z���k�(R6e�d�Fmˤ�Ș�!�'Tvm	�n{\���I2v(���EmǶ0k���4�D�����F\ɕ�Ս=��(��'��0Sb�(42�9��P!�V���,J? (-�a`4Or	;�*�'&��xDaQ/C#�Zf�[i1#K�w�p�2�O�T~����ǥ��t����@�I˸@�/�>� ���i?�BF�&LLx�6��w���͘��e��/�ِ6�5c��OJȀGǝ�f*J��q�
5l��]!���,8���j��D?Y��Q��@�5b�J��=?�Q�B�Uo�1�&N-<6�Y� �G,_�.5Z�N#-b���g�'t����@\-��� 0䎚1��D��Ĵ�'��7-�ٟ��I~g��.��]��� � H����hj3����H6��Q���#5���e,{�0��fm��ѣƆAxH<ɱ��E�Dc'�2Ĺ��aĢ#xQ�,8�/�[�`A��X��l]����XK�Yi&B��U��}άe(��Ȕ&`�i2�I���hΓ�Me
F�f�����T�Q5��v���{���[><�P"O�A�D�ǟ<$䠑�I�ՠ��>�E+���@��ɡ{\x@B��/>i!Bor�~B�	=b��H��'�o6
�abJ;�JB�	<c�n��C*J3� 0��F�VxC䉂e��Q�5+�.n�X;& Q�B�	�+
�� B��f�$����+e�<C�	?v�T}�àԊ$�L�0sM�P� C��7:�����,4pz�a�:��B�	�p���
�7��9i��ֹ5q�B䉀�0����Q���h�%P���C�In~�a�[� i���%��)iHC䉤^2<��OM�2�Wa�~rFC�3W�°�E�r�H��0C
;�C�ɣp�5S�1{^��j��C�j��B䉺e���e HР��G���\4B��{NR�hD̫I���Sw��Vz�C�� �ɓ��U�j>�[��)�C��C�J�K�%IQh�
�lC�= �,E[4�������=�B��{oP���-
���N��B�ɯ0���uf(4b�1u�Z��fB�ɝ(�<x�v �l���(S��C�ɑ^@�E�P�$�8��*4�vC�ɹd�̙sԨP	|��ĸ�Ȓr�"C�ɚG���%���	����R'GP�B��)4��T{�E�3�j�ɖ�QGvB�I�D�R1zvHBa�k�'N/6֚C�I�"�4@�g�ٽ6��zPJ̹LL�B�	��ڼ񔊞���!��ʵ_.�B�	q8�Lن�Mz�qh3/í3�ZB�Ilq��2vKZ��}Ce�M�5pjC�I�l�����7]�ִ� ��RC�	 W��]ӴoZ+l[Xie�L)�XC��$(,�)݃3��I@���B䉬�,L��lA	 ��B�&|��B�)� ��A���*9Sp�O;S�����"O@l��d�\%��#i�޹� "O�P�W������
4c�.qU�ɀ"OU����.�fݙrܘ5�dd3�"O&x["��\��53��G��r@��"O�]�g�2����Pc�m�и�"O�}������ւՎ/wԱs2"O�y�i�\8��b��!p�|P""O�1J�퐯]���_�^j�HQ"OVLR����p�b�,�8!gɺ�"O�E�b`6J/����7yR�m�"O�X�����ou�$�T�U�^�TPB"O2!��4T��+/ԣR����"O1�r��=�r���J�\ �"Oe��Ǝ0/oJ|#�M�OI�!�"O(�yNG1�R�����k3��Kf"O����}�T#���)d"O])2���'�"	��@�3zȼjt"O4�  �,8�]��US�1��"Ov	�r�XJm�dC�B��SC"Ope+窞G�lT�A� !(��s"O.E���1T��>����"Oa	 �E
!%��N`���"O6��������A$�t��C0"On�q%!�� �2��t�:E���"O �Ⴋ�����Z�Q8���f"O�	���V�B^"�5�D�5�g"Oh��i�%#j`ڷ��/b���e"O�Q�g	�9I���y�-E%d���P2"O��6��~�i�LKX,��"O�Q F�be�K�lA�kP�2C"Ofxc88�8�ptȵt����"O�T�^?���#v��m"&"O��!��"肝I��Du�z�!�"O(����5:"*�@� �$|�P��"O4q���,~J�c�T/���5"O>�x�L�	4Ru3E,�84����"Oz����6!���#)�-oD�6"O\ɺ�*�'g�fP��*ՙ64����"OT�8�&�$A�@��v`�Q��p�"OpD;��T:h%2�����Y�.y�c"OL��ЋW�!ɐu�,�-J�:E�>I�)f�����S ,t��*7�z��'�ў�|:lO%HH� �$F.`e�!�S�<�ƨ�>(L� �L��=��麡bO�<��%ـ޾�˲H6a�]�WBEG�<YR�@9K�Π���K=6+B��tFCB�<�����td[Gأ�P�:���~�<��/�)~|���K�cB��h�fNR�<�a˫/<��1�͝�~-����d�'�?%s�L�
+$H����
ǴEb��1D���C,�410�e���&���/!�'�ўb?阄��>M����l�� ���y�/D�kd�?H\�p7Ě�-�����+D��*�h�>0��j���+���h��=D�Lppo��sM��Q"
��I�tE�r�'D��׊R�G�� �P��9S2 qRE$D�P��m� ��ıa�åCr��#�g!D�PK���2u<8k���p�`83�
?}R�'-�2��$R� �.1jԩ�'D�(ÆĭC�R\X�	��+�'G�՘W*Ʈp��ZÀ> _�E��'��H�ԟRCX�LY8����'�9�T'D�X� �b�ǒ�O�؀��� ��)$ʖT� ��.�*T<�"O��.�ҥ2"MG�fD��Y"O^�ҥ�,'|��nYp�P�P�"OI�a�D BER�#�F���n�;�"O,��%h�	҅4�F�U�6��s"O�@`'�?tLtz&�/Β	S��mx���Eo،w�1��k�"I�f�	�,"D��ЌޝI.p�Ň"����2D�<�#�	~���y��ulEh )&D��x��@�H�� f�,"�8!9�k$D�숲FF�R��S�o�#u��y �$D���2���U��㒽a�d�o=D�x;�o��)���k��<(����!�<D�̣�	�m� (#AI���6-D�x�@&�?����FG�Sp>�JU+,D��9�7��"��g�$�*�*D�`�3��(����&!�BݙAn;D�8��L��dɗ��$t+2J�$;D��� �zΆ�C�2�"]���;D�Xq�'	&8oH�pK�4h�u 6D����N�a<b)�ע��-�iC�2D�H;3I�s1��i�d�x��c1D���b��1:e��"Cʱ=�R� �/D��QUE�;�Hi��a��J�P`�ǀ"D���,�8�Tq�e�
N�(��%�4D���#���简(&��!��I�G�2D��SG�	_%
+# �8��%Ҳ$D��)�a��W�z���!Z�pR��1�C D��I�T�`��Fأy`F�%(=D���iU$E���JW�Y��8�+?D�(�C�:9g�Y��߸;R޵Ju�=D��+vƑ�l�	%^�A�d��'D��+T�W����ka#Z�`|�d �(/D��r�JZ�0R�y�#�@�P�R�*D��в�N�ꐫ���}ub�)qJ>�O��]���� ��=-�-� �҉/�L\�ȓ@��� f��4j.y:���H!,���s�<%����(rZ�R�L��	�X�ȓ0Ҥ$��L�4P���ᷦ��Egb�n�I������aH%P�2@�	W�;��|�7��y2CA.Z��\C�+F,���A͍�y2D	:y(Q���(6t�	s��0�y2%�6]�����k� �290+O��y]�ۢy��8!l��'�)���+�S�Ouz�Za˚�V铡DA�|�@�'o����n�L$a�k8�tHh
�'Vp)S���!�Zpҗ��) T��	�'/�;�/S�-y�eGT�w6��I	�'8�y�r'R����d!QuA�|	�'t�)x�c��t�0()�':.m��L�Y;v��D">��H��'�V��%��>z��1Kv���7���'8�H��[~���R��4�$� �'lX�T@A�n�d9)Ӄ߯*�:��O�=E�D��j�t�(p�'�\I "C�2����J�?G�ݣ�AG,n=��Kp(��lxa}�>����"v�"�H��p�8Tp���T�<� k[>x�t"�A�,G����v�N�<%F� ��c���;��Ei���J�<q5+�v�<s�����F�(�HF�<ёOҊ%u.<,[��:|��cZB�<!�"��KzR�!r�oh� LX�<� �S�J*%��()`����Q�<qEkӺV��)�
U�5Sd��C�<� ���1@( }j�K��N�.��]:7"O����
�W��`���K����"O|Qh2m�N^ �+^�`����c"O��AD�rl�<�Չ��/6�Aȇ"O��F�A(�V��Gf,N���"O�@�"#��$P���$GQ1D��`G"O(���8W2��#��/�P�9D�lB�H>%;j�)猔G4�	
�`8�	Q��ħ䮭R3������@��G�n��A�x�r�c��ii�葮 �.��ȓ^+n���%A*Ŕ|�C��'Q����{.����N�6(���W#}7z��>v`Պ��hh�-��'�!g�	�']ў"}"&M��+XT��&#�
OCTQc"�U�<	c	G�q�L�x���P�*����P]�<I��>.��]#�!DX@��!��Up�<I�o�� �ď�Mq��w�Ki�<1A�M�J���'HD*{���Q@��i؟\��V4<�u!p!�%�#�K���0����(�`�$6�8R��3��ȓ+�ŀ:��(R�E �(Mx"'"O�` ��=?��FQ!]? �Y�"O&!#�U�>PDP�B�
a1���"O"ݩ��Y� ����/<�bt�c"O<�Bk�rxp�`��(-��D�"O�Ȓ'�O�*�N���A_=̶�p"O�X�3 �~\���m����"O.\s�o�'m�ޘz7��3eU�du"O�}3`��W��y5/F�!U����"O"i��2��3v�LN]���Ɯg�<q#I��5���p�(f�cA�6�bB�I�n}^�A�O� ���C�/�C�ɽA�� `�Ԁ.]��bEfZ�-U*B�I�t�X��#�-�����V�B�I�!X(�6��j��"J�D!B�I2t�D�+�HLLx��K�=��C䉠`*�Ti@�"}�L�����r�C��<����E�-.�L�9��B�pC�I��^\�@�
L�.��unD�_:�B䉉C�p���*G 3&q�.�>2�hB�	�>�T-���E5 �ލ�m�e5VB�	?{�0�/��wr�jǆ�j�B�5afnؚ���f�P[r����w"O
�uoݹ/à�s$�<=J��d"O�����"j����9@�|t�"O���b��Ip�ز����P Ѓ"Or ���<�hta�4Hڀ�"OD����<�Uk� ��$	�"O|1I���4*\�+'L �xx+�"Oz�:5�á7���Fk>w,4�5"OvE�EK�0/�5P�뒽96�3�"O���"@G?#�1;q���Y#\!"OXm���K�(��+�
X���"O�1�օ#�0X��
�)y�G"O�dp�$@,�XRbG��	� �#�"Olc�E1o��p  �r��"O��S��Nwje��6;ȖT�"OY��RbI�HY��Q�FO��"O�p9��c�� t $8�x�*�"Oؼ��%��A��A�`B�I�*\@"OF�֬W�ã�Д]�HZu"O$�z1�Ĩs��!���7�H7"O`��@��HFlI�Ł� �Μ��"O<�6�Y&F�͹4Ѧvؐ���"O� <X�B��~����Πu�� �"O��k`^	nQ����q�8+�"O\a�㙪PI}ːO[���"OXd`�(��T�DoX�`��)"�"OB���+S��`B�F ��="O֌(���g��lBo=M�2�"OꭢЂ8֙���ћ}�T��2"Oލy�P�<�� �-�zH�d"OPi��
�L�h�3/sd��"O@��c"�09%)�T7WT<�G"O8S���,{H��c܅��1��"O\@�Ό�$ ����C��z-0"O��z��	�w�@Uy��u�T��"O�]��f�Hh��Ж�_.g�Jq�3"O��pS�O�@���I�����"Oص
�Q�"�����g��58B"OV�ʣ�¯t�`�"0'�$F��P"O�8 c�8R;6A��%
M�h�"OJAt%��� �4P5��j"O
|q`��72I�К�ā��n��5"O����/Ѫ��$�#�v��"O^��@�ڮQC�,�l�#\��ᣥ"O�m��*sJ�RQ�]4Ppސ"�"O`�:�D#����X4�V��"O����N�qnɾM �$P�~�<���Q4~
�S�-ܵ6�T\�dd�{�<1�g��$@�A���	Yѡ�iw�<�R�]��� W����S�s�<�7�J��9�B$J#T&4��GKz�<���ݺ&ӆdhc�^^��iq�{�<)p�ݩ�ι��L�!��I!�ZA�<Y3C��2T2�MJ�JaFs�o@�<��$�:
���hJ�ZH!���J`�<�"�X0*�����\���2dC\�<���Œ^�T�!�*=Ց��Y�<���δ?4z,�A�dA�k�f�M�<)coa#�*�/�r��1	&t�<I�`P"v<����fI�q�M�t� K�<a��L?w.P e�Ž�DYQ`��a�<�'�I� �t�3!뗼��ers�X�<)�&[gNQ���5	�:�y��W�<��@Ցx��%)�~�aV��y�<!���'P�� �'+�!I���A�<A��ґ�т��?x�5K�#��<	�X�t��p�cmwV�Ca�y�<�u.Q*f&�H���ŔDNa�&�x�<�Nʲf��l�	�H<��k�|�<����f�Ԅ %�B�s<Li8�fS�<�� ��L[�h!�h�Ft:��Nj�<Y�A��`����R�t�$�D$N�<�ׂ �TK\ٻ���D J���G�<���+�f=�FO�L��;dH�F�<)t��=m�FȺf�W�V���,\�<)Q&F�UΝQ�dуmY�����S�<�J.b/�� 2g̷�x|��)O�<y����~��Wl.1����IO�<Ig�X8����Վ�,T��GO�<I�H�c���ZMǪC��cE��U�<1B����ձf���hQ��8�A��($b%Q6�pP�PJ\����m~ {g(���^P�⟏\��=�ȓ ����M*u��+��Mn�u�ȓdW��r��3F8��K<ǔ%��
T$]J0X�V�T5�3�U�%ޤĄ�S�? ��3�./N*,R�`�~&��{b"O�}@�]�����̈́�pE<� A"Oh;� �x��ӑfQ&O=r�q�"O`I1aj,��e��o٭D-F0y�"O���anK0<8��/^�|� �"O�dtˁD<�v�D�x4�` "O"Q:Ҫ9k?�x[���	`���0"O|	q�F��Q2t��4)�8��t"ON�K�Kێ}c��rG��\��cD"O~0�FlU�n�~$`Wd� �r� �"O�AY�)�&����$��|���z7"O~i��/B� �F̲F�M�J+����"O��
�N�|D���@q��"O2�����l�p�M=O��xr"O��!�!2X�y:㧃%a?0ي "O� ���@�ّ�͒� $^[�*O�(����|W�:VC����'9pE@��$8�5
vK�6
���p�'
}���_�F��Z�A�7�����'�l�C�.ߐ~F���� �
D��P��''hh��lU�Ůr��\�&8(L��'٪��C�T
G��A��M3`B	�	�'�.ɒ0c՜4�L���6
� �	�'�&�PB�G�V*�AӶ)ͯZ�� �'h�@�R獥u�KR�mR��c˃p�<��%��B�9�0��p�.���m�<�b�v�ܱc��(�v�W�h�<��ā.m��M�����&�d �a�Ao�<Aւ�!*�\xD��X��e�q�Q�<i�c�0+�Aң�,~�~��ej�G�<�C� >�� Į�1K��9���@�<�aCеipƀ�4]�X�+�H��<Q��,(���R�<Eti���x�<�eP�]Y�,[H�m:�]{Bx�<Y�eY�t��ūR��8��D����K�<i� Pm���S�Ӵ	����.�H�<�(�@߾�@�ۯe���Ҡ��A�<���K�f6���ɥ3��H�C�{�<y�T�g6���!i[$|�\�@3��v�<q�@�q:xE1`
��z��A���n�<�r�J4DM��P��^!֬!�j�h�<iV��xib�+���2@H<�&M~�<�u�8k�y 4�C�K�����b�<y�&<���ˈ[�&A���z�<D��9\�F$Z&�']��Aw�<Q��<RF���kȘV�'�Fq�<ё�U�lLACA��x��ðEn�<	ԏ��4�|A���Ȳ=�dT�l�<)h�8��dj��ˢ`W2�u�UP�<���{8�6Q)U��"JM�<��oǰq���j���"u0�4�kU�<�C#	a$��D�D~��p�X�<�uϖ10�$���,���ЂgDQ�<�u��okl1;�&�8H4����O�<�T�ɂ�R}��FDR��Dz@PJ�<�q�ݠW)��ăLO�^��`$�H�<Y�JL�&�\Ȓ����`�≑"j	|�<1�-�:,VLt�����eٓ#�}�<y�(���+���o����Hy�<9�!��L�$[�eÀ��<{ǫu�<)Va	�~ij�s�k%+��I���o�<с�l�(�z*��\2x�R��v�<�#nUzlū��ɇ{�d��!\�<i�C�G�M@B�=L赋��VN�<� d��$�Q�β)Pp�X���(�"O�E��8{S��AWҏz�1�"Op��!f4�H!) V,[��ݛp"O�`�$D�vQ��S Y�e\(��a"O��ڑ�ΛbB�ʤ@U��� "O�xG��&xH� /�F�`-J&"O�\��{(�-�,�(Öx��"O�}��j��F����R(Y:^���2"O�80&ML�A�5�w��Aɖ �"O�X���!LP` ��"O��`wl�� i��;��� L��"O���P�U�v�)�[�75���G"O�Q�4�	�,9�H��
|��"O>X�%�Q�Jـ0���X��"O� ��B���4q2�O�@����r"ON����RҐ��,Ѣ��E:A"OLy�,�<6�Ĵ𧉌�^�SF"OPaj�f�%$q����'P>,����"O=��+X1��Щ'gX�d��"O�z�mǙ^X��AӶ$� T�K�y��0��X�#O�4Y������y��#DtP����)�	�����yr�̴{n�Q�al�~r|C��T��y���+���c
T���2�`��y�/S�Ne�P�m�1S�iq*ߒ�y�̙�*�,i�!�r;&�0�iÎ�y�n�Ll�H���h�j������y�H��1x���H�[y��p�7�y2��U���(��Q�5�ci�y�,֨!]��1f�Bz�Խ��.��y�փi�mN�=p������y�� �6,�p�G��!;g��iP�M��yBNJ�]��G��6�2��'�E+�y�-Z2^��b���.t��W#�yr�I l?��p�dY�v9awB��y�`C 5�h׭2Qy�L�#�8�y�H˗ka<��WER�z����5�ybC2�H(��p(\�2�6�y���" �r���҆n��y W��y�!ُ>$���Pj�i{2��yB�W�]
�	���J������y�D6�}��%Ы4Xz�6�y"�y%�����-�"x��T�y2bG1��D(�ذv��,�p#���yBC[-�1	��Qgn�`G��y���0z�A!�;d�f�p�j[�y"���Y�|���2_�Ͱ����y��/7P�P�㛑U���;R�Ĳ�yJ	 <|<�V$Đ_��!e���yB�ϨlX~��!���Eh\rtjQ?�y��&ޚ՚�DY<�$`to�$�y�䜃m瀍��(C%3Kf$pg��y��\��,�b�(@�\��y13a���y�U�t��q�gG��Tݎ1c���y$P4H@�cEI�MP�zR���y2`��$�$#��=�p��"*��y��E�4��X6.�-O(�r�[��y�'ӸA����.Cy�P���O�y�.W�-qd���ei���y�!O�źA�.Fr�kӤ�"�y���a�萸@̓�L������;�y�V�z�4i�6��*a ��C�y2(Y�*v��3a3E��B����yb	5��L ���,��T���y
� �ı"�"'���q*̷> �w"Oh���2����t�W�J�c6"O�$�5ț�7(L0ԦP��Գ�"O�H;��[�>���Fυa���"O(\�M�:C�>� �Mg��`�D"OBA
C��cτ��!�4Wwl��Q"O�X���I�¤�:��҃x�u�6"O��`�#�ynl�!��=W&� g"Od�:�
��b���&V#g��"O�E��IA81�4��X]U��"OP��JV�Q�l9A�,��N<��"OJIp�-)���!E{�2mYF"O0Ma�a�����ηp�t1E"O<�	TH_�ec��A��'���1*O
Ҁ��C�^��-�rj��)�',y�q�$w��[U�<@�B�	���@���O��<%#�hרjj�C�I/ق�q0
�L -�!�����C�-`6���C�
�;Ѩk$�C�I#5z|hV�C7#L������C�(yx��� qi�M�3��-.�fC�	#<��@�0��9T�^}��M�sj:C�I$:�F��"����	%ewC�ɜ�4�Z��ݍ3NDH�d�#*��B�	 Ve;���#�`��7
�n�C�I��8&邎�8�p�e��xC�	)���;K!`Ya��H!���U$ɉ"i� �eR��3�!��ï;�QO�=����#٬Us!��ʛ�֘�iP�#��U#Rk�/r!�F�$u�AKu�F��<�p�@S!�V�T��� W拣!�D�+	X9p!�Ě�=~���@�ئxH��h�!�Ӏqm 3�չ'2�m�V��:Y!�dD�|�x`ʣ)��q��r�%�0?d!����t��L�`�k�c�8n!��eؔ�����
��1ㆢ(V!���s��
�X|��Xv�C�!�Č�|Pc	�:]�p�V���P�!��U�(H�0*�,NO����D�o�!��;��(��� (@��koT7gg!���Yi��N��5�Z ��9!�d��[C��BׯG JF�Q�=�!�䐳^
ҩ�֌ČI)ĐQ��!�d�0RB�=�c
N�RD��,�!�Đ��(�qA�@:2�MP���\�!��2TP����;|���a�.�:N�!���gx�$֦h�Р"v�ʃM�!�DX�I�� �/(�8���iѱTv!�ZJm���3�܆B��x�ȨH!�$�!!B�	)u�ŇH�1�ǒt�!�dAo��"w�ǆ$b8l��\&iE!���5������OL�����G-!�D�;��d*�Ú�yHxu����!!�D�D�j��5�̔�F�¡��4(!�$ο!txEڗkM�O��=��hٳi}!�D��R�|@"���U�
ln!�$��p�1� �	c�c�N�fl!�$W�-��ш�A�|\�E��U�!�,d"�8rB�YVЈ{��ݪ}h!���0V$��+�8L�L�a�!�D��4"��ão&=���H��L�!��!�)sE��o�ڱ��.M�!��,4��)��	i
�4	D@��!�� �����o��Ҥ��6j���"O�$�.ۆ&p�8F[�.D�p:u"O1 F&W9�<d�ԭ�v�h�C"O���-@���9%�x��|۱"O^dH�
^M��a��U< �@a��"O�����C�@��K�+�0=1g"O���C3ltd@7�¨�$�C�"Oj�q�Jچ)��I$*�4�R�"O�!�fE��{a�p�Aj0��|�S"OPIE!�Z�b��cfJ�m��=Kg"OD�0��ڃ6�n��r�G�"��"O�s5�Kj��0H㥀�C�>+�"O�4�K&mm����b�H��$"O��æMϢv�lԱJW�=�\���"O�-��m�>�f`����3�t��"O~ p	��c"te��D_�}}��'"ON���ގt	�T�Ú	`�h�a"O���G$Y7 �T���p��=:�"O�!Tg�t��iԃ�,��p"OdS M�gL�8+�nԽ0Qܙ��"O���E _�;��H�p�ݬN5����"O^�Y��,g���C��X0aU"O4q���/F@ ����!�`cE"O�Ag�
1	� I��S�6�<�o"O�KrO	^��z��d�İ�"O����=� H 场>Y�(�d"O�ɢ��@���z��H=��z"O�Ԃ��4'vx����*Y��!�"O�('�й ?�h�@�)=���I�"Ox:GCN2n�98�b0>6��"O�T�4k�"Jؽ �C�3���"O�,���ɟ9�L��i��S�����"Ov@2��(d��Tx��S�f�@�"O�`r��Q48j@�����7v�(�U"O��QA/�c�Ԫ%-��c����"O$�(�e`��ҏĮ3��A��y⫏��x��g�%%���lO��y�i��e���Hh����H@��%�y2d���^%���I���
�;�y)�k����3��
anI�1���y��$b1�2�5"0a��ꃞ�y2���������oQ�# O4�y��U8z��!�0�-8�QB���yfQ&M�")���4�@t�'^��yB�Z�4y����C}�����%��B�	�U� �8R��#�:��B�-�lB�i�T!�i�ꈣwh�y�B�I036d�Ӡ�%e�\��-�~B�I4_VԀ�����ihlEP���B�I�<��
�e[k�z�&ȗ�2�DB�I
��Xї�!4<u��N�)��B�	�gƚh�EƔY�^$!1e��v��C�	 _��@����	a�l�$`�=T�C�ɧK�^mkR�>!ߚ|�Ձ l�C�w�<u#���^%�-����
%��B�	M7�uA�@�5>�!��"�=}a�C�	�"ܨt��_<���Bi ~�C�I�<��3"�Z=�˃hޕ=U�C�ɩ%�n��7�>���c4���a�dC��7c���5D�|�b�h7A�d#�C�I�&�YW	��{P���KUv�B�ɸ
N*	s�C�8 L�rA*�B��<iOp����d� M!# 	V�TB�F� E�����6��>$B�)�  }�6Ä�:�><qB��0���Ѧ"OD��m�����D?����"O�h�ϐ�<��Wk\$�2�M�<�U^4s,�d�KW�\�������c�<�wJYV@����#.MD�Ia��y�<��� �H4b3�֪7�v�C� �L�<��+^!^�R���	�#����T�<�A�V)e�zSs*�<L�9(х�J�<!4�G�+��hc$	ݜc�h�d�p�<Y2��06`��K��E~N��dNh�<i�fM!t�X���ۏ:��h��C�f�<�e�S�2�rBBA oriʂ�	n�<&����"�F��f�H�C��l�<�&�O(���*�!jȨ���Mh�<���#i 8���oۻ)n�ѢUj�`�<i6ꙶY���5ouT�D�\�<�c�:lx�
K�2?W��
�d�Z�<��(�"w�z��瑥*�@A�ƄA�<���[;	���h���vL�*�C~�<����
�8��!\����w�<!@�,l!�B&?��A�r��v�<����McF
r��9�Q9��p�<1@ �ل��EmF�4�i�l�T�<)�H�&K��,ڤMGE�h�;���M�<�5'��3��|�Cg�	1�@�K�<�f`�-]�����R:$A&H�<�!�Gz�x���	�\��ᅋK�<a��[.:R�$�z3H,��ÛD�<Q �P�S� ��$�2���Jc�\H�<	C�<9�	�E%/WU$dzR��l�<�FcN,e���Q��(~�NE�bGB�<��$	, ���W���Z])�-�Y�<�G��.n�ܩ3w
�Qb��(�#�V�<��L�l���p	4~�:)`��x�<!teO�h� ��EQ��P�UB�I�<����`�ph��K�$n-��K^�<�n0[�p<���;`Θ�+�	`�<�A��y0�1�Ǹb�,$jd&X]�<�B��C���c���
�a[�%Kr�<Q���Q�ʳj�-3E�� _m�<�v�ljs
��b�bt�]�<Y��id�]����*xv=)���q�<�2�Ʃ9��a{�΋<������m�<��O
��"��4��Rg�e�<���-�2E�0k׶6�k�a�d�<�&�@3�x����2Ef"���K�<���Ō9��iy
^�V�:����Yq�<��jXH(��Z�%L�m�T�"P�Mk�<1DG�R��;сٕu���	�@�<官�_�jA�T"	%g0ؠ��W�<� ݏ1��A���L\
����V�<���Ʋ{��3L�4��e*�S�<�#�� �b�`����2vaj�@\N�<�E7b�Ȉ��5 0��@`�r�<qƁC7 �Z-��f�dU����_n�<��Q�r�E�t���s|�0Q�Ln�<�hX����їi��h���j�<�B��$V����BL	d�COA�<����Lt�b��A�D�CG'�|�<�`ϙn��8s�ХL��,W��{�<�2��j��xP �H�ı	ѣIB�<��M�@��;�-�J�ЙasIVS�<)'�Πf�����HC¡Bg�K�<���L�"��	�*)  �G�<� <��R�ر9�N�c�"�, �2��"OP``�ΜU
Ts�@�
%(V"O��ݛ�Ѐ3�.Zk�԰�"O�԰Ԧ �w(ԍbd��`�8]@�"Of!რ�.6ؘ���ڪ3��5�!"O<�)��{n�8E.��B�(���"O��Q��\�I�5�I&\R��"O^���1_�H�*�#�/JF �"O��y6��a��ϘNB(u��"Of���ə�}z�퐅w.$݁�"O~�$-ޠ"�a�o�����C"OD��hԬeE�����1�X`"�"OT��m�6��e	�i� *�:F"O`u2nQ�g�X{#˱}�,�@�"O�=�0�V�E�D�X���kS"Ot�(W�U��LUJ^xϲ9c�"O��"`�=<5��6)$ �*0"OBy��G��f\*|���I���"O�塵LY:z_����0����""OA�ሔ&&�Ф�AȊs����"O�� �I���T��,Я
�:��"O�H�q+7����P"�/!>6�Z�"O�<鴀�"_�.���@�K  ��"O`�)�̙%b��� դ^�nE �"O��[ #�=		��xǯ֠�bF"OV�x�B��Rؤ�'		z�>���"O�I���Y�VqĦ
8˂5��"O��j�fA <���/ӏZ���"O̩�6o	��ހ�b@
AT.3�"O l+j��<�th���= ���"ON0e�^!{j��[T�¢����"O���4,]�Pq�ЈDe	�I�P�s"O��k�BR�'�eJ�#	8�D8�@"OP�� fD��رqCm�0S�5�v"Obe�  �*d؉���,X�(؉Q"O~5�"G�'~�H�sʆ7��LI�"O��зa�>7�=m�����"ODA��o�9g42�q����\y����"OhMi#&F�m���Q�o^3,l�f"O�0 ��):1��Uo͝�<�Js"Ov��`��#p�|��;@���a"O�(&���f}0���hX4�"OH�ť��b�D�:F�N���j"O^�����dy�Ku��/�d�;3"O�]�W�E�[��E�eO�P���$"O>�����#u��¤ ��a`�"OR٠��V�)�������,a�"O.5s6ݩR��|��ɏN�^l�"O^P�D�8\,t�A`�.aЕ"O��K�jZ�K����4��:^�xD�""O�U	c�o%�i	'�8ό�qt"O��.g�D{��Νs�� ��"Ov����C&1S����ˉ!5����"O�E+� �,�l��̍5�ȵqR"O�-bтӁ[�L��#�׷x�2m��"Oހ�5�V>B~�)������\}�c"O �k�,i�*��!Jg���ȓ|�B�k'l�*�2U("+�+'XɄȓpB:@��!�@q�B0Q>FI��&i�,��lW.a#` a2D�H�ȓ��I�lG�~�L�R��9~6D��"k6��P"pH��6�م#3.l�ȓA�� (G��' IB��5@��C�Ѕ��$�r�.Y�c�н��E�9h�؅�S�? ��Y��4,nA�l	�0B�q"O*@թS�,�VPz�K��t�j"O���F�Y:��h��R�	�`�"O`�Y!X�< ��c�=
���2"O�ip�+Ҷ~ͼ(+1̆fzI�"OT8b�d�j�,�t��6+ˆ��w"O�Y�W��_N���f��r�8Q��"O�ڒ)�36 ���[	^�T���"O�qSg�-J x�1SF�G��1(V"O��ÐeU��d�
^���0�"O^U�TJ��Z�[�b�1�� "O����ί6hh�u�X�����"O
m��i���] ��!��9
�"Oh���;ږM(B�P~�t"O�`���6Ӯ��f�Q�ŀ@"O@(����R��E"1e�Z�*���"ON�H7��'J�;	�����B"O��S!��
;�Z���V"OB �A~5�27�Tr�f�:%"O:d���#:�"�B���v&���"O\3͖�"N��rk�Q�d�+f"O�q2s�B�� ��2J[i�Fa��"O���S��V�x��_�Xj���"Of���l5O�h��AX�&"Or�eJ�9�^3t'�b�E��"O�l�ӀK�[�P X��	 Z \	"O��0��P������%]���8�"O8�ы��Wu���qnU&%�j`�_�<)��I�fe�0} .��F�`�<	�&E�=��+ܥ^*���+�[�<���K��
���&�� B��Y��@[�<�(��#��G�&q��L�<�1ڂGd<iq1�Y8*�>���FH�<a%ǒd5�C��L�?Z2������<�Ήi���c �A	�Q���p�<�ň�/]Q���q�p�	���`�<ic�V�G��(åA]�Z����^�<�G$D�G�,3�lX�k��dˡ��W�<�CBB�YS�)(U	 4D�hq��S�<�ͺM�nA�N݈&hNa��@Ji�<��D3�J=ѱb��L���4eMe�<Ir*�*�b �Y׮HL�<��̓?3���s�̀?9��8
'KT^�<��Ϝ�-�}�"e�<S�1z�AY�<bH%dD� Xf���l���S_�<!�}����oF,d�d�!bF�<q4�ئX=�	q����q��C�<Qe�ϱA��q�#�=&��])�+Vy�<A#��,�X�T#�� ��x0#I�P�<A�f�D ��EI!uк���r�<�e�3����1$ӣ��Dm�<5/\x�z���#�� Q)S�<�3�O4{�L�`��.�ꄳ�@�J�<Y��1d!.�Oi�\���D�<y��7P@�ç�Ř8�놭O\�<�`AӢw��y�T�fz���b[�<�#OJ'Y�(I�1��	��Ŋv�Hk�<)J1
sz]J$�ا(���s��
b�<���_6D�r�ς�Ba,�� B`�<�g`��+,�H4�F-� (w'u�<)5k�<H~��A1k&�3fm�s�<!K��[���'��kDUo�<��l�:�D�ʁ�8<�
A�G�Ps�<Ag��7Ǽ��lD�qk���X�<� 8lho�% �JPKW�{�^4�T"O���!Dh���(��O�]�Τa"O�l#G��>,m��Q	 �fZ�"O�����Y�=~F)�f�L�j��y"O��a�Z?wl �,@?�聲'"OnM�WMiQ�(J�k['q�|$p�"OH!���0/�|�
1��Ѱ�9#"O�`�M��Sx9��6�R�"O�1�$ܬ&+�A�b�E�0�!�"O0$jv"����u�׎Ha2E!E"O����A�9�a�T�a6�k�"O]*���@��Hk�HE�E��&"O0�KQ-G�)������C��"Ob�
d!��S2�y�%	�i��1p�"ORy��� -��*C�%?~�ٙD"OhQ�f[2F�F��W@�\@�B�"O�i�Q��,i_d�Aš�.@����"O��H !;#tpÂ i�<l06"O��Ss䆝
"QHŏO �H�J!"Or�k�	$�l ��[�,�̽Є"O���a#�6��I`$-R�\����"O� (W![�=Ϟ����d
��Ӥ"O��2n�
x]�h���Q��P`"O�y�%V1z��P��w.�PҰ"O�x�Е~8fM�Ѧ�t-"���"O����m�s�f��$C��`��"O�A��(�/B^()!m�$.�V!C�"O�A��G��zI��G�p� �:R"O�\Rw��x@6�2F-˻f~`d�""O�5��o��Q�Љk�� eܙX�"Oꅣ�@=�l�uf��N����"O�I!`�"]tzl��D[�iX(|Y�"OF��C�U�j��4���Z��"O��#"$߬M20�#r#ՉJw�ȁ�"O��ѧ�Q�uj�l����&q�w"O�|bpo�;��IPS7#VjD�""Ol��B�@��/�	CK¤p"O����Γ̦�2��3��}b�"O�h����b����F�V�ƈm�"O���Dʠ4�B`:�>�U�"O4���a�;}�
e���әO�I��"O>��$�C~�� p�6T��+�"O($r�C�"N*��5!�?���U"Ob�C�ܚ*�� �rO۽W'��D"OzQ�ƅg��� ҍv���G"O��gc�$@0������k'"Ob@��;V&���܉B_zi	�"O|�ygD�[�f����Ӏ��	�E�<�gI�+O\�4e��$o�ʹ�@cX�<�	2U��Ƀ��Jopڵ��h�<Q�ȟ�D"���F�]�)�d�V�y�<����j�|����
~:̉5n�y�<�'ȇ=ȒM{�҄fTYiV��o�<��+�+0��xV��g�xkTcl�<q��Q�?Ω��
��j���z��@i�<ɕ�!}��`rB�{4WS`B�		�~��G��5�5S��C3�vC����M#Z�o/N@��l�?<>HC䉨_�؝kL��T��p���Fj6C�	&Șv�X�}�<E;�@3-4C��0.
(Eö�nH��#�
5+C�I�6\�z�+�g�.�Q�ۗj�B�		?%�l3��
a=c�S�t��C�ɍ��D���7Qb�<C�n�e�(B�)� �d��≊��"u�F �`%+5"O�Ī�nC�hÐ�1W�Y�7�TL)@"O|\�r��I�HH��A\����A"O��3
�
��萆a�%���B"ON�S,9���AC"�ുB"O��yfχY�"�@��ۯF��٫�"Oh���g�PX�@�[�a�"O1�À�%�� �!�4���AC"O���c�-hl2� V�ϖ"��)�"O}0n���r�mҏR��p�"O�l�oW(v:�wF�R�(�"O�{Rᐟ��|�b+ǖhݠK "OґI�.�b:�p��f��Tɠ"O ��6J�?.��i&㔯bP4l(�"Opx��(��Q!�!J���˱"O��q�b�$��wA�-m�u�"O�v�D�F5|�;!�]�p��"O�sB�A�E"����˙>�d��f"O�����s�P���%C
�-�5"Oĕ�@�X@^�u`"%��k���6"Omhd'[�S|}"uCP#SWX��6"O<�:#�P&/�T)&ޛ`�X�"O
�+f�� �4l�����5����&"OH�#⟦�`V��(v�b��"ON���J� �X����W���I�"O�Ah� �)_����I�%f��R"O�`:b��%x �2rK^H�T��"O}�d�ÚKHR,I`ꈡMOj0��"Op���c�=J-��V�' DHt�"O
��,W��B�?<E��"O�D��lTZ��� 3'���C�"O���1R�h��D�]�Q���t"O�M������9���.\�b�P""O�#qET�-�ʤ��C
&l7h��"OHᣥ�M�\�P��DL���"O"�q� 2�*�y���}��u��"O:��r�U2�Q��@8�p+�"O& �@�� H�i�.�*	��X��"O�"��+D�x��W�\���e"OZuҔdr��Ty��-X��� 1"O�H����\<�Ȳ��f�Ι��"OHe���_�r��Ɣ�֊��"O��)�NP�3���ץ�-d����B"Oƽ��*L�\R�@Y0���yH� t"OV"SO�!)p����h4�a	"O���M�E>% ���u4�S�"O�l*��M�J�V`xԯ_�v/�왤"O��Iq�;+:Z��"�H2Y:D��"O�4kR���"l(y�L��I�]1C"O��1�DޕX&���Ǌ=:���""Od�S�� J��ԀVրZ� hZ�"O-��J �b|sͿ4�V��"OV�!���:����V♸r����A"O��o� ��1�'\4J�H�"O��"��K��43&�J�{��0{�"OX�F����]�1��T�Ő�"Obx;�Z�.�`0�hԸ^kB�9"OD����i� agۻ~W&pk�"Oޠ8�F���SA7-wU��"OmA� ]
�ӱ&�h@��"OF� 2ǔ�$��������ak���4"O�eZD���.���i���:biJT"O,H ���BT5� c��P�A�"O\��coBK�d�W�]�=ϐx�"O� ���a�1BnMU�"�pb�"O�JG/A�M��\@ԏ��p	7"O��cIՀp��1�� ��M�Hъ"O�	�N�0��$¤�ڿ����U"O�l� ���W%�(��C	7�\p�"Ote邫Ĺ� U�)��hc"O���D��

d��0nJ�#�T$"O���&�?�xe��_Ӧ��"O��Rr�Ԩ���?��5;�"O�y��+�"�\�
̼0�^�a�"O" 2bH��(\x��h�h$�m�f"Oz ��I���[e"��,�iE"O��A%��2�:���*ܱ� �G"OF<!��>dlA��[�	��!rW"O�LKJէZ�*�Ƙ�jа���"O��1a)�6h�Ƞх�l��0�"O��1�kՌX6|y�Z�d���R�"ON-�ÁC�-�v#�+%�$$yu"O֙� �P�D:��$�׉Qs<DS"O؉���	@h�)G�B'uk X�"O�(�C�\���DM�`cp��"O\��2�?���K'*�dS�p�1"O��lĈ�,�XԨ<B,D	E"OR��R��(�r����S�2@�P�"O5)�dN�w)��$�E�y,��q�"OT9+��)J�.��QW�7�&Ը"OL	��ʪ4���J2Ŕ0��E��"O�HP�K�d+XJg)<n "�"OzT�1��/	���B�EZ�`�"Oέ�pǽJY�eP���A&��s�"O�;'����i�L>��"O������0�%.ZD�EcE"O��0�̀>��R2�,3ݮ�0�"O��w�?ED"�b��S8� ���"O8h���V�(ڮ��1KVU��l@�"O�{1��l�v�uOՁ!uDE1"OrLk��	4. �����mZґ"�"O�Y)���Ќ�j1c̗D6�"O@�ZV�ϠZ3�����q�L�t"O0��cS�x�nmK�B_�uY*t�0"O��{�@�\^zMh�Jx��XW"O�� ��>��ɪvj�%<����"O�0d T�M4D��G �;���&"O�X��P���\"G"O4��"Ǽ6��uc&I#r�ܑ�W"O���� G�h�!����6�Yw"O��``U<A��%�tn��whѡ"Ox���\0��JȒ,5eց�"O�=�񦊙\�h��̬|M�I�R"O���0��g� �����KM���"O�؛��\�p��W�+x��"Ox��"@30*��i0L��4�6"O�.�&R���i�	�p`�;�"OQ{��@Q\p!2c�Hrx�"O�E����N>pP{G��5G�vk�"O�	jA
5Z���^(L��!�"O$��"�=f(�\H�@eXRW"O����Kp% dCՖh⸑�d"O @�P��1>����;@h��cT"O&�8Q#�
r,k�΀,h0(�"O�<��DR8M ����1F�v���"O&� �eS�I�2�x��3�.���"O��3G��=��]���	�@�:�q"O�L���C�
����&8콩@"O� 4)3�9v��h�TlM�k�t�&"O4]����!R~A�ᅀ��4b�"O|\b��cb汁r��x\M�"O�0�cގ_���c�5z.5�t"O,�`�ǋ?1Zt� ƒ.g��d�Q"O��{B���,>p�h�с3�2-�V"Od��c�V��G��>�x�KT"O�[�Ϙ�V,v������F�418"Oީ��ə�or��� ��M�
l�B"O�d+׀J�b�F�;0�C�V��X3 "O���q��v�`ar�-Z�Q����"O��lY����%�O=#�V}ˢ"O u@W`ʿ$-4嚦�ߖS�a"O�D1I�'���/�l8�`"O0�bdZ�LEnhK��
/V��"O��  �&��� &��+鸄3@"O�x:�Խx3�9�ĒѨ��"Oұ�%aޤg.���S�<��U@�"Or
�	��	J�p��)`(��3"OZ�x��-{��Ż��ƃ2,�yb��B7*��P�A�����ꉘ�yc��вi�W��l��\O�C�I #9��%��-@�em�Q��;��!"w#B��� �@��R޶h��gmR��h�W� Z�F�?�����#bh-)å�%%�~�a$ER:H䐆�%�@-���8@�iܚy�4��Mz�PDƯ)�=!v��\]6���w&b���E�}�� C�R85�Z��!����vO9i<$"  ڴI)�X�ȓS,��*�4n�"���)E�V�x���T!g�f�~�p�:<�BQ��+�@��(P0��D�Fd��Ll����V�,=�7g�7L���Y���aG�=D�h;��ֶQZ\laÀX/��	��o;D��`kYN�jM@��=LƝ��7D����-N��d�w#�\o�M�V�9D���"@�+KdA�RF�2U�L�{Q�6D��#�R>P|�����lw@	@��:D�X�P��=��������:�0B8D�Ę�ѧ`�����>��C.5D���`N%wH�q�A�G_�H2/2D��ST��i��Ğ>�����1D���($M� S�원Aq�����)D�䛰�S] Y�`�+@�|��H;D�ڡ!'�d�A��6�dP���.D��@�*_/�����^��.�2l,D��p�BõѴ���&�c���&o(D��� hW�|֮d@�.[8Q?P)೉"D� ��'N�D��N�U�&q��� D����bQ�c��2�D��b��\Y0b2D���3��s�&�x���"3��Dy %D�T�G�X�G�UAc&Ѥo���wN!D���5(M�p� &�(K��2D�г@A����#�|8�0�d-#D�T���;���u�	�)���D%D��PuK��s6n�?"T�0�>D�tؤ�P��Kp_�{�F�Q��8D��A5΋�vRxyC��]X���*)D�X���*a���T�S3�u��)D��G���&KF��H��i/���@&D�����0q����+	�����%D�����46Ai4OL1���CE
6D������n��%���_����!>D�� 8(P��
��T��GS�t����'"O���ꔂ����T��F����"O��+P@M k�.�K�%F�'6:�"O�M�sA�lIpą&u��=z�"O�QӅ��v6���E(,|�2"O�d�s�݁B�8�@�T�6�9�5"O��8�N�T��*�&6'�qR�"O:Ԡ3�4�V!����z"O��!�ό�s��Y#FNB��$���"O@%�F�E�^?�J3+�%v�u`�"O����U-E$h�t��t�""O��aP�T� �ڍ�����"O|H1 �.l�]����)qt|9G"On)�Э�%	Z\9���5c�h�@"Of�`&F�f	�h8�BORl<�b"Oƹ��A�}��EbDA�<4��x'"O��ZR΂0s	�,
�"��q��"O6�!Ak^�V&P�E�4 �]�"O�!�
���H��I�\"U"O���`J�/c]N8!a�B!ǈL "OtxZ�N�{�t{ӫ/����G"O~�x�"��Rq8�0�*��h�JȂ�"Oܜ��(\���꠩�A�2�IR"OB1Pm��S�9{��ҌM���Q�"OVYPP(A�4�#�%E�JւaPw"OpPbgN����ՙs�
w�h�S�"O���wHL8�0��ëL_x�Z�"O�`�r��_�XV��"O��0$ʋU��J� �&/(����"Oe�D�i�"��q ŚYi�}��"OHE�4�Y�h�p]8B�H+X�`�"O����V�a�PE[4O�VTu��"O� ��--�*0��HԺo8�x1�"O(R�h1l��������t"O(��`��R���
{�ร"O&)`1IX .�\`���1ẖ�V"O���H�s��S�Ee8lh�"O
��!$��2��t��.kh��au"O�8zri��*�"�Y2ħp*�)`�"O|U�	��1OG4X���	��yҀF�/បq����Mn�=�$�I4�y¦˿1���8wKȾF�@U���)�y�	� $� � ���A@^)�"��y�V���� 9��i�眚�y��e�J�b�	J�e���@�!K��y��b�&tJ��	ڼ����y�b�/q�J7�� ��	�!߇�y�F߻D�@\`ӂ֬�xAօ���yR#Q1L�Y��T]|` � "Ӯ�y"�O1M����&��)$I���V%��y"��"yϚ���*!�4�:�cԵ�y��P�5*���ÄWHKE I��yr��?KI��c��_��0���:�y�`�h�6�B��FY�Y�sά�y���!�T�P(A�6�̛f� ��yRÍ�c��i8fo�?��Kf���yBl��a)�h��N�"��e��yl�!��|!�.��H�0=xo���y�JP#^4�Ycʒ?�&e� ��!�y����T�: �D�7Y�`{��D'�y��Vm����� )��/���y�)�G<P��%�{����ލ�yb�D|l&�6��)������Һ�y2�OwZrU���ȧt�SK��y
� *�񦏟^�<���-��w���J�[��Y���dHb	S��Y�x�0ZUk+D�da��@�a�@��Ⓡ���@�J�<�5hL�Z��%;�B�?]����BD�<� ��(B@�d�c'��)"���NY�<���H�Q�@��!�F�<�K�LQ�ɕF�a{�"�p���'�1�L북I,�y���I�
��wA/ �H�˳o2���6�O�0W�9��m�$I�/a�]т"O�yxt��sh�`�W2
y%� "O鳥�B}�20z#�Z�S��!��
OF7�M=>�ơK&��UE� � �Tg!�$��?�d��bW�J���uAԘ>�O:�S���ɂv��y�uJ@�4Y�!B�� =vB�	^�)k6!W�6�D���1`&DB�I-/3�5	��Y�d�,,xQ�D.�B��m�V�tLϘ>=b�"�?��\ɏ2�'m�7�L�)1"I Јǂ�(d8���H9�h�zM���g��-*cM* q��Zsh<1c@�j�J��dC�d[�|x�B	IX�(Ey��(f��A�\�XY����
�yRȃ%Y�I�%�I� ����������I���s�O�.���'�m��2�۝U/�		�'��5�D��!���#'�,{,(�ˎ}�3LO�y;Al�-oo�d�j�_����EOZ��A̚�Ψ�{RF܌?x����p�g�ЩӪ�6\�X�%�z���D7,O��<!5ϲ,<Ra� e�&U�G	`�<�o�6}��@�"�̸0"�_�<Ag�֟���� �ɜ^�N���m�`����>��
�'O��u���\EPP���u�<Ѳ.
 ��b������,��d�{y2�)�'b�qӇ��9D���X�oL;#Y���7�R��C�ˊN�a�E��>h*=�'�����<�s �JN8m����E�Wg�e��X��4�?QE
�\\� ��_6hn���u�؅�M[�����8D�4,?D�Eٷ;���	j�'�b=��-��p)�H~���2
�'5��h'�ƃx>Z3^<"�g#�d2�Sܧf/���ф��CK,�JG�Q�V+�l��_�4�Ə :n��rd-�2E�T\�'6��>\Of��-E�vhz2�5x�1"`"O�� ��$LU�$��"V���!R"O2�k�Θ����p��:Z��%�'e�O�UB󩈢N�N���	��Jp�s�U�`G{���Ƽ��ʴ�ևT�j����SkPqOأ=%?U�d�d��I�Ì�|d�	�"F'D��e�	p	a����c*���� $D� a��u�B�Q.��
�44r�a!D�ȸh@�(��q1A�<}E�k�kcӌ�O��IX�g�	�4r�0�j�.�(�qP$g��B�ɞ;�m�� �2-i��SVM�3SvB�	�9Iz��w�]%>K�����H3�|C�ɵI40�۰�S�U�rM�d��A�C�ia�aƮ_4���ʕ�.T�|��:�D?�S�' ���bB�2�|XJ7o��J
x��ȓ����D�c���C��b<��&�X��	�N�����0.� ѣ`Iy�j��1ړV FqY�*��������?M�␆�q��5Ȧ��cJɃ�.�#zi���'�ў"|C��7M�6�Hv�T:'j�1��L�<Y�HƳ7hʨ����>�c�"XR�	(}�{� �f����
R�L�����yB���=<�d�U; ��T�u� �y
� Z����1��AP�bQ�_}f��"O~���2������5���@t"OpH"VBU�$�Nu���V`��J�"O"���Wa<2L�1�(EF��Z�"O�H[HϤX���!���sX@a	4"O42���3o%���ICSXĠ"O�aVg;9G�x���O�m/���"OF(� `�-w��b��3Y��m("O0a��k�!$�ʄ�C��"
Rm�Q"O4�+tF@��jV^[Ҵ�Sϑg?���퓧3�@H���[�}��)s�\<k2(�	^؟��7� 4=ؒ
K;Oa� �V'3D����5R$Z �@`	Mߚ|@M#D����(�~XͻAh�Zgf(� �-D�D�$f�9}��MJªR$`H)6-D�D�'W�i��HƉO��T8�)D�X��/�,�3u�BI���Bq�:D�h��Uf4��+aO�]�|İ��%D���t%F`Zn B��@�Y9Z83O!D�DصΑ�P� ���"o^y8��<D���"��Ff�Ѣ�N�3%�"ukg!/D����ӀPL��A� _���()$����`W-mOT{SC��؍K3�D�yr�ަ�j����ƴ{�X!Xq"J����hOq�d0z�%�@� �JDn�&%j�R�"O�H�P�J$��a�`���M�`�7"O��%&�#L�`lqA�A�/�x���"O�	�p�|ƀ����ˆV�l��T���I�C䊄�pʑ�#(r���/�:B�	#\���F��0'�a9v���_%B�ɢ L`��/L΍�v�Ѳ��=��&�'-���$(���sĠ�_$��ȓR^6� $aR5^�H Q&N#K�L�ȓ��u��M a5��X�

&n_����zH$� e_�,�4\[��Y%xA�م�)�2�02Ά�6a�0c�Ƀ�Fh����4s��!!��"M@F���j�=���8�Sd��;�a��C��(���-_l�Z�ƴN�>Ȅ���W��&cF�[".W�<�����	����p&���G�8� ���b�^X�A���$�1������'����,F	oV�:��A]� L�ȓO�.�F��6�bG���=�,-��J��2�	?)R��@�ʊ$���'�@���)�ӎy�fEA֢H�e�Z�)3-Æ:D�C�
y�����
J�_D@�%A�2����j7<O
yk��\�u�pg
ڋt��e��'w
}�ҤOoxT��` ل�P��$��P�!��^8a�J����ױ+u ���ȩ��y��9��gܰ��G�y���T	(1��C�1o΍�&�u"��Z`���JB�I�G�^�Y�#F�	��
QhIk�6B�ɶ1/��	��_�z��|�tNFfF
B�ɂ��B$�ҐtL�8�vI�#/�B�	�p-��:T��5-�`T)�LT�[�C��
k%�@85h�u!dI�B.�K}�C�I�j�p���e�\�[R!�5��B�	��&�y��-E��E���{�B��#2<9��ݨeL*E��!ʀ[R�B�ə��ѳ�'�5&UF�"�͜#-�FB�<�(-i�cG�yy8�5oX$L�FB�	�lYX)�AN�bJ �Z=s~4B�I43K2xX7��'P#>�QB�>^� B�)� ��B�2lh���7�@q��"OD-�6�̫E�@�It��I��ȅ"Oj��r쟅�� ���U!,@�"O�8�#kıa�< ���D��)�P"Ore 3d���ӣO�%
v5Z'"O��+w�}s�8�,֊�5RV"O�a�$C��� ���i���Qc"O�	j2�X�;������"]�h�1t"O�aЊ�?��9:�L�?$MC"O��E�;EX�� ?`�u
p"O&t�tKR�Bd@,�6 �x�LRv"O�阖cV bF��׏ߤ*�T| �"O:�;$$�K=B�Q��v�عp"O����d��H{�ա&� IGNh��"O.|iA��l���pKX9e@p���"O�����35	��kiɬKǘ	R�"O|(��g��i�t�Iu��Ҙ�K4"Of�� ��B����2A�&k���"Oʝs����Eb�
�����"O�@3��9!}vE�QM�*R��9!"O��������Y$��.F�P�2r"O�@���<
$H㶭[�<�*�x""O0}yD�O�|8��߱k��D��"Od�wFV�!D�ٸb�+�] �"O��G��u��T�R�B�T�b"O�mP��3�0�Af��,&�����"OF(��^�1<X8���$�̹r"Om[��T��t3B珉h����"O2�IWnR4"`^!���&Y�Er"O�s��$T�$��wO@c1(�Kd"O4`�B�-<`yt.Z�\R�3�"O�DPF��O��$y�)�<=1�"O u)��F�O<��K�m�R�y�"Oj� �k�(m�j��H�p3e"O`{7IO�q�r5�5j��p�hc"O�1c�E)�h�`)�;�a;"OV��'F�'j,`	��ތ�ȡ��"O��zE���7=z)H�( ����c"OL �bQ"4�~�HG�?z{X$s"OJ��A:��-y� J�%]v��"O�Ũ��Y1_4ڝ�Tm��t��"O�Pb��C�g��K���V�~x���'�^uz�7��Tj��\��<�Ad#��)�`�3���&&�!��AK�x�̘�JQ\�a�L��0CqO�{� [rBr�@���]�M�1�њ�$B'f�aY�"O��W`T=���9����������+sN���I"+��O�A,>�y�@��jν%�>8���llq�Ɠ(���W���p���6&��P��-ޛ}1B�X0`KV8�0��� =tI:���f�F@��AC�5�O��q#�O<�s-ԛ1�X	{D
T�a���C"O�I����G�6X`JʒG՚�'"O~�)P��+�nĩcIA�^��SR"OE�$%S����
��Ip"O�gC|a�-
3�H3]��i�"O����Μ�;ؼ1(M�C���W"Oԭ��o �5�xMi�*H"mSvlz�"O.�J�H�J�c��է'1 ���"O�Dp�b�0*�L��#�(4���B"O��JF�ҏ~��+�ҩ"�p�"Oz��,�/WFЩ ��T�
u"Ot����V;t!K�.��j��H� "Op@� ��	��m��I*p:�"O&M	!��\�X�z�jL�p<��Ht"O^��ԏN7
dP�.Q�G΀�"O�  �7)Ig��Z�ƀ Ӕ�2R"O�	IE�Y^���Ȧ��!}���i�"OZ}�ՍƇp�Hฒ�I!3�"�{v"O�x�V��8v;<���Q��q�t"O��bd?!8���`Y�%�����"OHH��R�*k��8�z�i�"O+ti��3�H����ĵ	V����"OH����΂F%0L�R,���:Y0"OH0�d������̛*c���"O 4���ǧtg>��nE�NȌ�P3"O�p!�7zTȍ���I2�l��E"O��H	5O ��z#����^}s"O�pz��?EZ�XVf�F���$"O�ز�M�'�F��R�\�_���"O֬Y���A�,Q�'K�f��<�5"Oq�w.�E���pE[+�Z02�"O���ŭ�Zq�k���<��(�"Op	�D�-� ��R�E|�T��"OZ`2 $ţ�y!�#@\��"O�Izu'�n��yU�^�j����"O,,�� RW�C�H]�c����"O� �H��R�y�-�Y8�C�'{j9�!�Ѫ���a��$�����ph�*0��;W�~�"�&'�>�kX<�>`�-U���OV@��d�~N���]-��'36��b��7f B%�Sa�B84�ȓWȪ�i���PH�(5�ѵpK�U����8�ń��RgM�d٥V�Q?��G�^�-̒��6AԄ�`��Q[�<I�jt����+X(T�Dy"*��F��-P�HP^���b�%��x�O�Q�۶
n}�*@��C^Tmh�B"D��AN�;d@�@F�S�6��X@�4?9��Bg�l9'��iR�m�d��5"zbIf�0�Cq�Љ6�8}���!�p���t)"���nĪ"�Ds��F�<��h�	t�ր�4= ��*�ß�Q��j�HZ�S�8�BB�A�O&:)#�S1@زtjG�W�Xyre"O��j�D��!O��IW(/�b�;��O�qbf@J�Hm�$ÞQ}"GH2�O�5��Hǒfаy�S�
�f���j%�'{���٣v�VUs�,�_&
	:�#�/u'z��G#ʦ_�h�U��`?�+�?P�zb��'=���6O du ���ȅ<��'���"�`�.�р�T�z�)�#iTF+�)�ȓ�s�l�p�hD�`k��)�dP	Bے��ȓBҤd��B�R�<�Iq�ւP]Vp!�
��<\y���d=(���CԮt��"�I׼��&��<�B����L��Aa�dMx��������Iq�D��𪱢�"}h@k+@�Mw���O��/�9�'��#���J�(���]�n������nܓ`)X�v
ڒb��W�2� L'���/�"&`��VL�+��$>s������3����c��$�d�A'��'b(F�ₙ7%sr�w�l:��'p��"ӣG��F�҅�	���e�+1;p��;O��  ޟ^x��J#F��T=�B倉���EG*2�D��	�3ʆ-�'Q�y�6���'�T�V�@ a�qDe��['��q��(BP���D^r���BȚ�n�r��  `�e"4��Y$��(BR *v
G9E��}kE�A���0�8��Or�C�oxA�eZ)E��xG�9u�v�S��\�gf�ę'�F���z�-F�֍"�fȜy�Ԑ1T���1�x�yXw���YB���4fqOD�Yf�_;7������D�*ZXe!Q>O��kc�:�\h�唔�R�L������Ĵ(_VE-}(� [�H�qf�%�ML�m��Ԣ��8l�
�i�f�E�Ф�fk�m��0(���a���١�Y%1t�,%� ����\���h�lR��Z ��M�0{��(�e �8	��+D�}��gj�;\�0��$$.�1)j2�a}rn�㢶��9Y�|Y�hͰl�>�����M�J�1)��C���)C��-�TI3�diDH�j�$�ѱ ���YwR���)n01#� �Zl�S���Y�'[|�٦�U�j9Ku��]c�;��mJ���K��-=H={`,8/��S1AK�:��ŲB#U��<�# �^�����u�T2�4�+H>�S/�8,
7 [�g�V0Y��>�T��7� u�1���"pda���|�<�)[�f�^(abǖ�9�L��L��j��`)Xl��B&�ڜ��JW�O
p��R ��<��IM�0@������50P		�y��,j�$A�N�X� �/� �� �w)L�7M���-���= pi	�z�� jRaPg��E(�!B
{tvQ{ ⌲�p=����_��`s�F6���p�����y�3&"Dn��I A۟0�HK����:i@*$Ƙ��!�HL�V�W��IV��oz �@�Q..X�Y7�K�`:�)T�}�1� �%l�L�hM�0�9^P|�x#�"_�湡��"Vf\��N�"d�L;�v*��ĂYnȸ�A�E[ֈ����#U`P�e��H�,&���Ua!q�L�1�+\0�1'E8\�8JwnU���11NJt[b��Ł� s�@�	�˜��,A�e:X�� X���6��Q����}T���egAT]��kɒ����<,O.��@Ky�@�5�o?����M�
 ����遗Z��-˶�
jh�4�@@�z�
P�H}���"@6�24�"���~<p����B:q�r��D�  �x"��	�����M�������FX�1p�BX��]*�3͕!S�i��@Ubuh���'q�T	Ei�y@�x���5v��Aj��T�V�E��5sZ(,B�Qa���
�	���#+��y��f��5ۖ��Cc,�R޷Xf>]�AH��i�t�À܀Er�X�m�/1��7��9�X��GԘ�J3@��x|�D� �Ch�  �)����l��I��mA�j�_��2��k��u��f̻B��1K�%N�!|&�����;hʼ3D�1V��QRSi�HI2��
:N������2���aU�d����[��|�q`�>��2=+ �BUV��seh�A��}�R�;w�2�8�e��Q�d=!���,���+wO�VP��c�O��7�>q��i����K|Ll{�*� 'C�]A@!śo��"?�S�RAbOˁ$�H���':�a!�L�1U
-3Z�R��Ā?m��(3���-��%Ido�cM��F��3f�숱BHC�\�Sd��k���WA�44(H�LB�wc�l3��{y��I�
DȽ	cm��0��yu��	�<��T>����HS�5��(��n ؠs��.dF� �T�^y�6)�� Ï?���:�$˲MX��7HRk6��<�Tj\�:J�L��OΆ|@MZp�éI��y�$���|ȷ��& �"��$;N�P�qoz\MJ0
C(K��q���A�|���eO�##bu{��ѝtQ �ǄP"���Dq���GQ�������Z{h�0�Ԏlbhiu*��*�ۦ��L(6�ؘbj�?bڠ�+N�Լ�aCM�,B"A*$�ڠc;���2!?4.j��2�CƢrc�
-H�+#�ךXF*Q2D��7�4��G�I<*4�l�kN�%вuAc���y��۲K&��P��2�:��w��������:�X��2^��p�	۸Ly�-)'����Gp��� �f�D���V\�e�	� �l� !�-(�a9C��e�T�H��׫�-�b�ڕ4�b% ���d�2`��/.�Ea�N�B~�L�"�^0b7kX�1w��KU�ƹ���`���"u��Cg�;W-x�c)���
6��$�X�Б���o7�\R�������E�%(�ȃ��"�����&P�p�r��?�V`F{��H�/�%��/)X�6���(K#Dn1���3m�\���8���	�M�7�._���8dEС8�, ��ش`)��P�(����FNe�q摓y ў8¤�/	:����G��Q�f�DƠ.s��A�F#d�CeL��F|��7�zD��W�R�"��#)|����G�&b�����CԤ6��:��$y��86�*�D��I<�d[1�!�d�F�t%��੘5�ɲ5��j�)D�*]ĵ���_�^M��@#�.c�X0�*�dA���8��Mr�O|di��k3L�����1�>�C�ǖw(Ȱ�O�y0��)§�Z�!�� T,l<��ĄZx�� �NQ�;$b!Z�Z|�Ug�U�
�b C��S#���*��ӲoÀ���<Yz�p�'��ƹ�l��f,��+�5�H�qK�9H��贆��e�� I��x�Q�`ɎMo��dQ� g�d냅�e h!� 	�siR��7=QnM)�C�$�xP-&j�P�C�֕f(`��ΐz����L��P�p���0����
*D�@��o�$�"�30��Dsd��P�I�k��������`�W�،ʧI� ��W��^n8�V�b黱Ȉ(-�];uVsz����,����q*��z�X�@+�-I�R���R��M��ˁ�	�LŪ�	D�me2��jZ��"?Q��C� \�0���+2]Cd��A�'��x�G%Q��q���/8E{LO�f}4�Y ��"{:�5��#�?kC���q�K+�  ���j8��BH�i�����2�8ܫ���/�*�FLܣ[����<l4��"�R�k��	��y��όOt}�F�>/��p����y�
IJ�S0�L�*u���p+�W_x=��4z	^����:|t����O����`�j\���O�Ġ����E7\m���^a:,���1|Or��e�B ���GKT�C����Z�,�T�S'�\��c��Ѯ./��ےE:tPJM�˓A��-���QY�Г҅��^)"��?��녥5�T�3��!��L�G%�C�)��$��L�v*%�⅑��,}!�D��@�qAFLʴF�byh!�#|�Q1��P�c˺p��Wev� ���
	H�52�4p� ��]tx��7D�|[׋۽��2VÂ�Q��JW�w���[a(��e:2t`���"�~���8���R�	R���;:��{¡�C؉���߻�<��pO+f�z��@�0C����H�;���r���N]p҆�0< �#G�Rל��?�*Z�=.��� �̡FA@P�N��!l�)��H'[�b��ឰv!���3a�<Rec�)�� #\�8����P=P����ϘhH<���8J���U�T�1�C�K��E2D�a��ϖv̘���N�/eL��wK�`I�l	�}�v��"�%RMB����z�^Ģ��BW�)g+��;����9YZ��(�<@)btӵ��.�4aedJ#4���6_�x��$ƭWx�#�/m%��!bO(iQ�����F�Qt �ccT�l'1��9��T\s��,�mCr"O���5��J�d `A?v��%�i��؂�a�$�wP��6�1���Eȿ63�0(����p	 B���>R��Rl��Q3NK�I@5�.p�U�*��m%�İ5� �Y��'̦4���Ց8ٶ�ga�|ӌ�d�O�"~bu	�NAȋF�ڌ�,`�M�\�<� (�K����KOaB���� ��ihў"~n9W���� �22,��T�H*�B�I%����֩~��5J��H*m���d؟�B@E� ���B�NޕdJ���f +�la���IB��ۥ��<��;CF��0K�� ߜX)P�
5 .�ȓS��8� $�5Y�bdm�g h��B��'j"������V��'j�jQaf��H�Id�8�yb���Y�J��W`T�eB�ɀ�
J��y�јX��1Gg��]]�X�r!��y"g���T���ц�<�CB�@��y����1�ޠ{B��2T$���oA��y���f�@ԣ���H�P�C���yR'��nǤ2���O��K0��y�ϗ�C�yI�dZ�=�֜��ެ�y��)[Luӓc>i��X��&�y2�L`	�A$�$�H�匀�yRE�cJ<-(��	�c�1�ՠͣ�y��U�^(G�d�RAz5`���y"H�,c�ika ���A� ,�y��B�(�j��Ԍ�Ր��ÏO0�y"�A����0���= ��͗��yF�g��5�GMЛn�d��¯�y�s��d�5LV�->�d9�C��yr �|�j՛�E ��L����y�*u�&e���1'}���O�y����}z��ޥ-�>�:�%D�yb.�Yr���2-�#0�3�Q�y�-�m����(���9Z�E��y"`Y�/��UiDB�#$��0���yr�͘�e��R�K Ն�y�a��~����⇎�������yb1�������>�:���	�y�Y�F
��3Eڕ��E	����yB�+�v	ad��$��\Z����y"!J0<V��� ��0t�)X��y��(2� � ��]�sn�P)��?�y��%y�=t�_)Y��)ė�yBALx�F�B��[�D��g+J�<1�ᇁ*�� �c׿6��i����B�<��F�%e�Q(T��ҸIF�Jx�<ybb�C���goޱ(b���l
s�<Ѳf_�i�j��w
At~�����[�<IE�P�lCb%�s� R�̡��S�<	#E�
���!�bӉ$�x��Fc�J�<���<s2��Ȕ�F������i�<��˶ ���V' �I|��ïd�<��,��=�]�V�@5=�P�2�X`�<9r�N�bf��C(��w���hp/Ob�<Aqa48�)@ ~_�����Hp�<��䟼@��D���ޫ	�%�Fn�<YB��L�X������#�@����r�<Q��8cL!�b ͚
%�$3��q�<q�G��!��T@E�t�H�v�n�<q�ύ�"B}�ge��~�hX���`�<���A'q��8�0�O�o��X�p"O�Ay��}/�M���B�x�<��P"OZԋ7���Ԯ�8�Ǎ
p"O��ģR<�~�� ܡ-��`p'"O$�@ӊ��p�\��ʐ���ӥ"O��rJֆ;K�e� ΙRcr4��"O���+��m�v��t:o�qQ "O,Yх�)7��*��@�Ct�Q��"O�u 'X�bG��%�?x^0�"Oȩ����[���%X)	`��ң"O� N��*���e��u�8"O�� �Y:` ��2a� ��6"O,�B �\>L�([�Z���x�"O�1�p�ƛM�`]� Db��2�"Oܜ�S��:EuTua䇢F���"Ot�aӢއ.���Ì/V�8<Q�"O`a3�
ۑ\��Y�M�~��}��"Oh����/K���Q�T�?�z��"O�c֮�r��RM x̾}�U"Oֈ�T+ԃGV��GA�'���)u"O��X��$��*��_e>�"O��$F��`E�%���X�%����"O��V��5 b~D8�_���5�"Ol�q4�2,)�aR1�����8�"O QP X8jR�,��.u��rT"OL���ȕ$i�.i�	J5����T"O1٢iHg��i3��s^Q#�"Ox�b����,��%�ɀ:ye��('"O�I*w-
AQ�hv"ִkT�d"Of{�Jt"`D�'㘎D��)�"O�5b�Kܧ_�"Ĩf�ʑ@5��"O��4)J�;h4�f�8I(��b�"O�}[V�2Z�B�����;����"O0����� Y�N�Ж�? �a�"O��˓�f[� ���#%�H5�"O"��Å&�R� 3���K�Ty�"O��)"J�o�d��E��	�r�Ag"OЄ)����,4���� U�X�"O���P���J�բ"Lu[���"O��An�D������ �NY��"O�UqteH(+����T�ޱ-��ۓ"O2ٻ�HFr�ޙ9r@��4�b�r"Ol���M���� ^��R��Q"Ol1xu�@(&옔Y�bD'�UzR"O�8���(zXLi������"O���s�L=�@�)w��I��*"OR�Xu��K���d	��'�N��"Oʱ��,�
L�V4���h��c�"Ov�('�ҴD����5� �"OV��!�,:��Is�E�.�mrc"O����ٲw��1['�-c�%�B"O8�!�lJ8��9&��
L�>a��'�B��R�k(4��,O��H�)�x �"�S2)Ä<�"OFBHN�U��:��.�Z| ��0�E�A$X��� f��ȟ���aNS�;qn�P�
�$?�5B��'pl�p���%=�1J�'*�ܘ5.
�r<��9�g�<C�{�BK[�(͓r}�5�S�ͱ��g�tdnTAlU��F�Q/�DP$�,���\ڙ������O .�C�5Y:��� ��
y<���>2<h�E�����3�O��
!e��^U肧��VGؼ�AiL�T�̀!�u��s5$M����a�]�Lq��Z�SKܼ��������g/�MФ&��7W�$�uO����Kܺ19���І�P��'�hvʱ#��o����%]25q���Ƨ�:1:��fT�	'>�u�����%�
�w��5C�i,�PvT��!!ܝ\;��2�h10���e�w2�[G�I9�p���`e����qC���ɖepRС�|jb�Oܓ2�Ѝ�cD�0�Y_<�$�EIu��)m�	閄���_�B���D�"��S0�dMj%f�8�2��I -͈����.,���k5��>O�0�b̉����ɝ�")�%"J	u�b<�,�������7N�p��B]���Ò�٥~q\l�4LW
/)�q�a	�*�u��E�H�68s�)Ӗ���.
�q�+_ �h�bE�m�b��
�.ب��j0�|�u�ߕ+|>��0-��%(���C�\h�u���Ӌ�4���b����
�<+ʌ�Ȧ�x�� �%v�1����+-ĬY��	��b�����"{���"L!A���F߶%�F|(�#	�%`�䌂9c�Y+����`�������[N*(��M>�a�-���h�^<0Ƥ��蒋��]�~���
�dC����AP
.����S++b�O�B�H�HR�H]�榋����+s��C��hXn��le���+�yx��B�#W�o���r�M�T���U���3nU ��))N��0e!�Y�j�
q��%d���2�͈U���e*�:xA�E*
-w	\)P�?�z��e��D���`�O��ht5ѡ�*��  �'F*8q����%F�f��b���vh��3'(4�t
��,(�nB����ᷠK?�Ń�� G<�a���
;��'I����Nܓ%��qa��1l"Р�a�^1"L�	x(qC�	�R0��hل0��陵��-h�0
D!��EP�	�^�ੲ`��^(��H�6���%��h�F��l�0��W`V�`gZ�PB
l���֬�9y|�b�Ŀ,B�0!��n�<��'��.c`H�{�bf��F�ŬQI��9�!b���f��)5��S�8��P�bX���M9���jWbQĀ�H�A��<�D�cٯq- �	 ���Up`ʃ�L�:���Jg"�ٺƢ��Hp�L&1"�[q���}����S������$�G����O��j�xLJ�&����裍�z��K���g�R5��H��?��X�Ǩ�:a%nPXF�U���	�CmO��k��b�D�1(\(���P$@�?)֬�6ŋ�-�H��O�y��J�Pj�ѥ��|��% vبdI�ŗT���G�cT���BB�c�<u�O�@�x,+f�X�+  �a������ y�j1eY�����d��'��t�mAP�L���ņ�tŀ�#�O��y��xUjE
Qd�KG,�5�d�W���T�V��pEG<p͐�����x���CN@LAP^�a�`�u ��>���ŗ��:���(tP��M&cl����6c��g�,\�PJ&��8tB�x�L^9s~��r�'���|"��i��B勘I��hځ�؀F�Ԝ
Wf�z�����U����:7�&P c�Hr&͠U��U���D��id��3B��_Na#U��
N�ȝ��&? �X����P7W���T靺kb��k�j��YCU���h�Ɓ��l��a�FKy"�ܟso��rW�	"��X�G۹ug��GV>��V┟L��2s%0N�.t!2���D\�D�� 0W�1����'�(%���I��1j�E۲K�8X�<	��~�p�AgŎ�Z���=7�0툧-�#|X���A�*@E4��S��|��G�J�d�5�8嘠�
��5�U1��}���:�P��/�3\�N	#O]g�'�0z�����굈u/��L�x��cN��H�
���N�_�L8�T�iq��a)��R3��s1��
!�p�������	 #]�#W��:�j�;.�X�Xt��8�pm3����P�䐃R.�	CZ -�S�W�!S���B�*h��!«��/���Ed�].X��fH��$�DE���#^M���5Ĩk��9��C(��b"'��r[�	9C���B.ꄀ�nϕ���̅M��bK88\|���C�cA�b?�0gLT;g��6IՍ��e[�D\,'�V�+vn�m�Hݐ�Y5SC��*R�T:e��v�
��Y#�O
�qF@�#H�%3���	�L��Ԃ��c� �Ě�s
聫��U:H$�S�i��!�'��3U�.�pd&�!�hHʲb�	��Á�1Ss�x�+G&)&�1� ���(U���hO����鉘}�(I�Q�.^�ƽ9��܎4���kR5Ҕ��u\[?��d̾\����V�-n�� 8����D��� �F7@���s,��� � 	l�AD �S u����E�-��d���wfD�LPJM�N�.6��ٹ�d�OB��t�6F���3�Z�]C̝ꇆ>I[\eC��O����JN���%.:$����l��N���&�0i�K�1u�J�� 	)����=���ң"x��抆.#�V�SB*��4Rb�ݳj�j�R�ļ#��Sq°����7��I�m�9ڳ�
�S�`���ǅ��j˖�#=j�ɋ7.�D��A�Ϡ�!#k����3DQ�K;z!�H�+[���*�:N��DC�����%�-�
���'[�x`��I+z��F{����P���1	ϵ#���0��
����G4V�ڜ
�N�~�~X�A��
3ItL��I�W�qs�mԽ���`!UI&��d6d�T�ӱ�ͿD���B��Q�E�?���H?E[��۱v�Yi����?e�0��#�t�<�ծV�xS�Qw%��b�X`	4n�Y�dEڇ���rZ�� ����F��=�Ot�E1s�٨W��'��<��FEo�px���(1
�C0lI��� ��bD�1a��9�WƨY<��CBÊ�,M& #Vm�z<r��U#�9'0�<F~2��%D^8uD3�1�Aώ��(O�d�a�!ODk�$�1�%�1/N74�1i�F�2_��J3d�Vh�5�񀃒o�8�e�'��1x�.	/�Q��5�.�K�dꬍ�A�ߦ��t�/����)H��*�]�ϟ�J+C`��W��.��\���p�!�DպCg6X "<|llXs�@�*�X�#T�i�FT�W/�Lo�%�¥���`�`�D�|����Ԗ>�B�N���]�$���+ބ�K�"�v��������!!T@�h��%1��e*�Jǁ��J`�x[��� �Hq��u|Т�'aDT�6,�'0b��D%�J��2�r�_�Ը����Ho�b�IJ;��ӎ_��y��!�T,xRl5s�BC䉎;1�Q���u�H].��!���86��9"�Yr�Vi.~� ���((,�U������2X��6D�|�t�����5�P�ۦ,����RNվ��Ao�j�Q�"+���&��	�0�RT��*�6_����6�b
���ߙj�l���FQ6�Hl�0�B�|F�iG��`��p���5���P��p?��L��p�`,_�{���ٶ�	c��6��-)4Oط4+
1�4�Y<�t���V�E��5}h	��"�_<�b"O����ϕL	 0U�
�P<m�_�@�p�$`�1U��1��@�>��$V� 
G�W�$�ܩX�c�:{��B�&�J�$db\����φ=�z�xE ��~$v�qVƄ-��L�sI��������44���0.;�$�`h1va|�*C���+����O@�)I�`_�A�ΐ�c'�����bd�%��.Ү!�d��J�'&|���&�<�(Of�3��R�"�t�W�����Ovd��,m� 0e��j��,��'k2�e�	��9{��V�TiXx�4_P��w!ߵf�/O?7� L9�E��,Tr�/��dy�9R�"O
,��NS,y�x�0@ �A���3�V�p�5@ ��	ד4O�����d�,����ԅȓU�ԉ���'
������t�I�ȓjoܴ0�+ȕu�0`X��Li���ȓ�4�C��R*J P�{%��+"����ȓ%K����!�;R��f>!��̞t�h"aPҀ�����H�ȓM nx�&�נ	��١�{>&�ȓu��b�
�+-�UY�k�8XcX0�ȓSF���`�ϓ8< }��$µ���ȓ6P�� Ì"J���,�/�$��>�f�Ƶ1H5AވA� A��F���y�ƙ�3�b��/è��ȓ+�N�G̅jIH�xcNV�<<�ȓa������^:fM��Rbb^�0F���O�9�,P�~�T��W&Q�ȓ+e�	D���m[  ��W
C]&��ȓ[%����͕�c5�$�G�z&�ȓB�(}y�o�:b/6-�f�FGY��ȓt�ĐX��$!Y�N�;���*�>D��i։�1A'>L���J�V�0A�9D���3BK*Ac̀��j�=q2���`"D��sB��+<r�C�Wp_e��) D�PbS�҂<��훲�(����@D>D��yª1L�r|A��,;"L �l!D�0W�E�l�9��)�Y�6�cd�"D�,b�M�� v���
R�VZ$��#?D��I&Z.S|TpeѨnpZ�؄�1D���jS�3��p0�㎛=�t�5�=D����	��+�����=2%��P��>��@\\�O1��ϓYԀwi���=1Ꮯ\��y�UQ����䄿~Gr�)§|����,a���'i=�(�J�+Q49�|���I���T4�)�'X��@��$�~� ����Q !Y(����H{I���y��ɒ�_k$�k@�ȩz�Xsd���.��f2��].�a�t�5�|t�.Բ7���3�փs&rOl;eG
-����Z�O'�t�מj⌕QB"�2��jP2��	")f0'� d�a�`]�"�.UC���o�Y+�gJ(�~b�Z:d��|�՘��"���3�4<9�*�5K��ł6Rw�<{�h�c��'����i����ɉb���i���?ctt���x��'~���)	���*��>�6ĢQU�I]�'|~i�U�*\���O�vݥ�O3"���`	�P�<2�T=3���*O@M��� �R�Z�$�����*�̝�a��Q�1��HD*Jq��)z�E _���S�O��ab͍<G>����F��M��J_�!���+`��L~b�?�O�IP���lp�D	v:p
r��3lP7m2���Y�(��?�@�GP�S�Ċ��K�{i�؉�'��{h���'�'.�A�� 0@� ��.�LA`R8��dN�<?��;�4��S��OT+�H��v�#���|��1O�@q�O)�MK� =?�Od�O�p(� d=8#�h$\�Qu�L��lRf���d5�P1A �<֔Q���W�Q�꼰�,U��R�d�<���r>)"����z��_� �+En��<a�'�X�`�r��Oq���`��I�
*~Q�����@�[���Ue�6slp R��P$>�{��<�c���U�z ��ɀ&�^$��;w|QU�G��S���ɏ�2ͤ���E���E���X�'��I!�@i�S�'h 
L�ӍC|I�0O�>&�⬅�t��<�!�Z�{�0���D7u����"�"b�R�u�h�p�������9N��
'��I���c�R7l �����)��rn�\�3��fu��x�B�K�	��[���x��PI�zc�$2uV�!�Q�w!j�ȓ=)̰z$�� ~������"aZt0�� 鉇k�:Rt�@Yp��f�&�ȓd�"=�W��<H������UD�i��S�? ��Hr)�
;,����	��Ay�"Ox1��ԌF,6+)Y�	�����"O�C�n՞;��-��Aw�t
�"OP5�E�s_�u
� ^�<ϰ��W"O�05�ނk-�`��ʈa]��k@"Ox8��ъV9�����V�)Mx�:6"O�I����<��C�ې.@>���"OjDzF��)G��������?jL�T"O� �a'�5��՚2i�.j7ڤ��"O(=z��`D����B� \:غe"O�0ء�R�>���D"��"�
�"O� �G�C�y��� A��|q�"OyY�@�s����a�\�`S"O��g��^\��­-��y�"O�|롮�)B�����̀���"O:��B��54�	ƣ$t2"OPt�Ă	<� 4I�a�/3��;�"OlP ��D!���{�A@"O����) �e$l!I�� ���*"Oj�a�L� ((���n��	( LxR"O�QC� ��fW��6+� ��J�"OD�e�R8'm8��f
�$�d�G"O�Q%��v�<�D��:��4��"Ox����L:zH$HR2�Ӭt*��"O� 	Ӥ�SK�����K<��p�t"O�x�gĞ�I�D�Kũ��nW􈰵"Ol�*W>�h��� �P�q"O��
�g9v@�$�.2����W"OҸ�"R�n�0I �V.P���Z"O �ӣ�3�lS�/ *b�{0"OV @�g@�M��<[f��I("�""O�̨V��	M&�Z%��*�\��5"O�����ȩ��Z�X�DtF���"O|�@��<Z�P�'�]�]�*�"O��@��<U�a����$�X�X"O���"�A�4r�ĽYn����"O��Ю�z���p	pT�#"O���e�@�)����g��+0�k�"O�1s��D�:��� �f�q���"O ��g+�Q����1f���}�"O� ��%��<��n��⤽(2"Of��2ȉ�|�t�� ����ȃ"O�x��.Ǜ	�Pc�dQnw� t"OH�Y'��Gp����P'\:4��"O���d$S܀���(1�a�R"O��	�� ��
��W�>�Ȥ�"O�z6i	J�`쩆�Gp`E6"O�EPU��	_�(y%/�-_ʡ�"O��O�T�4"soѸYq8D8�"O� ���˅��"1N�?6�4��%"Or��ħ�.��03� �vH �z�"O���%J� �Y�#{2�BA"Oh)aeϖ�~
�� �F�qþH��"O.Œ�"
p"�ɇ�!M�� "O.(�"��e~����Nf�A�u"OP���jкh�Fm��9L�Q��"O�\��ȓ(��y��AM(Ϣq9t"O���ɋz�$Х�(?����s"O H�1��@*�y*�&ܰ��a"O<́�G�	Z)�A��J3+�y�O�������"?�y���	�y�AV�z�ô �� ��8�n4�yr�Ɩ��2d�_�v!���`�K��y/.���+p���A��y
� ��pk�<P5�1M+�,�"O�p���;&ּ���ˈy�6<�F"O�d�'A]9[o�@h���'ﴰ�B"O�ST�E�f1N	���'$�,q�"O  0��;�z�Kf��79�ͨ�"Ol���ɞ%6΄�j��)6&1��"O��ᱩD�[��� g��S"�@P�"O�����P�{�6��Ĩ��+���Y"O"v(��O�m�W��(+p�P��t,�5�&�[L*ȼgB�{Y���ȓ0��3��p�\�i���p�ȓ]�U�i��L{���3c�>���ȓvv��v�ޏ���HuL�:����ȓ �0�� ���,�ұ�7�5G���ȓl���Ȃ螎,�*LHT���v�P�ȓ+`���A
d�tۑF9�
ą�>j��0�:D�8 ��{t�ȓp���!V�x��g�8�2����ҩIb�B+��m���DU��m��h��Xygd]n�H��2LR7;����ȓFɢ<
ԭ��>�3���:*X	�ȓu�xܠgi���ڼ;r�+#�Ň�/���JΑ#2Að�ϑzXH�ȓ���P/<o��j���F@(�ȓ`72h2	�pRmz�`U�!f��ȓ@~Pd�EL��	����6Z�,�ȓ?��3@U�c�,%��
N"2�FՆ�a��Qbb�>-HFM��#N�W	�q��iM ��F��!x��Q�K�Q��U�ȓsJ=ŧ3wd�٠��I���ȓPNd��U���T�5�uHy��=��n�$���e�1fH��AB�%��M����2V���D����s���ȓ84�+v��P��T�e��2j���\���j%F��I+��	)_F���Z���aT]�_��bGA�p���UpX�۔��ji��Rg��i�~��ȓ;@M���#	P`�n��Ir���O�l�1��5� �V��0
�`�������)S$7BP��fN�S��y��u��aIE�?*6�Y��ܕg��ȓ�b,`�	*o��qp��V��ȓ^d��Pʻ[5��`u�\7R��p�ȓK�52��3K��@���4[2`��0�Ĉ��3#d
����!Q`��eD��:R( *H�J�W�!u�6}�ȓʀ(m^d@��B�ٟ^�نȓG��t(�Ǔ+-�U��R<���~�Q8��[�]H�`&-E�.WBY�ȓ��M��OS�Ib�0��C��tǲ �ȓ@L���>&�(%O�5����ȓ���u	}�d9�j�D����V��X�d�شF����F�K���ȓ5m�I�c��N?܉��F�`_@!�ȓ0�az!R3e���3E
� ��ȓ<]`I�R�.A��3IV�= ćȓRhޡc$�)|Ӡ��K�BɄ�x�Ё�m�#xS��h�j��#��\��5^f`�\�H�8I�%�� _rņȓE"�;��¦a�f��ë͈q@�\��,Ub���,��+7���N`��Kj&٪'.1P���aZ�zE���ȓ)i��9����a�1Oy�U����J��t��y��+CQ���S�? b\�.1d4�`ኝG@�|u"Ol �2�A&\겤ԅ\�c����"O�<h��� >s,��QDX�H.Z�c�"OXaQ#àu0�RA�I7�HP"OX����71V,�#��s��<��"O����R�y�fa��l�gl�6"Oz�&�J�e+	<tg�<�v"O*�	���2)JB8�@K@/$e�S"O�	kR���X]�W�>#a��R"O�����W�MB�K�;��@�&&%D��"Յ\�
0z�Y��M�B��$ID�$D�(����<0˶�R�"_�u)�t��"D��h��üD���G2P�f�c�� D�0i�)�O&H�r�͘G��Y�%�=D��p����Gx��EհVrjVc'D���$W�-�h|��;@"\	0A D�T$a �N$"#���F)`  D����	��@P�Ù"M�Pî<D��*t�!v\y�(�S}�(��/D�T˕o�Y��Qd��$IN��qת-D�x�e�.]qni
E"I7�r{�0D�8Za)ԓ9���X�
C,`I���)D�ܹ�A 2������MUJa˶�&D�pA2��!O���{�Q�[�0�s�#D�p㥀I�X�]�6N�	e�ʘ�+D�L�f� %	���qB)�(!����!>D������Jօ�&P���QD�.D�`��*�`�E2%O��*M<��f�+D� �G�}�`5���&ʌ��$D�@Х�]�/@f�A�iV��
�$D�����ޑa<�!Y72,���*'O$D���vϔ�;*� �A��*ٸ|ra%!D��0ؿ!��0�N>dP����#D�`�F[�:�m �ņ0����"D��R��m��qq�!L`ܬ��b$D�����(�<(����:2[�����4D��$	٥�v8#�0;���zD�4D�|�H&�Jw�`�NPW�2D�\ ���9/P�2�!%at2 2D�P��"���$����m��1b�*Olt��m�;rx����M����"O��&�Y�cC�����M�:5��"O.�v��Ov4�s��zŔ�Xp"O��m�<�, 9!lHy�"O��HgC�H�� [,.�2�/D��)�@v���{5�$P�$���:D�k�	UU�P�6	��;�
��� :D�x���<������m¬KPD8D��R ��*����J�R����e6D���S(�+s�D){rዮy��y�� D������	��O4�\XC�:D�����>�`XN�#0�<��9D�80�	v]Q�ϯ����q�<D��Z7&*A߬�*-�#�Hqs(:D�cĎ�B��L�f'�G֪l��b:D����朠�� ;@�	C|�2ɗl�<�Щ	�y.�K�a��\K��+R��\�<q��G��I� K=r�L|C�\�<qЎ]
���t�̓y���c�W�<�F��- @  ��     �  U  :   ,  <6  $@  �K  S  UY  �_  �e  )l  ir  �x  �~  1�  u�  ��  ��  =�  }�  ��  �  f�  �  ]�  ��  ��  ��  ��  /�  �  ��  + m u  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d�=����D��j��%x@�U�1��Ԁ�fX9�yB��-VI����	�15�.�8%@��y�EK�4� �.A�Q��ϖ��yB��)<N�C��	>+��7����ȓ�����	G�lP8[�)� WD���ȓ@鲕�oˑx��T w�&+F0�>�דQ ]c�o	-WLD��4�$��U��I\�D
*�x�gH�a���f�Q��jB�I'q� U���JD֚mf�S�%8<B�Il%$@C@�]�
����юW8B�ɥhvш	�&�z]�hN#6�f"|BsOC�g��)!@���N��Vc[wh<a���A�^%���6O� ��ĭW���QX��#U��[�T��S�]W
���F6�O��V|ȱ�hP'`$r@���bm�ȓ���b�r��)7��+G��E}�?O"�|Rt �3Lt0d�B��
��M�<q��0%�*�	�#���Z�� M�<q���*P��em�N�\�Ѱ%JFx��Ex"�E$^D������c�X)pS�A.��'��zҫ�X<�((�'�]�H(M���	��HORc��@a�ͷW��!C�S��!BL9D��3��ݛQ_���w��%:�)��4D�����d�e� �Q�l͌�B�`8D���3a��I��UM���F\ "3D��wǂ'�N�(�F-Q�f(-TfC�)� L]��"���SĔ	��"O����R�n��q �V$�ؠ5�Ɵ�E�Tf�T���A�:~��ڕ"۬�y�L�S��2��Z�4��Pf�F��yD�"I����B	�D�fP!�yr��L�`BWK��4̉͞����y���.U�"��C\�%L��pc�G���OR�rc��?P- �g�"p��S��J�<i�OB*7��M�e��|n���*]�<)���*x^p�;�L�8Թ-Ic�<��� 8Aq�3cRe^��	�v�<��N�#N�dc�O�)-����Bp�<q�8Y�H�#L�`��k Mk�	Z8��+��[֤hc"|>�Ӗ
?�Oz�p،E����r][�.��E����ȓk"l�m����yf�V�^ళ�O���$�� hc�= ��J��H�1�!���/��$�օ�Q%�Xȱ��J��9�S�O�|=tl/: |���af�U3�'������"Q���y`�\�*V�C�'l��'E��X��۽^������Q�(rޝ�ד�?i�4��$�=r���eI�9o�$��vM�!>a!򄖱:�봮���6 4�܅$n�O�=%>)��Gp�x�͔&lQ�Zd�,D�ث��5e�U��)T�Kcf��/���hO?�$�X�5 g��a"5H�"�\�!��1+)��vG�z"֟�BB\хȓN�F��;��@��;����O��=��R.��I<5�W��v�D@�<92��:^'��+�䛏:A��!|���=Yt��Dx�1"qH΢E<�@́A(<)"ȓ?>��#7� y�E���^�3.DC䉒q��)�� Eg��}awÉM�<�?9�O��>9�󂟹d�
�yaLj�����2�d2�O�4{�nӎA��ȱEGl�H����D���j��)�?�5��
9��!�%kI��{�,(D��#օ�nU��m ��ы�¢��lZ�.5�O�#=I��ի�r@R+F6�fP��+�j<�WM�=s��ПY-nyF�9L6�Qf�O��=E�P�#��������,���φ6�PxR�i�"4ж�M*;8����m�dZ�O4��$��{p�xS���3"� �M��GN�	�أ�}��%�ӘS��i���j}`�'N�"_hB�I�P9�'.N ���y��ʓO�."<i�`,�P�0��b���gFJ��2Ɇ���<��ߧCn�Сd%I$�<$�b���x���m60��ΫY��`RT�B,�p>i��-?ᦢR�w:�U9׈[�LVLd�b̑A�<f��)�]�"��K�hܠ�'����$�U-��Bu�R�n��D��H%����ȓh��)�9�B!abLP>FH�����hO�S<���V��.N�J�c���*s�C�	&�d0@C+~.0��@�;ihC�	�@I��m����k�e�.C�	b+v�a�'��HM�u	�Ò,��B�	�O�峇.L� ��%@�����E{J~z��Vhn�����Q,l8���I�{�<y�$�s��Q�C�Y4v%<�i4�J��ў"~�ɀ4D�OZnkVA
Wb�7& zC�	8;�+�*� m�s�<kC6�=�ç"w��
���r&x!"�`	���ȓm����(N8�T�b.@�r��m�F�����K O�R)Sw��U�B8K�`�:���)�S�O޸pbR>`�Ҽ�T��^�x�+O
���)� ��an���ܑ��*ȏu����T�>	
�-�
	�Ӣ!cC���gꋎr���#ƔA��P>\T$�5�[[j��ȓ;���h�G@;q�؍#7�Yt���(b�	����v(됬�6����wPݘ�*��LN�D*��ȐBw؉�'ў"|27!�5k��PЂ�+�f4 N�l�<9�̃�Ya茓a� Yʄ�(�e�<�$�H�YRsPA �mU�е�V��$�'����ĬeB��p(�>��Ik
�'�4�k�CR$e�(E��9'�X)��'�'
�NY�ȓNg�R榅�/�*�ȓGI��A�ɏ�! ��qi��:p�����hO��$�����!��#��{��H�1��C�g��U�r���j?N��"��4A4B�	�m�*�HT��C�L���	J B��S��!	�O�1�A�MY�>,�c��B5�'�� �cl@)	���90��F�Db�����8*D&)�eH�=}��A+և�e}!�DT@�ut(��_y�u�
�k]ax��I1K/
I3�*÷3<~�����5h�tB�79A��Ań��S@���@?"Z"<��w:��s�E*s1Texӽ�)�oA�<Q��8����'*T�tV��֍�����O���7,O�)��.T�4
0=Rrϋ�&rBl0p"O���"��JBt4�a/��z�,�f"O��P%Q T4+UD<n�H���'�Q��c�¶�`:�g y�\0 �/D��a�K�.u��IђnI*l�T�C� D���I��^�2@!%��f
|QR�/=D�p�#JN�x�z����VR.�q��:D��;"�ǜ���HbLN�DH���J6D��	�� ."�}����}	B!0�5D���!��8�PAa%*ȡ^�=��%D��H���i��m۲�9I �"(D��C"�Y�z�.ݙ1���=� ��F%D�H�c�]����@K�9JHTrb*0D��!��/��Q2�mI�.�a�cb.D���Gl��M�l0 B��'%�Uq�-D�D��� )�p(4iP!Z���C7D�X*c��u)��[R��4���:sC!D���e�m�l�0��G��^�Bt�=D�@��*�3f�=��`Eq_ 0�$:D����ꋠ]�v��N�h�)��"D��+�Jp~䁩u�^�O���P�?D�*�Ɨ.���pflׇ �����8D��9@�K8��`�Շv�$��G 9D��R)\�sR��
�.҇g�cU�8D�K4�\�We�	����,ŔL�,;D� �&�O�*	���(�Z�Ģ:D���7�Qt���H���+	L�)�A.D�̡$,��j5��E�@�<2�sׇ9D����	 1�"a�
`�HpU�6D��UEU�1U�#�7u�4���5D��XE�D�1�.0��O&�ޭ�I2D��#�� �Nx#��7SЈx��/D��PSmT1}��Qp�k��vI#D�d���]�z�����&-h�� �+D�����ќ��T ⥉�MJ(['�(D��IC��8����1&�{�t27b'D�B�B'n�-Ww<��Qh&D���ӁY,Ba0�p�E�K=��C0D�@jF-�7nr2�oA�v�l��*D���h]*3�Τq���-h[C�*D�� <ز�N�z�}� ��~���"Ob�o�'VAHPq󥂸y���"O��S�ƙUi��Ps���b��"O֠�Ƙ:Cy���b�N ��j$"O&Iƍ�72� �̨]�6����'�2�'��'��'�'�B�'��A6oXb*���`�ݨ �VA��'���'�B�'
��' �'�B�'�Xpx���B��� V@�0@�M1�'���'��''��'���'2��'�n0���q��Ch:	����'�2�'�"�'��'���'���'�N�Y'��>��q���^�D�y`�'���'�B�'.b�'���'�b�'��p�1@S�n��tE�t�Hd)p�'"�'GR�'���'�r�'�"�'�S"�$%Ԣ�p� ș4�N8��'���'5��'���'���'���'�t$����k��끣�L�ƽJ��'���'#��'��'���'��'��	:Z�|��E4F5�iQ���$�?����?����?y���?Q��?��?�P�W�Q�DU�)A30Ԩb�W��?���?���?����?���?����?��Cd9q��L�hk�,J����?����?Q��?��?����?���?����a���N.�uB֦�?���?9���?I��?���?��?����ؒ�G�{�h��NקA���ڟ4�I��h��џ���󟔀۴�?�T�}q�k��|BP��.�����Q���	Yy���O��n�g&AJ�����ڹ
w�T�\e0Axv(2?���i��O�9O�9oZ�a|�Ћ���fH�9�Q���`�޴�?Q�P-�M�'Y�,ֶ}n�	I��	���U-!ը�
ve=ې���'�%�1O���<���I]P*���s J�m�q3E(Z{X�m�=7�
b���R��yG��3P���Ԫ@�)X�B4�N�4�6���������`7Mc��AA \E��8�h��'����'{���UN��6�Hbk�Z���D�'���k@�Q�8��k5����@��'��@�� �M�'��k̓\d��F!A��p� �	�u�@�b�>���iBz7m`���'q$�P� �8w�t(A�xd��O�,
����):��@r�	�,B���	�?Y�Gޢ	�M���!?r(86���<1�S��y��f:�'�*;ޖ1iwү�yR�kӤ<�A����4�����h�p�`�tC]12�1��NW��ykn��o�ß��˝Ҧ��'$���I֢|�J5	AK,����qhƣ����@NǾ	ø$aQ�ԁ$躈��.I�L�{pI��(�-��2��4�Y���G&�JX�y�1L� 2�=��M��L��}��'������T�,�REe��#+���ˏ�(bf��Ō�)z@�-7.�0�J��>N>k��$d|X{3`DE��(H�%�e�:�ZR�X�[X�[�FM�p%
���*��V�Ĉ�Kr촩#�I�����S�Op��eDH�lzM1�)�%8����B!�eK�A��AﾅC@MG>BFJS�
�M���?�������|x�H J(<U��Q�]q~`a,nӖ�$�O��6�<�O.�T�>)�iO�7�8PtC��O��5@�"Eݦq+.��M���?i�����x�O1�ː�S�@������,Z��� �k��e8�/�<����?��g̓�?����9΀��!�H�P;�0J�L��-]��'6R�'�J��1�+�4���$�O�8#6�dc((�a�G�Qr�qg#�T}R�'>Z��h�<����?��?l��n'gS;�G�l�B��i�"��godO�i�O���<��I%)
p!���,N��
 Fh�6�'� 3�y��' ��'�/s<I�����O
�E��5Br�+���?a��?�+OR���O���r�xyZ���(��
H)1Ob���O���O<���/2�ȭlZ.�$�P����S��,��݀8���+�4�?9��?����?�)OV�$��醊a�.�V䎿b	�3���|@�oZ��
��^ӟ��I�P�	�;����ߴ�?Q��O��S�@V� ��Z�/J3Vf�P��ik�'�2U���	 � �S՟���]�v�B�
_�����I�=x���o����I����ɽj_XM)ݴ�?����?���U���[�C�/�~�S$_���ˡ�i��\����z���S�,���ܴ~<p�H5���t�9�6l�ϟ��1 fR9;ߴ�?����?Q�'�2�`pi�c �=@NTAVML+G��Yz�X������=��r�i>=����Q"4+�$$��E�� ^��+V�i��4�v/|���D�O�������O~���O�0�u�n}y��
4��Y�#Φ푆Ęퟐ�I|y�O��OK�L&a��a��PC����+�-�7�O��$�O�|RE�Dᦅ�I͟L�Iɟ��O�L`��˪ �m�����dӚ��ܴ�?I�r ��7"�<�O"��'���˥6�$ B�h�#F	��,�L�
7��O�lBWb�5�	ڟ��I��,��.���3|(�����Z�Rǡ�=Z?�7m�K�.���4O*���O����OB���Ox�+_DpP��@5s*����P '��eҢD�Ǧ����8�	ៈ���8ʓ�?���%ì �WA� ��]�C�	`ZPϓ�?���?����?�/��1��n�ئu&^�J�BUhuC��#�p�0�o��M���?���?������O��w7�k�=J�Cě�)����D>Y.���'�|�ȳ�'�2�'y��P�;�>7M�Ov�$�a�0�)�Β��0r�	��ux��lZ���Iџܗ'���mD�	s?٣ݻ(=T԰R��T�ĸZ�J��=��ߟ���؟�;� �M[���?Y�����y�q��,M#'w0���F�t�&�'��	̟$�Q�y>�&��s�� `��ʚ@+�ζe)XtC#�i���'� Q��AeӦ���Of�����I�O�(�(I %�*�	�11��)X��	r}B�'3��E�'Jɧ�D�~�%J+1�,c���[PdĦ}�dH0�M����?��������?���?��J�W�j�"d+וWd�`&`ׂ]ꛦ/�K��Isy���4��d5PrL�sLԲy-B�a��y���o������@`�+�M+��?���?��Ӻ��G�8�k�.O ,�$:g�ަI$�Pxw�d��'�?I���?�����R6�H)j줭3rLZ�p�jDQش�?I��	E���'���'(2��~��'�<��T/T����:cP����O0�A?O��d�O����O����OT�D�)NvH�i������+fOB�zU0�����ۦ��	�l�Iޟ0s�����?��fj�b&J��<�
�0� �<.O��D�O �d�O~��ޤ09�9lZ�����1Q�'�~l����>�Jm۴�?a��?���?�/Ov�ĉ�_��);��!�p�[�Vx�Wܱ��V�������؟�ɔ&I�0��4�?Y��f��DrW����a�-m��	%��%�M{���?������ORAs�<�������W��
�옐� ���Jc����O����O<�����	�X���?���n�#g�6q����&O��� ���M{����d�OL�R�ű<�,O�i���3-)�d�+�Լe�����IƟL�U ��M���?����:���?����y~p��%v`�a�*�b������� I�'��Sk�I�M�I�6ENr�X`���΂Û�b�n�6��O��$�O��	������O`�D�d���1$K�_G��z�G�R��Um��o�:-��|�i>-$?��I�3���b�J�=z�E���޺T6LI�ٴ�?����?9I*5>�&�'	�'f���u$i˼|���J��h3��;�M�J>1���<�Oqb�'��E�"mN�슢)E�2 ���nt�6��O�D(5@Y������<��şhk����	l̘���}���D#N�j��|�͓��d�OZ�d�Od��O,y����oq�9�u��8m���fPi6ʀlZ��x��ß��I��)�<��g�N��._ &tX���j�J/�ȊQ���<q��?q��?Q���?�� Yz��f�i�ځ��8+svE
�nTd�6:�fӨ�$�O�$�O�d�<Y��$r�$ϧ�|	�H�]�M��Toc�@�ǿi��'k"�'�����t�Ĳi���'�iK�B)����9֞`�/~�b���O �$�<���V��'�?��'��h e��oPx;a
^�Uf�H�4�?����?A�O���7�i]r�'�"�O
@M�Ff܌?XIu�?;�HM���n����<���l��"+O���|n�5o��Uz�g��8�8DK���q��6m�O��D�g�5nZ����ܟ���?��I�wc���`T>0S��ЗU�	a�OZ����8���d�O���|�J?�s��F0�����)2�ٗ�c�Dqa�Ʀ��	ƟD���?-�Sݟ��	Ɵ����C�%����b.ـ�x�A��M�s�R4�?����4�h��2���: ����J�'b����ԓ,ڌn���\����`	�LD%�ē�?����~r�շz�d��Q��_P2dc��Y�M�.O�d�v��?9�	ǟ����z%L�R��ɡ	�@E)��(z�c�4�?��ͅ���'���'+ɧ5�e/8�8��W�GI҄в���M��b�L	#���$�O����ON����2��0�����FJ*<y��W*/�'���'N�'���'���5	�z`�TK�e�0%x� p [$p�BV����ҟ<�IYy�K�2��S�M�����YK �"S�j�d��?Q����?Y�O�d��U�,KU���<i��¡B/~t��S�����p�	DyB�� e�^ըU+ǎnhI�'E')�����O�a�	e��ڟd�	�i����}�����~���͗M��H��AW�;��6�'��Y��{��ֶ��'�?����l�3��U0}y���l���r�x��'��-O�z�R�|��t� e��z���*�KZ6�haеi�	'81���ߴ
]����������V򠙒�R��ܐ � vC���'RdE!5�|��$��0I� �
��72_�u��F��M��E��
��V�'���'���.0�$�O�I�`�����$zpn� �t咓��Ǧ�B�)=�S�OZbNC�T��`��̧.����W�!6^87��O����O2Y(#��g�����m?9@)�s��Y�����.��Uo�6�'�ě��܀%>��I����	�8��A	�O|)5N�1J��ٳ�4�?! ��^��'R�'�ɧ5�Ë́:P,�XF�߬G��|,J�����Z�b��<���?�����%T�6�ՠ,���qR�&]Z�l�~��ş���\�ş����_7l��z�J#/J��zAxT�g�Ĕ'b�'��O9�Q���q>e{G�U�ER�جR/n<P�!�>���?�I>����?#��9�?�Ai%)�;��@�R��Q� 6�I��`�I����'+���"�J�V�tKD���  0���-�(1lZΟx$�T�	Ο��e����O�a�P�˝Rr��RJ�s�w(���'
�U�8��Z<��'�?I��ДAq&�c�΅I�XY��x��'���2)��|�����J�,_KZ�IGÜ�l�p�iV剘8��(��4-7���8��������-�v� M�7eͻ}��5�5�i���'�Dq��?�S�b��C!�Vk٘�`ק�q�,6�]�&��n�������� �ӭ�ē�?	%Z%."�Ԋ&cF�JF�2�^+1����ĺ�yBY��q������O����OЈ� h�qd���O<��A�?�%QS�i���'�2���#��O��D�O�I�L� X����&y� ��`�6y3N7m=�Ć=$�d�&>��ߟ��I; �Ѹ�h��y��4���ָn���ܴ�?�PHN�zX�&�'�R�'sR�~2�'Od���݂=�F�Ȏzꜽ{ܴD��LpgE�<1��?a���?�����I�q����jN|�� �ҡd��\1@�S����ҟx��ß8*��h˓�?�@h��&�܍F��	���@E��=L!�P�'�͟9@� ���f����B@�)*�E���U�P�S��;�y�l�P��)�ǝH�@�*�_��']`��6f���E�*:���E�Ԥ+�x�v��/$�U�&_19�v4�"rڦ�#SSe��es��E+F
�@��!�����R+҆��!%
N�vhb�	^
j�dᩒ�ˑBP�0siЩ�%÷	�!��l�􀗌bR �l�.G�i��-G�s�1i��]2s(�2�� �F,Stf�
 �4�H����9`��?��mw�JaY�N�4��� ���4=�wJ]����Æ�����@�6(XH�S��S�Kg�,��X� L~��Pd�l!�4�e 	�}��
l�큇.�:q #G(*�<�O�}�0�'�2��t����أ!:�AF�s����si݇�'�r�'w:|�a���tF��U���"|v�aÓ|;��Hᦢ_�^-���CY5�$D�&	��Mc���?��c��<�?y���?����sw�u�8Q��¬���U�ڥ��'�����'hZ����I��4[���!U��=!�{R�޲o�ayb�ҍL⁺0���Q�B
�̸'�"Iaϓ�\�!"�:Z�l�k�.�GVlńȓ[����/gl:�{�O�����'1&#=�'�?�(O��rnT1{��3�-)p��KMi��h����O6���O�������?q�OVr��)C4P�իX�h#��/B�>	�1&K-c�!P��[��M��n1�6X8���ڃ����,T�N]��q璀1�q 1.΁��-�ߴCC
\1a%7C} �yr!% ��$�tJ�6��-�!�C/c�����?�K>���?��n�8S��f����0eL�7�0>�L>��l6|[��	�	w�,��t̓f�v�'%�	�z��8�4�?����H�	Fǟd����ek�^7.�����?��.�<�?����d�S�'�M�m bV�$�bII��@��� �+���y���	�4ƀ`Nտ?T�CT쏹<�(� �W��PA�� P����{RK�E�d��%� [��O����<��hʩ�T��Ui(8��M��<���?������NNd��k�&r�,l�/1D|�|G{�O xA�1��@6&x�h��R%H���)�����
��nz>���G�Čګ4	roI�IZq�����
D�Qq5�+���'�D;��G��9 I�/G��T>��O��M�g� ��hx��gA�G�p��O
]a3cD��a�#=��"}��aА�A�	"h��W	�[��B�E��'��>���K���`�D�5!�P���)�ԅ�#��I��-�_�sG�'*z���	
�HO�)8�]�|�mSF*e0��Q �Ħ��I韠��,?֌,y�N��`�I����ɹ�u����������EƎ\#	����0�$n��<�7��-�dʱ�|��۹L�
D��F�>hm��P1��	L	�t���Z���@��W̼��□{����y�� �Ǽ{�ʹ?9��3HP*
�0e��9��6�g����
+F��Y���	;�Y���6W��
�#�6r����s]��(#���B�ɕO���\ϓ�?���?���hyb+��L�z���M���\����+�Z#�Q�L���'\��'�x�]����	�|�c��Z���;��g���'�b4�܁�i��E�.q��A�ay2���/*�x�PA
!a�N�Y�B�4C�45�⌇� ��J�RZL7m�;4��%�	s¾�O� �A�'	Щ2�ԟj��[�
ə]��'�'�����X�?���	t����T�.s>`Q�IJ��'�P0@:o����W�-?�(�S �>�I��MK���%��OV ,��-عkxȹ��0Ԑh��'��MFԯW�`Т��x+��Y	�'E^M� �Q+a6X��
:l�U	�'4�y�C�-w��$�F�Y��5D�dZ�!�1Z�d0EC��R�"A5D����YH��K��&�:�+>D��z�D�-+z��K�)?�l�0�<D����T��Z$` -ȩ\�4���9D��1���ow.�iaN�!H@�!��6D��Y�
�#+�4kBnA�e����6D�D򕎛M��R"�@�}�vɚ��4D�D��K��8j�I�\�)^`�n?D�����@V��1�X�Aء9�A0D�P�sń�HV�}���S!w�@��/D�� ]�#h�>]:�%�r)+Gl��"OL���\��ȓbS--T!$"Op�t���Y���#�O"'̍��"Oܤ���S��9�ҋ�d0��3"O��%��I|�h��*��VZ
� "On����r>�P���>Z��-�&"Or�� ��2STJ�QO����z�"O|��Ӯ�#Y�N	!��1 i@I��"O� �`�B�A�̑@)ϭM�Q�"O�Q�0 �F��x�d'Б-�F�a�"O�yZ򇕺H��|�$]��)�"O2DPǬC9 �2$ٕ�[;n��"O�b�E��k �Z�$H�Y��"Oܰ�p�۳>�΁Q�:k=�|� "O�ͣ����-��D�K�u��-Y"O��P�L�$(X�*�<��Z�"O�5+q��[���G�<�|��"Om`@��O��0�ČT'@GLـ��&FdP����Ƌm7:aদ߂n�l�����Cx����d)�g?�w0�
�� U �R���V�<�t��� �R�<E�4J��w&���΃�:)�V���?9�bA��0?�#F��F�!`[��X��RaQ8�$�r��٘���c���4jQ�T���^�U�RAj��;q�,��	C�W�a~���4v�7M� i}δ@� 
n�u;V��\��\+��ƥ�O�8�׀*?����t9R��B�T��?}�@Es�&T5���c��®n�ў��G�
Q����|�0�big��	3�%$�V�"�(�2�.|R��p�N;��<Һ�2FJ2j$)���nS�X��D�fcHZ��ӓ4�lZ�Ul���pӖ���-B�`h���0H<��t�;�LV�8��sە�]Is��sJdԋ'EQ`�\KU��u���rΣW��ó�ٰl�4]:��/lw�=x�Q��H�J��p�Y]0�J`$3]�.%٥�T�Iwa{�ƅd;T�-\M��Y3i[ "i:�(t�ħEp��'��uD{�	T�[�>,����fJb���	�\pA�I\�Q��t��I 1r���t�\qC�AL�s�9O�I��^���2Κ�9pL��ҵi9��K�O��3��[�9�b=�dсmL���xRl
5����Bo��:�84&���MC�HS���J�"]ƅ�۟�ObY]�Mnޫv3��QqN� ��)9��reWً6���u^�`F�(;�pzn���m��6i�;6�޹�?Ol1Z�.*}Zw7�
�g?�g���|n=�2�g�,�\�)���=?����'��k��Y���o���9'��"C����ʋ%)�b�3���V<i��W}����=�(��f��|p9�(� /��#�:�� kC/8ړ ��4H3�����vt��	%A�z���C���1�fQ�q!6-\-]�'mƄ"DA@�2�@�TnT�.̬�A�Oz�rA�6G)F5�+|�I&�i��]�� Ո&@��$z�$��b�'R?���T>�|�j�����ر�ljzAC��!���"�]�:��
Ǔc�ژ��bH6�� �$3FJ�9V��),��'挕�w�	��%���?��%c��{��B�Oy8�8
���G�U+���r �X��鲇Π.^�`�W�tb���V̦�붏ހY���9�b�4S*��a��,�&"�ў( f�X� �	 &X�0ɷ����2��W�!�&�Zġ�g��0��>�'�����< L��QlذI5pj�yBɟ!����1�j�Y��͍�M�&F�b2b�;":O��u��_�	�����s1�[1<݀`X�T�'��8e �.Wþ���uaH�Jt�n����#��
6��ˡ�)[�y���,}�bO<��?O�q.{����P�W<P�����)�>�����T�p,m��
��2Y�r}��W R���'�P���'#�']r|��G ����wܠ�Z�G˅.��C�:WV���D�.PV,��R�<a� �N+�ɶ$�Lxâ�Z���:uÇ
`b��8q	ӧJ�`mIFؤw�ڜ���=�	��U:g���.>�Y�����?�d�H�3�ʹ��뫟��!�/��	�
X�'C�=�U�\(�T�c��S�h#4!�0΃�΄�%FEfi:���	������/V(*���
586MҔr�b��'��!�D�3�i7��Sw �87��w��(��w��^8�������߱K��^&���!�
���Წ�4N�c˓i�\��mIü{��R�P��8�Qe�E�d��ǂg�'o�P!���'h�e��ϒ�<��ڶY�Z�Vf�j�����A�'wr3T@�-34�k�(F�VL�Ԁ�Oxah�N��N���BJ�I�QW8O�%[e����05x`j㚟H�0�+?�ԃ�n�֝���%x���p�����a͹�hQ��c[+'� ��	MX\� e��w����I��ܠӀ��%I�������4�Rֽ�� 0��u�<q�j��$o���r�"%S�gp��$Q�2H�;I��9�0-F�O1��K@eb�X,��4;�(Ok�ղh�b�LΧ�M�1��I��Ԓf�*u	�G*M�Ez���'=k�La bY�y�+���y�N�?/(r���E�{�|�څKP�3Sd��L̓i2�xC��n��1�����'$5ڥ%_4�
�D��v�BȀ����B��P��,X�$4lZ~~�������_8>�؁8��[�a2�KU�κ�����4P�tu�3DP�?)��[s)B_�'�N��*A6ER��֮l��i�4@��XJ~2�U���ԟj���N�>�f�f"8��#�Iv���֊ۇYᦘ��{|nli��s�=Qt��*���xFK��>�D����H��y��3��E��0� 2Ok,N�+^5��C7\QB�:W^�J���WHY��,�h�ſ>9S��T�u�ʮS�R;gX 9����O��8�'�T�� �8U�q�'R	9�`��^<�C�	�6n���^w����k�t�i�"��ly��O6�?Y�duϬ�`xg�M�����
x!��b#�7�~�Ӡ��O�ϓo��x2dkш�m�P$���z�(�̓8_��AZ����k�����DW>�ku�R��0�uB�>��Q�A�2�O�Q�B��rZܪđ�<�^�sf��W�v�"e��M�O�+2��Mq�b���~�!�	.�ϓv?���D�$,y�\��v�GyBg�6����T#Sa$-{�L��~r�N��ɗj��r�x���B�B�����4yR���y���+�A}��a��1Z���|�H)'�1I�okJ(;��H�uЎ��t
�$}�0�����sh��Z�O�����O��à�#s PІ*��A �m�L�<y:6o E�@��dX�@YE�x^T��F�͕m�������1O��GzJ?I�J��_�z���ǧ�,����[ �z�ᒦ`�y��;tf| aHO.j*��T��4d��R� ڔ(�'z�>��Ԍ��L�8I�PL܃z� 豑�O]�'�r��'�	9�p�����Guj ��O�v��z �iU�!EUZԀ�I�ZP 
��uAjע�
��h�0��@?�T3��f�x��&�3���uHZ#��b2��X�'Pr��� �V�nkLT��h
q7�P3�! -�p��T%z	�Q��:J1���8^f��pT���LՆ���X�Q��F{�.P.3�$)Z�����X$�ǇVj��d�q�>����VU�&.�9z:�f�C�s�|v�I5H��	k�"���S�#+*@ӧ�7�$)G��2��`S��+�(O��կ�w��%+C��>r�bW�O���,�*(�U��4Հ��5CϮ	��DY�b~���,};&AA ,ېJ
z�!] �'.�EkBE��8���]��n{�jN�f�P�E�C-^��d�U�Ɛ�~�g�'�x����$`U� �TT�8����?�1BFN� �KA�'� C�-Z?pnFL�U�'R�ę4�P8���O���1m�!`(��	v
�:�����)U>��'Z8�0��#ABY)�ħ(� CR ��ݙ� ��?��O�ܛ�(��{�|\{J �$`e7O����އG�(my�@�*9�<,��팢YG.`��k �Ɍc�0��1h�G�Tȫ�i��/��O�TS�!�,UP\���2���H\aR�@�Pե_a���'�(єR��O�|���ĵg&��E%�n�Xڧz+J]yb��9��P�d��5vJW�w:]��ǔ���H���K��y��z��ة�ox�"�P8�B��5�Y"{
Շ�	�0���p�cݱv�������F\+~H���! ��h����דv:t	t$
�e�lxؓj�#_wt]r���N�0�Ra�
fZODb���0`�ܔ9�k� �1�Q� �d���t�ó.|��G ��ke�@���'�Z*l΀aq>=���0� �L<��Ě4b<��34!�<j���0!��?!ħ,cS͡��'�b7M�)Dx5�c`2�ɢ"��d����8���!�/,�-(�_����7A�=R{���4更{�mSJA��Z�oX���*�E
��64�lŞu;��D@�]��!�ә��ݓ6N�kaxbF��%+�
�\�%v"��%8y&��)��j��zF�)�M[v	�0`�,��@U���x:�F��e�|0���'�pjK���i�>���K6���z'k��^�T�C�oð"hD���O��� |���UcP��4�:Qi��� `�@z�ɡE����d&G(Av��3А5�V˓\!�k�'���Yq`A�<�0�Gy"I� $��8 ��*q�����M�,�8GĂ�Q!&L�@���gI�j�����P����T�H�����&h�*�� �q��K�I��X_ʰ�Z������Tӑ!��P�-찌Dy��E��O�΃�3p,��I�	Slr�g�U��}�o	�w<�4˚+}���ƚ2��`
�n0p��%���O���3l}����� `Yq���K�2��0.?D,�u!L�6�ʣ=)���2�y��/Qz\
W�]S?�@�́"�P퐐F�$x�
 ��K?�b��tj$��E x�^q�u�Pq�'��E�&g�yp���C7��"ܴ~�����O����w�ֶ�Ey�O3�aQ�dA @�q�IR6��6�6U��,(�O���!��"#\lt�"�&���zT#�]�*(Dx���A����Ռ�E"��/_�iP�b�����d�,E+��`�b6� �LP�a��9��8���ɠFR̸�O,͛�͙N�O��ɷf.K5�^�c���,-1�2��7k1�8 �GԈO� ��-ֵ����b%�;G@ �ʄ2OBk%��'=|R���mڂ��@�P����O�B�(D�"�|Dz��Cbݚ���L�5=�$�D��#�~҄��P�z��5,:�hK�)���S�D�@�2�xQaA�z朚�.�)u;*G�5&����䐚Z��89��J� �,�TEzߨ�jP���ܮ��	����x"e�>9�h�5Ռ�QӁ�(�΍2ej�L���01f�� �agX|z�0�����pTx�'x����G�3&>��'�f�'6 �J��ҫ}A�d�	Ƭ��n�rԡ���1)����*ѸU���EH�z4t��&.u�
Չ�
zĀ#2Ș�X���u!}��M<���R!:�E|b-�6nHؘ���/F���ʣ��y���	i�:�`0�\�|�P��a%���S����a�D��@�6���Pv���D6��~R�� ��
��@�
|h Ó,dE�	`����?	����@ʟV@lz�}jˣ>�e+C(b@˓I�EuF�Y���e�� ��4�B��%��y�\s)؈T��
����� h����p��JE�Z̦��}��~RA�����1���+���=1�jQ#?�x$B���榭�egH�qlD!H�K��&&8k��0D�xʖ�Q�q#�O*��A���/��(w�6-K�=�>%[���H�i�Ć^0��)1�/D��B�J�V�и�O����G-D�����>`5>#�KH$J��kW�8D���`-ͲF��d3d���aW�*D�$��*Ǖ��X��m�=С()D�Xr�&�>@&��ѪHc.�\�"D��{g�X)Jat�CCņ;��\�5�4D�8�!�W�`G�\��÷\5�) d5D��H�,+4����@�0y�erk&D����L�(_H����^�F5L\�Bn8D�"�F�7	8��Īܤ�b]ؗ�4D����K��,� �D��
s�`��q�&D���J�	�����*'����R*%D�@
D� �m��X7����膣-D�h��C�A�b\Ze=6(�iSn*D��[`&��U�n��tK��p7��''D��z!
�.�֭a���.!�D��{�Tu���)Ƽ�'�D�!�䜱
���e�r���z�c�*]!�dF$Ƞ��D?9��T���/E'!���Uo\��2I��{��� ǁ6!�dE�=�`0�b�M������q8!�DW�^�r��R�*�h����Qn!�$3�ڼ �K����Վ��3!���MڍZu�хQ�:4����e!��8�,���8T|�qgFD2Hz!��^A��(��� &Z4��&9n!�$\�748����_�:�B�j?Kb!���P�����_�P}�$*R!��f'���*D�J-x��f�D�j<!�ΟMºa␈X�4 V���e@�zU!�DF�|�	Z6+�
nHL"Eb�I!�D�'��bD�@�v�NdyAA�OX!�Ā7�z��t��9f���sO��Ta!��Q��D"RD]��(!��?�!��8t@��t���H`�_iD����!M.)���s�|��u�_��ȓ~d�� �a�js"��J]�݄ȓ=s�q��/$>8S@Җ$��q�ȓ:)�hQĨց?$��(�h ��HĐ1p�������e��6�p�ȓk,):���	vPf�y��։�Hȅ�%M���J�	Ϻ%����:�8��ȓ{�Ui�o�PE[<:ka��k�p��+�$A�N���E �i�ȓK�
���ϴ_L��b�؃J�tЇ�S�? �`�7-�%e��|��/ȁ<B��"O衊aI��
�(Soޤ ��w"O�a��Վz.�1���
����"On��扇��]�)L��@�g"O �3TGܾ��K���&躸��"O:�C�fK�$�Դ�ү>�j�"OpUo[ZF(D�ԸM�j���"Op�(�1zø�����4�!%"O�iqJD�4�ܡ�T`I<u� �"O\����V�<�eLUd�P"O.��΄�N�4��FL�3�Ss"O��1��7)�r-� QUdL�Q"O�}�c�ИoF���î��4��`1 "O�`�Bлm �#M�4��U�"Ozh+'��/0�j�┋�Gr1�s"O(�W��gA���
5���2"O�Z��ʞ�s3)�)#Ŧ��"Odia
˼j�6�07��u��d1c"O�t���^C����A���I"O�-(.�#�E�������"O�4�&ŗ+WR�K�L�'t�@"OB�*M�>�:�K��NZ��p�"Ol��i�=��Ո�JM�i����C"Op�� p�H�%�Z�;�jDsV"O|H��ņ�uyl]�Q	̻F�U�"Oj�8�EZ�K_�đ��K�/�"�"O�M�d�����3�Ӯ�h�H�"OrL�!�?2��SB���쵻�"O��I�n���T��@��^�2%"O.`�v�(D�~��dA��X�k1"O,Y�I�1gdu;#0*�8�{`"O�u�cV�36�(󣄁O,z�BA"Of��P�p�L9�c�5_xE�d"O�Acr*�f�"����՚{��q"Od�j��O�z:,�T�>~�p�A���L����̥\�F`���|Ը)֮H Z+!�d�
��aI�J�%2�P��U㗺�!�� ʚ(`���?F�L �@��u�!�?zH��$�ѲjĮ����8�qO���L> ����@ݧ*�p�)u.$m!�d�.��yA�-Ӫ4�i�fh_P!��W�a�9(�
J>C�@a�2^ay"�I�O���j�����"�+π%��C�I�`�>Ě�c�=n�|�F�
z�C�	3Vr����dT�QQ�`΀S\B�Ɂ8���hA�0��Q;'K5vB�I�=Ԍ9*pn��K�nYK �ǳ*�C�I#CL��0��5ODZ�Ŷ�C�68p-�eBE/�8QRDNܬ#<)�	m �ȑ&��r�x�"�ȓ��Ls�E�
؞-򅈝�(���U��lY��X��I���7cP��ȓ?��:,�'2Hy��� �<5�ȓ4�L}��쎋nc��A�֕=@�t�ȓI�L��/G�rR��(�7��]�ȓXc!�F
U1�6Dx��B�o]�ȓ*�2E�ޯ�K��[���Ն�..����J�[LW3|��a��hC�|шI�GC�+4MѲ,RІ�Y�8#,��w��{4g�,p����ȓ7�"H�gK��<UJᤤc4I��b<�R�냒u�b2�D���D��X(N�
#hH�}4�)���_�	��L��L��G��Js*��2m£ ����S�? ��Kv�[a�l�ڥr�]x�"O82�E��a���s��ܩ.]�K�"O���F�ט00�Z&��"^k��� "O����Oܡ`�TM��d�8�h���"O�<�qƐM��H�&��h;BH� "O�I�(�y~dHY�n��V3��"O,,XSD���0�KA�D`�xc"O(�x�j��I���"�*T{\����"O��q�-X�&%ޠI%��?[YM�U"O"�k���(0��RșdC�	'"O��3��F��2ч�A.�e{W"OR�+��� o�1�	Ċ�z�"O��
���/h���C�pn�QQ�"O@yCi����q1Jo4&T��"O`Y	V�� 
����ʕ$ �L0 �"Od��8(Ry��D >`���"O(��6��'䒠°$6��#S"O <x�����rЋ'�,�q�;|O$x��*X�.pb��єn�""O�J�"0u2�/�^���"O�@��V��Db�'�6�2�(E"O\xr`��V��I����=):�p�d�d'LOfy+5�;��぀�8Nt��"O���(X*,�䩫��� �zS"O�t��!CET܀Ұ˔<!`銖"OЕ
tc�.b�4���a�x���"O���V-S����I�$1�0��"O��aeA&b���eo��hm�"O���T��.QYP ���w�h`J"O�AP�j��}��=�5�۝(�z	�"ORy��E�0�(��*��l�`��'"O�١�C��&K"���l�R�	C�O��xZ�G\f���/R�V
F�`	�'��䃓�Θ�j�i��x/��
	�'�$���S�o����jČnk�(��'���'��X��D���l����'�^ip#!ų*��%�a&��z9P�'7jF/V�\Б@�'SCf5C�'و)Ro�Q*F����5M��qC�'xPk �Ekh����2L� ���'M�$BBL�D��9!�,q|؁��'v��Y�"��:� ����ғY9�e
�'3Эp���P�Qɣi�(bR%z	�'�i*��)�p ����#S�M{�'G����	�
-ǀ��fIP72��'�6%�� /]��Ļ1�^\P��
�'X�+�O�nv�1���.�b�k
�'�M+��T�rB��)y� Hh
�'�t��+<���w�#o�t9
�'���!٭B�p�ƊaA����'9\0�B�� t^@`���/���	�'C�ZF��
� �É*���C�'����!�G�^���匘(�dz�'S�q�0mV�\=�𚁡C�i���
�'��zQ%� �B1����4��Ց�'��� Y-�,*p�ݷ){�q��' �M���,1Fb�����Yl��P�'���`�S�n0�!r�_�4p�' �����,D���h1k_+���s�'��;�dT���B,~�$��_�<�Q�5l��£I!K�`8Ƀj�Z�<�;2�n����1r�$���}�<�b��c���2�B޲/Be�Ј�T�<���5}h��P�̄i�^U�P�<� �	���=r�xy�2�;΂��"O�HQ��	�4�F�˜���+q"Oa���Ɣ����P[��!"O���D�^./���p�Ѭ8r��ʲ"O��i1�	1l~V,�l@� �@Iʱ"O84��"[��r8)���6&��sC"O�5P��kS�M��	��f
���"On)&'wQ�-�t鎞;�xI1"O�T��ό�t�����Sk�D`��"O�e����2HCHq��
H��"O|\a���u�Hx	�#�5LhZ���"OnE���SDc5��`�"ONX�Cu7�*S�B2@\���@"O@��b�T�oN��Q��L���S�"O����'Q	2�l=yR%_�5�fѻ�"O92�B�*��|��1�2�S"O<����^�&	6����s7"O� ����aEfKW�=L�BJ�"O|�H��V�i��N�*+��C"O��2�`�<�j�X�?$��@"O�q�%g�3���Z�^�4�C"O�i�˄�@^NA�l�7�<�[d"O���ףܧw����m�	:k<�@�"Oa��%3q FI�w�7`Z�pp"Or@`��"*��a�7��0j�� "O�p�-��$e� �;H���t"OL�r)�Y��K�W�
��A�"O���"ɜV������Q����"Oȹ ���$ENd�sgH�	��I�"O�@B`��iP���f�Җ��a"OV���@�L8�x���'%F%�"Ob,1׊�~Ū2�J�;�,`�"O0�j�oJ<�*��"�R��#"OҤ2p/�Q�<�j�
��}Ú�t"O������1�N�k��c"O`�@'�fZ��'(ϛ��1�f"O��A�\��'�
0q�>Y�"O��2v��M�г�W��%�"O��mC�/,���4FŮ)�&R4"O i��jT�%�n�!�����	F"O�,�'��/}�|8�
<�< xQ"O���3��'�����T>�&�1 "O���b閟<�^��	҅uy��""O�0�LL�v9ے��>+S,a��"O�,K��ɼ3��8�Wƀ|m2�Pa"O��۶�ؙL�ʨ��E�
gQ�|"�"O�%���
��� $K�2^���B"O�l�t,�C������9$�X�p"O��i���2��B���J1�	7"O8�s���tj���C���U$Ĉ[2"O\uB����^�:�He'rс�"O�u�BR�Ƶk�/u�nY��"O:�PC�/�����-I�b��d"Ox�J�䕥Y�h�ʧ��_Զ�Z�"O�rUGׇY���P�d�	�(� "O~��`#u�� ���E��`��"OT���BZN8v0���
���ч"O|̓�"��OE$<8�=B��{#"O8 �w'�Xf@��T��
8{>�@u"O~aƭ��3��I��Lbn�[�"OTq)R���Ī�.!�hS���y2a��C��A�K� �p��B!ޮ�y�kN���Jǎ���p=C���y"��Ki�5 d �'H	�t+�!�y
� �,�qb�/*\��a�ӥu��L�@"O�{��2�PH(�-S��)�!"O��9t�֍J� ��I
k�+�"OD���\�(	r&�
<v����"O\��U�p���9dnQ�vLp��"OLe��H R��d" D�)2"O�%���S�  �B�ɢ1R{�"O����Z KsY�a\�y��HC0"O��R�ӆH$N	rD�\���"OqA� ��X��IJ��[F"O~���I;�H�V�B�@�Q�"OHĸ��R
)mB��s�*F[v-c3"O,HrDD��J$�"G�L�%]~��5"O�-�%��a|�D��$]�sI���s"O�A���<Q�A�<~�̈��"O���uCO�xp�7#�,t�ZuCG"O��U�I�8]|���+S(rԵ�a"O�	
R�,r����b*��Rb�	`�"O8(��?;ZlI��.ih�+u"O]�cJ�!�\���-0P~ �B"O�,)�������tԨ3߶���"OD�����6/h.�H���R
�"O�CrO?]���J����)�"O�$��JK�d<r�
�n�VЃ0"Op��
i3�ye�J�=��5�C"O|���ۡ)�pyW�3�zA�2"O4�R�B_�0�1k#/`ٙt"O�q�BD �B	@$�H#@y�"O�����:k@ea� �^��Q"OP�����l
|��T&Vb�~�Bv"O`��D�#xbL8&ԉ i$���"O�A�B��b;DQ[�$I-)�>-"Oމb4bǴ�q�����rh�T"O���v��}�p��e U�z��hP"O�t��o֗\:Ve{�%��E�T��"OV�����%�B5���#A��a
"Ov ��'�.P�QE�!z���7"O��C����y�(@�\�c�K!�y��@����L�Glm�A��y�
�,t��0��ԙ@XD)��y��![�� ��/S^���2�yb*�'@�da�p�ծx�N�����$�y��/���8CL�q;��q���y� �w�0	3�~|ћ�O��y�n�<�, x���E-��X����yB��1s�最��:y�IZvđ�yb��1z�� �Ã����QF�� �yr!�4:~�� 2/N-b�0�&P��y�`� Xy53�
�#f���Ǥ�y��M�J�Nd��G��ncTdʀ����y�3
�^�j��\���+'� (�yB���1܂kt�( �@ٓ��]�y��9R<(�6A\�A{��ǡ��y"ѿ�@C׀�";[.t�6�,�y��/-..̛H $4�
�	����y"oو
����*�2��0@Vk�y"��l���!�.��<� P拟�y�撦o���pI��Z��ţM��y��n�X�rR�Vbf��c/�yb`�83jyI@"�;P���t+Ⱥ�y�mH�����JC p���*�yR�&8��d�Ż=�5�ǦK:�y��ф,��Ȉ�H	m�D��*��yRmS�{�.ӗ���16�p@��X�y
� ��-�kQ40R�ŲW��5SR"O�#�,+�5z��1g���a"OL�DI�Y�T.Zgf�Q "O�4��`2FE@�ᓒ&�v��S"O��%���:��j� � W�&�cq"OT0����SD���S�g:��w"O�P�a�+5�ླྀ��0Nn�ن"O�{�J-Tt���wn?>�NG"OBt`0��9��t�c-�4M� W��y��].�X���l��2�������y�����v�G6X�E�è�;�y��%���4���A��E`����yBiC6V�k���l�nI��BЪ�y��( �Tlx�l�o�>�Jg���y��_��E�A�>��ٚ'���y�쓣 �������HYҦ���y���-�\]���͵ ��b���y��H.K��ꆉ(���@d�R��yr��+�&���ڨ6/��k@����y���[(i	"I��5�0���J���yr��V�*e%D R2 �����y��J�P��'��ndtٚr���yR���x����250���l���y"�L�Z�B�@�.&��bWh߀�y�j�����6+�;%�J\[�Lǃ�y�FD�k�. *�@�{|P�$]��y�Jܮc��0z�AT&\�IS�ɔ�yRD�n �X��]����@�bق�y2'��R��5��;~�Ľ��a��y��J�ztb��]� |u.)zX��SG�a��:�`T�,A���ȓk>���k�N�P�Aℇgl�ȓM�T]�C��n�d\��Æ{$�A�ȓ|Ӯ���F
[����*��V�&��>OL�� ĜH>��U�Jq����I"�<z���Z :��p���O֐���v�P��B�L�X�X�Nŧe�<�ʓ{��a�ŭT�n�����B��e�^qc�` g\)�f�Xp��B�I�!u�ݙ¡
g���BZ(��B�� z��B#�M����
έ^�B�ɨ6q�E`g��O��R&�".�B��qs`�*`��9p7�tTI���RB�	
厸h!��KP
D%��(wEB�I�~t�A $�* ⮘�5G�!�D�g��1S���@��h�Nӛ=:!���z�r�"KLb��jB
4!��.xnKŮ}/$��,կLB�]��'� ���(�!8@0fJT�=��$��'<~,��V�z���Ń8�xݣ�'�����V���E��bKNi
�'��R�ʂ0-�u���M�Y��%�'��Z�F���b�n�/_`x��'���d�K�:���%__�����'P(DX�H88�x��� iFy�'01��Ә*�:�Nih��"�'7��C�ɲT�&4R�LT�hpV���'�xeC��1/�p-��N�U�f,�
�'����-��@S 9�r��M�B�
�'���� -̎a5�����)JlP
�'�xձ"��zj~�ra��xT`�A	�'ʦ��a�0�(\�0��u~��0	�'�X$ʷƝU��;�%�h��	�'�|�t��y��u��'S������ \�B�ŧd;T�sc�׷`	�!0"OBB�0��\��!T�c�As"O�s�� �H�(�:�Ə���y�"O��8�E�6gD�0����9�nP�"O�}��jL�2e��N8=BP�"O��Ԯ�~'�1"u��*r-D��"O�D!'E,{]jlC���E�b"On ڐg��F�<�qFK�5�2"O��A$E�s�0���&�|�D�S"O,���H֊-v6U�@%T���h�"O���6��- ���� BH��"O�!��X�
��@�f����-�s"Oh%�� �3Lq|li���#��i��"O(qp!�K"�ftc��Ж\����"O$h��C6�2|�!�Z3&�*D�B"OV}�֨ԅOJ��p$��q�x=Y�"O"�J�m��h��B�^�ҡC""O4u:��Vzt:���"ã&羹I�"O��g�l��%��F0ᾕAE"O BRQ�7n���d�Ⱥm �"O:l�+P�FL��M�v���"O�!��eY�BH��s��g"O��b�h�>UI�<A������"O�L�T)��[�� �!%����"O�Q�G�U	r�>Y���Iw�5��"O� �T�l�`��2w��K"O�w��-���ȃ�Am
�Z�"O:�s�*w���p�A�<g�Xa�"Ob	 �̿a:h!ˤ�Ð#_�	"O-j&�W3�ص��W� �g"O�Y�0����,QiT�w�r���"O&��ٗa���KӨ��l^��%"Op���Cֶ������8AM>=� "O����l>��$�.=\��a�"O^�ZDFD?"������cd�|� "O�\B�H\5FWb�3�,L�"v�P�"OrU;��%az`�F��c@3�'-�)r2�R�+��10���}z ���'����T���b��'�_�{�"(�'�H��A#gY��%i^%	@��
�':tE� j��Q�rء��	!J�%;
�'5,�S���OVF�3�G��6)`
�'7D�X�͔�a~���G�7v��
�'��f�7`� ��`�W�P�9	�'���{&�&nb�J3n�X�q*	�'���!�hD�?�(!��n�I��G�<Y!�Z�_�]#��a$̘9$\\�ȓ_L����B.\r�� ���1�ȓbYFɕouR1i�l����ȓ@h�i�e\�bE�a-�X�8��aR��a�*4��� !�֍;l������-�ࣕ>WP��ƄK�5��Q��t*�`&���]հ�zd��Eq��ȓn� �S n^%J�ώa����/ a�ݢEi�I�p)�ZP�L�ȓӠ� 㒘1�Ha�bD�A����YA�Mܹ�PMc�TØ@�ȓB�b��&B�]e�m�!��p�n���y�`�q0��jG�-@i]��Ԉ�����b3�K$p�>�{���d80��%���x��'b�R��EYN^Y��,�fٲ@ӡb셣��<)�Ň�۰I�h	�g��q˶���sBp��'��Bc��!<��2̕T�xT��S�? 6-Qt
U�e��t�@��p��"O�d�@FT>]�U�aj
�4|�"O]����N}���4,�3=�j(x�':�+S5|�ڜ�,պe���	�'o��ӌZ/Y��L���%�$8	�'�=���&�*����	�� 	�'Ϥ�$)��^��4t�2���C�'��P鄠ܪB@��g@�j炙��'�m���N"���Ë �wo��'�D�RD#kT��
�@?uG���'�Fr�H/v�}rP'� kr,͓�')���cNY7Vdt���mb6��
�'l������7�.(J7㕉i&(��
�''�a�HC���	�qdӀ`��T��'��yH��O�5�Iafް\{����'%�d1#O�3Y����-Q�z�Q�'"P!L�ID4��J:�n��'�n8�w���u_�q�  R� �|[�'�"�;����-�`���پ=r���'����0HŃ
�TQ8�n��qy���' ��+��Ȯ�8�e�,g~l:�'<�����.S�"iFD	�v��k	�'e05���?c{��{%n�Dʉ��'�\��F l�,I%��>"8��'~�x�ud�7WQ��\<1��0A�'q���낗�$�SB��!!?��8�'�j)�%T�Y����8Ep����'D�}q2+H8{'t��T��P�#�'%�}�"�yH�Q�.���A��'-~E����0ǀ%*�a�N�A�'�� bg�ҲR��1��n3>v衃�'	�mCT�7mളTfc� �'=6�q��˿2���IE!Z-�l��'@y
����q�J@5:�>��'k����,�G�pq�O?+c2�y	�'غ$�mT:��U邨�1�bU��'�`:��YHFH��㝢+�Vt
�'wN�`1��p��p�F)Myv�{�'DQ���2
}���H�?8X��'%�,b2$]��>��Β�4��`��'�^a�@0N�(�d)+��г�''~щW��(,h�҉<�����'��,�P���<����9[�PH	�' �sୌ'D�1�7R��<p�'	��be�͗w�������IA�e3�':L����0rg�- v�Q���	�',9�1#��3�U����2Ng^�
�'�|�x�+W�B��M����<@`$�Z�'W}�tŜ��ڹ𴪘�*~�c�'�N���j)l�@��E5+:.Ւ�'ަ�
g��z��)�q�,W6L)!�'��i����2h�+��˫Q� M��'���0���3 ������2_p�'�䳐'�%$�`�w�\�zBē
�'� �82 �C��#�բqV>91
�'}xQ34
������d�����'����� J�ȶ�ǩ\��qx�'�|L�d	/<s�(���̕���k�'�N�p�V4N�@I(r @+�����'�TൈD	P�عБ�@��z��'��ٱ���8�Rm���VR���'�Aq�Rt�d��(��t�Y�'v, ��MZ-4�,�QA>ԾQi�'�D��-����@T��s���S��� ����E
}��h3(8~&��"Or��NGo��t)��R5#m�"O��0�ղ�)����RR �I�"O��jV�ε T�õ)�B;�,��"Oܽ+s�@e3zȻA>
@�,s�"OV���\  �:L�᫈8+2���"O�@�d�9aL$���W4B���"O��`e
��O��%Bta�"(�d��"O^�y!L��2�P��@ \�B/�8j�"O
�kp�����b�쏌;0�"O�4X��_c�ˤ�8#	r	�"O��y �Qn*�,�Α4&���١"O��+c�;6�1i���p�p��"O*��W��
�ִ�V(�	$?.\c�"O�����+�^�W��5	�lw"O��P�iֻC�����5B���t"O��y�N	4��2���
��"O�b�l�Td:�`G��3Pl����"O�y��&#���
6�>r@�p"O(0����@pZ�K2i�!��X9�"OR�K��W�NL������ւQ*%"Oa$�Y>~�z��f5�$�v"O�(ą��x��dZ�W�W�p��"O�,��L05  H!�1H�� �"Onm���^�1z�l�r�wS��Q"O��B>ErLY�j��cL8���"O"DZ�D Y`<iъ�E䄨�4"O>�BťL�B��-Ê�Z=� �"O����'ؾ�\I���N�R:��3"O*X9�����h�%�5y�a�u�<��腲:�s
�!`�ج��Mt�<�c��0��<���H>�NA@G�y�<���Y+S�ػ7gӘ"��h�@�<!&
K��������~�$�;b.|�<�W%<q�@���A�z��Gz�<����Ml�SƄx���V�NK�<ie Dh8�Fƈ�h����Ş^�<�Ԏ��`z��*M ����[v�<oN�X��&�*�|l��
�t�<��b�s˔q��٥����Qm�<��f22C�`�[�����qj�<�7O�
4�`����+���ТJe�<yPEŀR1
8�@�0��#Dc�<A�)R/[?q�`�0�Qm�h�
���07bY9��Z@I�cR9r��X��F�z���F���M��j�9!E¬�ȓ�Z���T/�XQ�+�4]_���e3t��I5M� R��:Uxr���W���A�:E�6�¯��d��{,�ܣ��D�!f�p��]�m7�U��,��$y0@�@P�CmX�(��ȓeDѳ0/×����aC4z��ȓa&z�f柟57��c`��8�n���n�v) �+^%XO:�#e�.y ��ȓ*s�z&n�cFT�K��;D�ȓ+�hcPk�QD�Ѩt�Z'q~���ȓe�ʼ(��6@�~!��h�}�I�ȓe�le1e ^�\�$�]%n�T�ȓe�\�+S^��i���X%��Iŀb`mK4\*l��#_�>��@��Z�~H�����|8�Xq��Rh��ȓfy�1����Z��D@��ËI#$�����p�6�؋t��}�4��ȓ7XT ����� P��	E�_� y��S�? z�Q�k�u�x�c�o7O<��"OT��d��_0�("��ȑ~#�x�G"Ov��l@43܈u0嫐�+Bm�e"OT�{��0%]�E�&�>\;�"O0��
�.@�@h��UAR"O���GD(�|QS�H�Wۈ�8"O )��AŏR�p�3- �f�h3"O�t��_�mcL�@2B	�%��	�"O"lQ�F�&�l��F��b�  "OV��Vǈ�	��c�f���"O�ab�!N�a��c�)�R�(�"O������(�cq��uf9[�"O4���EGq�&iE�JpL)Q�"O�d�7m�&s-�ڶD�$_8D�"O�u��`� R`ĸb0��*~�E��"Oz�(d�Э)ט]�A6=Z��r"O�3b�;H�zX �E�U	�"OB�����*,Z�cãW,e�Rf"O.0�5.�_�xI�C�73i�b�"O�͓d�H+q���c���7���f"O��B���$gP�k�R+R倔� "O�4q�d��S�|��F��y��"O��
�Or8%���A�%�2H��"O�	:"��-;j�s�*� w��X��"O"`��˄��䠳��W�x��"O5�Sk�1�����H��D]Ƥ�f"O& �a"̄]P0K 	��#A\��u"O��R>g^�P�֪��:Uh��À	X�<����K�p�rp��9v�zX��dM�<��oI�[�V@dM�[�'��H�<�4LI�?��\J��MGh�C$hC�<��сU��M�T��aX���[E�<yᜀh�sW-רl����� E�<�QL��z�lPc���C��=��@A�<i5	��X	�yVte��cR�<��狌$F�PA� !Y t5�K�<� ��z�V����>}�@!J�<yPϕ]�Fa{BA�~�v9K%�Q�<A���7SF�1�Ě�	Č KЋQM�<�E�;^Q�����hksn�G�<�ˇ?J8�t�4��rHr�ۄ�M�<Yb _� 4�JP�ن/��i�2��_�<��&F'g<
�����?ږ��ŋ\�<��ԫ�҉0��^=.52A��W�<�p�5'�F0cGl�_����E$�~�<AǊJ�[4�yCR��>��Xa�gR�<饩��a�m2�:F`�5��k�G�<�+�'J��`l����h�"�x�<�c�n�C͍�?ڄT�E��s�<a��	�l����-6U�ى֦Cs�<���L�%��%�7�ϦRܩa��p�<)�$S�d��mqӍǼ��p�uEC�<A�iW%K��)�j^;"�V�MV�<�BK˅N���E�[ ���(�U�<y�C3i����
�"eQ&k�<9�O��8����)��p����h�<�B�@C��4�vF*r�n5��Wa�<if����9���U��+woV^�<��<�$��4�G�:K�{  
E�<i$�D �t{�K����6�C�<E ���� C@�e���{�<��p:�\����XG ���Bs�<��*��r�vࢧ�\%�f�2Di�o�<�� �q�N���왌ں�TBUm�<� p��PCA�&l�= 4��{a~8�r"O�h`2�N�
"����PK� T"O�X���';Ze s�܋I���D"OH,��`)|D��U�B�`/��4"O��v�^���E�^�*$&9	u"O.� 2!� ����Q�n�HJv"O�ʐ��h�z��4ˀ)>��a�V"O~Yz�	 ,����~��(`�"O�� �j�4vɊ�Cޤvኄ�@"OBH����2*FDC'��	2�l��"O�Q��|��I���?Ɗm��"O�	��dɉdY^�@�
��0Ī���"O�=��($����8�:M
 "OH�f3_}�
�c����)�"Oāʔa�h�j���B��[��| �"O�Yz��[m��>}�:��"O�8�JĨv"~ta�'�&Y�~̊F"O��0�}Ԁ� t��J��� �"O%HFO_�u�����}5T�I�"OF�#s�� 
���Ԋ�F�dPy�"Op[QF�mlAX���-��""O@�!j���)�c�$�V�X�"OI��S�'3�Рr5g٬�!4"O��T���*���!�Ȱyj�C�"O@[၁�R�!�����F:�5�#"O�	�5��K��UXR�a#z�:�"O,��3A��6�8H�p��,*�5�"O���ʿQ!�Kp�� r�"OxH`'ē�y���L0G�-�t"O`;�L�^��C�k��t�Fp
r"O$ɠ��v���W����Ar3"O�٘@nǿh��H����|F�@"Oz��R끆4t�08�h�/xT�	�"O�U���^�-F�x+�_�s[��j�"O�9@ҨD�q��q5���ܬ��"OZN�*8��h�E�=A��Ĉ�"O��kDjf����ƽ)�2�i�"O��>dR�P`gޘ@��e@�"O��W��6���Y�㎿�LLA"O�a����M�2 ���8��(��"O�$���U(gl���q��)xd�&"O��h�I_�}?��1�3w��"e"O(q"w���L��5�A� [�buɷ"O��@�߰xGT@H�EB j:�(3"O�4·����/��9�	�
�y�IH�hy
P�A
��de�Q���yB"�G ��C�ωJ�u�!C�	�yb���!!��XbG��8���8�"5�yR�����p�A�^����pBҶ�y���wyv|�#�i�$�������yBG�5���+&I�#hľ� $>�y�w&"&�S�^�v�� ��y���|��@�C�4U��)`�Z��y�������c�٩P���g�C�y�$�F�88S'ƺIS҉�'LG��y�J�&� hC��=PY8�%�y���2-䌽�j%=�z��#,Ï�y�T�=�>�x����F����
�yb�N�Ib�8�ÈC/���ç/Ǉ�y$�5��� S�?>����`��y"j� ٘�� $���g��y�!�#��ϔ����ቄ�y�EN��� �[����Β�y�AE��Ճ�A�whx�{d5�y
� d9#��� e�;#͂%`{^��S"Op��A��7(�C�G�bhҀ�A"O^mu	>8�I�1jDYX�l	q"O^I�H�(7�Uk􈜸f��uQ�"O��ڇ��W���Y��S�d�j�0U"O���(�q:
%�c�H�7�z9��"O�A�U�gԄ%�'Č,J�΅�"O��� K'cr�Xj!cA�bŜ Z�"Od�Hd�Z�Y�>9�Eg� %Hf:"O\1�k��c�n9H�o��"1�(�"Or�����o��k����8��`V"O�i7�7^��iӍPLH��4"O����(Rz<j9ڂ��=�<�"O:�٥�!� |��֗M�+mHJ�<�B��/Fdp��ET�?K�f�F�<q�a��VW8A�k��N�F���E~�<�ӏ�9lH5���F�hu��{�m�z�<!1b�p߂��KM��PX3 ͑t�<�LV6�"u���Q�0���Oq�<ѐ���(苐mN�eU��� �FX�<���[a�H��ldB\Ie�L�<�ף]03���9d�ٽ#%L�7oBa�<9�Ɯ�Nt�Q�*�QR�Z�<iB�P%mRz�343eڴu��a�S�<!p��<c8��soF�'���_7!��W? -���I�O�J��KԼ+!�D }��A��AD�9�ĉCD�=K�!�Ć�72<)2��;K���Z� !��١H�($�d�P�f�\�!���!��
�AȆ��u�ȅ_�>��$�7<!��XN�h�#�U=	�FH�'A�;4!�d�8hL�<*5��!Q��ШբR�Z!���l���G�4��<!��U�}�!�D Z�Ҥt� X�X��ar�!�$J!pўU0� sl �ᓁ�U�!�D���D
�ś"f��x�%�c�!���	Wʍ��n͔`����qN|!��i&޴�r^(?����GG�)d!�$ъX��mcQB�-Py~�8f�j�!�DR�4�p���O&<T��Pg_tY!�S*%J����X�pL��q�޻�!��M8����6D�c���%�!��-MN�ٳMQ�<J!(��G&!}!��61l$J!C�/
U��٪5n!��\�(��U �7N����K��:@!�*H�����L�$� �0�ݠZ3!�ۛ?5�� @%^�f����6�3b!�DV�{�A� �$������<�!�*8���:���%�@Y��"W)l�!��f�ph���ܝtP�,`U2Y�!�D���0�Y�΃� N2��t�-=�!��H�J�H�9ŏ3Rg�%��X&0|!���h�4�dD�/,E��M��!�d��iX>��M4_��9)�K�5~�!��P�BZ\��@J� �JU*�J*!�$�|K�8���&7��1)��v'!�D�-o�K��_�|9�	��!�D�2���#m{65�E��!��՚���d<v(�ʐ�Ɲf�!�[8�rɛ0���fr`��W=K!�$	4n'��� ₑ,S(,	�͓��Pyr�ڿ\���Y
u\�H"�B��y���}_���J�_Lf=*c��y���_��UYP�[�T!�8� �y
� �K�
L����3��	�Sa$�c"O�e"qӌ.�����;HzL8"O��b�Kɱhp��®Ҵ��"O� ��.Pl��R�H,�n}�s"O�)d. �nA��"-yz%�"O�U!@�2����F�Y: p�s"O�h��C�A�E���q���B�"Oxh�BG�`ъ�b"ЁJZ�m۔"O��V�5F�l%�u �d?֤q�"O��E@̷xܴ[W`��9.48�"Ortڄ%�h!X�Y�MŰ}I8��"Od�	Dߊ)���0��2͋�
�y�16{��4Ve�(#��\+�yr���Z|DR�'ۤVP��p $��y��Z�n��q��__x�b f׃�y��V�*�~pC��PR�y'Δ��y��K�x,Re��W0O^�0�N�9�yb�B6O���JVD'L�U���?�yr#	w���`B�>$��w@��y�F�m4��"��%��%z��Д�y�H#9���������Y�+o�<	c�C��{u�.���v/�u�<�R ��FF�9��jӋB����r�<a�B߹SAN=����	wԔ9�a�T�<� *ħG`���TCۉ.C�Y���Q�<�ҦP:�hU҈ʅ}���0@�B�<qf�[&b�l���R/V��3&d�<��`��l4t���  �}��a�<Yv���.��0B3�_��]`AΆ[�<y$�ʤ[0jU%Ș�<m$a�s��N�<��?zAt�iՋs��=A%�ZV�<A�JB�[i�|�ɊfY:��W�Ml�<����-Vnh��� �p0���.�P�<Ȅ29��� ?=��@`��R�<��#J�t�����Rgr�p�Z�<�!RD��d��E����BAU�<���(Y�a�f�Di��d�NN�<�$��I3�!{�K�|�����#�L�<Y��'/��%������q�ir�<��"��C�6Mc��
#RfP�	�.d�<���_0�2�a�ۢ[T�R��Z�<���_�lRD�~N4���_�<q����d��+�b&xД�[�<�Ab�	����l�i�t��X�<����^�9u�
	�EFHL�<I���;f�ʥ� �D0tY04�b�<��Zu��|8���7�DI���@F�<1��O,������5�R�
�BB�<	���b�`��$��H�W#!��0��c@|�ƹ��l�4!��"�6hi�`��[��Iw��Z�!��,&�
�� \-c㾥	�ܓ1g!�[�
H~�ؑD��ލ8�Ø�6R!�$�e�(����n�T=�%*.�!���1�9H�&U-0��@���!���Ԣ�j"$�U����+�!�P�_ي�駯��i8�ǁ�$�!���x�б*�H�|�7�<	�!��ծ"���£B�1zA��Ѫ2�!�DOrc���+7Vd !I�=z!�䍽$8�x�e|�`�(��b]!�$��:ͦ�2A����H���x`!��ϩ��5ՏT�F�|��F
�@C!�ĉ�9{p��e�,N2�Ҥ݀eP!�� �07II�b8B��K�HG����"O�a�w�E!9nb�c��D@�9c"O|�zb���I)$�A�iZ�G���"O\,(�l��4Q]6'ɹV��Mh�"O��p5��al,�D�
���"Or��*϶� Mc!�ޚq��""O !��K6�t�!�*�ni�#"O�sw(t~<����>,�HI`W"O�����SJC��U�E�#��*�!��!
��l�ǆ1��R�K�a�!�$�9D�f��u�ܙxhD��Ì�?�!�Ą_�Hm)�Ւe��,zR�`�C�ɥ-�T���FS ? �� �ıZH�B�	Z}`�p!LR(	���5��ȓg����Sʄ.a�v�s ȶ �j��ȓrI���%�P�
��·1�]�ȓz?�]"Bh	��( Y�	D��]����� go��r[HLA�͔H��C��Z��x�b�-R�zY���U;I&�C�	$rx���$��[n�HgR2F;*C�>5���1v �./:=�TIk�C�	>MB<��3�d�:��;��C�ɭ4p��DgѦ;�Pi���J[�C�ɏРY���r�lhV�/7�C䉅{��C���e@��Lܹc�<B�	l~����5}Ĩ�v��0*B�Isɐ`"S��6i��j���M��C䉖 % qj�!��Mbjxc�F�Z��C�ɳ Z��k�3y��ʖ�-�XB䉛kPTXi��� (��{0�I�wt<B�� h�&��g��T���ٖ��$�B�	�?�:�gߏ��Y{�ΛT��C�I$1���p��Ĕ�8�W��9�C�	����6��w[����]$$��C�	#\�$Pp@�ԖK�֨�vB��
Q�C��)�>�D ������Òuw�C�I�p�d �L�j�,  ��=�vC䉙 �81CQ$�� ��|TIк(�fC�	�>L��j�l�!U��PpL��H�XC�9*���;UJ_�:��S5��6C��	$��#�k�+��I�pA��:C�I�*Z$#RFB4޽��I�E�FC��i����	"Q�a�5oħO��C��z���-T/&�|yy��ߑ9�C�I:(p^�K7�O�y8����͞�{<C�ɴ����H�;87nP C��.|�B�I�E^�a�F��+&��!vۣ/�B�I�0�4��HJ����I�U�B�I�>���ի	�}(��E͞E�B�X|@0�/�}Sh�E��� �B�I*4s�-� �L�g��@�g��b�C䉟W�Dl�N�F�u�§{�a��<�N����Q�i~Ġ��'̺`�ć�H�|�b��(����I>��фȓW:��m[�X!ր�ѡ�:;��ȓ)���#m̢~��1��CV9s��ȓ`P�"0.��jʺ�Q$�3~�L]��Em�ѳ�O�dƨ�1�J���(�ȓ:?�Mǂó~Q�#6�����ȓ_Rp��v/;>j4��6�R6�I��b����� P('Tr�SQ�"��"��mr��� C.�#����\=Dp�ȓi(|�����.WY0lr� )�fхȓbȶ1�FDů"~ |Z7�L���S�? B��DHΧ[���hL
zgvH�"O�� 4E�
�9Ƨ��	e���"O.d�6D�D
.�
��>YmP�"O����8�p���/�+����"O�؛ѭ��!�zA�`�HXn��6"O����.�4jN��E���̙t"O|�� �z\�CFM4�y��"OR3����\�uҢ�6(��:@"O���4{e)1��ӯ[�,���y��L9a��i�m���@з�_�y¯�,K��@�ggH�J�|Y:&���y2E΅}�F`It�E�����-�9�y��I:��pHam��FBtk���yE�t�u!D_�g�ae.E��y��:x �ꂇ7�dH�풾�y�ŏ;���� ">c���.ů�yR��-�XE��18ன����y�؂NX�����^$@�V�Ϫ�y��X�Uf�F#����a���y��5%���ZGd�YT�Һ�yR�[~ �X�V͆B�Pۓ���yBO7Q��ABbE�m������yR��6Z�8�pk@�:|d���^��yB&KA���s۵`s�D ��<�y�	5.m2��)�(\��L�����yBCB<[�4��)+T���� ���yr�Ąpz(�D�5����o��yB�م%@v�hs��:x�͘Ѐ��yr[��A���83�t�ke�y�'G(�X�:=�	z�ԋ�y�K�8P͡�Q�6�4T���͝�y2��ud�j�.���`Tŏ%�yb'����5��*���p�J�y2L%�rh��E��,F���M.�y��.D!�=V��2����⌽�y޿O7&�cpā'$H&<S㭈��yR �i��)����s���U \�y�.D�A�&� ��q~4��e�C�y�"��=������v�μ
֧F��yrBQ�L�:B#��<�Dx�0���y҄�6��2A�L}/U���T��y"�Y�]�B����R�s�`���ʖ�y��F/~9f�G�P&;��������y�S_�|��P� �0�<�Q#�Q��yRς;W�=speW�0�������yr�P�F�8`f��謽�̚+�ybÇ�<�Q �����cGF��y���>��Y�O/m/��M��y� ���5�n!S@�*���'l�]pTn&+�LD@���7*�� b�'��7ܴg����$����`�'jL�:PO�g
�كK( ��ɻ
�'�ma"gS�V��2�!�� ^���
�'h����-J%8�jS�aυrƮ�I�'���B�H�=-��t�'L�:&zD�'z��S��ݜi����L�,����	�'w���H�nx%8tƒ�^�Ŋ	�'*$���M-�X�)ċ�DW�x
�'㨽��K	�9�P%ð��:İH�	�'$�RĤ�2WBDm�tJO<1z��R	�'gr3�n�R��ur#��-��9��'�TUb�*��5�̙�#�Y	 ��	�'���X�䋼i^��;���a�ƈi�'ۤY���J/S��H���`�z4i��� lL�և͸�҅�Aʁ@�@� "O ف�͸A��1fȑ)�|��R"O6�`�$�*m��Qȗ�Y�4�B"O���Yo`���V�8̝17"O>�q�D�Bz�Q3G�:3��iF"O,����%0���aw�4B�p�C�"O
������1{PF��`T�5R�"O�A�3/^�(Ő�kf߼ e���E"OP�C�勯UI�8𠄗�W�� �"O�H+�Ո`>zMPC6UM���"Or�P��i����b�3k�P�"OZd����/�� �c�3t��p�"O*��riF�s)�9�e#P8`\�Cp"O=(&j����{%�7��A�"O�E�B��4�����"׫Dp6D3"OF�D��*D��o�w��As"O�h��� ^J0]��<0��t��"O����޳X�Bh[QN�#k��Ec�"O�3 U�wG�UK�.@�>���"O��k�$��~��0���"� �y��S#*�~ �Ս�g�x��5C�(�y�̛�M��+��FYC�Lj$+�7�y→�6�mi��\YF��H��y�Ε�*�a�Re�1_�l�Q��yg��GnZ<�׮T1|/X@W�y�i6:���S���&oRV��0���y��P3f����G��h/�%����y�C�(�*l��݄^�Tp)!˞��y2��	��:���>,4H�Q��R��y"k<L6e��m�Xߎ��7o��y�K0������!{=M�'+	�y��/_��2���	w��!At���y,��.?�$X���v� ԣ�KO�y"�@
f�n89��C6bÜK�	���y2eW(u�䈛�C�3$X4m� G���y�e�0���"k��ܽ����yrMLc�p��V3���ta��y�D�f`����"��*�h����y�l�y��!����;j��eXJ�y���
7�t��`Ǚ_�f��a Ч�y�@F�@��Qk��F2rt��y��	���h£�>>�(4�F��y���Q8\����ث(�Ѱ�&��y"��3YiPf�)X��8q�E���y��H�4[HQ�r9Ǚ)�yB�^�"�� �j� Br���Iՠ�yR �9^��L��W&=��h/���y��)�� P�NC�
.�p�3���y�3 "�}0v� �rܦd:B�$�y�*�&Up��->	���A�Ձ�y"�Vڼ��<3@����_;�y��KC����-�4b�l(fc��yr"V�e�¢��)^�U�U����y���C͊�h��S�8���Q��y�M�?{�1&�X�J��i��G+�y��2v�,���6J�29�Á��y
ά`�$%ڑ昱Aq��b��_ �y�����D��@�??�֘�RmR��y��|x��Ig�M 8��`0�"���y�Ȣ^�����!ɟx���'���yRn�e�\�a@�m�#�H���y��^�]L�4
BE-^0�s���6�y�%�6*t��$$�V��<�Z��y"E^�
�R�!4��
����y
� ^�j2Iރ����똅
�XU��"O-�i��^{��q�j�w�n�"OeyRH���Ĥsc
��"ÎmR�"O�����F10���cT٦"O6�Br�ŮiNr��en_1mT\�b!"O@L�`#Ļe^����K��"O�(A//@�`����8.����"O&���ßj�Ƒ���֭~�x�+�"O!���Ȯ4��hRD �fd��"OBD�ub^;bo���B�F0�ݑ�"O� ����n9�u��-�"|@�"O��)G��Vt6l�ˑ?�.���"O�8�x���K�B�`UI�"�p�!�$�d��#&�8v���x(�?<�!�DR��\�*�͕"&r��D"%!��ʷ\�b	&�t4dx�@��v	!��ӵN�`YӢ�-1�Hq��U!���=�²G�.,I ��#!�$$4������Y"Ih��R�&!�� '�d��]�H6�X���f�!�,�. !M�1Q�ޘ�&㞳V�!��J=,Lt��s���4�L��$�\9R�!��D�0DB]1k�5��pTC���!�O  �&PC�%SL���9 ��E!�$:	"PXu�
�_�f�����0&!�� ;޺�@R%צib6�Y�FѼ2q!�Dôc���P�79��Z�E�w!򄉉6���Z4��@J.�15�@'Mc!�d�R�|��A�Å c�	���-7]!��0V*p�Z�i�1(W�t����6�!��إ{�����Wd�8\S�A�*pk!�d\ m�X��@��l��A��a��]!�D�w5���ᮄ")o�p�����RE!�d�
bT e�����s�.�n�!��͓E���F�R�%�^x��mO=�!�߉��1�Х�9ڬm��-��^�!���z����a�=Mp ��&K��!��>5¼X�V�6�"8S�F m9!�$��X��ؚ�K{J�h�$�7S*!�ċ	t���3g�Y�F���CD�4!��ȃSl0��I���1Hw#ݑ5�!�d�"ef���I�r]
��YK�!�D���T�����*g�Eke�Ӳ3�!��]�T�nC�ߑ)O�	���G�O�!򄙗c�9��I���ұ|�!�H+��[7(�h��;���",�!�$L~q���B�@�B�R��]�!��@)[P!����^�8l��+��Py���w� 4�7e\�N�6չ�bN$��O�#~BR���ѱ�Z�/	hy����R�<QTΗ�C=2���Ůn�MbE�Q�<9��	�j~NE���&�vM�A�O�<�6�J�D�`YGY+W�hQ��S�<��IK	8~��f�7�2"
�U�<AB��N����/š%�n�{�/��<!N<��O�O��I��9��
�^����,��X��B�ɋ-�N�K5�uH>���ͪp�$�� ᎝3����.=�-�Iۗ^
��V�ȹ�r/í �0���:�^D��L��|�S!�Aa������ܘ�<��4���$<j��_��9��W��z��ȓC
��YTFB�;mz�Z�dSW[��D}b�'>�>���-.!��T� )ֺ�K`c%D�@��[2��ɒ�.���b��M}��)�g�? ������S!��%#�!Z��P4�'B��YU�F0~��8ʃŞ�n���I�A;D��8d#�W��B	�#�n�Ha�%D�<ٰ?i� �Ca��>N\��&D��84$�"Xޞ<#)y���à�?D� %��*#gj9󃙩r Ε`�#�O��b�D<�C���!�fk�� h�̈́ȓd6�I����29��C&N�����8}Z��/kO�4�wm\ L���
�{�c
�"q�0`ؓk䞱��=	h!��޲��aK�m�tf ����?�h��d�FXRP�H�}\:u�uOP^�<	�D�_^��p�n��v��q�*YZ�<q���Zn�u�d ^!Xc�l�<�A%ˊB�H�P�*R�l��]�!�g�<i�B?�zm�D��;_�-C�,b�<A�L�**�
	��`vuA��-�`�<qv#_'OED����v��C]�<��b-<������}��p���M�<A�S�O�r��	UV��h���O�<��`L"���h�<<�RE��$WFy��'��X�e�ɆL��t�q�iA��@�'Q��:�'�u0D���W&bބ���'f����	H�JȣP@Jb�.I	�'��Q��߀0��d1���"愹	�',,�'�9�����N�P�}
�',���u��G줻��,�JP`�'�$X1��	�
�I�󅐿҄ٲ�'�1�b��`р�RlD�/p���'8 z��D/�r�P�̋��N,��'
�=�@c׫D^�A�%؎�vQ��{��)����|D@Ytƞ�X�c�͏j�!�0dg���g-�b�4e�לQn!򤃖n�� ��8�
̒�&cP!�d�;Oz�$���+tҤI�u$�.E�IC��l��߁5�d��pf��a-��K,D�16�+ZY
�[��P#�v��2*D� �%�O,�t<"E�,kVDс�:D�@P��8S���
�"�J
Π�u�3D��Q$A$v��,�փҤsAXI�*>�r���O�f���^3)��e�$Gϟ� ��'��<�c�ão&�ؠė�c��ta�'�� �G���c�ǎ�Tf ��'��
5 Y�w�Ba`	ٓ l�+	�'j��p�c	�}8�'Is���(O �=����'SveAu"H�/3|(2w����x�'�##cQ�y��AC��<N/����'U�f�<\�0 ���C�Q��[	�'{^��u�ޑl�<� ��ԥ �(�Z�{B�'g�\�EC�4.�lC��~�����������5�vp�t���4(���M+�'j��Q�F?&���e��cs������x�Oxx�O:ix��Ͻ*��Y���� �8�u"O��#w����ҐaS�Ō?|҄�R�>I�'-��c�O�t]�ЮF� Ѩgc�7~Y����S͔-��
P�^�ZAه�X1GV(�ȓ��\bRK\'X�z-�f���ȓ. �����?�R%Iu	�e�ȓ$�8P2䛙l��q�b_�.�ȓ��Mh�"� VĴ@t��I,��I��}�vd	Lؾ z'ˎb%���ȓd�0�3Ə��Y/Q
B�M?��q�ȓ<{�m(#��Ox䑈p���#��q�ȓz�BM�c���4����L��R�Ex2f5�S�� �0��f�v�Z�	�R����"O�KG�#
mN�Qu��>��4�,�������h��2ra5���&��)p B�I+Lj����j溠y�$C%FS��D4�HQ�ڬl��L4z�|#�8D�X��iH.Bs��JA@��K<��E�7D�X�����h�ˆd��D�;� +D��S헇%dH��qErD$́�H+D�P�p�m6i��'o$U qN6D�LQ�È*{�ۀriH�9���g�<�ү�'L��[�h�i�ͭ�hO?��"$&�8�EX
K����g�_[C�IMǶ�m�<!R,���WLB�B�I`"�d���
!Na�j֩,�f�$��"|zgǹq��X@��)M�2m"�/A�<�t�\���ʥd�=mG,Aj'Gr�I%m'a{��-v �պ�h�2#t �JN�ybi��e��5�	E�0!�B[/�y�4'���Fˍ����%L��x�!��゙���nqH�Y� ��!�T�/��DK�-RT��� ]\�!�DΩpIp�Yuo]'�ܪ���~|!��H
$XJ ����'@?bi�vI�!pra}�>�bJS�yV�P ��{�:��UQ�<)o�(g ,2V��#���b%Wx�<��L�$Q�`�����cd����DP�<�#	�62{��A N[��x	�@r�<��&
H��P	 À gA���àCn�<����$*�̨a��w����f�<��i�.ܒ�hF�T7wޭ	���,G{��I��l*$� ��=zTG�OfP�B��\�����N�?	�4���̇kC��Faa}��O�w�l����^�}���%��0?I)Oxt�� ?&�
��	1�8�Z�"ON�с\%+ j��\?-�(�b�"ODuqE͛h{V�jDU,d�!��"O����qmZ��્&�6@�"OH��5��0P�@x�����m��"O(}1����!n�]��^'��Y��"Ol�B`��}���Xψ�[���d"O�����٦]z��z2���$�ȈH "O8���B�,U��`W����B�"O�S6��&���A"����L��"OjH��툏nk`�Kį	���4+�"O�%�f�C�r���AS-I�U�R�b"Oh	i7E����K�'0�Z�R�"O�qP+� +-�D��)��~��8��"O4i����>+�� !@HR	iRqY�"O���J��\��U�F��x*���"O����ƶYa���6��(T��K�"O���]�* ���_��h ��"OVM�,����}Q�O$m��	��"O�Myd(� �"���"ʹ���"O*��@��HjX(�Y���(�f"Oꭑ3FS�p8��`�=�z�q"O��2&��{���3E���9�C"O��RgŇr�f3%�7��0"O6�#3�ŝ+��%@��C8*��y9"O��r�F�{��A1�E;i)p���"O~`��ǘ^v�us��8Y
v �"OĨt��y!�I#���42��W"OL`��P�r��dB�dùf떤jG"O`	��߃Ox�IҦc@8E�\Q�"O؂�h����1E�K"O� Ҥ#�ɋ$6���&�{M�hZ�"O�,Yf�E�6�gږG���"O���D��0= ���U�6�H�"O:	[�-�D���2��1&l��V"O�T9+4<y;Gb�.MRQ)T"O$��#LѬD�lYŊG$y���Qp"O�c�+ңW "}��dA�R僗"O�h�Q嘩=I0qSj�2q����*O� [�N�q5H�T�+�,���'�l�0���*�V�h�GC�?	H��	�'	DIQ �Ξnͺbt�6yl�R	�'wȽ#%��#�4���!3p��'�r�U�:L�����X�ݩ�'|"�Y%�Z1;��}��*��$�L�;ӓe��e��i�ԡ��)z%T��7 �%�"ERЫR*
�܇ȓG_�����^�T.B��է�����ȓX�h�v�I����j	L"��ȓ?qh,�`'��Pg֠Q7@���,���M_�`�C�G+��(�K

}�,��ȓ�����K�/**%B��_ ��"O��(�����2 H% V���ybC2�>xt��^�2��-�yR!�00���5 @�S��(�����y2�b��Z$�����1�'���yҦ	Pz�x��X��I�
�y�Y�Q��}R�	[�w2�(G-�y"�S�AM��� k�p�Iq�N5�y�&�nژ�C�͔{p������y®;*DHً !�~$�lڶ�
+�y�;<Lܘɳ������6c��y��O6\� uJ�+n�%�Vʛ9�yr)`%N�qF�	�l�ʌ��y��;mx�,C �ǈ_�P�!���y�OR����)1f��{��9���y���UD0`/O,}���"�� �y��P�,��0��r��J˹�yR�/pg�� b$�]�$؀cM��y�@�a0���A��]��t�R���y�JĤ?c
�2�W	������y"Ѧ}��bS�@.p�J�Z����y���PBA��$�6��B���y��1A�������6��c��yb��q�`(�V;Oe��Щ	1�y2�^�?ܐ��ꟆG���G�1�y����F\��r���cXLA����y"kK	�p��gD���f���yL�$)l51���xZ��F��y�Őh�TPx�I
�&н{V����y"$ې��H��ɝ�3rU�R-���yRb��Kz�mX7#��؍ۡB ��y��ܐИ���U�p䛠���yR��,� �"w�Z�;�-�qh���y�ym��m��:1�+\�y��Z*�s#��-w�i���F��y�b�-O0�Ⴅ�;�p=c5
���y���5�!AV��2��w�T8�ymD�>@���wÐeT��; ߎ�y"MR!sOfy��BG�_��B����ybh�	-wU��b�I�>IpƊ��y2"Y3aq���(Y�N3b-y�$ =�yr�ſt|���J�\�ɥ��/{ޝ��iIČjG�ʧo�~�9�GL�n3��ȓs�x�I�%6f�9���U�Dه�qmdBnݪa����K̶g4�-��S�? xU��IόEi4�J6Qe�a�"OT�k����f���3����p�"O( �)��95nL�"�81`"Or����#�бr�Q=T��"O`�
R�&Ya���&�x[e"O�9��t�>y��1�j�2�"O^ejf�=Uj�	��سE����"OL�:�g�#-�<��q���e�"Ot	6��*{(����hޛe�D'"O��1G�ל`xC�
�)�����"OD����	}��1P���4���r"O�-�瀔G�0�ڳ�C�Y�XQ�"O��"$ ��|,�SdH5C0,��"O� ��J� [�V�y�d��"X��[�<��kдi�D�C�%ZN�;�e`�<�2�L'ɔhB#
V���Y�k\`�<A���-.T�!�s�M�9m�Ps�`�h�<q� �4O��xC���L9��[i�<�rA�h6$���
�v�z��!�}�<)0%�M�]R4'���s�\{�<����1;���C6���|�傔�v�<�� ��J��EF*˞hO	� �l�<�UBE56LT�p���Mӂȝi�<��L!������G�Q��5��f�<���!e�>���HN��"p��/�]�<I4�N	M����%�R����c��b�<	��S����KT;���D�<a�!P�l8��#A/���EK�<A�=q�60r2ͅQQ�	�F��F�<�p�@�+�[PG��v���+*AV�<��!�<s�m���"4��Åf�_�<9�M�xi�@!k,Z��&�_�<�vc�P�69P������Im�c�L��w�ON�h��o���;@��$��:�'��	`j|�x@&ݰ�jl3�Q!rOj��P�3?���^��x(���}}��yf�(<��͂?db}���R(11-�|���cvQ��� 8�'IF���dŧ{��ԛV��_�X��Ó'(8���E5!)��R�b��<�^��Q�i��Y��h��o�<K�B䉢�䨐��7w��%�8UĦ�	\'��ä��,�ԍj��Q	ap�}��.�#:�cGK�|�6y�C^�<y���lU�f�ˢg N�w"�B�:\fY�V�ˣe@��bLL�D�$�)Dx��"R�	Z��@r�V�[*�}R�VY,>�g�
`�v5Z�ǋ�]C�DZV$L�/$�X���Sp��u�(�O�qI�Y��v9���ם�P\ۍ��.Y�8�Fl�}��؈KX/�����q��Hq�Q�=�5U���.��,��)��u��/
|��lB�oֺYgX]��]�O��Ԉ�Υ�|��&�-��e٬�4%�+]�2��M���U�*�t���!yDN�c��C��$Rh��-��I6�A�A�mebqZU�̢m�0<���ۖ4�i��F�%Pl��Cs?��-C55�󎓅  daZ�m����
�t�|2߫/��%���IP;b��Lʰ{�����o˯�2�S%G<TƲ4ӇN��yBJS�W4|�s�2����+V��&Δ����2L9+:�ffJX����k.R�Q�#&?|�:&���b��'䤬1�KM�x�~1�B)6g��@2�
����狗C���2�!gB�.b��.	/ �b)��ѱ�D�KSnK�V��Z0Mc�=� �:0�,IH��j9�L	2b�]AI0�Б��-��6��6�ݱ
#,��
�c���h�㇆CXd���C�O1�%z6�\�d<xXHd��5�*��t�\�f���0֣GFJ6MZ�_�|������;%B�b0�$X�ax]Z��ߓd=�g%�<���Se/ɝzl���G�5X3�]Y0���J�đ���-z�,P�]��0w@�F��+f�?q�٪qn
�sr
p�'�Ͽ����*�)'�\�2nA�~#6�?9���D 9�K��TCX���|%�#���AX���GG��cn`*��V)7��m�C�>+��iր�98ed�RC�=3������\�Gd<Ց���)vI���E��3ԨX$&�c�gM>Z�~��GLCm.��a&A(tO����(�;4pΌ04SE"ޘ1��F�Zn�)k��k�z0Kd"Mw�~���3�a{��GTY�ݺ�L�"+A���m�SKl�	e�ޮ:Ⱥ5��
3��)y5$�PT���sL��(G�����RHx�Q����Z�z$�[2&A� �Ӎ��=qRʁ=�mhcY8݀ l9	4��]Vr���eg�5Q�
�Cˠ!��W�'N-X�F�P�b1$L�XZh��0BT�a`�-i%jWD�V�;�(�$��E��2^[�1"�$K�:AV������*G��Ӡ�E�`��8����)yN�� � �������4�sE]�$�9"�g�t!@;_���p�ә&���h�D�#fddI[��40���9F��
, Z�&�7R�p{3/�gc�����c���W6Q�hKS�	dk����`C"e`Pq�KƆV���h�Y�R�y��Ec�|X5J<5���<$��FL�2If�[cB�6�6���!��Yi��䖸7"�	P�냩:<�f�2Ak��
�٥�U	��@��4̪ ���%]�<�''|O�I�e�(~l�8�gG*<�ƀ"7i���������'@v�)�(s�h�aZm^�QA�=�ذr��G9��fE��!L`��#I��]"����C�Z(XZ�X+e��&1���[�x<L�7bE6W/��J2�iάy�HC�M� �A%œoOQAW�6�$h�P�\,��ДUИ!uh!I���=�FH�/Ll�"BM��p��¥l���!"�>.l<Iddڋa�4`���H� �ƒFJ��H���m���@$�YxK��V*� �]��$
�EV���7�K;d�~�P�'k�xHBN	�,�h)@�DX~<�BD�L"�b�v���A��Am�`pB�I�(�t4DYz �2�f��%8�iQjJ#R�(�##I/�����������s�X���5NC�;;6x�b�8?X�R�J �Y�"��s�B4*XT�;QÄ(2�$�ծ�<4(6-�w#`�8&Te��A�u&C>^��Q�J�7D%I���� J����{�>-:FT�h�T$���J��M{b���=�t]h��B+l�>$�g"R�!*�؉s˗�w
.�ʞ''&� �M9�xMDx�-&V�D�b#�S"���35iW�
ߎ|*��U�1�&��ػU�h��@�ɥQ�Z�t�ĉ�\w�.�bl8-a6n���$	ҦSR���I]a� "�ŠY��{ �.��9���ɢV�P�-O,�+7��u��_����D�����1&4)<G���ٕ�� R����_>z!zEA�- mH4
�.�h<)1�N6L�;2%܆C�\���m��H���8&X�M ���Y�'���a��
;P�`<��"�M��9q���T1$�\��S�ڗr��� ���"�R9.ո;.�;�
�&p��ER�d؉b�.T9���97��q"'�8�O.��b�ӕ
�4}#���3�rl�d�B�, 0A� ��a�sI��O�0��� �&�d����9�!W�N�s��cM��5�d�t"O���qmױ �&aA�G�"m���凘��h)k�o�1u
m{���S1�,yq㇑�!h�ԋ�'��k�IK%n7b|XR���gL�I�2>Ȉ��(�=u.�y�"#M�~�D�I��'	�����-;� �G��C4&�)2@ًY��aE~b�ڜX��\��g�$X��w���hO@��g93� �)FiF9���2��
nxv����8b}�L��o�5->r9����{J���I	D\\ PB��-���T�M�ƓO�!����0H�ܩ8eD�#HF�1�_R�S�\tR�8`���\�d�H�FS2f�B�t[�jG�)&|"g��*B ��	%�#q{V�*����q���d"+�S5��DE�W��Y����\�^��B�U(T_!��ɩCD�{�J��e�,�(���(z0����=�ʄ#v(T�j��G�)��Br4�'��tZ�QJr�_�f����	�~��x�W�Ě:U�a(�1tk$�R��G2;j���cLc�s�"�OtQ��� S���D �#�@���DL�n0ɡ+S�C.���M�% �O�*lʶ��zL���2��-qC��q�'I�=���4]~��E6Z��B�ށM���9EƓX�^|Ӈe/�(��I�v�� F��o�Ra��K
��B��Q{��c�4^��c�3*����G� ;��l���P�40r����^�'ֺ�Q���=��9���{���ߓB��p�'	M�w۬��I� S6ޕʓIGE�1��%k�*u�'%R���KD�w~�Ô"�q`��3��̱}�\�:S�V
h����L(c��b����A)*�`MO'g!�D
�3�d)1J��?3��r���S����W0����CC�(�y�_>�.}d�g?��H�q��X���K/~��F��W�<� H�aj�,���F�B^��"ҟ ��I�|  ��X.���dN5(�褪�ŃK/B��WB�(10a|2j��J��AG�l&�9x_U
�j퀡�|���HH��x"��f��Iף���\PcQ�ٱ�(O��q��e���Q�����9��]+�e/zĲ�q�k�@ݑ��u��T��-�X�s�ٚQ�� #��'�$ �U>��O?7�]�o{��iD��m8E�Qb_~�!�D¼�j<A#,O�{�����1���0<���cp�3\O"L�B72x#�M�"O��Hf"O$�*ccψQ$4 �.&���a�,27!�D[1M{�!i#?S�졘u��!��ĵ=�>�y��_5x�6 ���5�!�$��a"���S���d�)�D�
!�ڙ�nD�lȍ'�L��!�~�!��bx&����,ȅYV*�$�!�� b��F�I���������a"O*Y��[\#\��_(IiFx��"O�ݨ`h��f���t� �4Τ�!v"O|a`��3�@	�4C�-���"OT=jp�P�{��%�`�"pL�C�"O8���&"��A�p司r�1u"O�b%�9VO@	�v	B0�(��VJ�k��'(45�G���	�U�y�H�'T�)�K�=3��!2�@�,�R8��'���c���FP�C.�lc�'U��(ç�8j@Y��$�-�L0X
�'��(� ҄j��q%aO:p1����'j�A1���u&R�t� Z��I��'��|P�,�'�Z��kS�^突S�'9��/L@T�W�<�X�P�����y��פeg����%�f�*��:�Py�IAf�tG`�zY�8�(W�<�&o��s~��c6aP�Z�Q�D�<�@٣n�P ��4 8���G�<����mWLm8#�@�Rl��P�U�<��ƟfwZ��NP�O���H"(�M�<a�b�h�r����6�Zx��D�<���Lc8�� �#�,����D�<����3C�p�aB#.4���z�<�7+
��b�K��ݖvj��Ć�w�<�jPS��)�fEҒ)�~�;�j]q�<�5���.I�3e�
0���Eh�<�qDױ^)^�Y3��H��ڦ�Cd�<�5
OqR�h�s�ծ}�D���	e�<q�jTPv�Cb�Ϩ'z�@��~�<� �3\np9�dG'(3�e�� Cx�<�3	
5
AjQSO��L��o�y�<�B4J2�b1��	RYddړ
]p�<)�BXp%�V��dX��b��p�<	Qi^W2��2���bX��A�s�<�#D�%JZ��aCS�`R���f�<����%^�օ���X'h��oLh�<�t��:�؃1"�Q�Xq�U�S�<I���0o�$����:ˬ��6b^N�<��)[�h��p�kX�B�$�1t |�<1�F���BQ���#9Wʽ�Q�Vy�<9���|�t�VNT"Q�h�#Im�<�7`�/�P�qa"I��ЀCoKd�<9�ƂG섅@Eo�Pq�M�A�M�<���ݾamZr���=+��XE
�p�<���ǖ+�j9��9r��p��+�s�<��h����Q� �;5 A�@k�<Ium�$����TK�!8��ʢ�|�<A�/;�,0#e�Ը#$4��i}�<i���F����I[�uyw&�R�<���O*D.*�ԭ�X8h"w��M�<Y��-�<�����*i�F�O�<9v�)�$����f�R��D��A�<	u)��T=��Y�׺��6T��!�cE>;n�*Uf�<&��sI8D��ʷ!�c~��Q,ܑ X�pfK8D��C&�'K����I6ek�5D�pc�Crhv�r`�7��
�+/D��* L�+������3�4�R%-D�H�B�3Z�`�X3�?b��P�g 4D���4i��&e����'.��l�Q�3D�lz�k�3+ EQbL/1�¸C7�0D�dy�NEx^�=Xf�ܙ��x(D�,D��0V��z�0�0�)$e�Y腁4D�� �eIS$V�D
Pr1C� f���C"O��1��C�}��̀pe� 1�<K"O�y�D�Am���ҋ�E%��2"O�	W �>�~�Ʌ�$*��c�"O6mt�^�O�<��!��8-
P(2"OJM�1�Vސ1����
5��`�"O��$ � �T ��º)����"Ox���˘^vB�s"	H�0�X0(T"Od\�7`˿?B��11Ky ����"O���/ڙG72�q`��;�؝1�"ON��c��0���aÄ�\��P#"O2M�r�	3��-�gD�/W�c�"O^a�C��X�Mrv�Ʊ\i*qBf"OVȺ`	�#j�`U�CA�#oY�9	�"O�8A�˕S��Z'׋Ae�!"O�H�Yy��	$e��h�Hy�K�V�<ɳ�� N�~�fEƼ^bH,��i_�<�3��ג�Sү�=X�d���W�<���N�XIb�,^>*��t���G�<qPFI-w ��U䛗zĹC7-u�<�52��]��󠽻C@�{�<�΢bqJK΍Èp{ӆ�p�<�.E�s�P����
	O��$Jo�<�E��4�i�
E�N^�%I�]�<ᢎ��u޲a�n	a�RYL�_�<�5M@�%�����=FG.�h�J�Y�<�M� �(�X���?nT�f�X�<Ab`]	���3�숟D�������Y�<1�C�8����!T�n~}���Y�<�dX�j���!�*°KV�<Yġh�|���+g.��@X_�<���J~�����
"��a���_�<��&ߺL��`��թl�Q3�\�<i��|�2�=�:E2�YX�<9���1�:	�w엕3�P"�R[�<�2�M�}O�����J(��B�!H�<i�lߝd,��ϕ�[�쬪��r�FwR]wIC�O�,T��I�TM�(�re�=�=��'MR�i� q��`�̀��]ʕ�g݄O����3?Q�C��rz��3kB,2o,�д!RN(<ٱ�Io>`����&�8<���ھ}n]��&�ji�|Z0�'�n\p$ъ	�y��ǂ~��T)�h�P\�P�/:����<����C����'غ���i�<f$̧n���m�0(YZ�a��f?i`�Ľnf�Y�R�L�i& R�w�O�r��e�'��p�D%�_��i �'Ά�c'�]����D#U�J�J�QU	=cxLu�E���H0^��D�՘���2�	�2ʁ�b��8;�Y�aj�J��$ѧF�p��]�m��Q(&�ˤa�ఫ��զ�t����]d>�h"&��{������o��:�A�@
5��%�+z�Zt��2�f�V@����ݭ�������+"��9+N<5�ĉSOMG�<�f�L�8ծɊV���:QBI�=h7̤�#��.l�XL)	R&����cL����K
O�,���^��}�4�E�x.�L�� �'	`�D�?D��v�ʻj/9�ǉ�H��m�G��jJ������"{�N���Oܕ}�� �6�
;�Ք�O����o�м��$~@�S�Ö� )l0r��EG8����(�<r�(�	N�eF��3���xTH��6���%���Dѹ:�¨��t�`C���*bI����L���'S6a�aF&8+Z٢A@ӑp�P0���d�
D�HZ KH�ڕ#��%�нP/꟞���KM%?-���փ��n�42a�����Hʣl:D����'r�uBQk}�� a�\����8'ߦ���gjɓa��q!��
fz�aZqK[�}��Y.���pVg_���5P'�?s��[EW�r��̓Ol��-�<��ψ�.x �x��,x�Z��!��� ���T[z���M��=�=��/I#(u:��w���Rc��xfrAΟ-�\���'���j���L�i���-��|B3cC0?�44��b��A1�����N�1?( �C�"K->�"��(��`zC��1<�8�O@�����^B �@���wP�ZR�$�[L��b �g��t�@X8�8���D�)x��bi��������׵ �dA�#D�*�tԓQk��Jjy30��Vx�� ��su�C+e|�xʧ�d�v1��I�TN.�*6�H${�P�	��2$��;�B�fz�`�7�E�c�hkBa?TCt�(�&��]��X�6�p�"� '4��+���<����T�!�
иf��}���!:���	�!��r��SF�]<��5�oJ�S�CW����I����3��pCI2�r0�e�5|O�4C�
Ɓ\�Du�0f����y�1��1fUȹp`�?8�,1H����3�H�����eɁ ��`X�%�d !n��J�<�w$ť���PI-�	��,��Т�>�$ωH ���Q�S
+ֱjQ�\�5�V9�t��%�XX�U��� ��T0Jx�\BI����<��l4�m#�ʿhi�����(x �C�5 ���&�۪����!�?�Ikc��=md���M��*L���E�r{�t��
´9ƨ�7Ú3��x�*�:$ѧE�3=�$2��X�(��r�B~\h(�`I�q,n��5�.�8 �7�G�:
�JwbWۿ�R�_�����I�).�F`���=�����dE8��L�X��@�������5Sj���ϏQ*��S񁚃� l[�G�K��dI�Z9�-�Q�|���1R�X��v(CU�A���'�b%�"���5l�,ɤA�/6�VJ /���l1}Qָ�Q���Iz�:�ǔ $�8-��̩<���t�V� xJ��Ix���
���*VX���U
6pհ�,�,6DR0ْe��E0B�������r�'[N�9�C��5wݠ�LΨn�	)�kĮ�0i�Ԃ�@u�B�ɮY ib�'H8j2&��A� ���u�Q�bu����'\��AX�ZiJ���l=8�k7�ă
��N�8kE� 1*˻)6^`�����{p4����M�4����lJ��%g�iW��~�&ir��:��}*��p*p�7�S!�5�c�ݦ`�=�}�hĨ6�����ʸ��@������'R��+ሐVb`0�Ft ����eʻ� �lZ�Ijbyi�券1��uRt�]=&��tF�e[��C
g��ʣO�#��T� kݹPc��@$kޠ?����������[��C��!�S����ĝ�2�R�]���fH:vT��d�P-Jz��x0�z�<�*�6L6�)0�E�p����ɂ4v�\Y��`�� ��ɤ���]6N 8�q�v���G����e�a�
a@䢦)Q�E�lL8���l���C�-��
�׏�tIJ\0v��PjI�
%"؜sc$��s��=�-�&!���(���2Mf9��s�'-�|A@ �P���Sd,J�+�����b�0�J\��A�H�fkgh{X�=I�ID)���D(
-\L�}�a���\�D5Zc].H�����$<�OX�h`&ϑ򅓤Q����/��`5\�H �qA�U"�(��^�t}p�c�
i� A��O ���?��_�L�C�G��$��F�^/b5!�d>l L%[��,B[p9	�J�#�ջ� �J��rd��ӦI)�D�?-CPdZ-A]|!9���~���5�:�ҧ��'�R|�@ D���>�t�@�\�E����OzL}S5��?t�"����̆b����4���R���;����|�p f�|�'D��e���$�T� �w&��ڏ�D_4�dQ�Af�+�2�S�A\
:��!	K׷n%b�y���:��͡Ԍ�_�]�B�[���J���;KS���	��<(p*��.�'��(�j\	#D"3Eܦ/Nv���.�i��K�ȱnTTPԼ�H
�R!��G#�|��)� hy��he��\�l
p� $/�L1�&��%UT����)
jy��ʁB+�(�3�U(x����I�>�y"��H�~Zf�Y sR�u
�
�;M�ީ�D͖"c�9Hׅ$E��������r�aѣS lTه�ȶK���	R�MAbMӇBM������B����:,�ĉf%�.d��I)1�'�pd�A*������'��h��\��{��5kd:l�T�
�U�����/����' U��D/�>y�KDA+_¨|�ȓ3^u8$b�)ʲ.�9l�(��Fo��I��X (���F��p����B$!�K�F'	nb�i��[�!�!��Y��6�J�W�ȹ��Vtz��J� ��%��M5xYh��9��&9:� ��2GPP�f�ݢs�����l0�	bgI� 2(����>-� U��(��3p�N�,&��
���T�7޿7\T�@'�N���?�bb\�w-]��Y>|i�������?k�Pr��]�/^��K�Þ�y(�k�lm��"��́G&�)��5�F��\#����Q�<����Ol-� ���/�"HI��GT�%a�"O\k���s�\���+'��e���'����T�Eaڷ1럶�p<�'_�$�d�X��ռ"�᳍�p�$'�n����=}4P���/x����#�X�f���'RZ �3eHGȅ�%
����Ѭ\WV�S��IE��4���;�M��kO6
�.���"O:A@��L�{ź�{�냮O�8�b��i
Z��7/X�s�|O?7�ʎ3���'έ0���RRI-&2!��K����y�M�o�F�y�O��	�4���1�%\O͹6�Cm�\2�ߴt�j�"O�eY�g�b�6-0vk"39�"O �䃝�Y�:@)Ω'��� �"O� ��	ֿM�Ь��G��4��9��"O�=�@	��=��A��c?=�b<0�"Ob\���Y�|nU���r�q*�"O�X��D�Pa��p� Ws`��P"O9��_�����O�VU|c�"Op*��θr�%�B�G�Iӡ"OE�t`p�<T��A�����"O�鱣�̎E�l���-=��cR"O�L���@�-j|�8��+�µ�&"O~i�e���4�h��(R�<�"�"O��B�O7&ӺP蕍)o��uۅ"ON�ʱ�X'�6!9 lX�v�>��U"O�5���Y�y� ��-U5/?��"OrIzA��FM �т��}�y:�"O��Ԣ�Bz�q�F�֥]<L0�"O@�X�B<|,1��,
��	"O��qD#�lC��KN��%�0"O|5A0.�i��	0CS�!����"O����䞡H�P9F�ʲ.ڐ��"O�d*7��>a�t���ǻH}.�;7"O���%��z� �D@�J8��a"O�m���Ȃm�͋��4���*E�'���%��yTX�Z��Z�)4-b�.�EŲpȵ�Q!Y�J-O����F�f!b ՆM����>%?U1�Y�vl���̔:1�n���`���1�l���@2��I#!՝*-@�F�Œd	� b�x"��%�L	�y��4��4F	�s �?b�9*�^��y��λ1���0>��>�t$�7��5�J�T#�<JN6��D��0J�V���S�OQ�T�r�	�z�D1�H�(�,�� �%/����yr�G�O�哋���	�CO7_�"�;0�Z.=Z<����O��aמ-���O�-�OW7��J���dty��'q��,D�2|A�`���x��O$���G� �I�V��f����m�� q@l7B�z����8�9�(�;�Ω}R)5�A&{� �B��'(Ll�7�0?!����0�գs�T!�U��NO�OR@��Z�$IE��Ox&?7���';��Qs�a\�1�D�A(-�K>9�A*)�ᓪ�f I��ݨ|{������SL�'��lyCiY�����ɴ>�FH���$B�1�%qu��}�M�!���=E�tF��@���@A��>$+'��'HgFe�a,�߸����x���<V�c��١u?�\"���]��>��R!���J0�y��~
�K�����cǚ n�X���f� o�P�f>yS�[)�j�O݆j�<��"�<G�ٿu���ش��d �4��~��&:O�I��X:V��vh��aiP�I!��C�
]ay���O�.�TYx��WMR<e�z���/ºP�ЙI��W/~�&��'�@&>-�}2Rz���h�lU.4Ӝ�C���#4�gj�>��\2���S}�Oqr�1&B�{��)qb��%N����O��[��K/�3O��?;F��~ҭ�nA�1cJx0����<y��[��#���o�Y�O�J33�P}�|-;��Y�NQ��J,�Aٗ�r��@ G�	�^�Y�c'%x�ǡ(D�XC�]�(�\i�@ON�}B*貅	1D����6(�~I��?��X�g/D�X(��R�f쐗�-y��qB,*D����JW�q�QE
�SM�� �F(D����HR�$�T#�˕(u��T(�*O�1	W�Nl͙Q�1�8="O
�IA
�	e�Ni"(�F�.��"O�sEnU+y)P�IM�%���YU"O
���E�G�D�ǁ�;\h��"O^y��꘴,Z�S�NA�xX�i�$"O:б��<�*`��]��&h�"O4��P�cĄ�Cƅ�5��*�"O�qy���121* yp�*vΩZ�"O�yR�mҶI*����	ƛx<��a�"O���F]? ���:�'G����6"O�`ЃbZ-�Ȳ��b�2��$"OƱB�^G;�L�u���)K�"O� �����/j�щ7%���=ys"OV!b%��AT¢� ��=y�"O�%���`�p��큩}2LI�"O���",�D�l�LƚNluS�"O�%�'#�	�F�S+��D�T�Rr"O�8#` �,m�������C֖�z�"O�RW)P�]���,�I�L(("O@��@jV�{�L� ��r�b���"O�u!�jU=R�ѕL�H��0D"O��k �^?9q���扙�6�r�"O�h�B]��q�
�
lai	3"O�`@K�lm�p��[G�:�"O��Ň� i��I��A��@;���"O�9c
ؙ5�����n�}" [�"OLࢂK�^�)�5�V�<`��"Of��'$O!P�V���O�"8#5"O�L;d�F���  �O+"�p���"O
�b���+h��{qI��(ט)x�"O�I��ֺ#����G��5����"Ot�I`H3D	�t�	%d��ay�"O՘��$d ��;A"���"On�)P莘,9f��hM)'���p"O~�;�o�"fx`��� b�:��`"O�s�Xx���ᴄ��@�� ��"Opapc��K�F���A�F�V�"OL�#`�R�Gg^�"q�� �V  D"O��yvm�0+���&�_��3�"O<���+s�J����ԯ_Z�)� "O:5�m�X��#�BQ7?O�Q�"O�p��"G�@�#�7)7�)cg"O�Q K�D]bg�˺E(0f"OT�Q��o���i��(9܌E��"O�I�a >b���R�߿~$`�¦"O�tP��!J�ѡSIˠo�ڰBG"OX,�!랹{�D���MJ�pZ3"O� ѥE�������i
΅ b"O�����ܰe1��Պ����"O�y"IF�s�8�0��V�6�|�""O��3K�M�.P�`�b�d�s"O�<��#�Hߠ�
e�P�Q|�|�"O�H(F�G�X�SŪ ^� ��"O�H��5n}@t����,��H�"O$ha����(����e�RL�US"O�Lh���Te��e �xv��"O���D�i\B�z4$�= ��Ȱ�"O`0Cl���FS)���J �P"O�<2���S$��BpK)o�ܩRq"O}[P�?	�Q̀7=����"O<H���E�q�0Ձ����n+4T�`"Od,4H�}�8�bJK�B"J�(B"O�Q2qfS*TZ�� @*9
��D"O�(���J��{��[���(E"O0` �>g/nx��+hz��P"Od��\�|�usP"�%h.�u"O6�B�3�>��@h�WZ��� "O�|:4lޝ&�����zY�JD"O.���i��d��4����@��h�U"O4����B�{��,r1��4)�N5�"O��S1�8{'N���>R�j�X"O:l��.�t�U�ִ�g-�F�<$E�71���W�O�"��4ڧHl�<� �$.��L��S*K�h�d��L�<Q���=����ǋec���UE�<�R�5��t )�.fb���a]�<� N��©4��Q���8o��"�"O��i�\"��Q4Iق XZ��&"O~��6Hٟmv,�8�G�2X��e"O.i��+^"nir���*j�qt"O*��̭:a���@;�v�&"O�\�0j�>�H|C򎑞:�d�� "ODt�r�X3"C ���d�5z8��W"On@���a�V8� 	(�l	�B"Oʅ�Q��8BD���l���%�e"O�@[4��!/*8��w,�	�v�C�"O<�b_�b����D,8XBa"OZ�1&�"[.e�t��5)��"ON,���U�CHt�1��=ri(�a�"OZ��b͢bO*�sB��15hL���"Or=�1��;n�TI�l_2�B3"O����w$`�� �	��`J"O�@���ݟ=�DI�dgM�l��"OT����^#ĠrUƗ���<�f"O�����H�y�C���@�XI�"O(iP��C���q.ĪR�[�"O��� ��S�d��'/$S&z�Pe"Op��2-�*9V� �Q��6\�P�x"O �����@�s�&�����"Oj9"eC+k��\�e��Q�,�p"O<�Jr��%_JR�ă��Iء1�"Oh=� �:[.`"��+<�L�RA"OH��6#ՙ#��9�������"OVY[6Y�/t��0���>���"ON  6�V�dfZ)�&n�&;��В'"O��QV�O��C��m�%&"OfU��٨8Ĭc4��P*v(�"O�� Ğ�>�� ��/�!C@vE1u"O��fCX�G����`�"6	�"Or�yӇ�'�h �
�5h�"OJ�{G�z�,�� �U���t"O`Au�I�I��@�ħn�~]��"O�LX!Cai�C׎\X��#����y�iE�npNx�q�I;Y���#	O��y�a ~N�x�!��5� ��Z7�yB�ӧ7��8	7��"y��т��y�K�S8��1�]�i�`����y��P�#*T�S���b{"p�Qnͣ�y2%�z�6 ��)�^7���ٔ�!�$G?æ0a0i�<��kZ�c�!�ę �>����,L��az�i�~�!�D(�!x�Dәq8t�����B"O>�cB`��B.(X��kO67Mj}x�"O$�
��
}z��j#��&(.�x v"Ofx�Ҳ5�y�r��o���Q"O�5�1bm�`<����8llD"O��(cI^�&$��0J�O��y!"O�(��ƥ:0"����ȂA�֑i�"O(�
Z�]24�Ab�a�()�"O���#�K"g�`Q6B�	͒p��"O��t�p���ɐ�ǕWYv5��"O<kҾ=�F@�"ʞ�^M�c�"O� �3j-X�pO�m�}I�"O6� �R�2�UQ�(��Va��`"OT�rUh�9Ȗ���FO$xT��"O͹7��_����3��8&�:�"O(<I#��
`��� %-IX��C"O.�B���T���s��
��Y"O`A�o�9o��:Ѓ@/��P� "OF�)�+Z�A�0$�E�6g�fm�D"O� $P0���y�r�����+r����d"Oܨ���G$d�`u*W!��s�"OH�)�/�l8q�H�':��"O�L�$�Q6O�4L�p�^���+D"O����m@<>�MKs(�T�2p��"O�bVlJ� w�ܓ���%�t�%"OtEB��VD�\��������E{"O�U��=qZ�3@�d���"�"O\�	U���+{��p� ��n�*��"O8�cfc>�fU5ià0��3"O��eI�-�m��~I�E"O��S�̓/�JL)�	��\��"O��)a`�R�� ���\_T �D"O��i���/���'.7_B.��"O��Q��Ą
�Ñ!�E�q"O��YB,L�X�����Q�#�P���"O�I���
��(� & 5��ሤ"O�$vЉ@,�,��e�h� �Z�"O�)`�F�,''65���.%t����"O�1�"B�x8����a֌Mg�$(�"O�E� �m���S��,d����"O�QR�c�nP�e��po�`"O��x��/�J��(�_f�`��"O��*`��4e� �i��\e��ж"O:ISp��a,�U肨R/I[�1��"O2�Z��	�8	�,X���)26Iq "O�E1ՅU���-�P���j��"O@\J@l�<!�8 x+U-@�j��1"O©y�g��Kg�� r���cG"OI����ָ����F��P�"OP�W��{o�g�P+
a~�z@"O��Q�Q�m��h�DF�Q"�aC"O85���J:�Zu���sk�)qP"O����8��p�nO����v"O���QƮ�5`��Է��EK�"O�u��&Y��0��/J�� k�"O�̱bߚ6��H�sO��c��h�"O��
�C�?.V1K!(ޓamv0
r"OF�� /�־١"�$N[X˶"OP�@1�T�;d��j�!�'B�1!"O�Mӕ�&X�e"�j�;XUR���"O@-{U۱��UhR�{��R�"Ol�a�c,�z��P�p�C0"O���������8���>@����"O|���ٳlĆīqV/z��4c�"O���6k9�P��h����p"O$��w�ɽrW
��D������`"O8%���N11��d��#/��QF"Od��.�6��q���%9����"Oq���
9M�����i���e"Of̐B��}L]B�p(2&"O24   ��   s  K  �  �   Y,  7  B  &M  V  �a  |k  �q  -x  {~  ��   �  C�  ��  ǝ  �  L�  ��  ζ  �  S�  ��  ��  ��  p�  ��  L�  C�  ��  � � � � 2 w" �"  İ���	����Zv)C�'ll\�0BL[H<�r�W��,Q9�	
l�a�&�H�<���@=-KD�ぉ�	�xhA�a	G�<!Ьѣ_�<Sw��U_N�F`z�<�bDI-J����Ҫ[�:�\`f�Hy�<�Àu�ꝙu���4��m�r�<Y䫐�|'�t#N		3 ꕋ5FWl�<A����z	���A�V��XBBGA�<a!�c�*�Cɒ,̰G��z�<�Η3���Qr��=�B� �m�]�<�p$�jd�%�RH�[KxH0Տ�Y�<�J#j���mŷKO�E��AX�<�W-��5��D8�5��H�U�<���N�(H�"�Ew��;��W�<�&ᐵ7x�X�^Y0���q$�<9����vƠ�Zϖ�n�<`�&	z�<�$k�+8*,}�2��\|k���w�<��'��$RPң�K�a6��ZE�q�<y��_=d��6Ȏ�.��Q�6�QU�<����:�u�9`�AQ�D�i�<\h�r�T7^��IB%�n՚h���b�`��B�y#`q!���
p���ȓf���C�
p#�YTN 	&%P��DY�uj�:�R�(׆�?�D���A�t}��E G��0m�2��هȓ7.�b���+G���P�ML�QP��ȓq�L,2�E�%�zY�f��#i�,Ą�?��e��ߵU��2vC^�Bb"�ȓ'TFP/N�gݠ����� �D�ȓi6�T8��	3>�ĵ�vH��W\���h�ic߳'�N1BKBo��U��r�2���n��3N�t)��M���ȓe0��D�G�n���EKV|�ȓB�|t"0,�*_֠p�%l�23����1�x@F؇�jm���'t��h�>Q�����
�y����!�ѣ^$́1��Z��OZ�<ٚO$ʸ�� K2A�8a	�cN�h���)���hO?a��e[�L�&	!�!L�c��j�N�'>Q?�+P���P����~5Tm�:D��H�U�,����s�B�rU�-}r�'S�U�2�զ!Q�i㋒4y�bDK�'�x�Ұ
X!&�|}!pW��z��{��'��(��c��[4R="7���d��'1X9� Rr򢀘�蟭�`��'�1O��S�gy�뚾��x��`�&4�#�)��?�Q
�<I�"~ʑ�ǒ�	1rN�	A��0P���'�yr��8G�� �����>�vȉ%����$9�O���*u�0��,z�600jZ�VO�yb�ɱ&�E�S�U�d)xW$�g�pk���e��%
���.X��u�t�՜/�$MbF���R"O�e�`J��ɼ�稜��$}:p�'#�����I�� �M�quH��u�ā`"qO��D$��5�ɀIg2�Q+�:%>�3�j�+[}dC�ɮ�������9���^� `c��o�Z�㞬%?U��K6�2*U�
��#��(,O&�'^B�I.x1�q�W�9"��eJT)��)B�iY�Ֆ'g��4�3�dI?C;��X��P_5�rc�A���b��(��}��ӋQ�^P�da7MbL%��*|O��9�K�=�Ƞ��N��f�̢��'P�h� �zcbX���yV�_�N.C�I�:�扪�̀�&�썑`�� 9�@\�~��'Cay�ܜ_OF���.E)-�m���Q��p?Q�O��b�8��X�慅�8�E��^�TGxB�I�3��ecDE��@Sų�Mg�0d�?��8�S�� 28��*�?���8f�_�)��B�"O����B�m�Q,H�ǀh�&Z��$��9��Y�H�s�\�o\�|+�08��3N#�O��QL$h`��N�#��q�dHS�c*J���	(�yR���y�&���/��Ek:������(Od76��>Q���1!�Qh��ӂB�z4Fyb�'j.$���auN�Y��2U�$ܙ��)��<��ȇ�%H%�ҧ�o�
H�moy��)ʧf�A�.�5$"��-�[?���h<��E"}����WHUX@�Aa�zy��'�:uʣnF����� �օ8��\���~Bg�8L@hHf��\�D1ɒ)�=�y��V"��W!�+Z5()�#m��y�˴5�n���D=Y�l-P���y����,`�.Y���Aw�
�'�t��������b�Q�ء`�'),�`Da\�@˪٨qDȍ6I��Z�'g�Y�3�)3�f���,���
�s�B�'��	�\"Z�Z�mU�o(�`��� j�B�	�'��㠍�#��y	T�����듿�� �)ҧ^J,�[@L_#o�6�2u�ќz��u��@��1�N��AI��+q'}]���r�\�ICh�K�d�[w�F�zD�ȓ-���g�}����G��:�ⴄ�<`&,qb틟W"�p��C�G��T��x���S"��9`�7z e��x����ᅖ4�4T��_B^��ȓQ�BtʵG �@�,���j��B�HF}B�S)iH�2�C� ~�2튜d����`��h����S�Da�����)*r=�v"O�ib,�2z�@R,ů=\�c@5O���D��ob���r�V3=B�8��^�k>!�ė�o*��g���*=DD��K1*!�F�Ot��I�(A�q<�9s��M��!�dE�Q�����R���� CM��!�D̝�  � �4L̔��"��)R!�D�'k4ms�HFj����� �$B�	���On�O�YRٜxѨPs�F�F`��+C�'�	�!g�����Y+��Q�v�U�!{TB䉊1 ��*��M
����OU�G�BB䉻K�&љ��5p��� F]R�,��{r5O?�	�En
i��kk���%�#g4���O�6-)�S�O��8��њ��`�� YL��L1$� �-�&1a�ѳ�N]�P�H6 0D��xb�į'�}�sH4z�D���-D�����)&�w 6_�$y�%��<�Q�19ۀpD�A�}U���V�VE����>��L�/X�#E��?��bM�e�<�K(z�����"GU
� e�c���~R�'��>} ���Anir�W�<U�c--D�����	G��X�qJT3b65[�,D��UɊ @�f��t�L��"�qAH+�oZmG���1��x��R���°���@�	/^R� ���aL�Y""=
h�C䉔/�\�x ,�01S�8�0O,�d!�Ie}����?�$�LU�u��l�kʎ0wB�>I��I�*O(��ec�X8�)Zf��P��I�+ڥK�
O�=��Α-��Ԓ�{�O�������Wo����D���F4bX����?��E�&Fq`�.�*_�b ��ePV8�Ez�C�$:��A�mß��8��ӄ�y����Dl�Ma�5���Re��$��Ĳ>�y��LJ�Lqy�Ɩ[�dH�π�U!�$��*� ��)�|L �z%��ў���)� �Hp���-ip��U�UreZ ��'����4jf��'�ƑL�H�3�J��5��1��' �9E�L��A
Z�ym��	�'�<���K�$J�1p�E��"	���GO��7��{���+f���Y�*0$�`G{��$�ڥ1I�݈��qZ�4
Ea]>�y��ԺLĂ 9��,f��k�M�5�y�@�l��s/��c3  8a�M"��x��B�W�pM�oŅc\��ks��sU!��L�J9Q�C@p	�e� PJ!�$̚^�H��'�%V�p 8B�N9az�D)n����ĸ&�T)�T �,ˉ'(ўb?�0�m)?~��b�E*�կ<�O�扠E�L���A�?3@{�b\�`2�㞨��	
bp�:��JB�����ٜ<�BO������O3�r%^K��`���۬8xy`�'���H�q��iW���(*��K>q�&��=��׍ �+�Y�2$��K+D�@µD�Qzl�s"��[�$����$D����B,<����!ATItN �Lo�3�:�{� ����T�W*B䉳LƤب���_B�xu�ʾqN�"<�ݴ�0<�1A�Tf89"�yj<4a�N�[�Ic�ht�ȵr�z}��(۽c]\�zd�,D�jC	C$��tQ'�؈-;J8i!j)LOp�X�A�q�@CBmX�9�v�g%"D��:E�٘@}r���h�Lz�3 !��lܓ��OV2�I!�ߵn"�	��2-ðԠ�'7�(
0��� �܅����7/���'=�YC&��[�(�;Q�H$O`0�'�V�J��X�6��z�@ͳ�a8�'�J�	�cR?ug�A8"�<�ĸ1�'��ɨ�a�<f�D�$O@�.�1 �'20�0v) +4�A*3%
�w
~Q#
�'����� N�����G�0��
�'�J�F��`YæD�k���'[n1�V\�5����G�$m�h�'&���Ͳ"Q��["��%� �+�':R�lQ�Rl��i�
V��'.�ȓ3�������	��<X�'��7%T�����^ m��Q��'K,�zV��*_�p�cO̥u��ݛ�'ª�#f�)Z
j5r����ƴ�'�aZ�-��F�h*�-�)��q(�'R�+�����d�C
��6���'��A#s�8t�>���jB�)����'� �%M�� z�ˌ�n�V���'�=� h M��,!5놥k��hb�'	T����c�u�To�;�V�h�'������WDH���Ӈk7Ф�'ꢽ�&F�9��HҐL�/x� �	�'^�`h+���S��1�9��'tJ8zV������A*,��3�'��
��O�3�|���Q'�~�3	�'��So׼
���)����8M��'f-)@ ɯDY �A&
ڳT��'��q�e(��#Arl1fE�>z����'��I�#�z�ʥ�Dcn
���'��ࢥ���}�L0�3ρ/hnR1		�'��|��ьBs�	ѵ�
�t�.�+�'s��p��P"�g�#onFx(�'��Mz3� �h�&}�׫ÔV�!��'�|4�]�A��+D[�]�	�''��*R���qֆp	�l���� ƌ:�&B�)ɪ\�&�	�k�Z 
d"O��P6�Ԕ[PM� �D܀p �"OLL���Es�|8��ÛB8HX�"O�$���>g8�[� R<I<��"O
����P��$�h�J�i��5ؠ�')b�'���'���'���'��'�tрQ��>����:�TU8��'nb�'?"�'���'���'�r�'̉cK\�D��C'��8�Jm˃�'�b�'y�'���'^��'��'��!k1m�%,r<)���[��'���'���'��'r�'�"�'�$����[�hk�];iN�Rt&]r��'��'���'�"�'u�')2�'���Hs��)�T	�.��;r����'�"�'���'���'5r�')B�'тQc��X&^�0�A&N�@��'Z�'���'�B�'J��'$��'4v����(0�<�S�k�6s ���' ��'��' �'���'L2�'X���&똹R��@���Ӵw��ds��'s��'��'�b�'U2�'6R�'}�[�냱n����o�""Ȩ D�'���'�r�'��'���'(��'�|�ywe��Kߚ,s��:i�#�'h"�'���'e��'���'��'f~����_�lx��-7����'p"�'�"�'�R�'���'2�'~���/\2V����6�8~fv$���'�r�'�2�'"�'�7�禙�	���U��2U�p=���A1
hT%�[~��'c�O�͓g��O^�D�Цm2�"ZC�i.�����<,a�q�{�ȳ۴n��)�O>�'!����'�6���=��@��6���S(Q9����Ot��������O<��@��2~�8X��`!`�	_����ˆ6`D�+��@P̓�?!)O~�}Z �I�}ܘX����;|+���m/����1��'
�8pmz�y3�#�6�ryك�ۯe����I���MӰ�iK�$�>�|� ���"�̓��r+ú:�6��F ��K�(�ϓ5�r�k0*Ҵh�8���4�P��>`O�{q$��<�ͣ��D��d�<N>q@�iI��;�y".��Aň芶@�$u`������o��O,��'�6m�ʦ����D�;�&�w�J�O�l�i�Q���	�<?ܥ��M��z�c>E�WM�+���I)ɮpZ���#RB�4��2�X!�'���"~Γn#����B_?u��B�V��T��z��޴��d�覝�?�'�l�����P��Q'���i�`e͓9�fp����\'9[$9@��T�B��*k�BhP$eK�y�������&�ý)�N�Z���s���F��ev�{�m��?TmP6ό5\����Ʒ=�Y�BÐ)b�\�"��$;̽Cq)�?��i�EH�7hO�! qE�>����1��3V�̰�'�	zLA���^1梵s�y��F��T��h�F	>t����.�g���Uj�ly� ��Nv���wjF�G�q(WD*\�D v-�ΐ�0 ��,�y��Ä�L[R`�"�G�;wH����)t�)t��!� �۲�� ��ٱP���Xs"�x�� MH֬BA���H�ب�qa	�a_n�a�c�4)��xR��6�O~���O����R~�h�;�j�`r��$�I9��B�M�+OF�kG�i>]����?6{b��2�&yw�`Jy�L7-�eS$�m�˟�����6���?)�4gn�%�'��K��a3���Ah6��S�&��3�ş�a�J[����x!�AwmW�M��?Y�P���Z*OLʧ�?��'�`�,9���@`��I���1f���O1O$PZ�iY{���$��䟜���G�X��Ѥ��~
B$�d@��MS�,�����x��'��|Zc���{��"E�ts'%/D�8�ȭOz)��D�OH��Oz˓Oq�D+���<7c:�"&'��q����E˝�fO�Or��=�D�<���P<\$��`a�8RT^��GcHX5�<���?i���?)��*D� ��\$r���,�J�ّ�Ń2\�5�E�i���'ZR�|��'[B�_G6ܴ��	s��	&--Dy�D@�Nx��'o��'�[��0�O���ħu�*a�2&�	+h)�G�H10�{d�i�2�|�X�4�&&��;0�MH.SL�� Q.��7�On�D�O�D��:;d��O.�$�O,�	��y� �.�4`3�8��Q�ijp�&��I㟐q��?�<b��^R���R�{�$x �o��:�ġnJy�̸zê6�j�d�'����*?��KN%�y�Ha��CN�͕'�Xш���60(��A�ˋ�M������L�6�K?>�2�'���'W�Z��O6P,a��נo���C��~�H $cӦ�Xb�A$1O>��'^G���GB_ !U�Ms  \�-���ܴ�?I���?��%�a��&�'"�'2��u_x���l��~�0�[�i@v�rݴ��JV�4�S�T�'���'�h�j�iǟL����*ݲmĚDb��p�(��H�R>��oZ�p�I矘�I��i���ҶS%%��p'����͠,o��QSKT��d�O��D����O$˧;���e�6F�H�0,�<)�6y���]�#S���'���'�re�~R(O���_�$��q�L�(Aܭ��L� ��A��3O����O��[&g�O@�ĭ|
�,L�S�6i�1YFU؆a�g
Kذj�$�*��?����?)��?�*O���Ζ4��	�(mz̡�6�H2����\j�Am�������x�I>���Q��nZ˟��I;t�VC#��
�r�X�XI�pS�4�?!���?�.OJ�$ǥLR��:}���	�!���1UO6Ds�.C'�M����?1��?A��H0���'���'���i�O�B��ʹ60�hA�@���7��O"��?��H��|����4��� ʐ�!�<v1�8��͗5�����i4��'a���PiwӜ���O��������O�	��ƛ�P���r�^�	Ӧ�k}b�'�� ��'D�]��S~���~09	b��2X^d؂�Z�F��&�� ��6M�O����OL�i⟆���O����!#R��
8J
��J�H�F�mZ�=*4�����D��������'ʐ��EF�% f)�M�0������lӆ��O��$����m�П��	��`�I՟�ݗx�6a�G%A�={!
�,�7�O��D�Ђ�)4O��?�	Ο`ڤ�HP��B�f^1*DD�:�J��M�/����q�i���'H��'-�꧓~�͜���0�4Շ8u�fH���� %a��d�O���O��$�O��'W��+էǌWr�����L4�hE�q�ʽ.~���'b�'Y�į~�/O���՚2�E
@G�$�h�Y�N I� P��3O����O��$�O��ľ|�@,t��/R�F�Fh��k�7x�θ:3�^�F�6M�Ob���O���O��?�pL��|*4bM(f��4S"G�c� 7NH��?q�F�Z���?���?�Ѩ�=z`��'r�W���\�a��6~r�l8u�ǁC�6�O��d�Oʓ�?i�dX�|bH�`�LD�3{����,
�.���� a���O�˓_>d�JR?����l�S4��ps��G��*`ò�·n�^X
�O��$�O<�D�H�D�O�˓���')a���B�
5W�=����M�(O(u�WM\�M��ǟ��	�?i�O�NK�%%Vu����j[�<A�]�����'�C:�y�#�~��O��s��T1����bO�Ui�A��48ND�b�i�R�'��Ot�T�'3�'���҅�$�v�q�B"UvM�աy�dL�4A�OP���<�'��'�?9@�P��F\Q%�Ο$F����JשT����'��'T�@�r�X���O����O���� ��"M:�I�IP�!D6(�i�R�'6����B �yʟ����O6��ދ �l+�m��X�d�ھIi\o�ӟ�����M���?1��?!Z?��4*�l*�d��-ʄ@Ȋz@px�O��;OX���O����O����|:�I>4z`��ϢVqH�����Z�܃$�i-��'SB�'��'���ODX�$��q�e�WҬR�~4�s��%{����O"���O2�d�O˧YM¡hS�iq�$[6�>�R��g��(;f���q�J���ON���O��D�<1�+���'iv���ҥ�#�vt/*D���2Y��A�G�,�I֟t�I�nb��ߴ�?��+]�̉3�T���}{an��SBB��ir�'.�U�D�I�Lh��֟���M��AxEɅ���jQ�� w���m�������T���8�e�ش�?Q���?��pz���2xW��[�I�2�
�c&�i��P���Ʌ	�J�$����48
-����4Ar�I���_(
m���	�RF��4�?y���?�'���=K��3���䨡���4��L��R�X���m����I������~�e�@/z��h�%E�##��ACA�Ħ���f^��M3���?�������?����?��k�v)�7���7!���`�)_��F��-
���'�i>�'?�ɷz��W�ۈk-ڑ�Wd�3i4 Bش�?Y��?�#^<���'�R�'B���u� s�a�����J�"���M;�y���<�Ok�'�2�:I���h���-&��*Ve	�v��7m�O,uq1� ��Q��ן�����P ��@�I�y@�5U�O�R��%  H�(�%6�Eϓ�?����?�����9OȄ����-i�"E�Γ�3F�p�d��G�6���O���.��<���yUV � �ֻg���Q����#��<i���?����E8ց�'B�=s2��=��u`���-YC�I�'@2�'v�'A��5J�%8�����&�(��S�pʔ�'��'�BV��ꥩ�>��'�,U:��R9X�y7`G�h�(�q�i��|�X�8�g"��	����O�k^�%��g�7 �7-�O���<QNP�yF�Ozr�O;�c�93b܌��c�<FD���':�<�«�\���	�$�P��e	Ӻe1%��C+(���T� c`���M#�[?��	�?���O -+S���*@�㏅�W[��Kƺid�	�`d"<�~2�̌�\L`x��S�g��L����� ��Ʀ�Iݟ����?���}"��!]̞	��ĉu%~|21e5�D7�ø)k�"|��F�
��F�L�ȕ�wA֛:T𣅸i��'�����y|O��d�O��ɵ,",��	�@�& zg˦u�c�2�h:���������Pg�Q��+��M�3��q�+� �M���/8ڌ�A�x��'�ґ|Zc���B��f��A��
e����OĽ[v��O���OV�f�P��l� ����m��)��!�s)݆j̉'P��'��'Q剻�x!�d��n��D����P.�r4l>��ן��	��d�'��C�8��=z�HJ�9��{7͛��� )��x��'�'剓���\
��D��=/���z��W#&�n�'��'�b[��Z�o�.��' p��"�NCCj�y���pִ�S��i�b�|�Z�,	� ���M{������L�s%ה'�(6��O���<��b�I{�OS�O[�H)%��*oV���fŬq�1än!�<�'Iv������P?PI"�cO������U��Z��P����Mc�_?�	�?1��O����0s"a���*6��p�Q�i��ɴ
\�#<�~2��2[��	��8q,|x+�Φղ7���M����?Y����$�x��'���Ybc�{E�k�*\ =� ���e�$<Ф�i>��ן��	ϟ\X� ���f�.�e��-��y��i���'�⏕���O���OT�I/\��a��l��2G�Mf�K�B"b�8�/(�؟,��Ɵ�:�tuI�G
dP2���M��;^T�Hw�x��'���|Zc�*0��n`Z�C"5*���O��+��$�O��d�O��;l��tf΀z(�8��7I��D�	-d�O$�D/�d�<���7]f}�FaӼ�YqA���8P�<����?�����D�V��'�&A�M�6�F����&\�'����E��byBf-��d[����1�ݰ'��V!7:��Iɟ��I�ԕ'�:av�6�	�$Po��q���J T	K/ ���iVr�|2[� �Q�<�I��A� Gэ2�@5�sL��k��'!BV��aeD�3�ħ�?I���ji`�h��H�E���=��i��oy�-�������O�i�p���z�&5C"�"Lc���ݴ���FF��lnZ��I�O&��f~�F��>��%U�s�d�U��:�M{*O�yA�N5�i>O�r!.µ�>e!��}�)�i���&mq���d�O����4 &��	qw�\�1a0S����哼7y�|�4$J�I��Ϙ'�r�Ƭu�������0|��m�|�R6��O��d�O��gO�J쓿?�n���X�ѱ"�0yS4�]:���B�$�3y1O*�d�O��D��;(Bҡa�`���@�^N�Z�m�ȟ<򒆖!���?y����;g�k��j�d�	a�P�m�\}Bg�%��'��'<�T��r�ㆅ iP�jR"ʨ��I�w�S$1�pxJ<����?�O>�*O�M`v(�2����˿ǔu���C�&�1O����O(�d�<q3��{J��K�1�\Hy�M(�^����{F�I��@��F�	{y"��"���̻V�ՁB0Z(ڱ1���3F���|�I��'��r�e%�Ʌh� ��O�MDH�,�pE������W�ILy�E���'b�S �J/2� ���P�D[�͡�4�?������Z>0$$>��	�?AS0'I��B��ueB�~�*�\'��O�ʓqtֹDx��&� ��_�ti�adeYg}rT逰i��	c����4�S��������d�1�(�b"+љ?�	"4G#9\�&V��JBB1�S�p��X�� yX� G�I���o�+��L:޴�?����?���-ĉ'P�'���и����K�q x1R�i�0����ٟ\��'R�`��A�kW�N~6`����M����?)�~VR��&�x�'|�O|c S3B,�ѱ&_�t��X��$�X�1O.��O���	�-O���R�  ��ÈC	N%¨o�����wj����'c�|Zc��ܓ�FN���b�bl�	�O̬�"���OT���Oʓ�����\Ar�-
5��s2"1U.���>����䓴�D�5nu�b�P�X0e@����Ƶ����O��$�O
�`i*�Z�:�6��$�	�:4��!c�R���'���?�H>�+O�5˂^��sB��)�3Aޡ1Er�3㢥>��?	����Pm��'>Y(�H5OT��`�Y�i���B�$�M������¿|��O���s �ZN���6`" ��q�i^��'��I�tjVh"L|����r("R6�Y s ˒W���A ��'��|b�!4� +WLo�,��@�&�M;,O��a�Ǧ�R����D���u�'��9����c���;��fR�0ܴ�PxB�ÿ&~��â̗A��h�&��M5#�ns�f�'%��'\�T.��O�5�B�ٛ�0q�^ :p��Y�l؟L�	�7ج�XT�[	�vQ�����h���4�?����?1��W3�'Ub�'����-r�$(8�@�=8���
1a{��'�B�'�̝�H���x��B4*?��ۓ�l���A�\��e%�8��� '���=o�+�E)al�LYW�)i�(�s����O��$�OL����;s���/�tB�bP9{�|a�BɼO��'���'��U���	柸Z$�¾��Q*�S���Ќ_�Vb��Iޟ��Iey�V�E�x�S'*��2V,
��ju����HO����O���?Q�9O]�OF��EdL
_��tSQ��Pm�9�O����O���<)7�D�)�O�pq`S!T�"�d]��Ʀ7a��q�����O`ʓ�?���7#Ha�����gP�����T�0�<Z�aL Z�V�'TV���kԉ�ħ�?���oP����'ѼE�D����j�b�P��i8�I͟T�I�w���g~��M�w�L��e"��;�=
�Vɦ��'ňA���q�@��O���O�� �r����96�(
���/Ƞ�oNy����O��>�cV��.)�7n
�Jz�x���|�x�A6�Q�����ޟd�	�?�H<���p�ܵ��ZR"�ex�%۱Um�-�D�i�t�bR�'Mɧ�.��J8����c�U�B�ڷ/۴L��Lo�ß��蟔y"��/���?!��~2��M���a"��I봴J�!�%��'�`8��yR�'���'u6��N���
 �E+z%����uӼ��$t�$�p�Iڟ�&��X�?vH#�a�>R�@1�S�E_���`�Γ��D�O��$�O�ʓe�� �5�V�с�l�3�K�,[��}�'����'��';�'��'^���'o�V1& h�/���:�� ��_�S�T��Ο�'?1�ŏ���`Q:o�.ա���x@���*���?�J>����?���<A��lo����7�����^�i����'<�P�� ��ħmo^<��͟�_��`UG�*^<��R�iv�|�'w⣕��y�>���29�L�IU��k}�uHg�Xߦ}�	ß�'�9�9�	�OB�	ŲD��@'��&��$i�˜�{�&�%�h������W�Kԟt$��'=26����>b�YiuJ2<D�m�Fy�C�TB�7�X���'���9?�ab
�7���jr��m���r���I����hH�Åן�&���}�C�ŸF�:���*�Y�.�A�@����cA���M���?�����x2�')Ʃ+% �8=�dp�W��9
(ޘ���Z�2��OL�O>��ɑ�%�pG�%B�m�+C���;/���a������	)����N<����?��']��
��2������jpb]�}�LF�k��'���'�"+��d(�gB%&aZ b�D�ھ7��O��1$�K�I䟀�Ib�i�9�!↛d��B5Kj�T@PG�>�ɐ%���?����?a,O|}r%�����r@�o��Be-�M%���IП�'���	П��'���Z�z��ѤG~�XX���*��	jy�':��'��<4�D�+�O��xSa�CT�S+�R���Y�O����OH�O����ON�Җ8O����3چ��A�m߾�Y�|}B�'b��'���)K���ZK|��,�87��KrnSf����ݖڛ�'Y�'�'*H�}�HV#!8ty�-�0���	���gM�}*��P�K]3HF
q���Y��B���0oġ��Ƕ-���`e,D��	�,�3�R�a���rn�M3�銜r�� ��oԍ[����'0_����m5�n��p�L�`K��t돖f厀2�$ߋj#`�XtN�hΘ�Q�3y9mI��ِ3��%
�5�`sW"ґ^K�]��E�D�(����
�mJ����۫p|��M�/(�'-�DXq����4j�4x$Eݱ�>�HU&�T�	ş\�ɗ�u�x�+U)vi�d�"��x�Ā��C�\ي1�@�/��ɔ� ����q��)��9���t �Cs!Ț����)ݛN��ɲ��qܧ��V�H�S���5�,yB�#�)Y� 0�������S��O{ў����� vpԸ�@��,f�8k`�-D�䲔�/��4�lI����*?��)�-ONi����C�eb�9-������$h�m�7��O����O�d��3���?!�O#Np��SS���$d!� �z�yIV�
ޢ��Ē;��8��&áe�f���@ ~���F��h��2t�a؞,M�;�ZQ ��fL�CF�4Sp����Oh�=���	�@���]�8��:����yB���I��m  ̄�'�:�'�27��O˓8t� y�Q?%�	b�E���]�0�Y���ϵTY`��I�4	�f�џ���|v$	W�����(d5��u�p������{����j�D=�1����A�X�0�ɆM���Eq%�~�^<���ߩ~�PX�am]fNɊH�)0JĨ�="���J<��Q۟��Iey��+M��yA*�Q͎��C�3ޘ'��{�@�=~)���$CK$����<�O�=�'7���9�b,�hI=��r⨋�pRX� U�D%�M�'�?.���ă�O�h3򣖏C�t\�g�P+#�D�+�O��D�M��S�I�2�b�r�dוt�Tʧ��� �I��5�#;*�N)yVى��_7�!31�ܩ ����OX#p���Dܩ�ʽrbE���uIK|�y����	;�p���Ň&��ɒvH���O�}:��ָT ��
ɑF�$R��x�'�FE��Hƽ=��hP��9Y�-���i>�i����q$��*�?	���Z�ilZП��	��y!��V�R<�	埘��ԟ�ݰ?����2d��+B�	����`���	�O�&�I�1��'�Z�%��8v���0g�e��9&�p} �+��O��9��׸��1O���S�ݹ�0��Oǜ+��u�Ѵi'n6��O���1G�Oq���ޟ	V$��i����[�3Ҭ!�[h<Q5BP�qw��qI��X��]i���{~�-ғ;�D�	PyIװ?�
���"J$�P�O� @T�R*� "�'�'��ß����|ʃBG,k�H��a�Ģe�2�Ӹ1�Dt�u�L5)Ш+��'�@��>;��+��]�#��Q�ԡ�� e~!�e�/�E��/V�{X�"q�IG�P��&��L���W�	�4|`pI�O^�D�O����<����'LX���̅�0�4�%�R�ܲ��
�'�9��C5x$eI� �/:��yb�yB�}�l���<)7�!u��'����*9���KA��AI3
(P��'54 x��'�3�M���f�Ay��3}�٣��}�����)I�l~НC#D��p<����4}�t��w���BS�W�0uꚥ�p"@��/��l]�����C�Z������	����'�P�C�0#45Ѡ�<2�^]��'���'n�O>�kfS
O�6�01�*򲐚S#��hO�)��� .!�l��"W��C�P��q���O��^F������'��ӚP��i��%}��e��l�b��,cd�Z�b�m�IΟ��Į)pZ���ѻJ� e��+R�����|��6&��#B��v�vl���]���) �]�1����)�����I7b�.P��f}Ƞ*y�e�wn���V1)��K!���F-}"ȁ�?�i9�#}z�'V��r�ѹIO�e�'�WD�4!�'7 e�'];���$�ݼTB(5;�i>����n�����@?%��K��P��amџ��	��h�Ga܌|{�P��ܟ���ҟ|�Zw��1�Ԍ�%���όo�P��;m���[�lb�"i頪�1W3c>�$��XPʍ۶����*&6�c��6�L|XrKV3rZRa��Đ�5<�"����$�1�p?�2lȰ	7��@aA��wǾii�O�m���i>�D{2� F��4xpˆ8X��u���χ�y���E����T�Pt U�@��y��'��"=ͧ�?�(O(��G
K$�$JSH�#`�ؐ�㐄Uj|�"�O��d�O.�$Bʺ���?��O^����� V�y0D�	"6*0B
�GV�hcE�y�@�0�O�jExT���T�'b�.�������2�0����k9��sQ�	no��H0�.c�2�uŁ�#�<)�!;
��Hᰃ��0��{֨�)%a�)�	� ������'�2����}i0C��D�U>f�зD�!��F���M��A*�f�Y�1O�هF�O�˓DS�"�V?%�	�#5��#5!N����<0OR�������CN����I�|�g�WR�:%ݢ =��3��_:C�P��gZ/	����JA��@ J����	���!��SGMX��G$�ˠ�8X����'�;i�h��� 8�L#?Q����S۴]Y�	�cQ��F#�����Xn�b����Dx����+��+:X�:�E���$M��x"�h�~�+���)	Gh��`�5��O�˓x���b_�l�	d�4,X3G2nO1:�)�q�B5A�J㦌ޠ9���'��Z��Y�^��ً��B*�1&ήq㘹��\>	iS	�� �(��b��
R|����6}�n��|L|�S51� �b^;�Ea�:+�uɭ��,"���?hRm�G,R9�Li �>�`�X����I�|��k��.Er��W�C$hk��u)̬dƶ��<Y����<��:��])&.� ,�4\z �x�,b���CX��Yp�شwR�ST�\��刄��O �d�O&���_-}U����O��d�O��;!;R	 +� X6�3'�ԆC/����%��2�j������F��u��b>�O���6g�7f���Ď��NjBlض�פm;���V�xW ȟ}�q��'���BN���2X�FюqʐR�}�n���@Q�c���>��?Yf��u�Y�A�%&�.�R��J���x��=?4�٥�I����(�+ޅ���l�'X��':�	��hl3�b��	���I���$h*H�*��C>1G���	֟\���;]wp"�'��I9�fI	�%\v�H �vMB@��l��8Z$!A˗B���I�zm��C*Ȃ#7��0ĝ,:��i��(�00���
cQ�2�܅?����Ǌ[ 9K>��� ^����򠄴
�"�b�ţ�n����?ᑧ�i�\��w
�"��$ɦ(GL�%�X9�_���cꜵ 8���#�I
�M{H>�`�Ի���П�qu��?QvM�%�G�i,���!��ɟ���BRf��	�ͧ>2��ig�p��DKty�L�?S��QЭ2���&�,�p<9Ab,b���m�+��!r%���T~t��SFA��������+qb�y�ўT���Op�d�OL�d���Tx`Ɨ>!p�u!t'	4�(ʓ�?	���)@�N���S6��mDݣԥ�
<�!�ğ�胨G*y�T�ԅ*��D�\��Iwy�	��$$����?�-�D�����O��B��@�6��H1��a9��!�*�O����#��mk�!�b�ht#��0�~Eq2(\7VW��'G�<�'�(qV�US�%Ɔ	�r��O�
5�Ɨ|Be��L���9b���j>fx�3�U�d��(x0@/BkFt��Qxā�01<�'{�����?���)�O��:Q�T�?�F����usB6(3D�lsʋ�Z0�CdD9��
U�Pi����N)ғN�0����	���� ^\���1ľi{R�'&"(ĸ7��	�'P��'��w��	it��� l����mچ4�И�A��o3�8�fv�j��`���d4`c>A�c � SZ�DG��i�5Íp�l����H�HU�DyMV>hA.h0Ī�  ���C�CG�Bѳf՟�ȹwBP$�y�L_ �����'>��y�
Q�������0��Oq���'�r����B ���2	��	�'#��c� �9n�C����k�'�b)��|������v+D<�P��"?@$���n�0slik�5x$���O����Ox8�;�?��������1Wv[U��Jk�Y����Q��j��J9bȤ�� 	kb�y��ƥV�0M��^'_�l�P�Z:��ȃŉޜKV�Q�vi�7Z�����$a�ў��7�!<��� i	�-�b��EΚ}��$�Or��4��K����Br���z��
��-R	��t���#�#~��Msӆ��N�P�<��i B�D2�� �8����?c|,�jE!=ت �"O��kWˇ����&b��0�,�ҕ"OxAu�-I2!c >"��8v"O*��
�#ظt��,$:&�y�"O�u��.�^f.0Za��IȪ�"�"Oh衊O8*��g��k����"O�Ĉr@\�%7�%aU�X&�d��"Oj<Ae�;h����GK�%sP"OR��𧉱>����� �t�p�t"OL���H,&ԡ�t���3PK/D���K9��-0
�$q���	�L+D�`CV�U&-*�æ��$l����,D�D;֫�:C�D���
�`�d�(�,+D�P�p�S�~|�sƩG#@\84�>D�����1.�L���*[�:����/D�01��$XMӒ�B�e��EÒ�,D�����u<�X�,��"P %Já)D��Ώ�b'�x1�!O��(���)D�� s���C�(�zeA�-3_4�3�%D��$
�9���0Ϛ�	/
m�>D�Cqkς������<%���K=D�lSڟ(��U@G"Cwe2�%D��ئ-�7���h�o	��(�׏#D�|3񃖨'��$��Y r�@��5D������*{{X�ǇA?:����4D��P�`
%�v0�); �����'D��R���h?�K���e�4'f'D�4bD�[��ȃj� #�\���k"D����M�+�����<f1h�I� D��
/N�> N����G����A D�4r�!�.XβyB��G%}���(D���c��Nat�!�/G��L��(�ɶ)����>I���?:��.@S�).�����B�P�(��R�>��'!�P����埼!�',*��OPT���Ε��8I��ʟIVB˵(�-��];����t�������ԟ��ZH��t����FS�}����KL����R�~���OD�Zf"�|�f���'����&	�C��X��C<EI� !���� ��PyB�?�P�A�f��y���{ i�E��/e��c�'�7!�JPGy��E� h�A�}��qi�GT��eA2�F��&�O��=�O���0�O|]�6d�)4&�}��O��j�F�JE�-��':@e԰A&Й����E������a	/��QZ�I3yќT+�K��d�<)�C7�~���"��ȉ⬪?e�Dʛ�.�,�xV$��C��(���:9���B�'ł��5L٨B*�Њ��,O��M��i�C��#p<�q�A&��<Ԭ� ��V?ᕅ�-r,l�n}>��q�X��V��T�#o��`�!W�7L҉iQ�O y�@�<��ԟ%�R�^�]��!� {��u"��A"k����b��J�R�<�� ;}�t �?�
�R��{Y�Y�HO������'Xў�'�B���'8T`Y�/!��YI���l�I��,UQ�)�)IQlў`|�1c-wl>�'�4�E��0 |2�o��&PX�<��DV! ��篓)E��� �@!2��8�e^�T5�P˶�\�q���%��j��4KQK�,�Ȅ��<ʓ��ą����j��k�n\��%)~��iW>ܺ��[,|���G�=?�^�?�EmQ�S~Z (�ںHs
��bD)T"<)��ԟ��ej���PYCU� �������=&v��U�����Z�t�]=$>X�Ӈ ��'a��Y0+Dy���5�S�O� �Ū�/S� �
��nY6�A`g�<��O����B&B@�#m\�mh��> τ/#p�1��,��SU�^f�|���)�Pe�r獊Zv2 �o��v��$B1��*y��B��T�Yjc^T����Xt���H	��Xd�BN �v�А�u�ݓh͒)�ON�#��gQ�$Q�	�,��b��d�_p`���cB�yO��(2�H�#��q�ē2�N��e̋�������\�a(��F�I�5a���(O����2��`�;Z��I'�ǴJ^�R&\�����Ie��`�m��5�eab[��3sN�6�}hO*�	����@��q��l���)����?mKP�ڵ9�yA� &�Ȗ�'�I=BY����y?xC�&`��iK�T�M��YT�(
�j_8-o�Y������"E��� +����Ύe?�g�'�R�B�f�4�Z5��mO"u��b�$EI?�Т-��� e>!j�m
d�HtŀS�	�1xŨQ8#Le���8a�b�1�3� *�@R(I� X�pDJQ#R��� ��+d�����-$�<�S]Ұ��$8�ҴS���&_����4>M6D��'�R�'8��'��S]���u�FY�^�)�wE��v��3"T��>�͜(�z,2�l�5E�d�k�	~Z剒1��q���/�tHJr� 5������@�'��i��x�]����X�"tZ�r/� Pܰ�Dԓ�y��&
%�@�
�-{�D<��Ɗ���R�V�0�'i�O  ��ܕk��I�s&�6.6D��3]�<`&�޹<[���C���s��#��'�
����N��h��F�^F��Ť0C4��<�O�`����y����Cܗv"���F1Y�(��`Ϛm�Q��I̷]�"���wG�y��ÀMU�$*m�	Q��� w��'Ja:�H>!�������:,�t���_0k�
&^�z.B�˃��Xj�90ԉ�?A�d&�@Q�`C���0HVd�b|PV��O��3#��Od�ʧJH����h*mAb�Q#;�l��F�<Y�t@�s+d�4�W��.��ȑ�D$7qO�S�y��X07FdE󢣆�|�D��P����I-yڈ�a�rA�J� �Ɉ�M7�	��|���95���J����~Y$�ʌ{B�R�l��N�O�Oz�@�&�VUBWmܸ8��0����+t�xa��fE4U���ݘ1�p�cD?�,ɣCI�-w���"�
-��Dłz� �v�|B�s���ǆ�M��#����~���Sb����'|��a�Y?[�6P�7���_���K<��I��~j2�{���k�zXA偟؟��.ә7���=�OWB����q�4��8A��\ɇNB�� �DJ/<���fݵ<h$��3g�+2ͤ�ʧ���[?C� &.>4 �jF����.%jŬL��x)�o����e�?�&�نF@�ū�J���ꜨY����=qqF��u�d3�'WE���"eF5M�LY3�G�<8�tpQ��m�fU��Ä�HO���9�4��wQX �ʃ�d��e�h�2��Z� @*<�JJ>Y����'���0xZ���Z�(�{a.�h�
q^�	'�8"lNE��a���MI<ɱ�( �.Y�"�h����nǦ�(g�>���*�)jd�G5K8��^csȥ	�H3o9
Qȝ���s1�L�`t0� `���I������[�)�./��=ʕ͖SR荢f/Y^y� �OLH�3���$�Vx���[���y��2�!D-��*SZm��ɝ�M�QX�T��b[~�������g?����2��g,N�UC@��J,����-�=>F�㔩MD�p�<���
�����5�&A�¬C�?w,P����=�]x�e��~b�ڗ�?���K?�T��}��'�&��~0�4qp"I�A�2����ӑ2�O���p�����J��ѩd�峟�ݭp5�1�Ȇ2�>-�2	��U�z�'�|Xtm2u+n������h� ]# Ո���T�bA�E@F�2��� ���Y�T�b��>�d��P�+#�� s!u�l� �ȗ����������5h������e^�@�$��M����xZR�E*d�ʓ.f��gy³���B؋X���`A��o
Bd��FN!>����A\@��<���/�Be��>�tPsb�X����@M4ơ��X'�~�O��?i4u?��I��'ފ�䏅+m�`2ef��'K>ٺ�@��;N�O�5��ឳ��������2���<i�ˋ�Q�paH0,J
,i�h�ń]<����!�RaK��P{y2b#���)[:���#�P���U�Bl�YFѤ,��;��;�P�*�.���?�6R�����w�.8G�C�\��+&.�8ik`�A,Or����$c������K���ܟ1O�EPW���T��ہ⊄]֐	a��Xd̓V�cشj���}n�?Q��)I 0qY�n��gTl�5+(�+�Um&�Dy��'�l�1#u�ISԠE����f[�O��p����R4j��~}�O �}n��p��#�;<���!�%�����V))�����ܯ4n����떧<��'Jt�X���*��h�2I��I��5yp�Ţ�����)�%y��N�.^�9i�<kh~0���_>vX5`󢁳&Q�������aӈEc�S���u��A4�=%�TL˄�+� �@�("}�	�aր `�BA�u���L����'�<��Y�Z�P�9B( 74�c�3�	:!G|��;p�?�Ip�ݮ	�(	��ě%�V���hٻD7��Ă� {0L�Gy��e3V���`i�uavEn�*1k�"��2�n��L7&��`㲦"�<���	X/9�~Tc���-�\����C"�Ot}� π( =��UA�9R�pU�x�Q�fXD�3�ǡJi �WdB�?i�Mԡy�z��{*��9B0�ؤV
`1hЬC%��ysc��l��uh��%lu:�R��wFH��b�J�F��Q�=�OX��)Y�p��%@�1/����Dſ8��'�^m{���?��0!�.Cx��R虷bCnY��j�;PQ��p�C��7��8ҥ�����R�.�bY
֢L*F�|�PD��QF��� �� �ʥ` �h��RL���睓w��UA�$��iTpѣnŻ�49{ I5t��O4�}n����@r�T/[��9G�(u0�m��D�*ۄ9�c
ٽ=l0�@1<#�'~l�1i�(A~��"h�f,үOD���d��&`�D�-���&_a��xԂ�&`X��bv ^P�r}���O�l ��
&��a �7�M;��uӀ��?�өGQa9��$$�]YB)��3��A/O<��sm�Tf�6M�����6�i�A��	W���(�|\��H=�v0� ��p�j��Uy���u�4��|�#X�r#�ͳd�X$x~,�#m�����)3���D���i>-�'e���y� <�g�ʃw��HFM�{� :��'���'T��'��SN���u7D�1�ԁ����̠�H�I� �Gy_CԀ��'CL��J�A��~Zw/�`��w
�R�n�>K\����d�K~Z�
�P�f��u7��W�B1
m^*,��!����S/6�8���� Q���#2Y|��3�jî#����?#<�0�L) fM�t+�<rU�T� �oLE��������҇���4@3&q�?a#�R�w���:dd·fǒH���<v�*����6])��'���6K�4�:�SOH���r ��+ s��Cաup��֝<\���a�!�J�>��xt��#}�X- ��'#�<��� � n�`/�`/�x	�I ��2^��˶�ė7ak��È�|��$�"E.J�	!Vp��	v�-4��R�C'(�C��|�J7o�����@w�РEK�E�:�2u��T銘rkK�v������,M���,�Y���j��^%�J �֬K�)@�`�'=�`k����p~Hl��I+m�Fy+q������He�̈́�Mk�E�/�.�В/
ya��ڶ�As���RM��kJ�n0�P
bθ���z�$�>���S�0=I3��Tz�X�$��(�ĠY�ED,H=�1ӭ޻!��(���8tk����&�T�2K� �JQ�f�$l�<ـ��O��=�� ��-b�6HVB���Gh�9#o
]�"Q�V��-XߠuPWK%�	�Njj�r2N�4N:�D�����0��'�Qq6���N!�#'e���/O2Q;�`�5��� ƗH��C%%�Ȇx ��Y�o��x�B�I/K1�a�"
?I=ĥ��{���+A�ҡ�l��z(���7?�*�4r2��b�H�Ԡ�)uࢀZsC�1'#X��$J�(�ڸ�"�Q�4p�ʇ����-7��m��p�T���7ʓ�hO�Ο�Q����0��.~�>��#�Zv�x<���F9o[n͡���X�Q���!�J=6xx=���V/�(��aߟ5���#�KCm��,���hO��c6��đ�O�:K @
��C�c�)	⬖=�v9k#��*�*c��r�Z�
�L�,������᤽����YqF�J� A6W~��#5˓�S.˓�M�A��}V,-��Eɾc�%Z� ������O�f��`6m"D�	�GC fܴ*3!�7��a�"JԽp�4b�E��r��|�S�'e��> 'xaQ&De�R���'S!~�r�@�1!�$P� �	]��4��#n>aS.Tb�+�ôj�A�N�0g�K6F^R��O� r�<9��4��S�IP= ��C'cҁ�@���S�����32��r4*-�#ҁ�D�Ё	����dB�PEnV<u���GA�V��?͋���6=���5�i��4%��6��@��X��yG��y�po90B(�l1�"A�n<( �S
/G��(�{/0AY�Y�a�myV�T��ό3:!��p��$" [U
'W�^aJ�;���A��� ���&x|I��ĜC8� `�-�y��������	�<��fB>|�DKqA�!h��0�����3�Q�0f�-~����?I0EѶ���Q��@�d!��k�e���lmڿ~�Rʐ�'��?��-���j囚<�Xa�K�2J.�S�A؏о�˧���0>����5H�����Y#sfh�i���A�<)P'S/�
��o�7p-�Y��z�<�CG(j�<d e"B>I�(%��j�<9Bo��	)	p���|����b`Lg�<��l@~E!vL
��e`#�\e�<��%��nӐ)���_g�X��b�<A&$�O��%�e�s�x��Z�<��A2|8g���fּC�`�<ٖ���U�֤����pD@˦n�@�<y�ǉn����2�
	�h`�6n@�<ic
=}�D���- bN^���EPb�<مk�.o@@���0� ���W�<1��ʿ(q�4��	 
$���%��~�<�K
�w�@�/܃j��Y{ӡKs�<���^�(��@JҤOnD�ȓTӼa�P䛫Q)�R�ק6p��ȓ-�N� "�V�U ��)f�B(j%����8FbY����3r�z`��f�<@�(1��\<��[F�E!t !eA=
�r��ȓ(L��rA�?#ܶ�J�G�,4H��d�ƩJB^
IB(ĊgC.+�x��	߰��r��i��p�!��+�X���$�2H[R Ƚo|N��	ȊB���2�-���������$�X)��"}|�*��V�Fv^����/>�E�ȓ%v��F�ޥ�<��k�}Z�܅�	AD���AQ+}��l� �ށ)Ƽ�ȓ&E"(�#�	�x��zbڇ(�v��G$D*#�ƥh;lQ�BM�Lx��S�? ���h�?5�
�2���Z"O����!]�V��P�mEt8^Ta�"O"��J�4|I�,�6TM��"O�؊`��6�0h�g�L�D�ԑ g"O�y2�cY�2{�4 �hH.!ƌ�6"O�D�$	���s���-��81"O��c�[*�0��P�S�"��<�"Oވ��(�{#��"��?�~��"O�S7�F�#��#��Y)Q����1"O ����s�Ll��d˩�h��"OX�H!���g��&C�/�r�@�"O���$ '�H����({����"Ob����>9����L��6�-�"OV؃�#v�A�a�F&k��a�"OLѥщ���GJ˼]P���"Oqa �E�[� ��k�`H�"O�+��V,D���A���h�z]�"O∃�dJ	>�����X�NCf0aB"Oĝ��*��R;bi0Va0|&к�"O܅�s�O�dU&�Z�@�u�l��"O�AX�qqΝ�����tA�/I�!���Dc����G ��� 87!���,Xģ�`� mpP�.��@�!���y�0$S���+�4��$[0]!�V2H�2�j Y��m�EQ	]K!�$�%}5�Y�wb0c�
e�!�$S�F��̣�'��`�4AzgI�(&�!��ش@�v���#���l��-�P�!���TI"h�
<=���A�¡8A!��IJj a ҧG9)���iW�6-!�D�3:8scfF�=%�Pq!�>7%!�d�W�z���m]�4���R�#�!���#������T�t��%�H	�!�d�!"�Ĳw�6��`Hdo��L�!��A(p����aJ	s*��24�.E�!��٠_�V�1TW�}8��tˋ^U!��̼e��q/ޯg�t� cK�qb!��K�Fᄙ�.ґV�8�@�P�DU�{��d�*�f�-B�F� �aƬ-?c!��J*n#���@OԿk5��IT+�rJ!�^T�pxK�/�/i��4	�D��B,!�T�|�li�$ �v�P�f�$Z"!�$��0�b'\.e�L7�4
!���\r]�$b�%P�`�w\�-�!�R�|�ЛDJ�.��0��D"!�7�r����P'jq�q@Ԫ�!�,x���G*E"J�r��'j�:Qk!�W�tV� �2h��Pȇ��0��ċ(L=�	��'�.�IK7���yr��88�.��Ɉ�G�8��	�y�/ߙV
�����H?D9��z桘:�M��'��L�g��7� �3��^��1J��D{��g�/n�Kɥ\��ِO�v=M�ȓ�|��C*(�)�ÃZ-�X�ȓ&�n9СED�X�� Q(��ȆȓSR	��k�|�J٠�G�w..q��Y-l)��A4"3�1��� �x؅�yh~��̐�g��%b�	d�C䉆.���2lO�\0��R'VB��۟���B#hh�@J�F��4�/�>	��db�m#4�Ա:H�h�@V����7�l�;�V	o5���
n��ȓH�v�rsMM;l���Q��v,tEy��'��A�!3
]�g��lI�	��� ���t#?l����Y�:����"Oʥ"a,ȍ vdSv�ɂxDA��"O ���:s����B^�J�[7"OŒ��OC澵��+����WB֠�hO?�	L�H��W�7k�����Ahr�B䉪l�)�>	�|�؂*A&Z?�B�<��2��	_���P��W�~B�	�=��qBK�B�����[��rB�I�F���:��!��r��X� C�I�/5�`���M&o�I��i�Hi<B�I�i��K@��=dh�a��L#7�C�6bx�!+f�I�c���D5g�~��D ��KV�R���L������!��7a~ҴiN�X�� YD@�\L��À�O!�
�Ht�r'�v������"���`E{����!+_
{�)"�F�/�L��g"O\���?ƈx�U�r�� �d"OZ��E�M�������()�L�"O�6��?�P!�7�͌��Q"rm-D��1-v
�s�j�b��A",D�l�6�( q��
��$.��S�'D��k���_טU��,ˑ0Q�}`�
&D�pp3���%�)�Ʈ�l��R1�%D��!�Bç\�(��F9+=��)'k9�$)�O�pՁ� 1悘�SŌn���p�"O&�ޤ����	F/f&:9�p( D�|�7�Z��0@�&ؐ�t��i>D�(�Ad�2*�d�hرb4�<D�0س-�(u8ހ�B������ń;D��1�����m;c�'R�`
ç:D�X�s(¨V����J��Y�0�`��9D��C��ۦźV�޳na<�Ҳ�+D�(��H�IXrEhЈ0o �2�*D��CG��U#6@[��Y�h
���4�,D��e
�Y2�r�J�p��)��5D��ƀ�yB�P�FܾT7�h�.D���"��7-���P��=NTm���-D��Q�!�A�	��17��}�"H/D�K%�W�J�+"�����"�	�yҎ(shHȉ��ڪ�Q铡�0?Q+ODxT@�r�(l���kh�a�v"O� j5�
�H�o���Y�"O�(k��W��#��@A�LI�"O�9�N@<	;: r�G�(.8���"Ob�Ƣ�5$<$�(%`�
?*�ͣf"O<y���5'�J���͇K�`B���P����eK��Ͷ/�f��DC@�	$pB�I� ;p՚T�ʶ\�( iiʔo�B�	� ���T�İ"؃��1}PB�ɡ%�I�AEǸcA�#D�G�4B��8��aK%�����kH��B�ɝ��P@�W%0�5�U���-O�C�	�|�T	��^�d)�Qd
%ps��I{����A��OUH��W��!`@�"O�=��e��Env6f��"O.�V�M��v�C?�h�x�"O���&D�+�5���A�"O���/#`6Ċ"�H-0a\�/�y����b\Ȓ.g�a�b���y�҃� 2Ee�
��mz�gӊ�y2cY!1�l��a�4��-��-ч�yR-$=64�#���2�\)�Vn��y#G�0"Z�w��"$R �aW�X��y���V�A�B����I7!Д�y
� |���J]2{���Ì$�:a���'P�'�5iD�N^��#��H8`Q��h�':�|G�toL���P)l��'v�����Ԝ0���ՏԌx�D@
�'� -B��h������o��	�'����Ɩ1�x���>�1��'ظd������U���J��-O�=E�t�ؔpi $@�j� O���k'B���yG0So8I2BN��M�(`����y���20��� ��zt���,��y�DR �%��0 �t93�Ӕ�y�6/ �(�7�8H8��i���yr�	]���9d*B=�j�HӦ���y�d[ �f�	\#8�ۧ(��y�G1O&�ɀ�ҷ�|3gD[0�yr+��9�HԸ`+�~.2m�q�܇�yR��N+�#�y&L)b���y���6��`��K�y:µ�aW0�y�f�� ��aE�4sk�q�ʐ�y���Ib�1m�	iLe���D#�y�![�?xQ�P@�;VF�$��d��~r�'�b���BR�/!��!6�>�>̋�'Q���wl|�p+�8��p��'�����NfP|��n�*���
�'
��I�(֟CL��F�U
#�m
�'(V�{�AG�>z�y(ř�P�	�'���aG�=/�d�`���`3����'�8袱fԓl�n��
&.˸p��'V�Hpb $%2�h	�Ά �4Qc�'7�p2�Z�z�P��D��x�J�'pnI���^�UP1� 	���L��'�ڽ[gb�(O|HZun��L�����'�M��k�ح鄭Z!-݈�'�0q�O't ��TG��oF�1D��d���p�Rd��#=Ȓ��0D��4(�=�剌�ڎ���*D���0O̪*�X���ɨ�leS�F)D�D�&Ԕ$O�Ҧ�<}0�3O1D�0����U]���Qf�I�6q�"D�(��$� e���D	�U���;D��c����)�(��ҽ|a��cë?D�$�R�C	R8�	����W�����.+D�p�e���6 ɷnO�9��l*S�>D�"��]�'����X�7�����<D��)q�Vp�dɪPMAm�ZU��'D��2��8{�!���^,T*��38D��Q�$D���*�_L����4D��{�&Ʃ4��Ua���7"
Q�E-D��R��N��l(�5���0���2�/D�HKB�*i'*@T����-D�蹶ၤ	�:� ��D >,��G D�x��W&9\`��W:9 6X ��>D�$g�E�޸p#��:0����8D�4�go[�r��4蔋�)��)�K7D��8&׫a$D�*J;p�a�*D���`@�0�!�{J�ط�(D�d�C�9k2y�cL�u�B�0r�"D��`7�0(��T���:��0VK#D��� ���O�-cV�	���Z�!D�k7l�/��e*̱,t��F`)D�L���ٚ6vu����>�2�&D�8�4��*g�2d2�#,D t��&D��YҤ6<����Ζ�v0L�V�#D��C �G&at0�D*J1&�9k�>D�� ��	6�ͿV��Cg��]-����"Oځ1�/��)j�!�"cl�C"Oؙ��j��|��yDaSVbЀ��"O������"Bi����T`���"O���
�jÆ�Y`�;FXp�""OL������b<3!)Ԭj��)a"O���P�ѱ`۪}��HϸQ��A�"O�9��MITprxГ&],�,��"O��D'�$*�V�2��* �*�h�"O.�:A��v�.�䞞Y��-��"O��y$�Y�r㴴����)i:�"Oı���y��-�cO)UL��q�"O ��Ə�����":�Pۀ"O:���ʹ)%��3m��%�"% �"O�,��#V� "&\Q#IS?�2yQ"O���r�Sk<�Z��̞4��qi�"OB��%	����!�c 9im����"OՋ� $V7�x0cP�5eJ��"O��+qf]3�J��Q! +;<���P"OČ�d�M$N�R���9<Չg"O��Ó"F����@�,�z����"O���CB��v�L� 0�1n=bu"O\�� @	����K�!5�m�"O0�%�u��q����~��� v"O�Œ3b�2�����"5~j��7"Oؘ��̖MQ���,A(k�f��"O~#( �QRf-s�J0梕*f"OtM�C��;�h|�#j�Z� ���"O(�w":O�lI@�ͲH�ڼI�"O�-�a�\.x�X4ҳǌ����!�"O���Հ3oYH	h-�a�f�RD"O�L��X4��7! z��1�"O.B�l��>z��`ӘYh�J�"O�\3�g�()!�p��Yj�X�"Oz�@�� t�8�U��
�ȕ��"O��$!���<�@�U�u �قd"O��Z��/Ȁ}� dˑo�Bu��"O8x8�O�C"���bآ-��R�"Old�A��R�v�#7l�kL9x%"ORi# V6+;�S�˃�qM��z�"O����`9�'Ԓ"����"Ox@A�юc���Y����bB [�"O���B2Ȟ�B������T"O�uc檋*^&�t�Ӟ��hI"O�H!я����8C�6I�`pR"O6`a���-KxU��-�4�D"O�Ta
��$*��Ξ7T��Q"O*����-Id��eEG�A����"OX0�䊟�JJ�x��v@�!"Op���	/O&�x8���m=h�)�"OZ	q��W�3���4DDD���0"Oha��n�i�TXU�5Uz11�"O@�"� ��
A!6�׹(KB��D"O���@�^,�Ċ��1&��8G"Oݡ�a��:Of9��m	�"�"O�t��B^�P��K��M%�p"O�=	�f�/`�B�)p��5�E#�"O~�`p ���q[���j�Z�@�"O����A�	~f�	`Q'�${���"O��PK�AQt�#4��D�"O80j��M'#�Ӧ�.%��-��"O�T����^�fT[�OG�Ⱦ	ss"OT�7�ϿB��*���=9����"OӰ��;L{�)����2�"O� �!�D�^	)��A(�"ϖp�r$�"O>5��۱Z,���`��j
`4��"O�\�p��nR�[ȟy���"Oz��G �
R���Qrg_6�H���"O(��"F��&��p�G�צ`���@�"O�mK�g�8
 j�L�9u��u5"O�9�@+ƥA=�) ���.z���q "O2��r����d��V}2�"O��X匌;	���PGM�.	X�"OHh�w
�:,T�1�%=��hs"O�mj�D��B���8f8M�$�2"O<)a�/ƴa�8)�W*B��0"O�uۓ�q�D��(4C�Č��"O�m�@
|xh��Ʃqƕ�T"O
��B1���� �VZ03!"O�9���̢9�0�;��.1!D��""O
�9���6r-��[S�K"p�4y"O����i'h�)�M�0!X^�8P"O�M���NF� @/W[>�02@"O�����#��k�.�>
�h��"Of�xǯZR�d%L�M���٦"OUy�i�u�}��*>;�,p��"Oi"0B;Bf�!�X�8�
��@"O��Z`N�r|��d�ݦ,ʢiq�"Ol����� N�L�&Ǆ _H���"O	2cM�`.���F���qt�`��"O��QbH��V'4<��S�f�=��"O��!�4\T�f�hh��j "O
���Ȗwf<|ʡ��%,Pr���"O���G��$T!�DV�F�9@"O�Y�3b�x�ʹѓ� ^�ܼ34"O���/#�F��a#�$]�2���"O���¡���ހ�@]F�\��"Oҝ�#a_�Aʠ˖�� *a��"O � �B��M��X�PN�t1�"O���I�+A8 Ȃ�R�	'�	Qs"OrPz�!�L�Cg�ўt��)�"O�P��cB�	[���$=����e"O艁�("�t��u�7h.���"Oh� ��|f <��+�-;��r�"O���BL^oN$͊6�̍<����"O��WC�#Q�:|��g�A
@"O�>�b`YqE��5�K�&@}�|��'/Xw�G�vr$("G:��y�'XN���d^�V�eJ��׫zr�ݳ�'�r���+/PtqPd�m��9J�'�����mДevPI	ph�q&��P�'��1[ ���%��=����;2F6"O�L���@V�� �EC)a#�4yP"O���ąQ{����:�9a"O��tbR�e��PZ^J��4���y"�N��!��#r� 7�H��y2M
o�̑���8��]!NА�y��ա3+���S4Y�ƀru�6�y���&4����,��=�X�d')�yB.L�MKbQ�썞Hy�C����y��^� xA���iwPu�@���y�l�>+�RY;�Q8Zf�B�-���y����A�`��/��ɂ��$�yb�ߐ8��]S�۹|bHM���"�y"U yɸx�����z��`é���y��;��Q:���%@�F���y��Fna��*��6j��F��7�y��	N�̐��#hF����y
� �E��
�+��є
�.|�0���"OH� �"ef��f �C��t�D"O<\9T�����C�myhE�"O"�f�U"-�P��A� b�uJv"O��#U�б����&�.M�a�"O�izc�(^�0@�FS4K9�e��"O�1���7���"3��u�$l�W"OrA��)V5d��R�v����"O���˝+'H�%ȕ�@�Hx"Od�D�s(�d(֧	V�y� "OT9���#NK�̊c�I�q���KQ"O� t��;`T��%!_�:�<)"Od����5�D��o�BF�L��"O6��D�&���QE��g&�l�T"O����F�!x�9��� 1>(��"O�؀'A@ L�����!��7�T�R"O�(�c�R�>�8RW�L�l����"O�����3.LQo�	��""O.ԹS��b����@NW�k �\	"O�s���/PS�0�ۢ{��\�"O�E�g! �4�쨹�J�h�0��"O�ɐ��ɭH1J,1���99���i"ON��mQ�q���� _h�3q"O��c�P-_T�m9�jK	~�$u��"OD�(�ƒ�Ilb�X)��n<E"Oh�3���64�R6�[�S�:�J�"O�-ȱ�F�0x
́�'���˄"O���u�-R�d����_� dK�"Ob�b0 ¨E�u T�-n���"O��#��b�Rջ�mΛ\l�I&"ON��;C���2��04�n�B"O�a���9�ʤ`���5�N)�"O �4n�;_KΥ`�'�P��=82"O�L�W�E�Z���AG�5A��m�"O�DHs��:�в�g^�N�Xl[&"O�t vÍ�D6��d�  {�1K`"O� 9Q�ޛ$6u��{��+�"O�r�$��P���%WE6���"O�Ux�
ĉ�8�g!SN+�0"OpT����5C	2'�#T6e�"OP�)�a��6銌�tL7K��ie"O�݁ ���@E��Bd�T$̡BQ"O�|b�F֦~�LE$Lհ9�r��'"O�ձ4k�����J�Ɂ @�`��"OniS�IO(��0��������"O��!��t<���e�wt�9��"O����₾\�z��e�<`��"O��j��n�iB�6wN�<b�"O�X��5�:�)�ƍC����"O�Msc�\@a��p�̧L�^�`"OH]�@�\
Sښ`0ቀ+rZ9	r"O�a���%Rq,�3F�6oL��"O�0�ǃ�]ǼX��̕)�|�B"OPph3F�@���2�њr�~���"O�ؠc�w�~\!��&��XK"OV�x3&��%b@�]�pZa�)�y���<R�8"'�P�W��Q�tl[��y��4Q��@���$�:�.���y�'J�N.�pP�G�(�$��7�y��B�I�x"��/�D��G�.�y"!��|��|�t��u��ao���y	�Gxp�*�ᑡp^��h�Ӿ�y�kP����X��d�j��'�]�yb�K�Dv��T(�-U3<�������y
� L�DIS9��d���E�$��4q"O���g�	���QBl�@)�"O�y��=���Ӡ	���1��"Ot)�5�>}8c�N 3����"O��!�ՀL%"d)lټZ��	�"O�j�Ш@��4²�P���z"OXЋ�?`�RI0��Ⱥ'��p"O��XQ�Ͽ����,���j�"O�,ڄi�3L�DQ �ھƚ�#�"O�ē���^vŃ��ϽA��"O*�I �K�xKR0��Ts�L�y���2�n��CM�'
	<�2�LO�y��-v7��@F��U`0�K��y�Y?�����q�)#��w���ȓp�DC��#�y3B��S�>��NT:��!��)�`�3�Mu����i@D�SHcV��>/�F]��{B�ɡ��%n?"tHD%J 4(�͇ȓ)�~�HUՁd���7K_"n�,��i���P�c]���@�&��5Le�ȓ4�`�3�m�'[\0���,~�0��#�~s3-N"�d\B�͞#6�*I��r2���"B�R69Jc�\
H�rU�ʓT�ƥ�Q�oa�Uk�5>�C�	�K,̥r�/��~�����A֭N	�C�	�Ib��eLm�xrӁ�5*,�C��6о�a�.j*�2g-Y�- JB��._v:qBT��/�𬓥7t�0B�I�'c��Ȳ`�LBr�pEh�A��C�Ƀh:z]sA�"H�l	8� �B䉋6�2y��FV+}��sp*��g�B�ɧ`�"mR�]�H�2�`��)�jB�)�H�1kٟL�� ��:�pC�I-:XN]C��$��Y0�c��T@C�	�oA�%	�]�S���3��j��C�	1\��UH�m�x���F�U6��C�I'w�B�A�ˮq�Uڥ�ݏXw�C�	�s��ًwc[�\�p�q� 	jC�ɚfo�y��Eɻ\�6��.�_�2C�	�%U[ƁK�!��A �$�jC�	5S��Œ#��tm �0�-1�xB�	�c�vQ(ˌ��]�E����B�-A���r5^=���	׮�
8_�C�//��i���*(���8c�R�`��C䉖p���1L�[�n�r%�Q6v��C�	6z�����
�X� ����
_Y�B�>z�a��M�x��@��R!u�B�	q^\�GB�	�,}��\6��C�	�y�x�C��<���!�C�=-ghC�	.,��Ёr`��Y�����5l,�B�ɨ�@BՋAAX����3��B�I$4��|j )ݾ>x�I�uH�S�B��3l����3�	�v��E�Tj�W�fB䉨��Ր�睶N�.88D!�8�NB�2#���c�&�s\5� ��9@{B�I�v,N�c�)�G�����	�A@&C�	���)�0h���Ka#�xD:C�	(%5����B�s������ۛ��B�I Y�.��B�;��+$�X�^y�C䉟U�����ܔ��[c#�"��C�I�*����C��.y��[�f�\2�C�I ~P��rmQ�H�򔱱���X�~C�I�S�������Nw�lXd`�WVC�I<B����Yj��e�{�0C�)� �<�C�XiF��	�t�t<J#"O:`��/��V�b�Cc�S�U����"O*@X�W(m�N$�t"
-����E"O�D{W�Ӡ���Ra\���"OZ!c@��$q�,�����#��$�"O����)@�\�֝c�Ä&��M�"OBtC�M�px���Q<yƠ4��"Oz�ha�̦X8Ƽ@,�p�j3�"OF���돻6H�����:?�:""O�e���_�s4QY@�q�H:B"O����'B� �1�i�_ljQI�"O��P�&O�L�ksI9�v�Kp"O.h�D!��Н`����t��q{�"O�5�Ӡ_X�(ӷ��L�Zd"O칦
!e�f0�����n@�5��"O����J�"XJ|�:���(6��܁r"O��j����d���7q�-�Q"Ony9�Ȅ��ɻoD-nM����"Of����3�4��sg?����7"OpZ�芢\[
����&J^��u"O�Yz�)\#R���O�hv ��"O6���
��{�d�jTNҠtS�Qkg"O�q��)�b�P@������8%"O����Ĥ"��ŀ�	+Nn*�"O:<+6��
-�DT�S)��0�B<�C"O8a:��E�@"�X�I�%,���1�"Op��n�5}�`�bO *��Y�"O����%Ԇ�@$q%ǦK�t�G"O�%()=l����9&>���"O�H�D�&��$�72)�t"O.�����$q�K6�{R"Oz,��O<V��Qeas<�@�"O�Q:P�<
>���FVX�$+�"O�y:3�&��S'�+M,ق�"OT���Ҫ���C޽5��`8W"O2��#�߹`"�z��X��QY$"O �5������6O��d��"O�̻F�ي=r�+��.3&|Jc"O���`�,P�A��M:MF��"O�H��f�f�	�2`δ`h�2�"O��B���KA��Ro�"���
�'Π�	� (D�06N�}12�
�'�D�hR�=-������/E �[	�' ��ԗ�H�r�v���P��y�O�uAvL��f��r�KΫ-Z��ȓ0wnAr��y��hSV.T�.��B�9�e�(��`�	A�M4�ɇ�e�\�hQ�i HEYF°h���1�����NU�d��Pi���8�ȓ"��u�uc]�%O����&-i�TчȓiZ��p���=��Kӏ_�>�j���x�M�5��(AZ��IW�:J9�ȓk��y���9%r�p�F
.]�ȓ�BD��ǥ>�|h��
��L����ȓ<} Q�R�@TJ�M	W��4l�~��a�Ĝ $K)Q����$(\� ��ņȓR]��a�$�$B�y�Nȇ�L:�, �i������9�*|��Uz��D]�,���R�H��@1 TCc��\2����҇!`� �ȓ$d�D�ɮ�*�剞O:�,��e:�&��g*��У�X
�@���L�6%��"*���%�<���ȓ~o��	X.SJ�`��Ƌ�@���S�? 2y"���_6�ɉ5��6|5ʑ`�"O��HN+gV=�`S�:� �"O>���J�)ζ4з��#X	���"O�X�-��0R�y'/ٙ2���""O����O�>�T�cN_,�x�"�"OB@�S�ʙ_@,�p�m|��aW"O>� ��0�X�R�]�HДLK�"Ojĺ4NV�N�`�*Ҭ��g��Mq"OV� ��֕ �2}�V!CF"0j�"O�Zw���Py0+FWԬ�I�"O���$Hk���z��%��!�k@!�d*;Ta�Eɥ<����Fb��-C!�d�)1ZrAZ�	Bg�
�@�}!�ĕ�9�����-�?V��I'`@>^!��8T�h�k�I,j�z�ōT3E�!��|��G�׿��h��f�E~!�N�1���2u|���Q�!�ˣY������>4[�S���\'!��jJJ9z,�S\H��@�C�0!��&_��H9�#�#3���"�/#!�D�"�T�D�ȧ$���he�ȃid!�D�}w*A`ob�X+R�JB'!�DR]���pa[.F�"���H*Ux!�$��pY�e���<�KQJ��0f!򄙄fe4�ঋ��xa���߂mC!�d�3_K��h��A$t� 0��3q>!򄁏m��p�kZ�q����/ݕs�!��	O�e�Sh�"z����Ϲvx!���ZR�C�畾M�4��v�3lx!�$��Q�L]q�؃SN\�;��X��C�IcXL"&)�"~�qD����B�I�W�ܨ���^� ����bD��jC䉓-,4]*5�N�<x���dA6�B��/�p��1#Z�)~�"�b_�e�C䉌9=ti9T咽ab"YR�D\�hӺC��	Z(d��&
JR�)/٪#z�B�I�A�zA ���-.6ac��U�U��B�I�i�fE�g%��q�"H߄K�B�I5P��8Sbn�8@��Eޥ3��B�I>㔐C�*��
6��q��Ɍ7غB�	 3�$)���P?;���8����b��B�Ʌ;;��ƪšf�� �W6��C�	.̀�sSǓ�LD:`!�+��Z[�C�		CTr�[��?p� W��2���l�����ą5�~|k��SJ�x��+uR�
Wn��>=�����j2�Ʉ�<j��x%i>,���G_)zՅ�
Ѻ���,�H�.�I�A�#sJ�(���j��@ɇ?	r鱃S�
����ȓd�plAVG�&��!��aU�(@��ȓR��i 6�F':.�0T��)�ꅆ�zxl�ra�	@ �p0�zK�ȓn ͘s	�C�l�*��QN��Ʉ�RV ��ůR1u��B�Ǌ�y��9��@`���5mE�A��j��Ŧ��m#�u��()O0���&um�y��1�|�H�@��Tf	p�e��D2��9�ty*�X��N`uDEA����ȓ��@0%�6}	@qX��8P��i��l	5ƀE� aM5/TՄȓ"�`��� �d���78�`��ȓhl5��͇�2��hҢ���@!�8��E�R��g�Q�|�:9"�$�U6�ŇȓR'�@�b����}#�H

�H���S�? ��E�[� ��ƌ6X��"Oع��C�i\Zm�D�<n�dd
�"Oµ*�d��n���k���/p�t�W"OZ�ccj@?�jT�q� �7s@a"O�	�ʉ�H�˕�_D�ha�"O��$�G&XrEʺ&�:� "OBPp�*ܣeDʄ0W�W�=pA"O4�����J�c�N.YF(�1"O�@q�^48	��KЩ8eq"O�M�'I$.��3�k�+f���ss"O*� HQ�s��j��E$�d"O��d����p���9*�H91�"O�U�T��=V|R� ��g65�U"O\�ad�8O�Ͳ`	¶b��PB1"Oz�듋�/9~��f�M���ԣ�"O�����W�\>y�W�P�p�	@�"O��S!0s
`�Ge�$s��1�"O�y��)Jb�1!��:�
qqB"O�Q��Q�q�^��q�ʧB��t[�"O�hiDƙ7b)}K`�7�H�#"O�yZ�,Y$ І�H��:�r�ӄ"O<�:U�Z���1�I'G~T���"Oz`s �
B<A.�&?� J�"O�9�k�t��%�@f�VzP�9�"O�dH���8���r��L����"OґK�W�0���I�p��c"O�u���4'�,9:bK����@"O

��
�;�jht,��[�D���"O2ukf�
h�~%ف
 C���"O8�3 	�&Xƭ����#F/�!��"O�u*��)gH��a�UxTQb"Odh�� ��ǡ�!p�-hv"O��x4��Q�H���\/ki��"OD�f*��#϶H� yTBX�t"O��´�L��9��N(u�����"OX���M�86��Fk�2J�zT:�"O 0I�%�-;���� �#e����"O���F�`�f$oTr��2�/=D��΂�lf�Q$i��oX���$=D�L��,֦tyr�xT& =O*�p
��7D����ۈ/�K������	5D����hv�f�x� �#4|�*2n4D�����Gўհ7n�,��`r�.D��"�߈SȖ�9�^1J���(�(D�L9�#�'s	��[��A��s'D��s�%ױ q�H���
y����C&D�J'�Ɋ&�4a���31���	!D�dK�t�참���2̎eఋ2D��ʔ��l,�0�Pi��B�N1�$�#D��ZtF�S�� ����r�=D���� z�*#���o��� !F;D�r��T�v���	��/�,i�A�;D�䓢C�$)�a9��0yLԽ��/D�0����!?n�`���Y3}%Ʃr��2D��� kF9�T��K�rB�5Y.&D�ē���QMʬ��
����ڂ,$D���6
�:?H�x)��� ӎ�s`/D�0�bOU1P�vm���8�}��-D�H��猊"��#g范2�d��ъ5D�ԫG/�5*^]�#�I7\%�4D����jA0y"d`�BB�-A.ݨJ0D��S�-��WȬ��%�AHZ�L(D�|r�=y�f��5��*�P�jE�;D�d��aH/�$�s��3D�ԋb%D�� ��įb[h�S���:L8J"O�-�l�?zf@��@
� H� �"O젺�\��0]Ӡm�'R��iY�"O �#'T�Y������~�f��"Of�M�'v����#?U,y0!"OTT{D�d�%2�ùX�L�8"O�sÇE G�ՋQݻ�j�"O��
 ��1��j��A�PN��"O�k�F\s�N]p���5q�I��"OhP0�.��h�R��Bj�(C�	�"O>����;��KEg�/ ZQ��"On�+`(�w
���Q�qZ�%"OTځ)_4�]�C;Sc��"O�%BCG�D,%ʒԄ7KlY�E"O|���Gވ�|�i�㓦k���P"O^Y�҉N6\��C�CĤ`s"O���$� T�$3aD�J���"O��{5d��^���d��P��4�T"Oxɑu�ݜ}b� D��b�z,��"O�8���(� mKf��w�V��!"O�|{0�%B�6�dŞ�1�"O����-��L>��b�GV��[W"O���``�#yhS��Ƣk0����"O����NQ"!��U)��,�4���"O4�����-A�T�Z9��ȑ�(�H�<s"L�:Li�'΅ �BX�@��j�<�qn
�z�`����	������o�<Q�#�!|+�p�$�Fj�(d�@�<���H�ZY�S�6r�rt��"�}�<Dݾ(��T�;2v)@ЫFv�<�u�e��%;5��4�x�m�j�<�禐���h�G�8p�U�p�U|�<a�&8)� !j�)�vc��؆�y�<���_�1E@�@����Ԉ@��_�<	F˙�(��iY3��z�j�2�YQ�<�-�h�:A�S�/vZ�,���
X�<q�Ö�E�@��wKS"N�:q�`KCP�<a�U�O�(q�4%�����q/�q�<�t��(N(��k�&�>�4�cG�g�<fj�7RO��!��"��DjCk@f�<ᧁH6D�Y�2�J�}x�Q���m�<��J��|tc�$՞f#�Iq��j�<��,S�R�h!k��de���e�<���/H�*���":#�2��+D�L��/	�Ш���3_1���(D�P����,;��'��LEԈ�!D���#�7�\�b��çc�bh�*OhpۄB��p�&��B�-�=��"On!�qm��#��	ТA^�+���"Of\K�i;|#~MSBܚ">�!�"O�H��KU�E�dj�aQ�a
��"O�`&'���.�&���6Z4�7"O��@���~�������#U"O<�Q��տ m@9r2EQ�p��"ON��2eh�@zU�Z);�FUT"O�勀�#l\��ǉ��/����"O�� E�	�6��6Tl��"OB`��ܼGB�Z'�J�����"O�(�4%�g�Z(�mNZL (b"O�9��M*���9Q�X�"O�Pu�_�-��Ы�H²}��9��"O�pPC� ��]�6�ڇ��e��"O(�bcMT�h#x�3g�ߺ,3t"O������&���2��K,)!v�"O� @<�%!�#6�nxʱ�ƆZx�<I�"O��g���l�#ʗ� ��"O@��w��$8dV�����&B.�!�"Ov�؆�,�D��ce_�b���2�"O��`cפ{�y��cQcɚȒ"OR)�Ҁ��Z>��0w"@3Y��$��"O�13V��7EB�ELA ���e"O�AcG�*���ė�Xz�%��"O|0!0N�3V΁'�]2yLq��"O��XpN�x��]� ��<oti�u"O�<���Wؒ�8�)9���'"O�`;��L����C,��"OZ�h�B�D��?�:r�"O��a�K3RGĹ��(��8ֱ�t"Ot�é�"�V��%��:pp8�V"O4�j� $76<��F��NW�x)�"O�,��fϤBx�l`&�ʉW�B(QG"O�c��4H�rE��L��B
 �H!��� N5��*�.���	�w���Y�v�@�+դR�l�l�[4�Z��y�c	?Q	z#C�%O�$��蚏�y�bЎY�h]T/MO���'昋�y�\�]���W,� e���y�AG�~�.��UA�7�8K�Å�yB�4q�|�J�7f�]�*A
�yB�<#8��e��,�FY��<�yG��.�Ι��앝/�Nh���y���%�B)�W�M)'�\�1.׽�y"b	9"�l8�-P�T��逑,��ybB��"��u�ì�"�ѐ3�ڭ�y�K_k:`w�I�Ţ��b�[;�yr��<�Dɇ�@x݆�K7��/�yĕ w@�Bw"R�s#�9;�#��y�	�V��D���!����؞��y�L�9h��I�4��]Q#��y�-��a$�\SG����Z�*�yb��Z�(��g�к
�	�����y2O�V�z��3��Xr�e9׌�,�yBkNyUX�봫��>��`�5O�9�yr��2R���C�é!����f�(�y"*;l����%óB�V�nMN�<�'�T9C0����j�2�R�)���l�<�AO�e�x�r�'QJ]Ή���Qf�<	���a#n�{G)��'�h�tf}�<�P�A:Ir9���	�n�d!���c�<9eBO�a�b��>9�s��_�<�b
:i�M�uI��$eN�v�S\�<1���-,J��![�;���E@�<���_(\G~��CX;~&�Y�d�y�<��-R�\�amI/&����0mn�<I����>�2Ѣ�*�8�Z�Ĉo�<Y��A~�"��B��?e���C��g�<��ؕS\:���0U�@IC��b�<i�E
�t� eNT/N?��7G^`�<	�F@�M����5�,Kͦ�[�l�P�<Q�@�8n���Avm΁n�x��F�N�<1�J�h��d�[*1���2�I�<ɳ.��]oTAr�GK�r
a��~�<)$N\~�#"kLd0�t�Qv�<�7�Z�Q{��)�A�|�Q�)H�<�soU�#�����P�k�Ɂq�G�<aW)3�fk& ѿ*[�!�A��J�<��eV=L��(X�,�9E���Щ�O�<�êT�c���ّ2sC"� 1`�G�<� ���g�
P��F)νoh���"O�r�mPh ��Щʆ`���Bu"O�L v��0`���C��F�A�Bt"O✒v��U~Z0u�I(
�"OFuKw+�!{���{S�վ'���q"O����OV�e}��@�/U�,��d@�"O�`����iyP.D�L� 4��"OF�9�D�%-�t��A+ݎ�d"O\�	[-=��3��	HΆ:c"O��t�@�dx�Uɜ3]�p���"Ol���j�.�Z�:�ʜ�F��"O�0��F�9}H<A�]w�(sT"OĠ��k��H�L����r"O���K�1D�=(Ej�~����"O�q�5�U/C�Jq��B��,�R"O�5ʓ��9YQ�d�󮟏��I#�"O�}���{��a�-��{���I@"Op�p�蔼D�
��܊7վ��"O�0��(��Y}��z�$еl���Q "O�X�o�@m(�����bB"OT!��C�b�>ܠ�`�K<��"O�d�
�.l��䅙+I�u��"OBy[p)(�B=ұ�X�
`L�Q�"OP�C�&!|��'Y�G`qJ"O�k���5O%P42���/9��1�g"Ox��͕Vz��a� ֫+��P"O��4��bgRU�!m�3s ��"OF���F5��ĉ��N=Oqp� �"Od)��Ҕ
�P�s�hh�Dc7"O�\H�bU8jüx9���)Ȱt"O !����&h��a�P��0�"O���b�YKF\�B��;���"O��QB��C��Py�$wC���"OX�Ap�ZZ�f-#�G�G_Έ:w"O�h*A�jD���ϝzV��"O8�j4���Vr�u�B@.v��A�"O�Lᶿ2U9���9��ဥ�_�<9��|o��"���^wƼx��Ot�<	BK���`GX6fQ|H����K�<��g�?2�����]���H�E�<a��3[�n]���&G�#%�QB�<!b@Y.��0�kH��@p��{�<I��/�x(�#"��(ԀŸ.�w�<!���+M�Z���C G�8���_y�<aP�a���W�RA�e��'�}�<Q&�t�\�!�%
��IB@]{�<��7O4���/d��ːy�<	��!C���
��E"J,h���x�<�RꘖO�"X{���(�\)� s�<� T�{��Y f�<���E�h�<Ar��W�>���KX�n�isBBk�<	�,\"u"��M	|e����B�<��ˣ$���sB��4�f<�Q��F�<�0��6x�u[U�ЀD4��{ �
i�<�ٚJ�`� ���!5T�ZV�Pm�<��bѠYx`��d�RP �%KKO�<)��ͻ>}�0(�C�C�T��F�b�<i%GX��`&�Հl(!�+�^�<�r@�1�Bu��: �9ѱ&Nf�<��I�,W��Bd�4����d`Bb�<	"��m���H�"�1!\h0��Ha�<�d�TO�Y
/��h�4���&�b�<!Ю�1m���aQ 0f�"L{�"�]�<i�}k��!BÓ�� �V�<� �0'����"�J���.~�!"O���B�ɁW�Y��^�R
���q"OZ����(pu���N�v�.!i�"Ov��ҩ�)J6�*��fr��"O�����'P�8���1'|�t�b"Oz	�f���|���j"�
}& 2�"O���M�-8 ��`��ϝ-d��ڳ"O�MYtGeH�\��
+Xe�`�6"O���D��!2X�YBj:�T�:�"O�j!�����[�ɛ����˧"O���u�Ď(��EØ-~F}��"O&��0�cs�p�vA�@O��I�"OH͸��k+��ʓO�b�:�r0"O��3"�1�6y��n÷#����g"O&X#�C�4t2X��,	T��A"O��#g	4	�ȱ8�-͜M�8� "O��)6(S8�x`��
a���"O��� �4eBѠc�jh`9۔"O�\���2/'<���׋ZT|��"O�:g���{@!�'e9�h�"Ol��P�#�hc�(Ռl&���"O�sD�)9$��cF���$4q�"O��x%,T�Y�䅁��U��"O���b�R�ҽ�F�A��t��"O�y���9Xg2t�W��|S>Ap"O��AŎ!`����l
&h+�K�<�2��� ��v��-_�&���$�H�<	E��#h��h2艴��[�,Y�<���S7^:Zԉ���-8�+�f�S�<q�͑<���ΏۨA��PQ�<S�I�V  � O@�I���� �[s�<�+�9 ]��z�����7��(�y�A�2p�=�dg�N�V�ѦX��y��\��q��Z<=���`C���y���V�� �OE�5�j�Qa��y�i�X5��B��-��9 ��y�\�_Y�&�% �Dy�.��y�jKe�����@ښM�H��r)҆�y���1^~�K��ZH�4C�����y2	���H�#ш)qfp�����y�
	BJi�ǧ�5#5@�����y�`�<�,�P���8�3�oߧ�y")�o*�(��kT	�x�p�����yRf�7(����@�Ҫ�����BI�y���u=̬�$�_0=��N�'�y�W 0��h9weɂZ��&.�m�<I�¥ՙWaڒ`;�e+%ku�<���C��A�R�Km�-��Cn�<�v�
NQNȒ�ϔi? ]"�"LE�< �4B�*�y-�]x�G�B�<�ď�k�
�w-��l�h @OC�<٧���l�U�J����H�ŘC�<9���7%"����\�d`ض�~�<���O�O�(I�M#o�vt��Zy�<�㨑�+l}�0̃�8�`����QN�<�"��<�
�R�B"q� 0���J�<�q(DC��iG�<rj51���`�<Y�!ڒ8�����O��!��lw�<9�S'1t�l��M�#���@a�W�<!wIX�,hPr��7�t5��(�W�<i��A�*��EkC�,(�i���V�<q�ㅧ QG���Z:��h4-�\�<�@l�-������q�!���W�<�V ;@lQ�� R�Q��P�<� j`[�.�%f����八@��[�"O�Aʟ�\1qwDU=@�ޤ��"Or�7[-z*��3u-8��R"O9J1f�/3A@�ˮ.�0Ъ�"O�2��#g�@Xc���`A��G"O$�$�����T �W4���"O>t���+B���1"��M4��1�"O*�.KWDp�`��<���jC"O���u���5'ެ���
AP"O�;$�X�0���nEs�Ք�yB�;n
,�KԬG�!���A��y"�R�ԠQ(�Pe��,��yR!J������w��0y��y��M�diB 5ʄ�"(�y�u����ydS�2��\���:(��IB�L���ybE�]*��u�2L:�gJԧ�yR�� �NP�a���@yt�b�,��yR�ץ?f�up�Jg����E E:�yr��yZ�Er�f�"�z#
��yR�Y���Yqs�P)H��������y�/X/L���ă5>�̙&��yRmR�w��$��ݦ<��p���؞�y�jQWW:��7N;���g���y�	�(t�ɩ1�1P���-ֲ�y2�� O��(�'+������y���V�h����r���V`��yBǁU �;�a��f���%mG��y�e_u8p��h�!UZ��:U�[�ybm� TxH�3�@ȗM�\��I��y��̕x����G̓?��	e���yb�@"|nri���	�^I���7�yB ��4�����)|O$���A��ya��]ꡊP�A|!H� �e��yr�lݣE��r��܀R�H4�y�c�<�F,9�i��rTZx�acM��y�OY tM ��ɟfL��w.�y(E�!�z��K_\��`�����y��S�sN�1!0��N(d��']��y���Gc|� ��Y-΅�3E��y�LL�X�D)ӓH�X.4ЁM��y��2+ XA���7|"A�h-�y�,�!����3��&C�"M�7�֪�y"�4�)�(�9�R������y���.%������,�H�#�?�y�Á�0_�:�T�Z�8�gC��y��Q�^:�hBb�(u��]�u���y�f�%�����mY�m`�4�U��y��C>.,Up����u����_(�yr��u�B͚���h�f�؃���y��׍k�T��Ş1bU^��cm���y�(KI�~�D��]Pٚ3C��y�B���� �� +N�()���^�y�e�1?��Ԑ M�/�<�Ї�y�/]#o�Xh�j�!M̼���ѡ�y��Xm.��6Κ4l2�M�O��y�����A��?e��<	#a��y��C�8P�`�(^�:���É��y�
��@޸h  &��aL�d8/��yB)�H�%��'H ]G���*�y��aN��a`ς[T`�xC�@��y�ؕRZ���KP�d����Bm��y��,��x۶T
a=��*[�ybB�*J�ƅ�S�Xi�M�਍�yR�׍���0���+i���
�y
� y�6�K"tIJi9D��P�:�"Ot�r��Z("	������z`"O�T& ��CV����\�p�D�"Oh�:e=�v])�߷4��� �"O��&��!����/<L��"O��KG&� X���2 ߙ{+4,
2"O�=`�BXHT��Ʌ��,ANH�0"Opנ�r�<
�@�[��3�"O�dْg�@���C�N)_�M A"O}j�b��*Թ��ʐ�9 ^%��"Oh1+�Gy|P��~mh���"O%�C U�a�PҥZ�Hj�u{�"O��8s��4��餄H�<�6us�"O�%��-�f���k�nh�t"O8�r�l�? d\l14�ס�¤�"O�(�sH$^��@�aρyT��q"O:�3k�|I�1�T�
e��"O�Qτj�5X�i1OH�\Z�"O��i�ŋm� �	��WOTaB`"O��awN���z��(�v�ND�6"O��pI�_Қh��&4J�\��"O���FK���R�N9"0�D��"O&$ؗ �^8�� ���y.H�H�"O��+W�tL����3|TH8"O� �T'�3����c��R�H"OhP�sAȎr��������"�`"OBX8!ȅ�.���/��u�"OXmi �۹{v-#�C��Va*"ObU�� �����A�:Z&��t"O��Qծ�R��8E��S���"O>��O��*���9�E
>��y�"OU)�C��.�X�I$*B0��"O�L�H~�|����lD<i�0"O�qЉ2f���@���z� E"Od�
��V� 0��jނ��xJ3"O%�2��@R�4sC�[0`�t�#"Oԅ#�o��L�lY,��Jsި�P"O>�YB	?0�F��E��*�B���"O>�X�c.��(�JI�.�`v"O�u�q B�B  Y��%x��5��"ONL�&�=��=0'���8)xE"O�x�Ӎ��Wg؅��ԝ}�b�b1"O:�1"�b۪(y@Ĕ+/� Dp"O�t�� 
n�R���!�c6�H��"O4(� %��5�ցڠ 
�5����"O�a'&$�Ł$o�2f>���"O�EbUm�J�r(����q��p@"O���Q�+��!k��˯,��+"O�3$�݋>B �b)*�X��"O�)���5� ��3�̘�L�f"O�떣X�(*>���%��	�"O�%R��5%��2Pg�6m�z"O��փܦa�Z�+���+?i"�H7"O��F��,K��E"��U6MZm۴"O����eȝ"0 X�!�3,B���R"O�0�c[�?,�k�O�*(��h�I�h�?�kъL�r��Kb
�%o��"g 9�IM���'a���Q���u�6����'d�2���Iؘ'�$����1>ͺ���j�(A�&��'�>�s��~~l+C�Fo)�Q�'���<���s���$��je%�[WP@��v�@-.�!�dl8d�	�aHp:C&�+u���Ԇ�� T��H{2B�8?|z)�
���C��,0�x=��Ӱ1����gf\�&a��	Y��� ��CN*F$(��ƤQ�_+��7�i_ў"~n�4���@*��A�p��C�#lp�����!��?O�Xkg@�O=Z�I����E+��)��1�S�S /|0�B���.i�$�ާ~2��O���$�7<����(�]	 �z�MN�7��{��$A�.���`^���h��&:!�d�3�����{�,�Ќ�~��衂�'z~��E�GK��Ƞ% �fan1R�'�H�i���q����4M^&)��'EV(��O1	VH��oF�Z���'�6��co��lh� c�#ޓKX�y�+���)V��)��$�����y�M�0ʠ$�-|ի!���0>q�'�D�-&h�@��3���c�ԸW$�'D��"~��$^�ܫ��Բ���h���*sv�	j��h�h���鎔��ۡ#�;�U�a"O�Q0"��,1̙��Ȝ�B뀉
�"O����a��Z#��	��U�q����00O$��D[�f�93�DاH��ǎ�	�0C�Iz4�\B��: �P�g�a��C�	��������?>S��ڇ̌�M�$`C�4���<E����r�HO-4kZ��e"C0I0 h��fq R�
(�Xr��E�$,���'5��I��u4��V[(!��HA��B�I"���D�l!�)8G��B>R��h؟T��%=	���h�jۭ-4�(��o$�I֦�ϓ���ؘC�H�3�dd����D �A"OHE�u�5?���ڕFB�!9>Q�d�JZax�ѧJ��u�T.�%â8Q�����O��~
AmI4@����T#�h2��զ��#���Y�!��	m�p��՝t"��ȓa�t��7�-��������k@V(�ȓ܎q� �S8]�p�ҥ�U�4��^� �c$n�7/(��B��3�J���R~R���HDt��B.q<��ъ��y"lG�'I��A�
�aZ^�Ȋ���O"~RbIU4W�)aۇ=�����E�'��y2�1�.��� �0�Y�p���y���&�Ơ
��ʅ$�=����x�	�"��&&.�f��� �+(O���d(�v��1�G�9��U�W6!�d�$,<�Pt��k@ �#|x��?��B��L:^�̴�:.�.�臯D�z�ax��	o�n���ۘ]�*i����%|#<���)O�d�`/-\���3�4}
A�|R�d&ғk-���.�6���'֜O�~0��IB��=w�^aӉE�k� {d��JԮC�	0p`�`	��tW!�e�K*tIL"<�NU>)�R)� ����3 �BM���!D��{T%ם	bdC`��$K�6�����O�Dz��)זh�h+s�5Lm¡z�D����C��m4�fX�!��щ�
P�1Az�$+�����*~�!��L4����&D�(2�.��3�&x�R�
�y�Ԍ�c�"D�`16�ٹJ�$�g J�k,رy�5D� Y�,$eQ�/��r���pB8D�tࣆ
.e�8��I����8D�D�5·�7Ve��Dʘ)~ڜ�A+D���r%�1s�nɲ�NS
SJ���ѧ4D�PJ�M�28�����"�d$H�ot�t��ɧf��2&j�Z�H�)c+W���C�I�2~>M��"
�4f ]�!��,��C�I�#n@1�M� �$�`�T8fC�	��r$ ��iR,�T��UZP�F{��9O� |�iGb������;:�ɻ�"O,˅�[6!�DQvaφM,�`���%lON��R5 ��t2�`�u�T����'���F4Mnz�2I�.�ވ�
�!�N=OL��S��80�"�Q������;OX�26��vg�S&샥1�� �"O��C�!\�v�I�R�F
$����"Of�{e��pl�}�ףH2!�)��"O����̛ZX�K�MĘb��"Opd`c�!����]1h ����'�剂>�p��G�'`l���	ˎ1��#?)��ię �`a!��U� ��P�f�7 ��x��ɋv.&�� �U\[`!TN�7-�aP�'.��gEH;s�l\��cS$(�0h��O�Q�'��'��.�d� &8�cW
�/Bڈ��"O�y�5��`�ehO4H5p*�"O��DY*y�����)nQ P���'q�dB�/_^i�B�ٛzv���@��#>!򄔒9O����E̗E����Ə'ay�'qO���q	"NFP��)M�A�N Y�"O�%�EÞt(��Ei������"O�i��Ȇq�
9�͝A��U��"O�1�ń�3%; � @�b}�4���'�O� ���)W��(0����M�4�y��۶*p=�a@ʫCS��P���3�y��Ϩ!m��8g�6.n�P�ď�y"���"�"�Qf0#,�����?�y"���&+4�$`�8RJ�1�
���?1�'/�p���l|������5>Uj�L<��*�z����GOfT��]�=�}Gy2�'ǎ�G.΃/3.�p�� (���	�'N� R�� ���pU�I''7���'D�;g�Y)�Đ��bV!
����'�]���I���qb�Մ5�$�'j���$*I�Fv��Q���%y�X
�'� P��	ք<���k�@ν���	�'2`%P�&ʝUw�M��T��	�'Q8���/��N�
���=y����'	�yi�kߧ=0�H�CC�:s�v(�N<!ݴ�O$� *F@�@*`�G�/3��PG7D�H����R�,,
Uʟ�g���iyӂC�I��PI�����G��A�挝�B!*�ON�Oa�Q���Ɗ-R��%Aٲ`5�܄�K�N��셰0�!�%%�,(Xb���g��)�h��qN����������ɫ@^�D�'2�
d�#��%��)����^�	O�� �A��(�� J"!��M��)-ⓘ�"����!u4����Ej݈��`"O��&�׊7�� næ�P���4O��Dz��� �}!�C6ʈ�zl�1�7,	t�!��Y�,�����]O�*��i �Ih���'>���N�X4~-��(*j�mJCL��p?��u��������H�J�  8��@��"D���b� ������'-���Sc<D���� 5�ek㏅=W*�qz�";D�801��,T~���M�+�z�b�%D���`��!m,!��l��m%Z��@#D�<&�̺~W�\:�����=��.D���Ql��*�8�KF�Xad�ɂ(>D��: ��~���KF=tVUص$0D��v��L��i�Db<
~�@�9D������p`��AB­aA�P�$5D�8�R��(.�҇ ��4��ീ4D��6�^�9��h�����0�6D�� |da"�vy�o���"Or��JN�z�rX��nF�U~�PX�"Ot�tiZ1>+(h�.�(ux L0u"O�=�V�����cfM�,
��l��"OZ�j�� 3K�сA��0朁I$"O�l��+̸4���w�� �j=r�"O��u��09��˔n�T;3+d�<�6��r��\��'B�!����,\�<V���d+G*�I��Z���Z�<�C�eQ�鰱�	wĬ�4�IY�<�'胋?^"�
ȚY��da�p�<W��whd��H���!�!Qk�<y��X��\�T���a�����\o�<��f�$��x�WN�:�� �ND�<��m֙51fu0�]�f������Y�<��jE���}+��V)��h(�H�o�<Y�Y�o����mN��JA�<��h��=���1���>td��ui�D�<1v/��4�b���8�:%b0j	Z�<AAdI!?O>�eN�N��J�HZY�< Ņ�#�:�K���7��T�L�I�<� c֫B�D�
I�MY��P���j�<I�O>�z�*�F��C���eF5D��&ъj謩I���T�,�0�2D��x��Q�݂��6mX��=D��[��L.;���Sg��/��Q��
6D� 2p	#a%N�;GeÊ�:@*.>D��c��،e8�e�Q《��m�E�:LO��Ё���y��څ�ݐC˲E�'&�x���� H(����"O����j��B��=�rF��bш1�W"O�i �L�^��ب����r\�"O6ԳL��<D����{G�L��"Ot�Б���^���HJ!ܡ1�"O�kl��~��0QÃ�h��0"O���@�L0Q�t�R�U�!)P,� "O�Ex�'K��x�i��I��xk"O�ɷ�U�߆}�1H��.����"O��;`�ȦV���b�"xN�A�"O4x;�۔Z�����B��hɐ"O6q�L�$��)d�\�w�la!"O(T� �,t
-�Pk�6w��)�"O�4j�� $:I`��S��3D�����"OV4Sg�@�*4��uE4���a�"OH}P���"x�kD�f��pG"O�	�G�O� I�,��C�k��A�"Otム��#9�Ȃ�B,X�D�S"O��q�$a�n�"`�s��ag"O��*�Ǆ	V{�Mr�/F;��9g"O��{5��'D�LRQ'��+a9j�"O>��uf˔&N�u���Q6"J���"O�Ȉ�� $>L���@�]A�"O��S��W;
�5`B�%��%�"O<�Ȗ&DV�T�S�+��1��"Ov���ꈂ1�4�5�� .�	
�"OHmPq��V�"�E3E�
�r�"OPh��-���Z�DL�v��5��"Oh���	=�dU���IR��H�"O*,H���-~WTi�Qk�'�@���"O0���ΌN���0����o��٨U"O,@��������J� ��K�"O����Ht�VUb��6Y:�"Ou���8,뢱�f�Z/	���"g"OD)���0�H�B2�΄^�(��"O��խC�?�6|��`�U��:�"O� ,��.�4+�T	 A,Ƚj�Ɣ�B"O2�Y�P;��a�#Ͳ?�T"Oq�̐<pA��1h��=��"O����!ؒ?(ś�ԼA�j�3D"O4u�$��>4?x�i��V����&"O�uPal��Y���)8W���"O�D��B^U� Ir#�G5\\1H�"O�|A ׳M.ȸ���<:]lM·�'�^�a�C�xv�ܒ��O A�5��9u�t�B���4Ԕ=�C"O�p�r�
�M����}��� 1���C훐����qP/_,XE�䌕�*1 �x06n���aV�)�yª�Vw�<J4:d��]I@l��t�"�AE�I�E�K��^�^�kO~�=Y�,ە6�4EX3�T�*tл�/Y؟�3�D��)��q)F�x���L�}�@�b���hp�Ǭ��P�Ƞ��	&�n,KF��W�䵉B�;�>i���fֵQu�ޚ+�2��qO�'�l�y�+�����ؒ�C�{� �h��(D�0! �0-oJH3����~1��z����ɰ,mNL�?Y��?�l� M</��cEI�l�<�3��F
4��ka�&�����'|u���Z��L]q�0�8���~6�`��b���'c���'7r�s���6Q��y%ePb�壌{r(�1�ay���
r��jQ�Y�M��cF���HO��i@�%�'9.�yz�'�i����5 ѣZ�b�i��F���L�f]��1�D�i�t2�!Q���˸9��O�)I�)qOB�&kO�| N�6x�p����IrJ��cm��	0�yQi�J���'r�A��OK�I���'�~2M�"K��̩����,��Ĥ��>IR���~�U�Ԃ�`q�V��^h�4cW���'�n�zݴVG�<�S�y��%�'� г E	[�#=�r.��ը����"��,5��C�&Z'^W� ��.@L��ɹ��S�O�p���EȔ<MH���ۦЃ�-&@!x7�t�"~n������`Q���Q&��-h4�(!=�I��M��'���������N',�1Rui� ���PQ�h1�(+�hO���d���'6���Pn�����O19ŖQ�OڀFzʟ��	�L���8H�c��cB�
�UO�a��&�I|����"
�
�����H���w�&D�(���N�I�2@�C]��%�s
9D�`�"��"��Pc#�}�xU*J6D�i�J��\Ȥ���B�'�.���)D���Ď�9Op4����@�n$D�<�c�
%UT�����4pl,����&D��{�$�-Jg�a���� 3��rG�"D�L��
w�DJ��n��S�� D��(N|��ݸ�����Nȋ�L>D������o��w]'	�b|��>D�� ׭�ߴm ��=p���;D��a��"�~hhuC��y�t �-D�P1@dM/0�|��Ï X��r*��p<Q�G^�_���W�E�o��t��,�_�<���m'\<З�X�e�&�c$k����V��Ȟ�r5��� Ó)X�
؅��_ܓH踁f)֯K@e��hM�~��"+hը /K�DU���G)�@��;8
�A��[�+�̻���8N�h�ȓh��1�i�54��%�D�?V�̈́ȓ"��d�:�b�2���,����e������ ����R'��LJ�Fy��'I�<���I5�,Ջ���
�ʨ;�'mP��L:-��RN�'<��aA�F5$�<[��G�W�h�#鉊y��
fD/\O�b��'�V" &:))f�ƈנ$�3� D�h��O��7�x�i1�Rˠ�Z�K!�L���'B����Ъ�b�r��ڕ+͆M��v�&<Zwm�o'�tc&��'�v�Gy���� ,(;����L��:��?v6@�˖"Oޅ�$gu��<;��)���#"O�`��O�R�����-	V�p�C"O-Q���&5r|���	92�jG"O��enб��q�&R,\@���<O�aȝ������t	�
ZY����^�B8V��c"O|ų�"ֵa|��h��Z-w0�<�"Ox !V�*��r����I��"O�����0F���qf��S@P`""O����T�g�P���һ.h �x�"O��t	��@ꔐ2�K
N,$�"O��9`+2(DuJ��]&j�,(�"O�XC�	�9��� !À%(��	��"O�h��%Ƥ,��pB���\��䚷"OXt�pΞ"5��K�&z�`��"Oj���.�fv 1)��Q{�<I""O�����c�ip�z����|yצS�����`�O`�2)$��ت$���Q�4	�'{pdb�,��g�СDa�N���˃g�&G����I�Jҵ�4��?��g�r�֐[$�زt}^�Ff�#Y�T��	�"W��Bn\C�<��"i@�g�* ���;h3�eTN-��j��'T IЂ�+P��q��� ��T"���� Y��AEj�#�Z��@ _�K&����R$�h+"J�0f����M�.!�6������5{��p� h���?�D�q�Q���&�~���G��h*dg���h�1
1��ط�˾6^!�$�X���C�v��1*A%!G���%���{0�Cw(\�R�� T?�۠A]z�_��i����p
W@3�����	-W�4�2�@�nr|1+V��4�d1��B�DlU1a+�2ab�r��Vh/�AAP�'�Y����J7�� kKSPV�#��DE��M���^�N?�8��k��PVZ� ��\D\݋��B}čiPbQK�n��'	�����]$`�,IG P�@'�H���[�]2�a�p�B�?������$a��y'n�CX�����vg}��NΤ�y2��O)�X��m>mn���DI�n���̔)���A�/5"Z���O(�T��́�e�'��ur�I]N2��a`�3֙���x�I�.�'�.$!Ve���H��ׄZ;. ��R�g^���)���rU����"��<�DCG�`z���"d��<@��$�M]�'� ��IF�H������/u� c�I͚9�`��$�V!k�f	��Xm�͓����$P���B^��*��iP�鉐"M�L ��Q�s�bq�Rk݅C��8qr��AX"�O7�9�޹bs�U�B�V�ٰL�4�h�	"O�T���ڼS���� ��)E�nK7O���)J��E�ХU g���k�O�����/\_�'��ÖYC�pK��)]�XYC�5D��*�e��`���C��D��+]CfL�"#�Y�"܉���&]9���e����<�s��2~��l� ��F~N���R�'��Dq�ڪa�RA����%�䰰��&~��BF��Yg��J֯Rn�6H��ǘ%�ў�bVY�O%$AQbHUk�a���ڴ[FhM[w"�'�X��!��^t�yӵ$�7p/4]a�U�i��y7L�`�b1��OT�U��
���M�1�������<E�ܴ	-�%i���J�,��埈\��� _�b��4� �]TꥨEn��|z&.�H� �M>�S"Ǔ">�!�d R�`�D��V?���0 ������/"ɚѥ�EB���Y4p2�`�$k_L�/�T$�@/�v9�@�D�_�M�"<qÉ��g[��h�4SHH�h���q��!�v(��~z�TEx���(���BQF5w��2m�".���2�ɩ��U�sj�(V������H4���#�6s����n�O.<`�S�ݦ��!���ȱ�"�B��4ȧmK��pϝ�, $HQ�Ӂ~���y'>&,�!k�eW�4r����ֈ�K��Ȟ��|���'�~A��(�){q~�I�剷@~�����\�����\�dKd� ��O�Hի���K̓NʚM�V�S�C��P�(ٜ����p�� ��%F��hO-���9��)�@e�b��IZ�OҰ@��i�χ+SH�6M\��.�1���(O��1bc.T@7D a��a9��25 �X���`���#B�1w뺄���Y�w@�K�n��1"S7��`����Mc�u ׍-vS��<qg�	�n��]3��],���A�
X�|�t|�6G���
K�U������G6jux�Y�]�-���E��
A#:��ip��c���fWy�f'��)p�2�y���ip����\��Y�-� ǜrSG��mYf0�E�5Aٺ�!"l٠���6���9ӠU���$VF���2�U='��H����Ó'���ڧ!�^i
pD4U�b�	�@l:rj��DRHCa1�O�(熩pk���� �F�4���	85H�Cӆ��46=2Ԁ�w� @�	f��P��9P5��=��A�"Oƈ���	J�DR�G+Z�T�ԙ����hW�5����X�Oc�����y�b4�ݯN�<�
�'*��X����tՋ���&9�$x�	�'a| a��'1NZء�H�+;&~�B�'6��'��5+XH��ek��'R��p��y`�SNW�`"��[�'ު�d�̻X��L1���lo���'JU��f�#1&���D�Q��{�'	B���Y?`@�Z�bQ�K���	�'�TPQR��ahxRb�|ư5�
�'kja��J��	)H����ۊi�Ah�'�:q�F)נ}�� B�3�j��'8p�c�S!�]�v���#Ee��'�V͓�G
;BҹF�ǵjs�R�'�`���;o���V �!fZ��
�'d�������z��EPcݒ\��'Iތ8ЬŒ$����-�
LDEC�'����6KP9�.��Ϡ)e����'ȁ�c��741��Y5)����'�~��F��.bN��å"�����'�p�V�U�3٢M�4�^ �1�'k�xA�#N�E��(�$���'�Py�O\� =b���`���'�0\��	���$�E�F�J��'VU1���M��+"jވ|��m3�'�����ڲk�:`&L�9j��h��'KV��CK=D���D��h�P�B�'�������*L��bW٭��y�A	�NuA���5sb�I�^��yB���vn�б/N1/ъ�����yr�ѷU��1+$J�i!�`rj��yR'���=ʶ�Y��J<�y	�8ھ}���J��@�ߝ�y�'�/۸��OR8�ҐI`�6�y�*����s��5%��)t��:�y2	�)]5��A�
 IX�����y�+��_�2�p���?������y2 R�/�����7���(t���y2-�<R�qtN�6M*�`�NR4�yRo����$v����2�yRD^9�j���㊜c�>8�i��y2���, � ƇK�����'D)�y"% 	4�ܪ BZ'J4Z1kX��y��o�4�s�Z���<��:�y�ɒ�{�aH$+�
�j)j����y҈�(z�~вU眾��) �A�y�A�0<�<�(�%Q�{y����	��y"��%��Ҧ��Z�F%{R)B�y"�
�TB\��p*`#`9����y҄��!{:�ӂ�ft�ae�+�y��
b�y���g����Te���y"��#t*�ŦàAI:�R��Mp�<y3���:b\��͘��p]���s�<Qe��
P�8�1�jFP3��3P{�<��n�5(a��w�S�p�8{��v�<�J-[f9z2M�C���f��q�<�wf@:~�$���Z��j9��Ks�<����6l�v�P�=�&�0A��F�<1�ȫX6��6o��t�f�Yώ}�<�T썦d�~2�oY�)8���Vb�x�<��O91�0�۷K='^�U�� �]�<���?,	�t+�=K�j!� E�^�<I��:��L�B�@� h}��U�<�  ;�lB.�K�cY�nx%f"O2�ە��1:�@`LE�mު=��"OL��7��%Sɺ�b�ES�R���"O![0\�s������٦�H|å"O�#a���8���@��U��K�"Of����^��	:�m�8XV89�f"O��
$ �	[�05�Z�^*y��"O0��B	@;� �]eFH��r�<��ςU�H!,x�0�Qb��d�<���	|nLU�ፚ?K�h���d�<�UJݕYLU�@hW� f>�ab��n�<y�k�;3 5�pO��_`>��S�<�!W�[���� �� G�]�EJ�<Q�h�A��y4!iI�pGB_�<��B�,��I"�h��>���@#��`�<����>�n�1b5ZR�B�d�<����� �+��^Y�����M�<�q���n��P�Gה|�pH0�n�q�<�%@�5�����̮>��Y`�`VP�<�ro� ���c�
X�<�x��H�<am/q��q�*�+L��l20��D�<�iZB+3���њD�mH��y�h�
D�eY###?����Y#�y�̎'�z�#2��:�pѬ��yb��q�f]Z¬	'���(�"��y"'Ӄ#��j1
��ͺU`��y2�	2��q󇎒�h\2B�+�y2�O��`b���GC��A�@̻�9D����TG�Vm�ơQ������J+D�T�w�C�P�r͓� �2n�����2D�H��(�N=\��$�+_�v�� )$D��:�,��L���G�6����!D��@-���r�"֣O�d�ԨR�/9D�TX� �	�؁3�a�1r�f� �H4D��1'%\�>�C�LɇP�DH#E!D��`G�=V�:�O�d ���;D���5-��l/� ��2BmJ%�l:D��Kg �0�bV�����ۖH;D�t��E�B��H��b�
**Ri���,D�`В�Q�\�`᱃�@;vxz5�E -D�8�q���T��8�DB�o�f@�L*D�<8j_�T58��ύd�T<��+D��C�!O2{� ���ʏ@ V��%G)D� c�F3�0���B�'0)��$D��#'�܂#撬ц	�!BkrTI7�"D�@��-_�;�ZY0D��!7�BD��5D�խC
Y0�-�t��.-
���G3D�l�V��31��9�Cɯnt�����1D�dr7��8#z�rb�|�|U0��,D����U[���
;4li F-1D���U��Au�<7H�N9�\q��=D�xBR)X�<��!�<A�n��� ;D��(%V (8P�f�ݹX��S$D��y�ԟW|Yv�Q�Hun���"D�p�߬#���� <1�Rm��@7D�У����u:��vk�J�\e v$8D���tk #z���w���
�#D�xJ��[�ukƝ(���,��B֎"D����&(놩��3l�x�$�!D������f�����hY�5"��q�!D��5f�-����5Y�ι{a�>D�,�wn.(�� 7��&\n��"#D�0�g+Y>b�h�҉܄^`D��J D�|:���=��YC��BaP��� D�� bhb3?�j�;S#S����D"O$-jb�A�m�6s�S)��`w"O�!"�o�R}z��!��a�#"O``j�g�u��O݉b0��"O\���"��o��s���2{�29J�"O��HP!=J|z�/�#f>P!�"O��B#�����q!��b��g"O�uٕ�B�!�� h4N	Z*�H�"O��S�V�^g֍�am�1!-ޜ�4"O"H�`�69j|��� L��"O�І���'��wX��b"O� ӕAN�T� ՊCPc$�A�"O��SU&�-W/�[��W�k��؁"O��1�D�H�n��d"�G���ې"Ok�`G�<��W�A%4�:�#"O$�2T!٨c�@�b�W(��
�"Oh�i�JP�?,bW]�<�hmi�"Of�
�R5��c������bA"O�9X��8�ny�t��Ƣ�y�H 5I�I�V�
'�`���y2F�:�б��H�J4�q���y�O
�#bАi�	�H��Y���y���1��(y���5wl8�JQ��y����V~�@�sEԀX3 t2��ɑ�y�%����Xy��TO���D%���y��;JL���ՐC�d�A�BH�y�H�:F �X���=j�A�r�D:�yϑ
(4����U�2�q��e
)�y �2\�6�)򦊢prT�31�P��y�nU��I�T����y҄�J�Eb5�Wf�]��+G��y2L\W��
� XO�Dy����y�V�_$D���BK�<As���yr)q������E�b��#T,�y�N5J�|a8�C�d��df*��y"�,V���Z�O�䛅�З�yb�B�@�0|��<�0�rI�9�y�a�Ys�E;M�$z�^1�[��y�R�$��20�G�da� �˻�y"!�ۚ,�d�LX�\dj�_��y"蒺$��m�7��! QT��'���y�ʛ�b�NUqSIE˸�ӦL��yb�4Y���3��Z*�IN��yR�@�aR���V�W6�����y2hyA���'��7��#D�,�y2�K+�Z!�4K/`�R�%@��yҏ�^=��n��5ʣǊ�y��M�k����#�
6�2����O�I� -�'_�RɓS�̜Q���xg-�8k&��s�bк"��4]ʹ�u��T�!oڌ[R���V�+�)��Z/M�b<�tÅ/zc5CD(4D�$i��_E볩,$����@��� Ҁ�Hn-���1J�X}��b��4ZH���wP���$��}IrӾ��m\�0��˦��+t���c"O��#U�F3J�x�B�?d����'�	�}��P��d�O >���`��-�� 5a�0-8���'�8-��J>J��P�����9�]� ���) ���O,ᨶ/Y�[="��0V���"OdL:3�Z�]	 - V�O�24�S"mO��D� z���pB"T�CU� � ��T��|2H�>ON��t�ik`|`N�}��"/��}j\���'��#@�̗6Z���E�6k���y��DHT��s0�,�']��#G!:9\��$��X�U�ȓ��-	FG:��W1a�0n7$�FDj�'�)��� �e�V��6�>�@�����"O��&#H�*�f�A���/K���⑟ĒîY��p��+�*b��C@J^ M2X��a	$D�
`�Š���&(�"~8 ��e�#D��b�G�P�����ה2N
M���?D� i0�d�Dh`	A�A�
<!��:D�X�t'O���I�f\�f��1-;D�<8��J�@@Y���v2���8D���R�ء.2�ٳ?�q���%D�D��A?�3!��`��c�a'D��xBD
?hb0��*O>~Q���9D�`���Q+)�б��#h8�� D����;uj`$Y♾���sЎ(D�0��ň���p#)�:����5�3D��3*��0����L�Y�E�g-D�@; �OY�f�ƸB�%K��)D�C��%�H��nS�x�~-�d�$D�����)1��'�B
P2��7d1D�p�B��7�Z�����D��A1�5D�P�%Ñ�x�np��&�+�:d�d7D�ȑ`��y���a^�	+��h2D����\�'��!Ɇ+ȟl"ܕ��o-D�Hj�(���.�q�3fN��+D�cP�>i��Q��O�����(D�<�A�\'OQ��(⋋=<!<LR &+D�`�p��t9H�S�nB�Q�2���*5D�����ԽrR*�����=Y��sb�!D����M٨0��K�M�9ȜR�<D���*�2Xv����I�Լ��1D����Ч:���!�6t��0E�-D����ƀm����+?�ʅ�9D���чˎ"d��-۷J��Aa:D�(9���>2P���/��u�D=D��ٱ��l$>8�2K�8%�6$p��>D�@#H�-{� S�@�[y*�)fM8D��r ��[���P.9�ڰ�u�9LO�]����Lc���7LW�w�J��i�<-9�[GGiX�����iR"�G�<��'�T�'���|�IK�h(�2�RG"����ʫ��&}b7O^����7A�<�g�Kդ��g�6O��b��E{J?��cY*NvT0���Ck���L0�$9�Sܧ�.\�6��O��;#*xݕ'^ў�|��3#s��ǲ��橃ٟTE{��i̓!�~�����9"�h���b�3eў���Ӆta �S�W-�E�ä0���dD{J?��@�d���	a�z+,P�*����(O������K�@u ���i� 4v���T���)�'`<����RSB�}�m�Q��)*�'=xʜ�F��
7��I�I��	��ؓ�������O$d���OƎC�d�	v�"�a�j�>o@�qS�'N����V��yb��B>����� 1�kŒ~����!}"&�
�(O���� �mK2E�e��g@0@q V�,���)�'>JT�b�؟E$��Yd	!vbDmZ�J^Q�"Jé����CBG
il�ۃ
Z�'ia��`�!Q�>P��n	1�~|�����'�ўK`Z��1���ns0@�'�_#+
r�!q+��?�S�'�����cW�hh���u�U� ݢ��'�ў�|�T�K*N_��&�3j"��S`E���F{��)�mEt��ah= V�#�_�`ў��>�K?%�#n˻6#�(�	޼(���vhB��s�p�S>�%X�-�"��׭P>o�	�PI�>��'�(�m��<�O�駉�%�/r��kW�Űy�����\;,|��0�<v��~�NѽN����쒘"�, I��O+�y�%�.R�lP�d�����.Ǵ�yrJ�,r:��v)
3����,�y
� J���=Z\�;���R��:#"O�Y(G'��~�J��c�5#�:aAS"OV��#Y&Yϐ�1CA��K�P���"O�dcK�����1�U�V��5"O0ea�(M:0?�h+����h6�A��"O�� -�*��Sf� $T�P"OtD:D�Kx.�2�Ҵ+��A"O@�0fȊ�$t�$�^	P�{G"O��P���$M༃�f�v\9
Q"O<��%�J�oh�	ڧ�՛Ei���"Ov�`2�&j^t�ZDFإN^��"O����쎜R}Z4�b��FT�@��"O�
'&T�)X�l�e���H�@�!"O� �N�$Ur
��t���H�*P�	�'��$���6Pn���I�y�1�
�'��y�gL��`��"#��~��Z�'E�@��V4/�����l��1K�' @y�/;@� �9 i8L��y�'<`,��홢�L�`�@ĜK3P��'Bb��%0_$\����C�ʓ$����B�:�ڤ��ǚU�q��!�0�7�	0S�TS����r%�ȓ�p�F��6E��%kQ)Ւ?����s�$���MT�qEvq�$R��n��ȓ/^d�@��rδ����ѓ3c���4f��G@6}�R1�Rb�1�dQ�ȓ��g���+x���P��%C�K6�ܔ6�,(�T�XÌ��ȓW����A1K'���Ӎ�HZ�x��s�48��l����'�l��o[<	�$�X����B��V^֠��S��FX���$Ӥ	JhX�ȓ8"2�Є�Y���(B�!�ʰ��/>�ᘲ/�98�"��6�Gj�H�ȓ#�}�6�ʾ�M����`���t\��v�X�Y�@��w�F/*vՆȓr��P�d�G|�Rl�҆j
�'U�����
*w(�#����Ĳ	�'��ܣ������� '�����'b�b�6Nf]�l
;#�00(�'x@�kuh�6&�%��T)G!�MP�'@�ܣ�ԩ>\��S '�'S�Dl��'����
��#ì踇m�߲�@�'Z��gK
���7�E"y�'��� �׷�(T@�C�(=o����'	r���DV�Y��u��iU0%�JT)�'�2I`���qZ�p�fb�*n 	��'���Vg��u`�ax�eǒN�(![�'���Kp+	�Y��,[�˃�B���'�Q��^w�\���ޝ2��a[�'��`/B�x<��w�ª!��d{�'4�<A�T(W�Fyf�ϟq�6���'�U�6�� 7i�X)�.H�m"�X`�'���*�b��Иpr�Y�#jԀ�'v�d��l��/�d؁�е?L@�K�'k4��ӫ�=)��pJ0�I�G�v�x
�'�&B���W���*���Q���'-�!iO��U�®�M_�h�	�'�v��o�w�n�qW�<u�	�'�V���Oh"@���2^�<u@	�'��'��=������'[RR�9
�'�,����
.� �E*TNO��h
�'����I�5If�Ah�M�rD9�
�'���Wi���Lڤ��1]'F(�
��� ��#�����eх)���p*�"O&(3�Fۜ2,ٚ󁅝��-#@"O*�(��ļ7����G�G:Rx�|
�"Oh�ӣ���^�.1A�Ǖ<^��F"OR�Ɇe�(W������/5��p"O������%���T?�� ��yr��h�P�;$h\M���x�
�y�aY�n>��S5���F��F�ϗ�y��%�p�@C�"�晢vm5�y�E��0iza)��Ł��c��y"�(�1��B�Y��� ���y"	�1y%��k&�6W	��ÒE��y���Mxv��b����P�y��p���B�L;Y�> ���yBذ��A��(��P�(رbȞ�y�lW-�j�a��=JD���	8�yb/	�p;ĩu/�3�*��
��y�c]��i�a�#�"!r"/��y���xU��9G��sV��y��זU�`�@��$,޴2�� �y�ܾb>s`������SLQ1�y�¥{��#�jAΦ%��m ��y��F.�p���������u�!�y��8b�P� ��O��D�rM6�y�!ړ=�ʒ� }��k����y2�ŌqD�@h��%���F���yb����
|��FZ�"\B�3�N�yR�X8$�!���
�k�ȅAc-�+�yg�:G6�E��,_��6KO3�y������s�,P�WƤ��k�yBG�s�X��4�N�%�h�B�A��y�nR7f��t#�B�My��J���y"�ܙX(�`n�;L~�l �-��yBc�,���X��ȎtMĝHFnݘ�y�M�e �$�Q�
iB<Hf��5�y��H+�=�gK+�H:�Hǿ�y�a̺4���M�4~0Q'ǅ7�yR��k">���)�l86<����y2K;����gV�z �Xd�R��y�o��M�\�UmArc6!xC��(�y  L�|��F��*2�������y��&b��1`4O�#k��a��"�y�$�	k�����������Q�y"�7`x��a���({�}� �M��y�� �d��%AaM�"��40P	��y�I�0n�=��-�#	̌rbG��yBퟴ06lHY`d�={	����L=�yb�V�V0t��H\0lO\ ��e\�y�D�V�]*��Z+`T0e���G�y"�_'|���[�隚U�����ŕ�y�'~�E����T��g&�y��Q2j�=�FT�E=��pA�\��y�v���2U���:s���@D'�y���h%����?���ɂa��y�.��Cm8,у��0Jp	r���yBC��4k΅�T��..q���y��M
=�8�c�HvSر�2���y�Y�)�vT���ۘt+(EbB��1�y�!8'�Py�0���q����L��yBˏ�u�d��C�|ۆ�P��y�ę UG����H�u2�ʥ�O:�y�b�J�ީ�G�R�C�<Jen��y�㙞C�ژRT��9���RD�T��yҪw߶q��I�,*̀��
�y
� N�q�b�=~[�d�A�R�R�8���"O\dQ��B n�2��@$Q��R|�"O:�{���6+�Tu�t��L����r"O�țb�؊j�:�"`ú��"O$�7ə�"X�����<Ē�"O�٩"Ȕ9�bT��!��egLq�"OD,�db�(X�
x��A�4_Kt�"O8�d'ˍ�t�CV���E���+�"O0�[wW�P�p\�$�U$6�@"O����>��0҇�R�v��"�"O�Y�fGږ&��;�ꍜqiP�Ǻiߡ��U�P���>�!0�v�!�$�,"a�mK���lwX�� 3x�!�Y2*��f�1}lt���\�?�!�DG;<�`�����0T�Ap¡�7�!�$��K��j�PK���"�?`�!��NP}B��Μ>4� 8smċV�!��-�$���N�r�h�QmX!�$#Զ�;��βW�H@�(��!�d�0c$���u)�T��0�Ӣ�!�D�>$�,�WЫ !Q�`Nxf!�d�*�Tkw�&dN�3a�g�!�$ b}��h��)|�{��΅'�!���)fC:��S%G�Q�r����<4x!�Y0J[~̳�C�#� �[$NҚkk!�$I����rFv��!�d-R�;@!�D��x���b�)!�X�U�4_5!�ę(O�d�����&�P5H���>!�DQ�u�r5��'��h���K�!򤇋j�6PҵǇ%KW@0a�AC�z�!��v�H�aG_U��³�9#�!�d�(a�������+TI���dA��z'!�H;x�QGM�>���c ��M!�D��S��BB�|&�s��T1
!��K�n ���z�R��.�!��A< �~��FF�UB�ҫQ�z�!�6Y�fЃ���?g�̱�I�<y�!�dH =b
��D���J\Jং-��$�5g�T�c���+�PAc#��yR��z�'Ò�nvHe�g���y�
A 'i�	�E�ap�����¬�y��3`�)R��ku���%Iٌ�y�EE0����&��l�]��%W�y��$������p$�E띫�yrAH�&��0�u��6�SR�C��y���
)qB�ze�Ю_M�y��i�3�y��Wxf8�8֨Ba����Q ˜�y��R�����O�`�p��rJ
�y��(~h��O?S���!�$/�yb��!C^� �~�VT �"б�y�Ñ9�	��L_��lEzᨓ��ybϗ�R1c#��u���0�)'�yR�ΘZZp4�@(_
V��5)�y��l��1�b��9Hi�l:�lԈ�yN�('��0UI��qt���ueݕ�y�L_<e�L�HB+΃omD�� ���y����j8�� �72z�l����y��F�8�I ��{dX��!5�y�닃3�05��؞�;�ʚ5�Py��R�:��U�j���U"�U�<�1`=M��Q�&Q c��V�I�<a�&E�['��Z���4_��&�MF�<s@$�<�3�� �q(���M�<	��㪉����;����̀_�<� Ȱ���]43��]A��+'(~�0�"O��u   �!�� �I�[�N��9*���-Ƕ�q�"OT�&�L�е��ԢB�FX�"O��9�l�-PD�)4EL�k��`�0"O�x"s��6b�� dE�L��TC�"Ox�Uj[�p��5q�C[���"OXՠ��t�Ju����?H>�u�"O> A�n�D�>��W��AF��A"�##W�$��L<�@�]�n|���c�4yu�ܐ�d�J<�`��97��9���̫r����&{��h3�^�/����$�-RH0(Tb�4nn�ܘ���%V;����c⁡�aS��F�<G��<�����������Ǔ�?�\B䉁3RqC�<a`H�e�6Ml��I
Q���!S�
��yzÌ�A�O�^�aa�ձv$nQI�`��h�L0��'κؘE��¨�1+�<V���[G��L���񳀅���3��.)�x�Q6�J��OXO����,&�|QAG��9Y��aW�U�#��1W�%.��%Ȁ�t�X-3
�>�~�b2�R�Z��w��G|�G�\Jhp�!�׉Tˬl��zr"ćU��k��*��e9��q�<Q7�F��9�,�"y �
N��pA��O@���y"g�-D�Z�{�W�O]tp@�ٔ3����O�i�F G"O�|���H$"�`���郔�vX�R�jـT:rm�
�.l��6.��u�'����G�#{�.�!$#�W4�i
�W<�Q��ʮ|y`�k�K.=�֕(��>@3&�KF��9 ����3�	�0>��C�,-���bc%lF���D[u�'���8�ʉ~��䠓�4�28�F=�L$���_��*�R2hP�F8:X�R"O 4P�f%W�<Y#�@�#9^�!��'h�AZ���w\,RB��v�
$H��SC�t�IA�r�%!P���^ �ȓ�켁§[�Q�x� �oӛ�t��g�O�*x���+
&�"���ɆK�D�I�r�Xn�7D�Z�R��Q)u�h�?AP�l��'�N��'C_�d ��!��i:HI�&�U|t�q��N@��#T$oa|Bc��F����T,��"c"�
��䏵���r)Ol����ݳ:�T�j��_aDhA�OC�-��e�1'���4(�D�E��'��ZԮ�<mvȬ;$g��>/$���'���6G�;Dpp@����
*���O� ၁EK�C"'�x��mH�΀�������?1�NG�AI��h��1���cš�]؉s�6R�a�'�^a�קW�u��[ϟ�O��p$O�@�B�!��4Mf�(���I����"p"�ɲ{���XT��-g?&PA��~��0�%͊��Z��������0~��h �_�(�%U�5����z� )}R�	!X�ŊA@_PQ�O]+u%Hz�d�ku@�y����'DTq��-I��l{��B7[j��O$���*˄n��"N������b�tu �%A�{���K]?3�豇�#9p
K9 S@ѡ̚�5�;�{rm�p�c?O*|�4��>f&t�BD)9�9� "O��d�S	T��$�'#S�ՄKc"O��@E�Zd���d�)|�vd��"O �+�K7
����C��@&�d�"O|���E	]b���D�,˸<y"O
���(��B -
�Ԋ�P4�"O��KFN����ѠHI�#���s"O�AT��%`�dT�Tǈ�^rF�"OJE�!f��G9Ԩ+�)~n���"ONᱧ��iw�%�g�/&^D�x�"O҅S &��8M�5���bG��A"O��˴f/.���[,\&���r"O� � �J�^��E*h8�a�"O�2����%�n��u�^�5@T�0"O�� @����a�!���,���B�"OZ�����f��<1�a�f����"O�bL
2@�8}9Af�^4�9r"O�	1Bl���:� e_�EC�k�"O����o&�!�s�%I����$"O.U�)��0HX0`p�@�|f�"O\0IP)J?4P��;'7j��i!"OjY+U�\7fL2�s�ᐺb�^q@"O� �����߭mh@��@���b�ip"ORD��617�im:stH��0"O���Q�|��j���[i�,	�"O,X�"a�"�f����smhm�u"OP1�T�U�z�Y'��$B�Db�"O���J�x�VQ��*�WPd�Z�"Of�I��ǮOQr4��I��T�0��"O0��uQ|���(r��tޠѡQ"O�<���+fn&��6쑓�X!�`"Or�t����ˈS�H\C"O*| "E[�Ns@��5��@�p��"O�H����90����ro�8T���"O�I1(��j�%-H�w9t���"O�0��٤}��-���
-"#b$P�"O�,���θ&r��K��x�i�"O �`��լV �� �I�DI��"O��+�"�.��L�cH	�q�d�r"O:%+t����ܐ4��F�ab�"O<aX�$�>y��i�oN��&���"O���l�}
l@z�N�����'"On���.3<�5�cU{t�p�"O����ő�a�\l�l�N6��S"O2�I�&E(-��(��IV(�
9:�"O���A�ǆka��B��-l�ʔ"O�e�1C	1s�"]� cU���t9�"O��J�x�4y�tc��<�R�"OHa�&mǯp $CQ�S5f�����"O.�a5GΓzp�L뤀@��``1�"O�ʴ�ڮ	q�)
�l��+| \ر"O.���nχH��e�Cs���س"O�L�хݑI춤!���@�"(i%"O���cL	�c7��C$�ܥW���t"O����Z4��,ˇ�U8{f�5Y�"O�i�gծu;0-q5�T�nD �8"O	r7��H����2#�F�4�� "O�|z�o�&f��1�@Y���e"O���b�p3���m��ABE��P�<A�k�4;�$�6J�5.f�u�!�V�<��(�;qT�aa��@>(���i�<�`�cJYBhD+J�PP|�<0`�s:�(F�]�:��%��e�<�#�ΦJ���pH�G�!赨�^�<��KΥT��#��-r p{E�\�<���B�(>�t���E���r�i�T�<���ì�0�+�d�H�0��s�{�<�ve�%{��<�P�Z�L�TP�%�II�<ce��{I�0��d �m�UK�@�<��c�?,���g���q���<a�ԋ�NP�׌�u��(��^�<�D�͉6Z�4�
���lhafT�<�WG�fp=!�B
gv�q0E]�<!C!��o �H����T��1��u�<��Z�	�	:��܁iRj�p�h�q�<����hiQ��O�����f�<�t�RkΌ���"��� ���<	�B�x� �*���_�&�#Nx�<AVG�����1X1|_��*��S_�<y�B�;�z�5MQ&;J���� F}�<�#τ#@.��-T�gS��;���}�<�d���g;�=�B��;�0�X��{�<�%?H��تցQ�\r���t�<!���x����ĩ�.}
��E�v�<q��^48Y�@�ʎVmjݸ�o�<���x�PC4�^��0؆E�u�<� ������r�V!��"�1�F��"O&�!s�� r^���!�Ĥ���8�"OlX���L�Z�`��&M�`���8�"O����g�L$�:��M�W�hd�$"O>43pD�0P`؂��ƅEX� S3"O�hh5G�1A�8e&��>��"O�A%*��~��xDER. �<)�A"O�=��\�4+M�<�dz��c�<�7�ְcvX�W�'R��a%�X�<aR&�z��h�$�	-~tiH�f[�<��FN �.�u)Ϯv@ ��##]�<�eU0k2<a N�/:Jua��\e�<�p	K�@${!!_�r�~!�$ot�<��P�p�����B�{�$=��^���Р��+��S�H[�;>@a��S8��po��������5Dr�ȓE����W���/8:�8�
D����ȓF�v�"��
.Ф(����"Ąȓp| $hs�2ߊ���O@�t�ȓl�����ô�����@���~
�HX)^���xԬ��,��uDI�R��_BH�DX0Dܽ�ȓ����@��!X�A؂�G1�\��ȓANr}���N`����9{}����8�4�PB�@/K��m��N:jU��ȓ �0����O��	9�ߺf(��U��$S� ��i���vhZ�ba^��s�L�+! C$�����* ��H�*8��ϋ���u`�R=G�PA��|�Ve(��\J��R�.�;G�jE���Й��	� Jh���.I+S68��2�]J��ݰ}Q&Ua�q� $�ȓ Dj�i���z6�%��h��4�4�G������a��&]à�ȓaONq;GA��J�� Q��_�|�ȓw�����B�7Ax�	�U��( �|�ȓ|W>{���.i�  ѥ	���E��n�V9�͔�<��B\�ń�>�*��vF��ߊ�bP,�?_(\�ȓhTR����44q��gĘgF�4�ȓ$⪔��,�e��$��jH@L%�����:���i=T��GbL{;�h�ȓLr<��`Z�-!����G�%�v8��7�4��ŇDǤ�f$_#q�~X��$��H:t�&>D����hĤ|�Nчȓ	`��G
�9����DϤ"�RU��:o"�y$MO<5��
%�Ot_���ȓvv ���4o�*�#��Y�0�ȓP.���C��?ROnXÕ�/L'�ȓI�ƌ��[�8Hz�P�H����ȓ��zO�SڨV0-��(�.D���k��>I�=;�β?���S��/D��p�f�		�xii5�O;b'����/D��
Ů�%j�`U`!�Q;Yr��Q"�9D�,�!�C�:�`��LX��0�6D���&�3^%Ȭ+SGK�8"e��`.D���$N�g�V 	F/��7�F�z��,D�k���	�Jt�d�F�C�l횑�?D���r�ɺ%�蘂�� 0�JU��./D�`�w
��8���[4��c~n��)D�ܪV�Ͷn�D��sa�`����E2D��׆��u@��H���64�H�3��1D���R�˳M��A��7z�2y�E�#D�dc�M6NA\ݣ�G��V鰖$>D�� :+�ڸk�|5�.&���"O��7�IpD��r�2Y�bUAW"O D�`��k� ��D��cڪ@�"O��큔t�0�q��;��a�"O:���u
����'N�
���"O0(�Vhߚ=l!�7��(Y�� �"O�(D@S�F�X@���K~�x�"O|�SB,�	�&�r�.�elF�1a"O,�
�"A�ky8�(2���7D��Ap"O�a�!/.�������'"�={""Or��H�K�������s�bVm�<��f1h1t(��+�1���Ns�<�$�$�ܬ���ο��x�@��b�<Y�)R;=� ��^,d��qq��f�<)� �5pĴ�@G�N��� �j�e�<ADY�ܣpj'MJ,UCg�c�<�tfHMBh��_�9gDܙe	�[�<!��[�����p�6K�,ÃǆL�<1�NM�)c`D��	��"gt@q���J�<Y�<p��I	�й"P,�[F�A�<A�c�"oe^��Kc.�y&�Ig�<aQ#�$e����MIfxK�WI�<�*F�&��g*��q��k5�Y�<���:r��C�䂖)86fj�U�<��a�N5�UQ0!L94�6T� �P�<!"��9t���� ��4vE�<�ǚO�<����&��2�+;�|�Ѣ�Q^�<�%�,-�X�׌�)q7���)�Z�<)S�����"t��$Gތ1$�GI�<���:��@�򆖍$j}2%i�N�<!�O�+*���gLO
j��("E,�r�<�bH�k��рAJ�����+�B�<)��Tu�dkVb �"�^\9b�_y�<a�T�\fv�Q�U�a�L�u.Y{�<�bLYѐu���@l��P"Ys�<)��M-(���1o:5�VZ�,Fn�<����#�b�����a�hdLj�<�'l�}��ɢ`��2j�z�"k�<q��-�8-��$�>�n��'�Fb�<Y3�`M$ 
ٶr�^��v�T�<��	Ph�j=�RD�;F��Z��M�<��c�j�0X��2J�0գ�q�<���Y$^���e�?�|pb��o�<ٵ�_+J�����<[���[�/�`�<�e/A8f��C)�>?�V]���Hf�<y�܄���A� �6.��â�Hc�<	�/G�
M�q{��B&nWL����Z�<ك�*w���B�Z�6��� @�Q�<y�����(�GɶY茩B���L�<�E(��JX���LW�p_(|U��b�<q� [9X~B�A��� ��m���b�<���*J�D���w3Jؚ����y2b�n �=�@m��7ONL��%�9�y��K�P�"�[�u�H��Е�yReԑ|VQ;�%������>�yA�&�<A����x��ar���yD��6,�Hbi�&-�$mӖ���yB��\PLY �ܘ S�p�UhT��y"d�X�r�2pd��e�GM���yBÄ~ V��EÆ'�K'mQ��y��O5%J�:RgɊ����Ƣ�yr�#�p]*.X �%���yb�w�z����I�zښ5��]�y��ִ��ua���.E�N ����y
� ��L�D�+��<�p��P"O`I�j[�b�D��K�)�R$��"Op[a�D�W�z��d�#�ryZ"O)JW�R:���ѥ��=�>��C"O}2s��M���	�h߳Ԇ�@�"O����⏣Z�P�G��Icԑ�7"O�� x��D�#�B����"OH)�L�X���Q΋*;����W"O�u�Da�+N��Q͊=`���H�"O���bB��D�
�X@���'�lL��@L]���ɵ�r�|h!�'��JV��� �26C�%�t9��'�D�ZP!N5<h���Ŋ���2�9�'m��5Eȇ]>2I�P��x�\���'��i�`e��uJ ��9{l�)�'�� �e_Y8,�2"�_�$m"���':V�hԫЫq:�ڑ�	().Q�
�'"y�qbҍE��������-��'��љ���)G�(�f��'\�mX�'iL��Ψ!/�ab1)��C0҄:�'?^��/�~�$�Х�,T�H��'(��7��]�� P�
 �@(�'@��)�m�ک�G�(v���'P�(z��}��,#燘%u�ȣ�'0��Bo\*�"$�Ơ�1]G���'���'K.&��=�a
�V�`���'�r�����8�P���� 5��'hNx0���\|����0��'��I�� H� Ѐ��	�$��'V�HSM*'7�0�c!�!�AK�'#�����iٴ��Bƅ |�1��'��e��&A5] 4Q0UkCz�&y�'v��P��cA,41d��M�����'��H(��5"�ɡ��s�|��"OJT�@H�S�:	P2�K�_�:�Is"O, �a��q��Љu	F���"O`09��o�1!���
UZڥ�"O�`�L@�`���)AE9DA���b"O�<ɒeG�>���;j�9>� %"O��3 �*<�
Y��\o)�|��"O��/��BԦ�;1�Q5 ���"OT�$��/&jPsc�J"�est"O.��p/�#ߤA�VA�]�Q�"O����d�6)�c��K�"O��S�я��jEIFD�Z��d"O�e:�NF�\�e�G'�h�T��T"Oft�F���B��I(�'Y�K�B�HW"O���ś�":~�J�GG�V��@��"O�T8�P�'��ePG�	�
�t="�"O�� ��JG����Ҳ%7��a�"O�;p�Y�0S��g[<,��ˇ"O�5�W��u�"��G�t�v���"O1�f^2V�Ȉ�u��	��HE"O�A��jɦ�����ƣ��-k�"O�H����,I����� '�(\��"O�d
`d�%n�Ή�@��;&z�}�C"O �3���S��%�"�G�z�"�"O�	*СT�u"	�1�	TR��5"O��Cd>"u.���O^�੐ "O��� �֤y��QPD��XM�"Ov	�Ő� �̢#�7`���V"OZX� �Fdq)�-x��:�"O����H�j��ad'ٗy����p"OzPk�@����BV暻(��|��"O� ��s� ;�P���pAc"O|[�������#��m�`"O1�RA�1�ȬA��\�a�� "OVa�7�V�K�N`R4�@"�-+"O�]�#�G�F� �I�	�V-�%
g"O�(���8��t�^5O<A0"OΙ�V�]�wc�x��w��(R"O�9+5�W�p+*�v�SGN�I"O2�B���S���Ѫ��=��"OnE�GR=e"�,��ڞW�d��"O�e�Q�G#:z�KUEʜL���[�"O���.�o~��e��M�f�xU"O��B�)��c�PX���vA"x�A"Ob����ԀeH��Q);UA\ͩ7"O�l�@-b�q)g̮KRP]��"O�(+��L!+������P+��"O� �$Ġ2��:!���h�I�"O�5��╼Q��U:!��}$�0"O�8�5#��r���V6Xt"O.����0~��ai�؞>���#U"O*�������$R<�JIj�.U�;\!��N&��Y��hZ�N`����	)�!�$:_���gd�#�5��IAK!�"	ԐH���Q:bQkp��=@!�d��NU鄠8X�!Y�� o1��˂`��2%�E�]���R�]'E��|�Ó	-0�J�`ѳ�HI�G]�J�u��F<[ 9�Q����x5��Χ>zQ��^������ �}��S�W��Ě�(�đ���Q>��7eN�S��ـ+<e�e�sǋ~R����`��C&�;�r����-�t�r��&4��X&�ո�V��.|S�ѺҤ��ʦ�g�"�P�h#�ф]����+:�� 	6cI�eo��\�����	a�T�J)��yp��T��FY�d����n�V(�@U��� o��@��������2��3`�"`ũ��ص0��FRA|���bD�8�>�fU����
Y��]��`Bx"iC��5*��a��+�@$���Ҷ4oa�違>.T��WĈ7��b�M�-�\��bվ~D�|+]�6�ڐ�
�'!�n�  %L�DOr����ϚL������ Q��@�W�n|����x�O��Y���D�(� {A×�{Z������
N����`�j��Ak>����W�<��7Y�/�F���_+_��mx�s��%#�%�(r����S
ڒ�
pj�@v�)˖��! [��i�L����e��2ܴ��Y��g?I�MS/�{�l�|�Np��o y�<a��]��Ͼ&�bi�q�Փe��C�	����š�/A��0���w�C�I�.F8�7!�5{���6-3W�VC�	�I�n�k��q�����L�LTC�Iu �)�KT"9�D5x��H$
�C�I?3�D��+�:,ȽK1�C��B�<Kf�{���5w����K؎lc�C�I�5�pD"���0�=B�+ ��C䉉<5:�3��E������g�tB�I�;�H��B���&��2��ϗ(HZB�	!4$Z��&�L�yT�d�bBA��*B�ɇ.�T�Ѧ��ix��yr(ݡxX�C�	N�:a������gő H�C�I�~J�ɘ��, ���R�`�=�HB�I�d���!�f�T��YT�9K��B�ɲ)�a���R��P�r�B�C�ɵ|�X��X�^\\�zA8܀C䉥_�L��
9R�d��F]�7AB��$I4��@CG�mx!����,>B�<Z4|�!H��D�2�Ӎ0&B�9���[C�1C4��	��a
�C� \�8�I�N�O� B-D;4!��ْ;8��#�ƗI�Dd�G˗�O!򤗿�V�*@��k����~G�A��"O� v`@��mqh�3���/*2�%�P"O4mr$��
`Z�a�&�C"�a�A"O��&kÄ}*(L�#�mf����"O��h����_%�I�+(W]����"O�TAFʌ	�����>K���4"O�`���7߶�C�kR�a?:��"O�XQԡQ0n�P� g$�'�Ug"OA��JܝT\L�scIORL���"O��P֥�f���􇔱Z�nY� "O��Rh�-C=xYH��7�UF"O�����^�Z�1�4�C�L��9�6"O,X� �ǩ3� Pz��ߘt�4"O�T�AʅKHl"� R�.V��#"O�p�S�G0J�L(� b<*��P"O�0��*��vz�xA�R<93���"O����;��X@Vj&x2��"Ox�{��	'�=��A��f���"O*<$G� ?u0u
���r�x��V"O =ru�@�A��r)W�_�|ٗ"OTdI�i�i�b��n�B�"O�hI��3N��8�b�9p�)��"O��J�!L
�����Z�`-x�"OH��Dd�"n��ı�l]�j���QR"O�}E��.z�ȕ�X>b�И�"O�$�q O4	�8@�ǟf#Р��"O�,�T[@��k�G	L{b"O�x�0��2U���W,	nQ�8j�"O(�KD�ͅ6��� �na�4�Q"O��@���"D�j��_�"T��0""O�h�"]�Lt��ro�	 <@E*W"O�Aj��>� �q���e6���!"O� �I�;J[��۵
�C���'�|�3��T�P��ɂt�X�T��'��!���̌��U}�iz�'0 a���8�a���6���'��<I�����ar�8#����'�=����R�T)⭇� �B�
�'�^��fȀ��j,���`#
�'�n͛F
�2!Of=QQӸ_@�:�'�bu	Tg�:j20����#L�8x
�'A#�ƺp��K�����	�'5�)��P�J�4ǈ:v�\��	�'I��3eLE�`�tC�L�i�fA�	�'�:����W(,J���=j]�T��'�&<���Em���c������,��'纙1��X<}!�|�n�-\L�X��'dp��ς�5��*�c��Zl�@�
�'�����;$tz�ʏVn�
�'���D�r��ڲ���S�xq�'s���CI*c/P}�FD�U��T��'q��r�+� k^$�Y���U��|��'��eڥ�Y{��xEOŒpA�'��P�o�6ߒ`�Ɨ�	2��'�&�"�
q;�i�D`��y�ј�'�"��!-�*�>r"��'$�ǅ�>\�F�S�D;�,Ȫ	�'�x�'Z���GK cv�q@��'��E����P��0��Ѐ�'wv�w�՛H"|��Ȁp����'��
Ď�u�������6�����'Ub�:����MF��/�N�r�'��]X�n�;V+��y&�,:���'���A�(c&�af��#$Ġ�'������h@qd�:!��
��� 2IRT�.���"�� �6L�a"O*4��A���Q�5���j��"O<��dA2���3��%!��u��"O�
'D���lh�#I2'lPdK�"O�̹��/v��;#Ixe,#�"OR��5�LVdЉK�=@$,�!�$P?aI.<ڗ�?�b8��}!�$Y�c�Da�rE*d�@�ġ{k!��M&{a���J��<�޴Ag*�!��L�j��� ��4z��<���!�ę�>��$�̼.��z�cK3�!�䖣%$>DB�h�-&���W� 1nq!�d�0j�R�ٰM	�o\�E�DJ	X!�Dǎ6T�3`�� s��3@�R%`O!�d�=D�6�Njj�	��+�z0!�$+1���E,�9Tf�i����A'!򄅝\�ʜӀ]�wXf�Ý�8�!�$VKp
�CM�	<��@�شD�!�DC0U�Iڒ	įJ�<,��JT*!�D
�\����Ʉ�k���@����!���X?��x�A�,�������Py��N	�=�Ss7��A��Q/�yRL\� xԘ�J�:k��i 랔�y �1�d���#?���$� �y2j�%0]�fcܢH!��Qb��y��`�4�i���<�a��ݫ�y��#Z�L�۷G�0�d-c�I��yBf���9��C��B�RpM��y����1ۘ,�`��0�x|H�
��ybC�7 ����eU,)1h��?�y"��{����sM'�0��l��y��	�l0+��^�8�&%�&���y¦�'ꮐ�'Aj����k�ڈC��'8����,U��-��fW�4ݬC�I; >��*�e��=;ލR ��4��C�;Y.N�ɱڊP��$�w�M\�C�I�G֖)q�\<>���@�1�C�ɣ/Xh[0$V*3��\�ǉ[	15�C䉽W��q���uĨ2�ڐ6��C����-�,R%j�9F�W"
�*C�	06P" �e�¬p�>L+� �$!C��=�B	��F�T>�����'BB��b".�*���}r�0��i�&NW�B�	�Vc�	y�B�5���3��|�C�	�}���Y0��)s�N),�:U C�	.%9�R�LƻMu�@U+N�C�	g}� "Be֬M��uLӉ?SPC��M� ���k�AتLi6샶e/HC�I�<E$�&yЌ��/���B䉓�K�/"�$�aƪ@���B�I�X�@	���BN���I5�tB䉧)��u��6Y���E�F,n<�B�I&ڒ�p�+�-�����?<TB��%w��@Z i+�H���J8�dC�I�9���,�;ԩp�Sj.C�ɧMp�1�i �kո�(%�@�r!�$�9�4�#�ᆺy��E8ĄT�!���	R|�W�ƃŨY�B�� t!�R3�:�c��[�*�h��KCsX!��@�遶�P+l�Jd�Ip!�$�"1��P⦠L�~j��B�MV9vH!�B<�RC%+6Zh(��a�3�!�D��
�نʆ22��c���A�!��6:�R��d�Ơ�#�r�!�� 
�h��Lĕ�k�K��<y7"O*����4(���i��)���iG"OV���
���!H/B�5Z�"OTԫԨ�G��0���d��Q"O�5�
@���=���@�X�Ҡ`�"OT��B�6j��S��ؑbJ��c"O�hc�a�>.���k���%sP"Ol��f�9f9<�yb*�:t���b�"O�Ҁ-N
kDA�牋�X>�}"O"B�'KKY4Dp�����"OZ�#����
l��%�'>�XA"OL�Rg`0C�BT�G(�n""O�e��E
(ke��Q�޶�^,h�"OڴYK@�H����a�+��%�D"O�\CՆ�Z��@"�K�P� d��"OhAq3ǦxAB9$n==��E��"O�l��	n=���P�n�I�"O� �)��Z����_`&���"O -P�fvɛ�Ȧt�����5�y��5Kj�Wm.t��Ia���y�ɘ/e��-r ��s��YJ����yb�W�,���8�*B�?���3�+���y�EE�D���Û*:�ά@�	�y�ꛤ-�,j��+[D�˦��8�yR,�L���86a�B<*5NJ�y��Z#r��!I���	%�H�����y���lD~IY#%W���Y���?�yR@�&I�02����FU[E�[�y�L�9����#ҲR|�)���+�yR$�*<���c
�{�J�����y-�i�䠐P�߉w/�[����y��������RM;uޑ�y��*s̤��R��B!�AGܿ�y�\k"�!��=W��x�%�*�y��Hd�����\%S4���y�)�I4*���/^�ٹ� M �y"���Mb@��!�7kC�b�Oځ�y���$4,x�ΠK6��r`@$�y��^���R�M9G����1&N�y��A\�h���=��Ғ��y"�2Pz���؛d�ƀ8�LZ��y���I����[QB`ecClD(``�B�I%>JE�&dZ&T�b��ᦖ�>��B�	�w���#�,rPI[ʒ�y��C�	�D�J��`�:o�@]�7gܥ}WC�	�cp��:Fko��1c�Ā��B��"�c���5�1e�>(�C�I�v����!~��ieȜ50�nC�	�j�f(D1Gb�91�)�z8C�I�
��	W-�>'r>5��[���C��r�v0�5���B:-k��Z�df~B�$*�~��Ud�;{F��p���sN��0o|d�S��C�`�Q��m!���;-p�@e��u¤���5X�!��'W7f|�G�A��93c��e�io�C3�<�W����?a��?����N�O���s�4�`�
�^� ��Ũ!��������G�$d���1o�R��p/ho4� �LB�l��㟘SE�ˋXK�9#g✢0k|�I�!�1oc��y�]2E&�5"�Fʀv��݂\���J�Z�8�OT�ŉ?m��M���۰=�Z	CѲi�<1B���?ل�x��';��xB�Ԅq���2���"���=1�Y�d�'������r?	��7M�qz �/	�1'��pA�7-�OdEo�şD�4�"(� � �Ҧl��^�KI�r=���I�9{��i;GΓ��`�	�(������Iޟ�j��;�$�[�'Pް��SAU6`���Ӯ�BzR�#�Mţg�ْ�4oMEy���_��iD*דtW`�faK�1�^<` 4/q0T{p�W�Vhs�!��ѡ��=ޢ�OD8�5�'Ǹ7�L.�{�#�.h7¼�〞!�xkN����ʟ(�?%?� ~	R�D0����bc\�m��ڢ�>!f*G~���
�,�{��^6�h��Fa�:?T*����i�6͠<Q�o�z��'{�Y>]�!�4k�0��.m���N�2�`�Ißd�	�g���0b.R���I�Y,W��E�O���N����S��!ḫm���C�O����!R�+'�\��H��|������j�d(G�_�ACPf���H�/H��'��#��rl��.}ӎ��>�^�|Y�V ��B#����D0F����?��S�D�$<K�Ȑ��ܱI�^\�K�=��z�Cq�&�l|}""�_�Yq��C�oJf� ���n"J��vb�T,6���Op�4�b���Of���O�6� �C>�E�'�1�~m
�J�8����8Q(%�D�O�;�)2t�E)U>i�S���JD�kB(A��ks/Q"�M�7G������C�N ����K�s��+�8����y'���=�Q��@ԋm#,����1a�<���O�Ĕ'ƀ�"��������]�1����K�5h@�t�	Ҩ	*�' ��'��0Y�%��Of�ۀ&Ðb��sL�4��9�M���ig�'1���O'��#���4��h��x�
`���^!R:��D̼O��+�j�O`�$�O����ٺ��?ݴy`�5�&�ĂC�<9�B�W�yW�)�����W�ܠ`�H��F<Q
���yav�ye����']� ��� Pl��F��f�����;b���W�Zk*]�$G�u���Gq,��ƩV��<���$Ey�\�H3g�l�ƼoZ�Pf�dͫ]iF�%���ɐ�u��x�eET$���K�,#V�r��=�p?�O�	�qaE?z�@����Ñ3����Ǟ��M�O>y��i�\��h dG�M[�4rf�X�r	�{ݔd���Ju�}!�'h��'��	@�' ��'����˚�6j� �FşM�
(�,�,]JZ���B�L�荻Gz�p��Ⱥ�(O(��NN{��M*i@�-���t�ڷ9[Ѕ��O4 �d�B�LN� c�6�r���r�	&%B��SѦqIT�^�a �� �������<Y���?Y�������a�~����nA�d�A-W|r y���g�O�����# ���Y� T�>�>�Iѫ�+�4���?9����M�9 *  ���c�%�y��Fgf��cm%*��C���y�JK(1� �ȴ&�d�cr$9�y�!� \Y����,� ��Y7Ε��y���T*�#Ђ�"nht�q�`T:�yb C �))��_�b�}�'E��yB��<B���a g��_�P��G-��y���G6��[`�������y��̻X��%�R� ���K��y"���(��[�蟰D8���ի�y�ў#"`��lR�;�� J,�y2hE>�£�Ҿ7`,�3��y�̕�0��X�q&Ŷ{��I)�h��yBӰ#�a:�$�w���+�.[$�yB�0�pə��Z� 9ٺ3·��y2�āi0İô�)����q���yr/� i�2�c�	X�
��I���ڐ�Py��_�t�v�z�jJ�E6����UB�<�t�]�%�Z��B�_:��5��F�<!�E1	9v�w�Ҡ9E�X�<9Į[�G���q��P�<�`2EDI�<t+�61`�`	��6����RV�<�g��4rj:3�}�|��F�x�<���z�Vx���$&X�ԸA�Eo�<y �N�%�i��!H�~F����i�<�P�wk�] 5/R"(�.̓�\�<��R<���a&V##�8�!�@O�<�1G��@۔1eB6)�P$*�HW�<Q`���|�sL/ּ���JBR�<�����b��'��8�H�w��L�<�wS�."���1���%��S�<i���"jɫ3 E�(����o�M�<���1@XzLА-�,nLtp'�F�<� �e���i� ��P�H޸�c�"Oj����"`�"�B�~��A "OV�sC�
}5�pH��;Xȴ�!c"O� CBJ��
��0���	��8@�"O���w�HP�Ƀ���+0q��"O<t�DÙnpu��"((�JU��"OH;J�1�X1�@'H�yD�"OԠ�n+<҂��׋�L��7"O���]<@�ZQ{�+�_6�1pT"Oبp#��@��m�֩ܕ*j��&"O���m�oL>����ӉK@���"O~|c��#*��BT��2����"O��Ѳ�T,�����Z:��v"O���Aۻ] ZX��J�`�Z�"�"O���bC�Nɪ�{4*ϳS�u�q"O ����p�̨�5J��p�;c"O��bb@��[^�(˖�A&-�Y8U"Oz��+@(�R��Lk���#"O$p�P�L��B���	�3�&r""O�J�ԲL���7�����T"O^\P�k�5�y�F�Ƃ���2a"Od�:��%��<5.�S�^z1"Ox��#�Z&.�ت�FڲK�eKQ"O$��(�,>ͼ�;g�G�z@��"Oʕ�%I!!�0.{�Q)%"ODx�5-�1��U��GĖ����1"O��Y�L�?�ΐ�ƊZ���P�"O��6fD�!�*8�E�bun�V"O�[���9A�)j.$��8�"OL���Of��L�en �q����"O<���mx����5	���a"O$�c��C�i��u���U� ���8&"O8$Y �2^r�9�c���Х"O�;t�Q�����	�Nw��:�"O�b��)!�Rp���Ⱥ'��9�U"O>	��#C�s�24ص�˹;�<ġw"O2q���I8I:�b���:Sn���A"Ol��E��7o�p㶨�4jc��"d"O|�r�'��b@���L�DO���Q"O��q3�͋��(��,ե>]�|1�"O��������݋g��<94"Ou:���<v�~\Ȅ��P��-�"OrA� �z-@t2u$Իcb�r�"O�=c�m�����Ƣ�)�9S"O�L�b����=�bB��2k0"Ozs��\x�	0 �//�(H�"Oh��f�G���Z%�;�z"O�,��+{��d�\��B�H�"O�Y@��P�R=���,v��E��"O��Z���K��Rq�j��0iS"O����H�I�0y��cS72Ǽ�sf"O
�q��ٲT��j�c�!�n��"O@�C���� P-��_�R�"ON��b�ҍ����7��		�@qu"O���֡/{���,��cb"Ox��ș/�bّ�R)�ԉ�"O�2�̚+	4�b[��b�(�y�'�2F��x��� @�izA'��y�m��CpRl�k��e��Ạ���yR�A�v=�S-��@ѷ%Ƶ�y2���I�R��C�*Nm����	��yi�{.虅�
�<��� G%ˏ�yBc�H��dB�#4�X{�D���yr B*T��U����z����oT1�y
� ���j�5[�t�1rn� Y�
��Q"O��w*O�N~�X���.n����"O�X�� k�D�3��E_U:Hi2"O��p��M$����ϙ	N�#�"O&j�Đ�)5�À��hJb�"O���+J�Q���A2b�2!P*�"O�!R�- B(I�@�r	Ѥ"O�|��9Kp~�Z���s��� t"Oxa�4��U,�b�/\$�ҴR�"OZ$[���%&��s�2Κ�s�"Od�B�E�nn�s A�5?���e"O��4�/"\�Dc��[?i���{�"ON�� ��(xp퓰Bq��"O:���у 3~��눘Y"U�C"O9xbB"�U8 $��1oh� "O$�*wOY�M�x�"�%f���h�"O�3Q%ֲ&��r ��/, 8#"O@�f��?N�P�+ ��.5�]B�"O���ئ{U�4���Z�؆drd"O2�i��Ơ
e�us3�W?r�ӄ"OV|�`��0q�*�C���:b��"O�)�FV�(Z�`J"�Z�|C0Z"O��ɑ�#W>�qd/�<��"Or��Oԝ5��!�gʴg�iX�"O����|����F	8{
hu"O�%�тA6��;�e?�p+�"O����h�BV���bdQ�A^��"O��rW@�{`v���?"z�j�"Ob@�U�9sQ:���~+T��y�_�s�$h2@J).�h8ɇ���y��d�0'̕�V�*��@	��y�'��lzL�%	�d��Q󧥚�y����v��,Y���
`���"��y��\����q(�<��c ��yR��_	x%q�B�"�JA�bm��y�nV�y,d#�k�8�@-����y��T#2��@--�0$hU��y�L׾n����Ĕ<B5.��C�T��y���2?�ʰ�����#�Xu��GY��y�L�0� ŏ��T��3���y"���my&��u�uR�Ο7�y�E�w
�أ�M՟~X(ŉ�i���y�ہ/>�y�$B:�h�3P�J�y��ޫ4�����.�t�r6�H��y"�M���:b �7�2u�U�;�y��D1aR8�;F�t\�"r�A�y2Ή�a���sc*W�	/|T�!"��y2��a_�����
�\x!!Ԑ�y���J���
��/?�j�D�#�yr�ϥF�~0�բ^�}�L� q�Ɂ�y��ʥ;"P��	W�hX�1����yB �<\\%���$7(����y"�� E䰃�
��7�K�y�N�����H�&�($-P	���ѵ�y���"v<
�	#!y�M9��[?�y���:	���k�\�Y����y�C�1A����B�b�^�QD��y�i��L{��R^�X|
d��.�y�`Z�r��`�IQ�"��hC�7�y"8E��	���C��]q�I΋�yB���Z3~e�,C�u���_�yBJM�{a���'#��B��1L�1��'BP3�e��?����ADϢ&�"|��'#,XVφ�$̼�
T�  ߖ1[��� �y��/�>�d���M=S/��S�"ObiBf��Xs��"-�p
qf"O�M�ƚ�Q�q8��؉QR& ��"O�x#��?�l�'e�7pX��1�"Od�r�J(*�bGm�4$A�1��"Ovx�V�^�:O��QAn�**6��A"O����	HQ�e�D��(Iw�U�s"O���E).8���ρM=���W"Oz��]
r��3��)�&"O��굦�7&n��J���0����"O|��B��
~:���%��!�:�"O�!�7�ǵJ��"���8�t���"O^uр����j�����"��"O|���`7��Z�|��M@"O6m{rg��0�"B!�2)+�s�"O����ƨ|Ʈ��oO�R: ��"Ol��R�ߥr��\�An�){�D��"O����.�np�c.�>�*�A"Oܑ����`���80��y�0\hG"O~!p�֖`�\ղ3�ů(�20�u"O�w��~-��j��#pzDP!"O|q�%�p7 �W*ʹd�å"O��
�L	4O@L:��N�H)��"Oj(Ň3�2�X��B"��y˗"O$<��*ۓs�M� �Z�}+�Tr�"O��D�_�Q	�1T�J:+&L5p"O2���IGJ"T4��
�BEp�"O���[p؂1'
��|�"OPa�2#�)#ᩍ�u���"O�bfA�	24���'ܘ5"Oİ�L� Sh�M���W�H��D"O������i+0�c���m��q�u"O�)*�τ4��t�O�#<�N�[�"OR��dAHB9S�Mڞq��=�"O,��j&Q�8xZ��^�0����"O0�L�<������R�  �S�"O
5�v/�"2f<#�S
6LX��"O`�!��Cń5�Ʃ������5"O*�H�aM�`⛠.��(�\Q ��,D��S��+L26�ޏ,5p��>D�t�o3j_�����&&X���;D����ΝLm�&��?v�*t��L>D��k� �$S�0�A��"mN��!D����Ń�1�\��TJG�p�@�cc>D�X�RM�;tB��"Y�T�4�<D�p�2J7$.��V"��"M�3$<D�t@�e_�<u
 �C��Kl
��щ:D�([$�H��lIƁP������8D�Q�˅�0��8C�A ��AI��5D��Z%NB�ZwlH��ʌI����1D��G��f��m0�M	,|���;D��W� 4J�Dm@u�E�Tة�,D�d�ggR�x���������=�k4D�p��@�O�F��J��G�E��'D��Q�� 
=�V93aÑOޞm��$D����-W���Ѡ�����j�7D��P�Bx�H�K�8.9C�0D�Kt`AAƪ�r�H"7��Q6)D����!����;���S��`� g'D�l�F+\Е�A��g�a1�)0D�,ó#	�(�-Kc�D�j� D�"D�$	�h�O�d�)�Zyh��!D����Ði��P����vX���4j3D����βA)���Uh�-(�U�%2D�� �`��<��B"�� E�Jh�5"O���@�- �.tȢ���9F"Oݑ�F �_�h勀^�{JH�ڑ"O6q:Ц*J�V b��C+T�0��"O,��3��S��q���]�y�"O���@�IVi�P@b����j�"O�azB֋����&K����"O�89�,1*�8*������B�"O�X�#'�i�4⣅��~�ZbC"O���u�]�4�0!
��Q�j��a"O�� E`_�b�H fl��np|�h�"O��F-�
,�2a�c,�l�T��"OE���Z��+FK�J��h��"O��RbI�l&��0]���*T.�%�yBף9T9�C`#c���)��W�y��V!qJ��G#�o��r��5�y	�)$\|"��2]��A���X	�y�<i��iKOt�9���:�y��@�|��!E�>a�!
D�B�y���b��Li$n�/pҘ d
��y*�<�ܙ�@�^�0).�{�	O��y҇F�M�bq �Y8v��*��ǃ�y��Cn��幁�D�m7���B�y�C�L��e��K�=T6�p�����yRN>(LLA��[=j|y+A�O��y��/Q�t"lЯaap%�����yb�ƚ ��umJ)Sq0Ɩ��y���r���թ�9Lۀ,ZF�I��y�AE.K���84NC�<�j�X�GԢ�y���!SP����1�f�Jح�y∓�2����vJ;;��E�h��yb$�\���7'(-k�r��y���0-�q�dCɕ<9bȓ�Ƒ�yΐ-US�����%j( ��,<�y�n�&�dm�K�D��qqK��y�
����
�#�2c)
%ȐjE�yB/S�I������&VA�1%CO��yB��7%I� +���Q~f)��*�y��=ttI"�׽Oj�=��)M��y��ƟG�f�8 	9�x8�(���y�-��-�&�h�) �6���!�jU��y���4�D��f�	<Z��-�j���y��Bܠ�aK�L#L��A@H��yrMY�	A�<3��.>n��5�*�yr�B
��@kw@X�)#��Y�c���y���B[`��t�<Y-2��T*��y;Wi.�@�.�%�]KuϞ��yrJʟ*;Ġ;GeՁ��Jp�*�yHۨ+���(�$B��r�͋�yo��<_,HC�[$섐%Ȑ��yr�-�hQ���P�)M�ـ$���ybf��Z}E˶���>�!�K���yb�G�p�Q�d�rу����yB�
��ySF� �* *�$���y�e�8��D��O�A�6���L���y���7E���:Dî=e8����'�y�X�{8���v W�<� ����yb@^?v���ߟ/�*	 �D���y�$ۤ.�1�A��Ux�����y���
1��1��ۻ_��˂���y�\�yk��*���8SI��0�#��y�c�A=��R"c��JcPa ��0�y���>\ �H�JY��jB'��y2��<\��!�W�
?���ǝzcZC�)� P]4�)z�ڰ`�iΉ"�8�a"Oj�ZPm���අ�(�0k�"O���s�8�8�!o�8h� ��"OJ���" �=�tj��QT�L�s�"O�9�mS�s�X�d!��s�\D8p"OzM��ھt.a ŠŗG)	��"OĤ#�猐�8xP2���Lrl�y�"Oh�����5n&�툶O�>`@Q��"O���7�9�k_�U�ܡ�T"O��"R�R	PI��E!�>���u"O���E<rM˓@вn>�@f"O|�0$�:݄�����"||%�"O�,���A�A��`b4�Ǚ<󢅘�"O�D`�A�Mءqw��4{�n�A�"O �P� !з�S�v22yJ�"O���n[�%��Eq ��%-���"O.�X3d�<X0Xe�&?$|�Q"O�T3t�; ���c�TRp@Y[�"O�E��͟��32��=x�XC"O,�'`Ҡ���ɍ*���"O�ض�ƴ����\��j"OZ���6D�X�I��E3k�>���"Oح���]�4f���ʍ�.}��"Oތ�g��7ͦq�G�I ����5"O(|��DR�AfXP ��SzdE�"O�*��7c��% �d�'l@�x��"Ol$��]�5�x�!�"o)F��"O:q�D�B|�:E��m�I�4"O|y8��#T��ٹ��2U��s�"OD8�#T�F.q �G[,�p���"O�E�t��%8J��R�B�@���U"O����n�'1h݀A녃z)����"OP��&�Ip�dӄ�O	r�z��$"OD�)���ԂA ��-PX0"�"OP�b	W'Jz�a�(�j���9'"O�a1�
����5������yBc�+r���x'�٧4��{Ӡ�%�y��G+�Z��&y�x���'�yR��9S���Wݤ��}��̵�y��_�u�)�"�S��@�#�T��y��T#9��@	� C"AL�,��y䙛y:<|1G�S�$�@�c+���y�F|>�e��Ƴ!^��B�y���)͢h`a>.L�`�a- ��y2��N���0X�uP� ��ybNH9`D��pA/R��Am���y2f^�eD�H��w��ɐŐ�yr�LL]�, ���o�hT�^��y�`�=8����df�R�0�ۏ�y"�U�mǺe�&���v�� 3��]0�yr+�7q*�-�V�˒W�'�ω�yd��.r(=H6�`T���.�y���kCh0h&��V����%-� �yO�Tsl@ 1h���x$�s�S�y��6":��W�-xU\���ֻ�y����zD
y�0)§�$h����yR�1��Z�A�?�XR4�J��y2i@)k
°b$I�xv&|��-�y�혘"� &iنd+j��&�D/�y�C��64f86g �q_H���'��s�͛�Vu�Eőp��=�
�'�6�y�a; GF�@��@5n��5�	�'�b�ХN�!x*��s�kIl$p�0	�'���K�n^���͡��a �L���� b�襥��$)�`��!O�6��t"O�H�vhǆ\�j�7ϔY�!	"O�-� �Om��۷��)6��i�"O���	He\q҇�ϩbpfe�"Ob�3E��%�&43��Pz5�T"O�<�#�ٛSQ\��s+�:"O���ۿj�~�:@-�:��,2'"O��s�*��"(�D����Y5"OZ�B�-��6��t]<(Ǭ@�s"O�qڗ,��/��(���>M�����"OX-��Ǘ0`�<�`���le�Ј�"O<��T	�}��rΜ:tb�V�U�<���٧�b��QJS���[e$�P�<i��2�ؙ����3>���1 G�<᧊�3�m
%o��~�"7�LD�<Q��B�d��PG�~R���UW�<�2(�S���ɗă�1F�9!Ai�<�V��}_�����k�4&�h�<y��(�`�9��ɪf�ER�C`�<�Q�S�m#r�6.��6~�	B1�r�<9���$N����aG�*-����OV�<�qe�8ή{p�s��i�[�<	�*	17C��{���6�@�K�U�<�����#\��[p�(��&�J�<���>Zh@%&�]�A��l�<�3%��3���eX��^)eJ_e�<1v)�8s0}C��bJ�� ��d�<I�e��I�j�a�D�q(�v�<I���t
�]��!�3�|���j�<��:vR���B[8x��ʂi�<�f(�
&^�<�"��<��W�I�!�D�<T��$J�9UȎ`8��Q�0�!�1mĸ�Ԋ�$v��}�Ba�p!�$	1NdA0W�D�W��q�mO
q!�d=k|�,z�@2s8�$*�L��R!򄏂A~�#�8Z�\���� T!�$ύG!4�x@O��Tj�A�c�ܰz�!��V?9I��@⨊*L^�j���a�!������Xa$�~?
:�&ne!��� ��%���M�_1H��,�46�!�$	`Zl��NP�(�`��Л�!�F,I]�0cD�*�4bT�d!�d�"7X-'FT;��0�+�p !��ӑl�Ti
�=��e�u��CJ!�$�r�����fY����3��B!���<���� kΑy�'T,%!�d&A�@,a�"������ &!�d�5k��4��,i�&�!1��3t�!�%k~�1�faU,m^"Dء�Z�U�!�D+4�]b����Cة����']�!�d�4/�$董�Z�%B
-HU�Vc�!�٨����4	��n� uJ ѻl�!�	�Y�4��\�Tw�]�"eۃh�!�$R�er��j6O۝2����\"�!���7	p��#d�lD��+�[�!�P��(q�.��H��ڗĝ.V�!�D'�K��:4{zi	Ɂ�Qs!�-r��1(��^��z�H`c!�[4�8bR�8��I�DHۑ_!�dU ?����
)'�pi)ч�3=m!򄊷zF,�S�� ?gB\@�:6�!��{���r�Cܧ+/%�f o�!�#cx��݀#�ф��!u3!�d��,�l�:'G7b��	�F�ĜoH!�� :��Cƽ-nN����,��s�"Op���֛�0�A��] q�8h�"Ohܘ��L�)"��1�nސ�P��"O��JB�φ"����&8O���"Of�!Tk�{�a'ŕ{1�u��"O汹�F!0�b`�U�Q���"O�����-
��T�,,��"O��n���3�&; �b�"O�lpf�j�&e�d���,��"O� u�\�)����t�Z�[�"O�c��h���Q��U�2�9t"O`�x��5SD�qMJ,��4:�"O�MR`0ec��M^"���"O�eu�^7D�qK��^�*S���w"O��gϮA�������4Mj�"�"O|���Ӳ�Թ9���
F�{�"O���l�>gl�MѤ$�2Ή �"O.�pW�ƄGY�R��&m��k�"Ox�	�b�k#*�C1kSZ1"O�XwCħj$y�$f�&��@�b"O.؛5%ܡ9��d�eB9���"O�X��5L�E�W�M1j�dqab"O���6�]l&Z��l�.1�t)xR"O�$�$I��}y��� *�Jx�9#�"O@M��$�
}N���i� kQ�s"OʝR�%�W�1�ei�*g���q"O��Fֺc�b�[�S3QJҷ"OD@��u������)O���"O�A�� �C{�����lHzL��"OZ}���#t`5` ï/4�@��"O@:u�ռP����n9=uT�r�"O�q���Z-B�#��_>7f̰��"O
}�2cF�#�I�բ�MfJ�˗"Otܰ�O�g���	�G�b[B�3�"O~u9�-F�ei"e�"B�1?�A��"O8��@��'�J��惂&5,���"O<=R���)_*��v!�</��u"O��VK� 1w��Q�W�A�$�C"Of�2Ǘ[.���A2L%�3�"O�EDI+2�p�ن5%l�0"OEI��V����,V�E��"O����X�"Ӭ�"��1`y�"O�,U댨Ac$���ʤ&�8��"O(�(0�X�Rd1#o�1�CE"O��p� R'E0�]j�͈q_��K�"O�)A��9j�����Fy0�C�"OV�C7�Bߊ!;RM�n"�³"O������+�:�Z7�O�3b)k "O�x�A��F��y�êPVh�"Ob ��G�vO�����ԬhP���v"OU�R�$QĤ�cq�G�~1��S1"OȐ��f�6Ɋ��c�@'���r"O��6�b,8�e"ݍ,	��Z�"O��`��
&I�	�����]��"O��#aO�&ƭ����>}H�P"Orԫ�&�;u���-�T��#"O�����[�k)��q,V8NN>��S"O8��i	�2� ���'p�ܺS"Ol9����d�����]O~�� "OD h�ҬzHf�1�*A�Yʥ"OHI�r��$70HJC�*2R��!"O�2��82�,#��O�0�F"O��8�����Ǉt���	A"O�e��T�~�8�'�eט� R"O�  ��ņ;G����� G�T@��"O� WOE�cl�5c�hƹ�*Ij�"O�����M�Y����ö�׬.����ȓA�$JgCJ)X�&Qwb´�(1��HHAP�dE��`s���Tu����E=�,@�m܃F[h�˂C�l��̅�2e��IF���P��m��#B,hyj,��Q���A"�(z�Z�)A��(B�� A�!�։�H�z��o�(Z�X��ȓQ	�q3�Jٰi =��c���ȓeh\,�GM�WʙJU��Z���ȓ\�D��K6)rL�(
׈�ȓ~��u�n�@�N�s����-��*�,��0\�3�h�(�|I�ȓu��%
��,b|�p���+��=�ȓx�\�TΞ�R��q��Re|Z �ȓqS�|�#�U9<gX�¦2��]��8XĈz��
y�p����B?�̄�f*������z�J�u��&R`��ȓ�m�5���E�ݩ�m�z����ȓN�P g�W�va��g߲�>a�ȓH[�(C��о~A&L����5e�����3`���ǟ)i�8)�N/|yԅ��<��`HV�i��aq`�5P�h �'�60OPc�|�=�v˙�l\��ɲk^(��@(�y�<��'D���1"��2�QQ�Yy�<�T/T,���B�43�v5�7Ywx���'� `���L�B�^ly!$�2t"T��'���cӫ^1}�҅���#�l�ߓݘ'�R��%ΏV��1�"��<�\��'�f	)4o��WmD�!�/GhF$�ڴ�hO?7�Q;]+�ux@R|ahL����c�!��1Q���VB�� Ȁ�K��8"�������m�b�Ti� 2BaU�^oB��2 �RL`��t%������[XB�I��t��fL�{dV�"�-k��C�	?#�ȰЈ>�>5X�D�2;!�C�ɢd�f�胪�-{�x4�_�(�lC��
��,8��;cќXۓ_Xn�C�	j���eI*s������%�|c�X��I�4�� w͆ur~H���N850>C�|������H�	i#�.w��C�I�b���*��SWI�v�B�I�j&Uy4�S8��h"r' ŰC�I]@D����U���2�Љ)C�C�ɫ�>����Z�K��@����U�B�9۶L˶m�=9��h[� Q�! ����������bk��T	�1���X�5��p+ԓ�yB�КZ5+�gB ����;�'IIA�- =�QgȞ ��R�'���G���<�7)7`2�1�'1�}A���2pF�!gc�7��x�OV"=A��)[�rl�p{ӊT	xಘ�H_8#�!�^#aB�`V�S�V���pd�7��'шIEzҚ|B��(��3���_�}�!F��yB��!-^n�:���I3�	����IE���$�<	�`ʜ{B�3����ǭwy��IS�O�=sD��V���Ж1�$���i�����,n�TE����Dp�ؒ����'t����58k��kv$�U��Q�A�D@!�$��.9ht�6�C90��81��S&w7!���r�R�	�X<�#%��ZW�x2�		)�=J@JG'Br�`y��ӼH��B䉡Cb(���dB�=vt����1 �"=�#�π �$�F_w�&p�"@
NOB�ʔ"O�(�@��P2�i�TA�$�� T�����*�j��X�f��,�"�)�F���y��C/J�����	�,|�B̤�yr/J�I�n0���8ȴ��K�	�y�H�7�8u��cȈ0x� {���yr�Ǭ!����ED��D!��o���y"g
	L1V�B�h����z�팔�y�j�;1T��3�#@�
�p��瑦�yb9�R%�`҃�`*㍜��yAȝj$4Hǌ��ZHa���B��y�KA3j��WH��q*qС�	$�yr�"P��T��T;����`ݏ�y��ŀ�f��i�E�� #đ�y�AD�m�*8b�M�C���"
-�y���f�|Q	:I��Y�朔�yk��|��dDܿ���Ň�x��'mv� ��H%|�H�]����"�'�B�е]�~ŀ��+R�Nj!gۡ�yr�Ǽj�Bu�!E�6��T�����y�ݸz�f{�R�+A�ՁD/�"�p?a�O�	+'$�v96Dّ��-"O��c�H�=�\���E46���c�"Ol���<��U�'�k����'�����L�#�Ҡu"��@϶7�az����X�z�j�'8[2�,)�.�i
�'�x�g�2Zph*�D�DL��'����A�֙U�¬�v�O?"t����'@±c�ǅ�<W|�F���x� �'��Y+����;2��Y�|_~��M<�
�i�qQ��%_{��@�@8����}J��o�<�Q��K�=X�U��`s�	R*9d� ���\:C��E�ȓ��d�!A��{��壳%	�5�m�ȓ+v����ي[�hE(�T���Ԇȓw��i�r�ͺd#� #�	5Y�ȓ�n|s���?�X��1	X�^=���	L�غrDF0Ab���n�,R���3h�8�P3|��) ��E JՅȓ/|$��f��C�i��=8��ȓ'�pRa� =d�51�m��r�&4��ThBy 1��(|��S�@Ҫ���I�)���Fzx2(]8VU�Lk뙜L�6B�I W� ̰g�('���$@V�k^*">)��I�
���!TbA�9g����<5!��<n�*ps3.��b��)�6'R�O��pG)ǉNŤZ���1��k`"O�0�7D�,B�rM�ec8$0ra������I7Cw��򊇶)��gA�I��C�I�[��Uk1Ό�s2p��p�N`�C���2�+�gĵ0C*�c�N*�@B�I:bY��)��Yl�*QQw�2B䉻j\x��©�,X���M�&��F{��9O~�Q���B��r@@2?�@�W"O�y�@"DC`%a6��-�&�C "O�1;��C�flنL'M�"�3�"O�]�M$Ĝa� ��-/�}"OΔ�U
bsȽxWH�)c�r��"Ov%�C �5 ?��IuĈ9;��!�3"O>tP��
{������)�"O�` g� p7b�S�`��xQ�U"O��B΄�/μCO�.U�nŹ�"O���R�c�^]�rL^8mb�Z#"O�Ix!�O\� WI�_u��ѵ"O� �����މP``];�b��aR�7"O�H2N΋.���Ț.��%@"O�t{BmC̜I�JL_��"O���g��,Ei�����N�1w"O�MC�L͋""���pcX;����"O
�a@lס���)�:!*�'��O.̑��E��F|5�҅a��6"O�j���3B���x���j�v��"O�%�L�=�� �ʜ-�j!R"O�4�۴�t���H6���9�"Oք�ӊǺv�Xq0�P:F�X�k�"OLH,VI`鱦g�#��И�"O�	��X�@D��s�'Q�%����"O�Xk�ڠ|C���rjFX[""Oh�%�C����*�ʔcF�=�!�d�-T��<)�FP�)Pw�,�!�ۨ�v���-�<)`� �ԦI~!�	�W���	4LˀXV��$�Pk!�$ĈI Pe�$`?�H��%��1�!��oN� {A'��%����!���2\��rh�2X�-`�vB!�DZ?&>^;t�.l�%:�!��V&!����6�ʄ(����JC� !�$ ���
� ��sB��6�!�$��&Q�]�1"�k�^該�_]�!�Ĕ�0hQұAˌ.�2��f`��+�!��]^��LxmBx�m"ao:<�!�d��H���הgr84���D�!�$�7<�"I'�O�Cr�5P��V��!�:F|.�i�_���))kޣ%�!�$ 2~L��)�\��d�Lђ7�!�$	ECj]3��#X�8��u,Nc�!�$R,Q"��ř=c�) &l;!�!�D�~��|)�Aѫ �^aI�Ր)�!�$��|l��(�l�乓�IX�!򄆕t��(�`%K��hI��ǒ�SJ!���e��$S����jtDc�O��V5!��.CP��Bb�5W�\	1��!��Hʆ#�zn��[#�O�#!�L�!�ٲP$�-	�m 2�T>�!�ҩk��a�甐B�`��_�;�!��úe�"�:���x������G�pj!���"~����/A�T/(�	��lg!�D�0.�IÜ**��[r�eM!�54U`y��B�h�L�s�k+!�G*uLu����Hx��ȳ4!��Y;4�:wO���Cg޽ b!�$�|��!Z�$B4u��h��d!����ɛ��
bR�ȦC��_az�芆6�DX��%(a&�`p��)v���G�	&&L=�����PyRa���^\
�]Z����`��[�<yb�ٯ	P@�H� �	��hJ���[�<i�+V�C���˃��$%p�rǀV�<Y �عg1긙� 	�&��yQ ��R�<Y6K�*^"��-��en���"[e�<a4 �*G�0RHQ�'4�0���Da�<��EX�`�X��랱'��i�Bb�<�tLl��1G�� j�t�&�LX�<��k�w��C�"ӾR>��O�m�<�����5n6a���AXw�<)���]�f=;��k��uH��E{�<���B��D;��̇�:�:p!Jz�<� 5$I< �̓37�%ڗfZ�<��Ϟ�Lw���8�<��G�U�<� ����7] {Q#kZ���"O�i�Ԉ��t`����M*W"$��"O�t`�A�O�ezs��AJ�W"O�a`)
1JL�(�d��tn�A��"O}��Y/g2��������(�"O�����F��do�(�9a�"O����"��Eh������f�i"O�aX� ؙ^� 
2�#3���q�"Oȳ�� �����NO�y<(�#E"O�P�����i�.Y��� �"O��V���!���(��%D��Ç=8��t�D�(Jm�A�"D�X��Y�;��򵪟�i�=���>D��r���1k��x�J�)b�����3D���r�ԕL�����X 4�\�*3D���s��%Q~��dKB{�>�pr�3D��˂�/y��i�u׃�Vܻ��/D�LR(X�����*՗8/���k+D�Ly�JR	ͥi�,���NG!�D�*Uor�X��� r���A�C�_?!�D�2yԸ�з(��A��!`AŦ49!�D� W�L{�Obc�����S&o"�|�/�N������)����X�֤�tɘ�0@�m�ȓ[��ЙF��!]�dy��l{�f0�?�@���H���,ҧ�����&�����9�u�ȓ&�,	 "�<fW���T'sD	s �'x�{V�<�>��o�>K�����W�b��H��Pr�<�w�N�H8j@+r* X�Y���}V�x��c�5!�N� ���Z��1 m2�蜲�lB� z�X�(4\O�4�p���.2uD��T�D���O7rj���DR#$�*N>��d�! �:vm�Έ�� �`	�p��0@�OȎ8"$Bf�dH�=,
ƥ�2%��+�)��q8�\��Y	�hD3��I�8솜�cO��q���#x�̙�(�3��	�8�z ��C�v	ןR@�dأ+�u����`�Or�e�s�<�0g��^r�,���)c��хnη_
�e'�ji��*��J\��z2*�Wf@k�䂸2���U��d@�F�3 B4�{����0��	�f�xh�ƙ7d��ʤB����/U�*b��΅S(����܎�0=YWG(^���F�z�$���רu�>(a���'jؾ9c�!��	�MѺi�,A���:�NV$��^=��I�|�0�ag�F<�<���Ć�>��AI�I��=�M3�9.��"B��p��\�u�øV��O���b�)�S�]���!E�ϹM�f�����"9 HV�pq^y��/Xo�B�����$S� �W�ܻ?�ѱ2���b�����F8�$�G�b ���&L;����"{��m`�@9c�x�SYl8���N�'8T�h�!j^(# ��TI�c�}��I<QB(\�U�����q�$�#:?�+'J�>��UG�1j�ay���	9~b����`<�,�A!�x��`�65�I�zD�E+��ܴ�8�u�pExD!3hɊ<�8�R�d�+&�2O�e���z�S�5b"H� o
f� D���еy��@c����x�*�<�3�>Qu.�!�p���툵V���ʎ�U��k�`Cq���g�L���1%�`U�K��P�	RP]&A��ax���&ye����¢$�~�i�#���|�ao��le$ R��':�D��<�G�F�	].0ÍǉV����M�J�'�h��%�0�t�@����t+��#u��1fk�%'�B� wh��yR"օ8n�Q��ֵs�]�v,B��y�F4?�dAs@�l�.T�r���vl�}�2(V(�t o�>TVB�	�r@�t 	P�t6�hK��vgD����j�4 T�8��@�|Fy2oBLSbհU�V�0<F�bA���>i2���d�0��BK��
�S��M�����A�Ȋ	+��@!���g*����Z�^AZu�'J�����C27'ў�Xc� R�Li�$)S�g����\?Y�ǈ8N��x����
@�c�� D����fJ��L���G	B�����O���W�
��ԍ	d�E9j;�����i
h�X��b��w!D�4cC�@�C�	�kC�]I���*O69�V ߮[���F�ڔu_���DR�o
���U��|FyrG?:c`�H�O���bT��ڰ>��(��-�شh�$i���p��� b H��!�y�m�D;���)� �ѣ��H� ���Xv'B�M8�x!�&���F�	#'��� �gC,N>��O�%�v�V7m4i
P">s����	�'��ѳ���r+����k��=��ٽy�P�I���2E,��Y����}��?`d�B�`��͐r�Ȥrg"O��;g�T?6mH�mR7P�,̑a�ar�da���a�<A{�m�-��	
<�`���8��Ȱ+�{1���dï_<��w�5/�x�׸�� `���]6 ��"�ʥ:Fx��	�W[��H�ʙ�;�
�!lI�w�D�?���K����a�T�.z�1�#�XR��_�71BT�c��{��RfY��!�d�!J���K&%���+v�ɤ3��b�Aԩ;]�X*B�^<f �\:��SY?镏 	}�l���ğ*� ślt�<�2���XNP�p��a�蔛E.��(�
,��%��~5`�n�:_�@��� �j}^8��'��*E��N�Q�HT��I?_��a@��)J/2`�"��VXh�Tg��1�ƈ,K������~D�7F�PT2��`1N�i�����a2F�Qw�[>vI�P;����$=��2vc�Z�i˜s��L0P�ߵDj�����3x�!�D��<���8D��+����$РҟtGV����]=w��@1��\�*T��"���G��=�<q���Iȣ<���\#���W��Ȅa�\ԋ�.�6e�����K�7Q��ܐ���?��];v

�O�Eken��Z�R�G}F�3zC8$���B��{F�Tc�0�wC#b��;�O�)ȇF�5���P�r����c�M`�������;dڸ+��U�U�uH�JV�9���Cs|�r덦3<�R2Ϝ8Iw��	�,��tc�/"�ҵ�G�D|b<�«�$6"�R"\8Hv���0�a �/Z�X{Z�@�ꆎ�T��$���T���^b(p�(=aR2P�⍎ ��l��bK�t�
�kօBf!��p��"��1�H�}��C�(28���'wƝ��������QbV�T�yp�{"KI+�,���E�@��ŘdO�������9�@����\��i���az]�:��U���_�LO�H��$R�����<�R1``�@��iFx��ć�`�F)�C�$�<öaE�Mp�fԓS2fp� LR0lXD�P$Fg�Za�#G$V���b��0�t�ٌ�,�Ac�R���B��,�O�!pɾTՎT�F��1p�Ј%d\$���;���n ��`�ʌ\K�8��H�Rޚ|��B��	y��E�%��P����EZ��<iHm���'��ݙ�a�U���3��<(j=X���/>�q���ј!��pS�B�V<���Y\|�Q�ʴ"z!h�e-8�m�'���Ĝ&z�$x�U��|����d�j���=9'	�5UZ����Շ)��8�Ԕq��M!c%ջI�R-��)�%�.l�T�B��B����܌ R6�\��G��Vu�Daȍq-�P*W�H�4t��D�*o��p'bζF�l���-�%iF��faIt&�|K��N�*H�䐨i�� '���r"�e�J6������eE^q�m'�O�����:MX �"��,��@�2��	��ą�,�,���ꏔ/��ٻ ̎;IT<��ɓ+��t���\>�(��-�<��q�g� P@��'b���_�x����M��D�3y��8�����sB��ܦ��poՂD^���SzF��������HP��N:,�7�k?�r�1C����H:�3�ILT�%ą���<(�%
4f��g"t(��[yB��!���a�Asd��v�Ru_2urRό)�Y���i�<�h���g�'c�,:�&��GQ:� ��g]52��Q5��mw
���郌y�aK���8nl�!��L��\&�}Q�N]�z��Q��/2����b\W��x��<�z�ү)c��¥	���a�C!;�I8np.l#ԊZ�[Z�$C�e��!"���B8q���Cab�
b�*��P�p=��BX1� �P$�L�z�ڭ�TH-� �2��n��]���>yD(٦����=�䑰��̖*��Z#ُi��a���O��Ƀ�ʤK6nQ�6�BD�nyT���}����O��[[8aʁk�6V��ǋ	 �yr)��{}R11���Ms�8�GG��u���'�ԐDDP���I�|y�a��XP�'�v�AA	�r�6	��k2hNn�jAO���P7�R�H�L�6*�l ����>�E2OV��G�i�4���E�gZt�R�� �_�� �P/zP��ə=Vj|��(=H�G�"Z�,���Eǔ>��ࠩO��ݴ;Z~\��40v�@t/�B�tu8��
�1s�=��c�<<&t��V)��xIZ���ɉ\l�I�qA_P����
)L�z�͖�6�:���A4W�h����T�u�`}m�w,$��[�[&��e�Z/)`�A"g'£n��$�,��49�@�Ht�p˦�ڰCƱO�e�V��y�fԫ	�_2��͛�o�5���o
v����M�w�@�i�bM4FH�& �m���+�jEs �#aEj`�>��J8���Y�[(�0���@�	��\��� B���)�8h��AjL��?`��,�"�� `W�?Q�].|F���C�
w���u�Ƌ1"���W$,�OH} 3�ɓ�l�A���e�!�S�Յ3�,!@�'Dfi�k>�Fa8C^��9r��_����w]�L�Ѡ̇����҅��p>q�/�Vc YyÁ�,���yE�Y�meB	��Кe��Bo۝Q���F�] ��0Ǝ�)��)�A�-nbLّeP[yr��g�dPFC8C�Tp��.W��HO�虇g��}],��ݢd!�E#w��	V6�Lu�6hYb�{ۗ _'Z�<�!ۡgu���2lM8)ax�H��8��M�b��)	�����?��l%%$���b@̏i,va�G(_&=��aJr��(���BVx��A�s�Z)�� ���+$מ�ٵa˛s����^�a��
�. �=C��).�����\%-��5��@Y3%�޼�R�{��cƆPK�j�<� Bqceb�"v��蚖�ԥ���ۀ�'����L�P+&Xؤ�',͜P�˛5��0J'��JŦL�",�&6���8��Ȣw�<�?�g_5HB$y�$QT��E��]�'v���MB�1��Ղ~b-��{��Q"���*Nm�Q�ƃUu�0�5��$A����D��ko����ŭ'b��1d�z0��>XN�2rA��N������mb���C��$f�ތ0 &Y�H掉`ץ�>*캥k$D���G��5F�;���m3d](F!«�nAI�Õ�%� ��&��g4�rD�mBэ����d�	~]IT�����p�DQ2C�~�� !�U�Xf6���/X�� ��\�4@P�NR���Q���Q.V�F�UσD�'0z���cR�~@��JT ���ɏ���6o�����J�V�ݨedM�0@L��'��M��m�4j	 2��y��%Z�x~H��s<�[뇶l�")��xr�(�'۰�k (ȥ3L�����J���-�������x�KS��lP"�]�woLp��"O��ڱD���0�1�ѐ}ObRQ�O�D�a�N�[��d�!����1�)O�!j��O�pX5���]ƨUOBA���O
 `3bK|�>,C�aZ�I�� !� 7 �J���C3����­8Y��j�@'_����C�z��}��C;x�$ĺå\5w�N1#�ʻ\��=�sk�:��Yc�'J�y�r��Y���(U�m]&E!��ɱ.U��b+@��0��,�LxN,�P�޷$=�ȓo��tk�k٢#:x`���ʰ!K����^���#�}�S�OuByH�LRL���
g��-��3	�'���j�^Hƞ��O�z⎨�'Y��P"G�]i�����&q�p�'��yՀ�3H󪐫�*ˍp P��'�4a�u�^�x���ҔZ'�}��'VX���:.䈣�U��IY�'S�y���/1�<�/�/J ��K�'�V�3g ��v�RÍÀL�D��'��C�cӢ0�S�ĠD�I��'��407dR�����Ӥ0SJ�J�'��H�$rH�y�雫*��(��'�c6�܀gf�	���v�P�3�'S�1Tʇ0`W2`�.�;>t�UK�'�6Q��
Ƙg�l�vC�&����'�.A� �B�z-9�L_�)���'LDl�`E%-�~\xFeޔ�����'}��2��͢@35�D���jIQ�ȓN j�񎖾���0�뙭�<��ȓ
�n1`��{>x��#+U��	�����o�4j�9V� vx��#��q��)08��5��7};T�ȓ?; ���'T9<�\��`j�R�L��	¨(�N�y��	�E� �	պ0�ȓr�*��RE�'zI�q�P�S�u�ȓ��J��K�J��p�'R��H�ȓ��C�Y-A��X!4g�"d��l��!����
8:=A`��������L��t0��Z���-��@hw R�<i��?%&��8�Y�p�:��F�Uw�<i��\-f�0��>G��S���j�<9���\󆐢r'�KN`%jd�IL�<��靈8h�-XDE��k��Lʑ��M�<�(Np��0!-�U�A�S�<Af�s�� 4��W;�B��D�<�7,O8V��ؑo�Y�(���J�<�E��I��)�C�٥:� e���<#H��P��K�!����w��u�<���Q$L��E�֝V�q��E[�<���o�kQ��Z���2G�[�<��]-�6�I��;�T�Sa�XS�<)�fՆ�&�"�+ ��\Âh�J�<���
8�X��b %�>�A"&�O�<�5E]�'�$�� �.��|9t#�G�<� r� H�vJ]#4�I5t�ԹK�"O����W>$�^���hY.i�кP"O�\V%ɇc��Y�Hʧ!_Ԁ{"O�xW&�DZ~�����/�ҐC5"ORѸ$璃;Mp݃hĎ5����"OL�����O'P0��.�3w���"O� �#&�%Q	�99���]�����"O,����J����a��6�j��"O:]�b
M"8V\B�%E.e��	$"O���s������~�(W"O�-�#i��<��Q '�U>\���"OZ���k G�Y��YG2ЬI�"O�j��P�%��cWCؖ�P��"OP8�bᔶNmZ6�H�<s�"O�В��N���� O��'8P�!"O�A�g��Tr 1��J�l�[7"On	�NW� E�)�� H�rZh"O��ؒ�vx�SAN�D}���"O��#i�.Ej����ΧLSJ��&"OָK�3TоQ+ǯИEQ$Y�$"O(�3c��lBt��|D���A"OD5
¬�#4��L�����!:���@"O�uj����_��Mc�E֞:=�+�"OR��/�,6�D�DW2c�|��"OzXqV&S(I]�-���T�.pr�"OZ�����	+���aJ6�q&"O��R�Q:F��K��UP����"OD��%��)-b�*�	=�R��0"O��d�O����:�/� �2�"O�ģ�MH�rqh��F�+n�*R`!�$�J�t���[�g��i�$΅%h!�����������"v�^X!�ė�K��@��ҹ`�-�.A�!��=E�d���,)����p�^�!�d�*�r���%R����w�U�!�D�4��Ի���&%�4�1�FҊ �!���)	D�7
�0V��7Ǎ��C�I�$�Qh� 4STt!�FB��x[�B�	~v~ �r��>E�*��b
�T%zB�	�|��	��;}\=�2*�8S�@B�I-|/��rq!ڳ�,��&Ƣ	_XB�	E�)I�֬@0>��qd�!f*B�	:c#P!@��W������P�!�:B�ɚ(����JXl����;dԪB��EC�f*�'at���v(��8��B䉔u���xe�O��8@d���]�B䉠D���1���!�*�R�a�6}��B�I�{(b���.�$S�#׬��nB�p/�0�ю��&�,���h��S'FB�I�$^�-;gՑ,�Z�g�V8HB�	�Fb�QD`��� ��$F��}��C�I�S��8���z::% ��S%��I�pB 5�N'?� ���[ @M;�&� ��YfK4�Oh�Z�c�7����b �_@X��C��c��8X���.���>].�#3N]�\Ί����E'�Q����E�91�������v���E]/Y݄� ���?��C���\�!��S�(���K@l�Kݎ�I�#�4���(Z;�����XV�O|<� &�;Jje27�@�;��Q�'�R�$�� C���p�����5s��B�8dˌdP���K����I�c��S-ڛ�f�y`%G4����� Լ �fZw� y��
߸F�Zm�%�@	�(Gn~���c�������K�MAO'd$E{$ �{�n+�N,@�R4���D��H݀SC�A����P<�dq7 ��yK�?V�Y�%ǻlAh�䘗�?�#%]4Yij�c� �`G�e�F.�'�� 
�x� �H�Т�ٷ�!�F"O�\���N$�H��Q�Vd�C*��k��Lr�ԑz��5�G-<��3ʓ>v�diԭE;M�@+cM��Z.✆�	��P�qeg+�ʬq�.�8`\+Ah��s�!�1��P��C&�O"�i�	�*�Nْ7�'4��7�	y.�)5iЩ�T�ʇ��$2��O��dۧ��$N��F��)D-8�'I��zůFi6��
��O�7�Ř�D(U�z���#�(��@1�Oڍ{J��}��1ݐԻ�)� t("$�#o��B�I�p��5���'��財��1(�h;�ޣ)�\�9��_
(T-B��?�=Al�?�L��OC�l$"��ek8����K�/�<#Oζ5��7g��2���B�jy�@� P8{qa~�	� ���b��5R�	@U�\��?IEJ	�1�B�b��Ϭ!��x�'@��Ӷ)��P��ω?9��\����#R\!��L,��9Rؠ_(A�G��4h���ł��C�l�ubP7}Yh��+�'�~�iU!~���C*�u&�ڰ �>�y�&Қy?����)׸~h����#�#o.���[z�`��w��(6�y	�fZ�'R@�i����;�����/�����_���;�(@�C�VQ��j��CB%�d(�3j�3�-T�F�8�S���O����d��H���3�O�	0�a��H�.��'2�q8��	 *�4}�)�TA���p�����^��#U��VK��Y֎ߍa�\C�&+n� H���N��HWnߨr�A�RF� Q�L�@��q���:gN0��9|�Ƒ��:������R����Lƽ~��#=�Ul�t�����	G�8�� TBl�9L�9G�Z��B*��D.�t��a̞��Ʉ�,��0D}�KZ��D�� �O��R����P�C�n�O���x�&�h��� '����e�V��*8��\%�`�sOݮCy��G�����=� 4�/��N��в~G��ɣP�ȽC��Ġ6��P�:�> rUo]8�P�a�F���Z��Ů��p7���;O���dS��� ���!؂��t@5��%Ξc��2��(6�2G�0Q��A�H�.e/�x����o��������(�'����YG��I�!�AG��H�{��� Vr ����$� Ҵ`����ƒIp�	񫋈��aA��f҉������ �(ؕSf���F\
(+�=Q1*�j�$���J ��lJ�N�0�&\����l4�(�!�j�J�a�U�]D�ɵSԨ���p �9�!7E��Y��V�w���BѾqȠ#����b�cg�'���R�HE�d��i�Y��kX+'�.i�ɤ+�����j���:"�� O�H�"Iؙ]����+&���,E�%�Fy0��O�\dl�rדP�<�c�֚\��e�"��S�x�1�MP�6���
��̬�ՌƘ�aC��,�$]a1,[�V�v��-P�5���r*RUy҂�7/�){��=���A�����'������;�ET�W
��NN��|| ��ڕ�4*�cW�$���!����䭳�#e5h�2b��5$@ٰ�:��OfA�&��x&����DN%0��C�V�k����M.HC��	��ʹ5ha��gJ-}-�����"?��3Gוmu��b��/�d�e��*r!���K)5[���I�5)쐃Z8(���ӋnR��E�0$��d"X�8���fE�Z��0b�:(�<1���`L�Ӆ�L�4-�HwS����0 F�	%@��n+\O��Ec���j�����K"|�ۗ��z8y�T��.8�J8�ܴz�Z ��"�'O����'P"�Z��O�#$�T��IZ�(�'x���u�7H~Q�$�:b���R�{�0WvL�����,Dw��9+�GS�=-O$�Y���$#�iӷ����|݀�/�EFtJbNZ�{�bmcaK��>�1��L�t�jLy�g���.�i`�G�x�ΠwM s��Q	��b��gM�z�'���qg���&�:���+؀ ��]� ��#np$�0BNS�:��~��.lΕ�
��U��j۽��̪6G�x��X��w�� 5|8����mL�KPYR(˚a�vA�A��q�z��.^Y|$y���6b0iD	T%v�8��k��E���z}⩍��MÑh[�^�s�镦q�"��ƒ��y�u/�>�d�'��ջF��4~Z�u�4�=+�⇊ݥD��9�M����c�,|�󄚑Q ����!�95$��w��6Yɺ5q�B=ܤ+��	��@��l[֨O�,�􊜘X�ܝ�0˘�w��n� K�ҽ�E.��]g�N�D���j][}��z�(
7�`Ӽ<���ۮ���t�5C���;�m
�]Ͷ���+�A�d���HD���J�n��	���7L�b�ˠT�|��i'�i��i���S�Vo�x�K�Cűj�頰��x9�IbW�1�)�|i����IM�bNP�Wc�#x������> �t��D�0�҇[�XF��۴d�F���X%3M�\����=q, (I�+���I&P���A%�8JϠ�� ���:W|c� {�e[�V��D�3�>���B1"P�p�%�'r��7��c���6b
�"LEh�'��~�a��̓h(����UUy�E}��4��=�`@E���I��slT�l�N��P��+�w�����`��(	A��vfbď�uk�qBC��, �9�׌<wO�j��Xg�� S��Q�b�TAr���2��%A�/U0Q��`�O|xc,�R�N=k�@�>�'`��`����:��Q����r���ƈE�)�'xU��D*u��[���.n���*�b����� �9� �L��U1�N���1a��"+~�����e���(O)(�	�y�,�cD��!޽{F�I�;���4�N;n�Yb������h ɀ �ѫ�
К���eMӪO�N|	�A��x����O,^�<��Dk1axb�q'l5P �B>d�|� �C��?7���6�;v(֏W4��y��ǃt,z �)�e�x��Js�l ��]�5��bR�R-f� !Yƭ�>2��Q��g\6��ϙ�&����&.D?0���[�%!���*a��*�Y�D$I-a�.�1s�<��+�|=���ŒŦ(�Qf�Ox� �1���['�C1g�,G�pi@���:m�b�49'�P�Hѭ
Ǫ]AI��+dY�S���x|$[�M"dh�đ�"�Lj��=���� h##��;~:���R�/}�E��H�$Sz8ȱ��-��S�̳�JT�'/�P�e��B�@!�Sm���h��Z>P��Ռ�$1��o`"��8a�I����2�IŪ#��;��I8��#E�%�0C�	�G8E8&b���3�$�6�!���f)�D:�-�8cJ�8)0� ���5���<a�G��7af�D�Ѽ#���t �K����"���$�g�Ę<}PUd]�.�4)�� ~�^��p���PH���nR3X/Ģ?�`�GG��t�ҌG4�k�F�M�'��4�F!x�h� �ɜ:0�v`�3��<Nb�a�VΒ�PQ��1Ci] 6N��Df�V��D(&(��Q�$0���]�9�B��<��
P1bl1��<�!RT U7��8U��df�1H��)
�b�F�V�zf�	��y�@�
��Y�NP�<:�;�E<��� �q�a����S[����Ď�Vy�br����1B��T @'��xR,R"iX�u�t��'Z�PUI3�݄(J -��eܧH��a���7$�]���'��0a�lUXl̰;��2
��ı���Ё�ʊ�T &��AȐf�\Pj3�7i�ICA �](<��'	�Gr��J��E� ��%[F�'��(���N^��c?�˃��+�p4HE�#Cپ�8g#D�x�F*<@oH7���m�՚P���rC R� Ǟc��}��0%�x��ԻN��R�p�<) �ݒ>�ȧ�65Kx�R@ Y�<	�A(@�	�.�R\��S�<�ƌ��=�n(Jᬒ�P*��0o@O�<��O6F���*�AW����Q�<Q��2��m�dC$t�Q��Ot�<7��7�N]S�iȵ?��L�.�p�<���~�+c�O�Nbd���_#!���uW���¯��i��a:��S�U�!�Ď4,b����Y�g�H[�6h�!���]�8`��N�N���0b��!�䊮;��p�+�s������\�!��5�0iH��c'"Db��ެg�!�D��T�A�
-y:�� �2i!�d�:�P}��B�3irh0��L'T=!�D�0h��C�$6 V�QK�cs�!�O)�n������U�z�W�]�r!���9�!:/Ө$zmB���i!��Y�M	��H��4Wc�?0�!�E!c� ����.0�@��Pc֒U�!�dB��"�G��$|�xE��6�!�J$KHa1�V'L�Ȣ八S!�_s������~�&�r4囟k!���RB A�P��m�ju�7BH�8V!�ɠydʁ	�OY/����cȅ�!�L�wQ��2Tͼqݒ�X"�7q!����-9ڐip�
a�j�1�ݮ}!�d\H�H�H��1(���3#C'#!���ƔJ֤�hHA��i	!�O����˓iP7Ѷ8{�RQ�!��O4��E΄�E*�8
��X�M�!�X/ur�����VJ�+��azr�����en�	W�d������L8H�bQ*�Q�D����~(��>Q����'1�xҡI,U>���F�(n��C�>���ͶQ���;��i�~���@5x1,\@t�W�/n��cT���`!��_$P���>%?���"رr�� *�n,
4+�
f�Ԍ�I�w����φ"@���S�O��)�Uf>]��D��s:�5r�#ۂXd���U�O<��S�S՟��O0
8�=0�
s#wdZ�� *�$٣ +06�dF!�0|R���K׎1�6EɺQG�pHW�Y�U��i�d�X�nR��ItԞa�g�)�� ��tb��v�p�0��:8�<i!�xr�-uqz}�6b"���ǃ��YZd�S��D0(�BU�-Odm��o���HM�"}����8(� �J&�D���]hs���5V$\�Ɯ@f�>E�T�g���/��`��907�@�V���x�(���D�v���H�O�t#/ʻ����Ʃ�
iyE;e��OA3��DR>�l${)�}*F��;S!~���@ۿn)��g?���qק��v�1vDX��� #���0|����T��P�&Y�7qO^,F��E������B�M0�y���M[�!�B�>��~*�*��s}Zw��4��[q�؃��s��ϙ�KqO�����65p`��6A�$�=3
��=�r�ޙ�@�D�DNQ��&Q�2�M��(u��ē9�6�A�V�5y�>�	)<&�������̹3Ap5��^���G���S�O���:�--���"K/¬j�4^�A��C���S�i0�S�Mdq�"��*P<�ɠ"F+rt, �T&Q�.��
��>�s�O�n�8W��?#�a�s�{�p�)�Ɇ	sx��O:�{�Y�O��t˙<���+p(P	lxбc`�U����OHd˓�}����?&P� �@@ v=X�$X$h`.�Q��'��	�O EcI��H�;��8�#��f������5R\9`!,D�hˆD��%��Т޽z&8Mqנ>D���޸K5�D��ʚ�:���Š7D��!ʖ*(�n9�v�[��I  ;D��1cKJ�n�f��6uJ�,K�9D���'ɥ|+��Cҥ-\g^���7D�ȓeC�*-�����l� k::�k��4D���pL�:~��@3���D*��k2D��Z�Q����Z��`K��/D�lC�댦p�\9qaš[���S�-D���%Ά�6e�(D*M$t,��)D�dq M�i��yY���x[V(6�&D�L�b�̟a��R��ƻg����#D��6��6v��U�P'�y�B&D�\�d�����3 �/}ڱRt�"D���H��d�ZHqF5*"�i���>D�X� B�5&��X�Q�MפQ Q*D�<�c�лx8#�ɅA挍ѥJ*D� x�/H�AP���d�\te�d�+D�@�ō�D�ep��G�� ���+D����C�����}��X�#�*D����e\�X�*��R�PT���@#'D�lzQ.�=*J��XPd֔b&�qA�/$D�`Z�́(�.,�rj�>|���Y��>D��4�=�X8�fRcG*�Be�;D�d��Z/��l/���0'�9D�H�܆�.��w,W(Q�m:�:D���eړx0��V�$]�8RB+D��@�B�5�V/�3�&�c�	)D��+@,�,�0�Q%�>C.�U���(D�:C�ʉ#���{�d�Q�t��@%D�$���I�� RjW�k�(hc�) D����)DQ?~�MU�Kg$$
��(D��@@��%�` �'��B<���+%D����,���aC�&P�u���"D�8����?�څ�a��?�ȡ@�;D�j�d�!ָ�r,A�j�N�He�4D��×�T�]BpA7 �Q6�A�.D�|��@�/��I��J�~�� -?D��22��X�Rr&$�;�d1@��=D�@�C��S/ �R��S0�BY���-D�lj��E2*�Bt&r�$�3`,D��2 �K��h�֪H�cB���)D��rd̎�Y;��U�5���3�"D�l(AU%N�1���BS����E.D���`"�5%�L�p��H~t����(D�9�M6HH�KY�R@�A�&D�� P(j�K� �<X�#���q�e��"OH��g�6���Fh?l����"Oh�ɳb�_�Ca��5-��X�1"O4�&�Y�K�Z��iG7ײ�p"Ob��D��0@=I�
L�� Bv"O����ڰ]Ml(�&���d�\Q�"O"\�*�,*
b̉�Z
��0d"O������r��\��`�	M��$
1"O6i(� ۽]W�4���&|�x=2%"O�����j�Kf���'�Lc"O�L�Fd��Hr*�"��!(�\���"O��"A"���
�J��I*[Z�K�"Ol�a�F�1��1ul�A�"O�5H7�P�|�r�{S�.08��"OVQH�^�[�>���_�LA�"O����\	d�F��B&F��Ɖ@"O�Y����8g&p P��ģf�I�F"OB��$I��4N.$ۆ�O�PAZ[�"Oظը�;&`Q���Lm��"O���aHP�N��\����0=�"O�t��)�����W�W�_�pAc1"O�q�`�:Y�f�lJ�2\9�"Oz�ӲJ]�x�F�a�k��F��	`"O*!�#�/���TJg�m�7"O��Kf� ������7-	1!�$�V� ڳ���8�ɋ�E !��ej΅����2����g*f!�B;̌0H�+�
�"�A0�c!�d��s`�����$`���V!򤆉~��YJ4CNoY���U�ʮIB!��A�ʵAS�3K
�{���~+!����jCb �c�؉�&ˇ�M���'{�6��"aӬ77�Т�����y2�@#BZfDK�n �a��jEOQ��y�(ܼ1��xb���J|v���>�y����li�7I�0n�ӯ��yB,G>g҉��!�*	�J0p��і�y��н'ôdC'� ��s��^1�yBjK#@�Q��Q q�R=y�]�y���,u������f`���L\
�y���){� �K6J��L��-�Ǥ�"�y����O� ���S�:�ϣ�y�̕8?��1�pLJ3Z�3��>�yB�L�+�\�Y=y����͓�yrlL�'z����ۢt�`ö͟4�y2�ݻWdE:�%W�n�h6l��yeϒMk�,[P�ƶLj��j�����y���'<ك'�ןKs,c �W�y"#�!28�1�
�0 ��q��#�yR䁋Gd@����<lX��VhF��y2G�iS>Y"  *;�θ(sA�y��Y�r(�Ɗ�7HDp|�I� �y��� })D��W̭G��4bL�2�y�jԋ.tT8��/?������*�y��	<W4L�ֆ�GjT1���3�y�����)r_%dq��EE��VB��^E���"�M���;�j�� k�C�!nq�I@� �F���P��6��B��/=6<�seh��n�zv�� M+�B�U�������Y_r[��F�"8�C�	�n�dЊ� ѭf@���7�7Ja>B��'w���Նӕ*::[5
ѼV�pB�	>X�=�'�16�h�eh΅|$jB�IU�
����#<����ʢ@TZB�)� 4�xf�?sx�؀Ɍ�NT�,K#"O,�i���x4<ls#��6��V"O�t�Dn) �t�[�b:vy���'"OvUx���-�,@F��<df��3�"O�F5^R2��f�X�JY��9'"O��PkS�H�Ą@�-·OL�C"O،C�ID	�&�cG�T�U�d:s"O�e�0oڟc���H�g�32�"O8H�ס^��k�$�=,���"O���� (��I���v���"O�L�ÉΕg�5x�ӭ+j��"ON4qe�%%�e��N�4�Fœ�"OT�e4��Y���(?�k�"O���R(ӹe�� s��b�(�"O�5�@H0��$�+r5 �q�"OTЁq˟�!\�i��k�2"lS�"O~�aC+D����j
59�b��"O$��mS)L�`�p��Gr���C&"OХ�GMGX<A��L��n�z�"O��[���J$���b�p��P��"OĨ�KJ"Mh)��C�>��5"O�BÂ�H9:1�ώ����"O2`藇ݭv�J�a�k3J)��y	�'	| Д�B�:�c���]��'�Z-���h���;P�K�`d�q�'��,+�<�4�H�ʓ+V����'{����Ą'$��	g��Gy�1z�'��4q!B<<� @j�`��Ca�P�
�'�P���?�$T�R�6K��`	�'aXx	V�ō^��a납0�؃	�'3�1!��8ٲ-��'7R(�	�'``��Ѯ�O3�tA6�GGE4�r�'�6ph3j׻��q5
֥;�N�'��L`�N_@� `���1B�'K�]��I�	L�Re���41��,��'�| zьŻ5
���V�[|��3
�':����mT q��*� ��?vђ	�'dj�@w�,CaZ��D;O'�e��'��TI`��	�(�P�<o��'�X����!�=¶�%7�Ek	�'��x��_11(�����+;h���'(�37�����e��J�; ���'t��X�lғll�Y8iI<�>0��'#�|b�])a��T��̓�z��'rو��6G�,��S���8���'�A���+L�\� R�4;�'� ��ξ
Cd�
#�N�AmDz�'��dr��9=ú��B��>=���j�'�H�sS��x �!� bl����'��8��̝-gԂ�&��+Vz�ɺ�'� X��� ����a?N=���'�ĭYpiF>xRz�j��[q�r���'��-aY.`AA�=T ��"�'ې���[�dP@�N X���'�h�bPǓ�UPf9�wg�* ��
�'�]�0�\�P�@t(�b09�'ՠ�y7#C�<��p�#cN�6<h(�'���p��AS
$�o�#]84���'��!�&�
o����� Y!4��'i\�H���J��y��	�x�'�p����	�`ur5�32ȶ���'g<Y�����( yK�2�FH�'�H��l�s����p�U�0��iR�'
6آE)�\5+������I��� y�%-П�V�3�ȖO��"O 	B�L	"�����#4�P$��"OBH�eaU�%a�-�殆56KR�Js"O�ThT�o7��8�{�B��"OX|�`��4��!t���O�.��B"OD�����;X�֑�E�֭\�05�"O>UB�$ZV͠'`
9��!�"O� KAg����� �i�.!��"O�y�b�/�`y��X@r���"O���@ڡ  �����(q�ڱ"O"Q+1ˎ#S$AStICU\�Ѫ�"OD�(�ˁ���0Ҧ�)?���v"O�-h�j�9f�4�SDہ*ؑ�"O�
���6"���L?}	$"O���tIZ�^�z�S������	�"OJ��礄:{m�82�]9~֪2�"O�J��P7���r������"O��b��P���P2^��!mK�B3!�d�>g�i
E)fA-�C�H
�!�Eup=`�k=C��7`��!�$�D!�P�5(7vנ��ST�!��Ŋt��x�G��`�b�h2탲1`!�$
%` �  ��   ;  6  �  �   �+  �6  �A  'K  �V  B`  �f  �l  5s  wy  �  ��  ?�  ��  Ę  �  I�  ��  α  �  S�  ��  E�  	�  L�  ��  P�  ��  ��  7�  S  � �  �  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|E{��Oh"pPC�}2$�����x-+
�'D8���$9���0�]V����	�'�6D
�/�/%�a��jA7Hb��	�'����R��/����.��@�P
��Q�ܙ􇈘�HД$K�_�D|�q`,D�ԑ�� |^eqQ��\n�#e �<a�4�OQ>�S�GEa a�v���`%�tR	'D�<�E�sY�u˥�7�z�[�#��w���	����3��A�%Ι����F�$D��x���u�,�W��p���#D�D��fG�k�l��8�FQ0T��>I����P������0�&C�,�ȓ@R1�ׯ��I�F�3��EǪ�Fzb�>�U�	�"�rA��?;��h����0L!�D��.3Py'/Þu�r���I� ��)��H�0u�ӕH�*}D�Z1t�0�i�'�ў�}���
X�z4�ʇ�RX�&�R$�O`6�<yc&+S̊��s��)���˦��U�IU�@FP6W���Ї�B"	���3g�)}��'M�D�:o:�2⋒)�ec��N@��y�	�0�`�H���YN>EKB�ԾdD���� ړPU`@��F�c��IZA �$G���O��س@��n�8=�E�$j�du�$]���<E�����K�t���rr��"�Rćȓ9|ڬ���5R^|ĸ �S���~2�'p���B%��tHD3`2U���wL�C�	*�e0f�D	c+� �e��� ���hO>)ӕC׎7�>����IOB���O'�������[W�^�_�r&f��x�80;��d�)�(O�O�I�ǣMAn\�B�ėG�A�
��� J����0lBʙ��OG%%���`����Ҭ�mn�qB(<:���f��y��Z�X��d�0�D �T��?��>H�d9F��||����]M���V�#�㨟�H�N�����U�T���K�"ORh �E.JYЃ��6S�O��=E�t�Q�����M�
ju���,N��yB��a��ӈ\������T�y�A��?�ڭj��BZ��U�ߘ�y��Ӕ0���Rd�֏􅐷J�j���O���DP�tAV$i�(�>r0P��Z�j�{�';�	�&��2�T�C�GC<BZh�5"O��E��9(��]�-�Z<Jv"O����-�*>�ڗ�N�+<0LI��IC>U:`�V�Q0�dI��j��� D��	s+�{4@D �/s�$ّ�":D�8�i�4}��Xf��C���#7D�887���mH�7᝕v���;�`�4��	lܓHl��r׮_�r��g/�b�rՇ��y̓��x�B�G�(UYfd�&w����ȓ8�va
w��I�L9F&,-B��ȓ]J���R�J���(jNS�%�^�'�̆� ���8]
c�\[d!�|�x�'� ٩����	$R�0q� m��e�b��7��{�!򄈸t�L�Kac�: ���'�P�����<���'��'�噆& 6���$�c,��	�'���[��P�5��)PF � b?A"	�'�n�����,R2X�� @�p�`����ēM#�)�'<Q��Xn;xaNBH�&j�.  	�'t��A�.�����Q���f�LM��O 6-3lO!AH�=����Z)`+�0-�І����yb�Α:|�=8P��MM
�R��&�y�/�7?���SeՒW������O�0G�$�þ3w����	
����d���y�I�7��B�/��7 dP�c���y�/70��q��FʠG�z�B�,�6�y���.���1g�V��
懿��'��ϓ^�F�{3*�.�X,2���r���'���9�1JŶՈd!4[9���7D��*�W�6���ʶR?�,��K7D�K�a�(��������XXЂ'?q�O�O�gyBg�(z��)���	��b\>�yb(�?��-�ҩ��ļ;�jč��$�O���d�/	 ���ѹ2�l�'g-kI!��T�&*�L�5l+`���G9":���'p=�����:2�3ᄭJ��`�'azR�|����0 f�^t1�U���O�'G�%?qq�qC�Q ��"\q��edӪ!x�xB�O?7�֥l6����O�<,{���3e�	H��H�(	�!ʒm�Z	�V�E�&d� 2��yb�D(�0�]����L��%���4�'��n�P��x"l� f(4⒁�	��lA��'4�$���Av�҃�ӳb��l
ŇXO����<	�5M0P���b4n����T����?٠��Q����j3xzB��dh�<i��X8(�����H0>�E��[b�����OY�D�F�޽MҮ�b��,YI|�
�'��@K$�F�A~��c�$[b��Ɋ{�k�m��uG��D��N�)C0�xQ�� ��L��*D��iugH�o]�5�q(ُF��0"J%ʓ2��x�	�3=(L�+EF�M��Z�L���O�"~�B�˔R��Y���	�@٘��Ѧ��]Ĕ�f���L:�OP����ȓC/�4*�}#�DZ�hv�T=��S�? ~�"�.M�	�H��R�6;��3�'y�'�>L���-m�*@:Rn�~|�9�'1V�����T����1�U�{�����x�B��i�>e��I,�v�j&l�!��=��{����|eb$P���V�F$�Rʘ��y���� �I��ןD|J��B�]9Ǹ'ў�������3 řl�~,��'W^�<yT�_&*�t�A����C�rM�Sj�D�'���D���kd���1ڮ�j2��$CbC��R�<<��H�4���D�#��C�	���H!���*��t��2uZC�ɳ��0͍�C�BFU�VC�I?.W�{V+��(�D@V/�}�B��1��~�	PD�"z:!��lΈY�ȓ!��Р�>}���&'�U�~��hO?YД�E�|��e���U%��H� -:D�d
�/Fy��89G���2䂸8��4D��!�cT*�� 6��6O�nh�f�4D��´��O�1�c �(�:@�D�2D���a
�nM����(c�H�)��0D���1�KtT-*Ec��1����.D��a'-�l)V�� ��8<I�e��),��'�S�'�T!�Rų\�(�a��1Z�j���j���p)_��n�)"�W),��x��9<щq��i�(X)5mM�l(���	���7���@�,RC�蠧F\?x#��ȓV�a�Ԏ�9 �����lO %��">r�:�jyr�#�رr�*�����5�⡆�b�	�R�E�1�=�ơ�>P�<�ߓ!֦)�T��˜X��c���u��ɯG	: �ɒG��8���ԟ,ȸq����(�C��=l��C�U� P!�W�Y���=�V�p���}$�3@Wf�B�*z�|�*1iYV�<�"��gg����-
wTi��aWI�<!����p_��
ՍI~�r�ه��F�<�U
��ZN�`e^��ά�u�V�<�T��^B`q;f#/]lL��N\�<a�ګrd��+�A���H���Z�<�A ��vc�N�C���0-�O�<!3��7\-��ag��q�ziX&k]L�<�5�4<��P�2Mfa�a8�!PE�<yU�̔tjYВ��) �=('�I�<���	~���a���<�|��&K�z�<���SW |<��a:xr�%	@ϕa�<1��*@ ��
�ϒ�\��Հ`�_�<��H~�M����-\H���S]�<nڄ�)a�F�V�2d!qZS�<��&����R�Z�$N��tnNP�<Y��M>#�D`��G�1����W�r�<��S9H#��;3��pw0rwn�y�<qRc�b8DQ�"e߂
#����d
|�<!�l^�Y�L(7M?.|0ȹ��t�<�@ͳk5�<��i�?eI.��Љ�t�<�͵KD��3�ȽU8�M�&n�e�<��Þ�쥨F�O���Kr ��(�C��;�vt�E�W�`B�����*��B��.1ض}��7�Z�9������B�I9sঠa$�S0ɈV�)ueB�%128��OO�+���� �(xS�C��i��My"ĂNيQ��0��C�ɟRS4��-3xe ���C�I�C�IYڔ���+R�1h���"!@�ejC�	#�����ݬg���i���)=PC�	�F�������[���BS�\���B�)� � ׀����14ꐠ� ��"OP�z�g�H�i����31�.ˤ"O�t�I�(D����肚A�e�6"O*$Jt#�?b�(@�uJT�X��aa"ON�a�cV�u'4����Ж4��8a��'>��'���'���'2�'�R�':���]����h�i�0Tb	"��'���'���'�B�'���'?��'�.x��O(@�����\�s����'f��'RR�'�2�'���'i2�'+1����7���*���*��+��'���'���'���'���'��'��R2�	�FQag0^���	�'���'���'�"�'���'���'�BpP�M��gR��E�Ժ$�*%XU�'���'}��'��'l��'�2�'����W!R�H�P�Ej��`W�'���'��'���'�r�'��'�n�(U����t��p��2{�h!�w�'T�'Hr�'�r�'�B�'���'<V9�(ɐ <����\';	���V�'�'+��'�"�'�b�'��'	2��k7�aC��SXy{�'�b�'���'�R�'���'��'�t�k���R(\��o\j+����'�R�'���'��'��'!B�'�N9���:%8��čU�����'���'��'(R�'3��'�R�'�2�z#�֭&�ٳ`!�tK.5�'���'m��'4��',�
r��D�O����ؒ$ut� ��r7TE�A^Xy"�'��)�3?��i�*]Y��Q� r���y�*�񦭒���
ͦ1��v�i>�	�)�g��=(#�<�u�⅏2�M�r���@�4���yK�U1ւ��ӱi.2�"�]�,�4��W�)�b�0�	Ty��S�S�2�0V'Ҧ�P� #/[�T��4�L�<!����'
��w��rn�n�r╃.0�Iҡ�O47�c�����s@r$y�4�yR�Ĕ3���y�H��0QJ%�"E��yr�K)tݘ@�Q%�> *ў�՟9�d+g�Xt�U��p�Y`G�`���'e�'��7��/l�1O,L�w�߂)��U�ǯ��HtQE��O��OX%�'
B�i��d�>9w�H�����Qzh�K�BX~Bʋgg�Y�N�	ҘO2�A����H��I�'cdl�S&�PTA��*X�,!x��'��	ٟ"~Γ+�.�8��s\���(Z��X�2�v�!���[�����u�i>�uF�k����P7:^0����X����!���8�r�l�[~2�0���+B�U(�����b�T�)#��+�bC􅇒d�$t��؀��x2��6JKPx�&�G�L����Q��?�2��r��C6E�Zd
�)���fSf���C!Z/l� !ށS<�<�����#��APy!���?m�И/44��O#a>����}d��B�B�(]�̑Rg>D�q�?8r�*�&�7In1C ��a\h]�`�Q�ԕ��&����7�Ɂqޭ�F�S�9ji`��	s�LXPf�}�d�82#�	�民��̏I�MQt��U��$p�/��[됤S����&�V-E�Y�F�����	Ɵ����?}�Sɟ�;BLُ<5�ʇ��'����
�#����OxA[E��O���O���1�����O|�)�G�� F��{խO�sc�� ��SƦ�aF"�4�M;���?����Z�'�?����?�$�^�M�t��B<����u�6����V_|�O_�S�ɐ&�����t°4�M��7r�E)�4�?����?��B�T曖�'F��'_���u�`�y Ή����M>J�84ޮ�M;J>)t,��<ͧ�?���?9��!��ybD!�N�J��DPX�G�iD���Yq&7-�O���O��$�d���O��$�("HP'�D��Ad�im|9�'A�y�'���O;2�'�哙7�%X����M��Y�EE88��@H4�\<�M���?I���?	�^?}�'pB��P�;�n�$P�^� 5�J> �
���O��D�ON���O�˓x8=``8������4P>�xcw�^/?���e�iw�I㟴�'v�'��g��y��C�<q����9M&<�!햍4~� 0�)���?���?�梏g��6�'
�ʓk�N��L�?0Q /4fϔ6�O����Oʓ�?��"��|:(O�`���� �p����!bg�����R�WG���O��$�O�lP��Eצ��IٟD���?Q�r(Vd��4�o*7\�芖B��M����d�O�LAV<���$�<��a	�%F�y� �td�SU�C�NdӸ�D�OuR�*_��	՟����?�럈�AgnIBp��jDP@I��G����?�W����?�.O���S5�*�O�<��E�^�"}� �1f8�8Q�4u���sv�i���'F��O6���':��'~��v� 7W@XT�f��n���Z�%mӸD��(�O��ı<ͧ��'�?)D��*w� {ql�2w�Ј�`8/����''��'%D�{g�uӴ�$�O����Ol���h(r�f(����f4a������iK�S� �g�m��?����?y��8���N
! nz�H!/Zқ�'Ȃ�X��m�P�D�O0�$�Oе�O��dC. �n�s�)��uiz���L�~����q���	ԟ��IΟ�Iv�=J�$i""�B`���3Guеi@,�M����?)��?	�T?ٖ'}ra�(|cf��v��\���c�	β ��1��'���'��'LBY>������M3c��d~Bሶkli7*A�.�iq۴�?���?	���?.OR����e��I� �d0jc ;D���0$�~.p�':�'�b�'3rOX;Hj6-�O<�d�eD�ҢY@<�h3`ԑV�ΑlZş`��ǟp�'�������'��P�?kܭ�0*
�b�ۦô""���'<B�'���A9��6M�O�D�O8��͚*�Y�f�pWB��`ۻ���o��0�'��C����|��M� �8�p�
F��+w%עg��{ѷi��'(�p#��z�*��Ob��������Oܝ!6+[��ވk4g�i߸|	e��_}��'vJ�i�U�`����O�N�%[���"��%	D�X%o�j���z�B7-�O@�$�O����P���OV��� wﲠ�P��l��5r���n��)mZ%~�VsӺ�D�OԊ 1�ܓ���	�D�r ���!P����fE!7��l��������Z���M���?Y��?��Ӻ{���I��݃"[�G弤�H�̦��I|y����yʟ��D�O2���n9��X�N�>����,�5%J�lZ���J�a���MC���?����?1�_?��"�
��(��"4Bq��H2Eb��A'�O��D�<���?�����$ԭV�8aڴ "	�E�c
^�l�>�A��f�I��|�	]�	}y��گ9dPВ򩉽 *��d�
{����y�'��'��8,��8�OO�1"L�0q�nlѴѱ(��\حO��d�OΓO��T>,��'� PR"^j �d�X +�1��O2���O>���<��c�T��O��1��9C�\������ c����?�$�<!v�Nd�F�"0�d�ΗBv�I@��ˏQ)�el��L�Iy��B:`�������b0CH0R��أ'��
�%A�IZ�	ry��	��O��>Q��1X0�At�e��.w�6�<I� όE �6e�~����2������}�Z	�#ȑ*<5&�T�l��˓ s�YDx���IU4[����[+I,fyqw*Ö�M��ӝ5��'_��'t�4J �D�O�٪A.�/�H@!��6�d�c�ͦ�`�7�S�O���A�(.�E���֯g�])g&��k��6��OV�d�O����^����	N?����@x8Ai�)�/H ����I[�?����<����?����=�O�t�h����(Drֲi[r*RO����OJ�Ok�ؤ{�,�H��f�	����I�:H�	��t�I��`�	�@�O����$��"�&}���;J��kT�M�I��O����OԓO�ʓ:�\ʰ_�OJ�L�҆I9M��b&�c̓�?����?�,O� aîW�|b���,x0�Y	bH�:
��ǂQ`}��'��|�^�l���>�Q�̝s��639r])d��X}��'�r�',�	�E�| �N|:sGF�%M�(#eD��U�l�)䞦l9���'��'���&{�b�trs'�(5bA���Q��JL��+e�h�$�O�ʓ]$��������'�t%φ~�-�6NѝTi9�(�t&O�ʓ!��Fx���<�2��g��ò�E�}L@Q���$�$�D<mK���'����)?Y�lİi�T쩓,����F��榉�'�:�Q������4�Q�A"8E���δ$i��!��-�N6��O��d�O|��I�	ҟ��!#ƫx{tq��J���D*����M�2k^p���t�DW��J-)5�C�!5��8C��3hx�1mZ��x�I���V뎌��'+"�O ڡ	��Y��C�ٻF�4�B�d�	?1O����O�D��f(~%���ྔ+�e�F�l��p!��%���?������C��G� �q� B/4f(곢	E}2�����'���'I"S��
�&djځ�/�6R��7�AZN<)��?�M>!*Oٻ���i��F�Y#hV4�1�̑X�1O��O����<q�I�GD�1YÀ	Ѣ&+���(��;44�'�R�|R��v��>9w�	#;�$y�U��s
���ݦ9���P��ʟܲ���ɦ�ڦ��m��߷UP�W�C�>�Z	���Ϧ��	b�Iqy�]���'�5ж ѐ<������Ɋ�qj�4�?�����=y��e'>��I�?����� �Pu�n�~H$�pM���ē��ٶ���'HA<%q� ��@�@!D��VdR�l�gy�f
�mG6M�I���'>�� ?��ˌ.���E�S�(����Ŧ��'at����4��'{��Z���'�Lq+d�)�R۴4��B�i���'���O�XOL���2)X��M�6BUc���|�m�_����?�g̓�?�t��u�fH��6�4����Q�F�'���'"TZ�f"��OD�d�O�ԉ2� p��"1�X�sRt�0TA�{��*��?����?)��?����8V����FI����c.Ϭ���'tY��4������_yZc�� �DÊ�V�&�S�eQ�B��
�OL�p&���O`���O��NC�=�en��qxZErR�0+�y�.�9�'T��'S�'U�I�YP�,���;0�#=P�P����\�b�,����P��}y`X6X�t�%Jnz�{�+/��D͖ ����?	���䓡�$��yB��[OzT���H�f	А�7�I�P����?i���?�/Oxp�',�Z��@�5ڵMB;2�d&�<�5۴�?iN>a,O�Q�������x ���f�
��r!��s����'�\����ѵ��'�?������S�Ȟ)�̤��/0Z����5�xR[����b �S�� g�6�I�"�����8�oM�M,OD�����������������'�9�g���j��k@����ڴ��D��{�b?�a���jA�p'k��Ɉ�1�j��4��-ئ�	�����?�K<��U�8��*����� ̏>
b<S��i��s���ڟ�x� H�'�+j���,��O�Z���i�R�'���O]DO��d�Ol�I3l�@���g]0dv�lEk��M�Rb�4�C�>�՟��	� !J�2��`1��!K(�+�.��M��0�n���x��'�"�|Zc���x!`
(D�Dm1`�"+�� K�O$Z���O��$�O4���O �$�|z��z�Be��o#��zT+'kڨ�G���O��O˓<[J\�u͐��0Ƀ�a_1�J-�˅��䓡?���?1(O��	F A��X �"��n��3C�4��cдg�fO���#�$�<�4Fy}+�5�"��	�*0Ӣ}�@������O����O��e���2��d��@��&�%.����'� s+R7m�O��OT��d�6b
��Е�5JN��S`�2Û�'�RY������ħ�?��'r
�%3e%��t���)U��G����xB�'�(�J^6/�81��ú���4��$��Z~�oڲ��	�OZ���~"��B���#�61$�I��J���M��'�8��!�87�`|�5��\�����48�)2Ҷi�"�'�B�O��O���XA����կj�)�+Q*<2&���I�,�,A�\��Xaj]<j�I+��F�M����?��s�<�(v�x�'fR�O��2��ӱZ����L`�d`��'A��'Er�-n[!*�n�z��P�?��7�OJ8᱅m������	Y�i��3D鋈��+��oC�ԛ$�=��?���?*O@��7��0i�hC�ڑP����[�N\�T%�<�Iן4%�8�O̱����6u�9�p�O VTh�����O�D�O>����A�<��$[q�E.���wfč;6t��&\�,�Iߟ\%�(DyRL�PQ�Aԯڊ/��r��L�����O��D�O0ʓy2iƕ��+�`�L���m��v���"F�`�@7��O��O���$�h��0�N�j����	@�����'�B]�0�Ӌ�ħ�?��'x���#T�+|;� ��Ε���� ՝xr�'�X�YG��Pkp@�G��8D<=��4���H�}�m�����O��	N\~�
(��D8�F�eU@� �.Y��M[��?���P$����L<)��<A�l;�*[�o���ߦ}�pn��M���?i����5�x��'�� �ɑZ�,[����sr��V�i��m���/�i>c���3G9��A�'�S&ʡ%I��tA;۴�?	���?�EmS-d�'��'8��z�;!�ӗ�H�c��A�	��b��U"�I���I����������m����J�M+��:��u�d�OX�Ok��*�ԭ��D۶����5�����	�f�`c�D�	ݟ���ny��\P�U�e��8�<���X'{��a��J>�����&������p!��߹
nx �t ��6���8�m۶q�ܙ��sy��'�b�'��	�R��� �Oy�AZ�a�e6*	Q3����C�O^�d�O��O\�D�O4I�TU��8�O�&>��;s�O�)W�� gi�>Y���?I����DX9Jh��%>��� z;
�����A�F�1��X%�M�����?��1%�����L��a��4X�x0��*sJ�7-�O����<�I��u݉O���O��s�#C� �%X��"p`b<���OF�L)`�t��Y�(�
��\'d����fɑ����nZEy��C�L}�7m�n�t�'��TH:?�&�^���j4��QB��o��!����̉e
؟$�b?�xā��Nd:ݳW�F==��)�d���$���]�	�0�I�?q�L<q�d��qF��1^���/ϥJ�r�J"�i���'�ɧ����͙^�Re��c��G��\[���,�0m��H��ߟ �f�ē�?	��~RL�-BX<����i�p�6��M�M>�wMۚ.�O�r�'Fr�P/m�p�X��T����0!�؞X�6��Oˠ 	q������IV�i���T���e� 5���d@�>ѕM_ �?�-Of�$�O��Ķ<Il��xߖ�2r唳.� �p�G�A�~uK��xr�'���|b�'��Gx��U�F:�*���CV� 	�c�'��Ο,��ޟ@�'�hQU`p>}��rLX�P/�� �R/.��OГO����O�yJ�2O�ۤ�Y/
���bΎ�*S Y���J[}��'V��'U�ɜa<�yjJ|z�˅�s�!BV��?d�$��A<F����'��'���'?��!��'8�y�5� B�Q:�sӈ�
d�*$o�����	Vy��ץWg��>�d�>5i�d܊s�BYh���U�\�@�[m��矼��"e����i�~��$[N`��WI�Ӗ�i�%��ݔ'q���l�D��O���O��>� ��׹d�B�)u��
\'@%m�ߟ���~�h�)�9�t`�f�frf�����u��6M>l,4�&ꀒ �J���);O��H�O�zd$a�$�1L$�"O�*��¥ )�T�&�ߘ8"i��L�(*,�RL�dV�=�2���+=��kc�ǯ4��+��ؖ$7R�Z�I�<N�3$�0̤-p�)3��s�d;I�Ƞ���mjr!RB��<�As��$����ǤR%)���0�.]���Zs�@'�zD;4��J�(�0B@H���2í�Od��O��������?��OO�-�F ٹu���!��N�ҁ�Z$6=T)U�~9|l���q8����� ���垸mM��<
�~d�5��T�Z��М��|��K�msL,i�3�%ob��E
�;nT@�PGINkX*PH�"�П���4P�'M��'��Ov�I�F�;�90�G��3`�1w�'��'�$,���] M3�1æG6Kg�i��yJx����<qv%OB�������M�����n�1�� G��I�-]V��	ǟ��'e�"@�1cQ]������"�M���9M�"���I�2�\<
e�N8���#�� ��r �e;t%�3�]^�Dzt�S����u�P�#$���iE�t��pf�No+��}�!��џL�'�IZ$�1t�bmS�`P�&�a�y��'�"���*Y%�@�C6�u;�'e�6���Y�j�D�[�`۫GS��<1Ea��F�'R�^>}�����4������F�8\���[l������Nh�*S�|�f��%C��-˛.��˧��h��5N4�(�*_�tM2ͤO� E��*W�~�����w5$Р6O�_�eSՉ�:��$��e|J�yWc�9[ϼ�ӂ�_��s����F��1+�4�?���DED��X��׈!�x}��X>Ә'�R�'>�	�3�L��%��˙�8�6�J��i>qˌ��Z7cW�C��+��Y6ōm�q�v%�O~�$�Od+Ҧ�^Z����O����O�u��4�,�� �9-Î@��/Os@HPgƢJgp6��Ϧuj��^@I�b>�O(�D'R)bC8	(����"ƴd@��^%wt�-5f�P�= ���eh!R!��U/��S��f�mz޽qt��22��Qd��p)�	���H#�MKV��[q�Oq���'wRMH�K�mH��
�|KB�E�j��<���O�$�	k�I�2��I!�HO����O�˓`�4�6��EA���g<g��y7�ނs��\)���?���?&����O0��Lfy�1�ף+�`�Jb� 5E�1@g^�"j�����K�����9*l(�JM�Y�t� B��L4@T��3��u�C"�}�r�J�t���Q�m@&k��D�Ywy�	�m(�(֎��]��YIZ���Ek�sB}�Qm��Ȗ'g���U�L@�H�UIm���`F�3{z!򄘞w�.��6�Dq.a9�AZ1O�z-�O�ʓxɊ8�c����d�O����`E<T����`�	%.D4���Ov����2[����O�擬d��%Y���<h������ym�l�낊.�N�rp���Y��|ڧ�'ix|:�̙5$&��0z�l��	"�ɚ��ŵw�	�1��L8���'�O���<�(�
D���H�)Ir|��<����?����)K�c�0��T`�y�<L���ٍ7!�Ĕ���K��Sv���VHDh�iE���ԕ'��Q���>Y�����&b�����^J�pb����|%ʋ��r���Oj�b3�[�H�b����,~-q��|�*���`Cݥ1i@	��B]*�ؐ��>!P�H�=�	 �!Bw,��� !�'5�v8���5<���0��T��4�OVE)��'��'>�I�ZA�tr�ō3nA�!�e���1O��/<O���D$��*381	EA�(lO�@�'>*#=�i�?`���R4g�Mly��a�#��&�'�r�'D*���'��y�B�'�B�'^W���;h��cC2{�½��$�4kuP8���jF6�4�[
=N�p�G�I�=:*̣�'�N�s�����v����ܫi :US�ΉW�4("ï���OuȑA����q��&r��(a'!9��x��L%�M�c�i9�	�+���,O��d�:y�(��K��p�䟛PZLC�=k�ށcǁ�3o<��DH?w"����ʌ���.���d�<�U�K"T���q�k
*z��ҭU�A @��@��?���?���X���O4�m>9y�φ la�)cZ�7����b���H�d fFӫ!~�{sɅ5"�X���H�UQ�� V��'�P�B�/<�U���G�i�5ʢ�[2S~%�s���������?�HO��Ф�Q�@FX�	�h�6|������H�$��uӬo�埬�'����q��djU�)�4� s������X�ҵ�C6���q��1>+�@�<������?	-O�2�Zn�t�'��!�A]���@q'�LW�V��s�'���q���'G�)��$��1o@t�x��'/��8�k�z� ��I�JڨJ�lO�cl�?b���a�-`����ʖ��y�1 \�N�8����)OL ��']87�m}B�33����g�f��U��B����'���'�DRĪ��/^p���D��l�	�';�7�ǔN`��D�9��}��@R�*x�$�<����DA��O�\>Y��̟tAU�w�,��iA�i��ԟ���#�lq7�}�`���O$�.��ʧ'�Dd��PY	T�8t�"٥O�-#�.�$`�ła�Б}48��1&���ra��S�	o5��!:)�1���?s�l�9WM�+7��Ɏ~��$�ЦE
��i��"��Â�3�H����*y��s�34�Ȃ �� TV	s�k�H��d�)Oj�Gz2�&tU�p��J�u�����"iF6��Ov��O q��0t����O*��O戬;� �!!h�CR���`��^0� cD�%�<�0D�p�*��2m=1��'��]Y'���i��J��m]r�'��V:I����R؀��&#�k�\�p�)��)D�T2�T���� k#��|������ձm�Hpj�Y�m�,O�a�T���O��O���ei>csn(����$�61
�"Olq3%]B�FE���)T��I�.?����(�M����D�h���RǍ�Te�I�KG�e!�֍�z�j߹xI쐫�)�=YI!�?	6tH�$���hqo.i>!򄗅0=�e�� �5B�>�y'N�1'�!�D�-0Ƅॆ�m�tѼ!��.<��9��o�	.�DYW��(�!��o�yX��=����d�!�G�D��#f�<�~0C�X1c�!�ē&EFdkЧ��F���o��6�!��ڄtC|Ur`��yD� ���fi!��D�%y^���'sJ}Ђn�#=?!�Ć�m���j��V�!�D��ph�a1!�X��¢�˒m(��1.6!��zj	��W�M'̭2�Mƨ&�!�d=N�t�{T�ۻ]����ҋ]�J�!�Dڣ�2�Bb�Е.�Z��KO4S�!��V@����c��y�J 'WJ!�$��7N\*'�T�$A��b��;&!�U�⢽:����r���U!�ϕ,�r4���T�x��e,�!�dЁl��!��d�9�#*u!�D�	^Ny��Z&=�,8i�"�7f!�$:Ҡ%�$hց ��E�fH�!�ެ*�,�0�ȁ�	�}0Q��]�!��Cg:e��!J�(�r���A�	"�!�d�G��a�gI�q�`�RoV)�!�$&� ��kOg�6�E�^�!��A@i8�_�$�PV^5!���D��u��,"�"&~��Jv"O���l�~���	i^�Ka�$�B"O�H*��F&��0��Mx_�TB"O������o��E�5���^��<��'�z�����=�F$	=���观#�Xu ��p=��@сCFʩO�M�Ӎ�$Ψ�y��	��*ذ�I%B��U�r�		�Q>��.��R"N����V�`a��&�	�m�ac���.<`Q?�+c�K2�4r�"ؖc�6A�e��rv��#��Xw���A?!��PW�b��4D�b�b#��?HK6�z%þ<��O~��eG�7�� Ȉ�d�/l����3	��bc�J�z�����Op1b"�u,�\&��'������ S��s����l]d8�r)pE�,2�G�z�'N�tR�I��l��.}XR!
��H�Rx@Գt&�,n��!Ӄ-�<)�L-k'���$��L<	��og�H
�*FXߦd�p�ǡt~��>�u ��aþ��&!T�X�`|�����<4�éIR�E؁D�/!S�����"Q�<�-Q�=D�6�[�S���r=�%A�}��Y�ۿRB]���U�RJ)��)�5o����$-�5�^4�%��X�Ïl��\���-���;D�D��B"^���y�A4�<����H�,^�hU�u�X�H?Zi�?1���8�
<;�P4*\��@�oR3H��EP�G�"=�ā�-9��Lh\w�Q?I�F���z��		��Z	Va96Ɛ$.d�9�c⋰P��Gy�'I�V`;2�`��12��VJ�ܘ4�2AȼKF��c��cٴ;�0C�'�S����ϸ�*��� |�Ը0�K8]�B��
[�9)Ф�Ʈ���HQ��D��u�'��,i�M�Oĝ�!+�$"d��i��RV@��L̹_2�O�)�b���k���@��AG�/�4�dN�`���TM��+�t�6@ÁfT�r���U��M_�OC�<��B� ���|r�í� �c��������q~�@E'/�p4xS'�-#� u�1h�OT]1v゛EF����@�k���0K�5#���X�e�Yu�t�����3���0���Z�#1uZŰ�"B7@_�e�R�W�I,K�"u�Fz������[�N}s'˄�@(Q�*_�_�~�	���F�"u��g�I�>��"@�.B
@��Lk 둮Dv�'�Ҕ�B�V)����~V�I���ó-�/ �
	�5ʞ�{i~��.��)�B������OV�k�iw���)LY�6���X�a,�"�J8xwh|1'	�R��d"ɒ�l����s��73`X"��Ҭ	�$�R��}2!�'.��yܘ� 5$K�J��t���J�|��I����va˵ y�0�0�_ Q���+ٴ$��#�dZ=��yJ���{0��#�`R�6yK���O����ʧ$�v`r�ԙZR��ab�H"%Y*U�gH��!m�x�'�%P��B��yF��'�PAvY-d�����̡�?y�$G��ӌM1H�,��'�6�!�9� * I��8G� �M�;�����	�?rTB��%0� *� ��'J,��A2�A�eq����./��������4�';�e���K�c�lI�Dp��+N?��H1X�҄� �2�}�R�M>+���!']y��#�Fȷn%��i>����5���q #�V�R���bY!'�]qe3Or!iQ$�:��@u�럴�s$�I�&D�	2g�k3�h)�OW_�UkFl��\�%\�p�'�(]�~�ҩF�=� �҃@MX�&�Ǎ��mj��� B}�ԣ>�gB�?\�ͻz�&�׋ظ)Ø!jb�3-j��	Ay���!hO�)�ɠ����d9ֺ�8��.����򦎺TAL�Gx�"��=�t[u �_�5�]=�~�'	�E��&n4%�as�T�'��	.X��Dr�K�;	`Y���`8aj �
�o� sH�<1�p�-g��UA@��C����h�8-8ԗ�c�!����'#�66�s�� �)[j�Q��L�2$Ad;O
ј��֮P���ɰ$S����Iv�'=~�0��´V������C�\���K���(3�.Mi!�x�\���GO�'%K\�[raŪ=g.��VH�s�`P��E�e�V���� ͓�9��a���H4C��q3��V�	r!�E�'��	��&-��ħ�?A��\l�r�"f^�Z�@��Q<��u�>ғwN�7'Q��``��>u����ݓ���+�.e"�_ U���TY�Е'U���i�
��F�B|�R�'
����xWbmh�%M�3M�?'�L��s-Ʀ&��P��L�#Q��q�¤�ֽ<�.O���r�ȫ}��8` ��	E�p pN�L?��#94N)����3�da;C��^�'!.0�B�[�/n�͘��
7��A�#jt��dy�X�|G��% v4�Q��4�A�snX�J��eO�=E���G~���3C�T̻!i�=�4�Ē����0�E��!�O���?�*O1��$ưtl�YhEH�8R�d�
܄&�N��H#c;h�Ԃ��1$��f�I͌��'�M����H!3ïM�pp���X�(�'��.K�4)"���v���b��n�j�)S�%�a�D��$�]鶇Z�F2�YF�	tЩKV���.����I&T�0h���/f�V��0♗ 6�">�|Y�oӨ'��B�� L��Ey�h�$��唤%tRP�b�(D
�<B�'���f�'v��{�*���lh���J>!VZp`�!�P�'�,�aK�����N� �����mK�$YJ�A��Qp؟8��LY�U@�F�倉��N�pN�؉�D׮l_*!I'
K�2@DKa�D�B'�ɓD�Ă��>o	(���c�4vR�>I �Xh}0��	�vpKg/��$��ϔ;Z�	tU7_�Vd���pӀ��v�P�yn���CɪLT4H ���\c�@�r�>|d ;ӫ�2Jq������$ɹ��P��M]�q� �=����`�̉����Ҁ(��c��Y*�2�'�0y!���	8����@��=�Dhz��72,��7�'<����e���Ql��f4�pp�7gs�ш��?�O"��#�W���1eg�w�8�(�,_)9��Ȉ��W��򙰏���;23��hs�Y' f(��.Z`��O �����N5��W}NMRd%�krfYJ&�i��(�GӉ	
��seE�IĜ�Ϙ'�N%ZB��Pf�-Ĳ%ke��*+P���r+n�"�%I+�TX���auў�r�m	*V��ዖ�z�6Aa���
W[���h�8Y>h�PG�Ԋ@y]�mEEI���B�$�V-Փ���&��x ѳ�Z��#^��� ��l����.��O�8��]�'ݜ�a�jԋY1�DɣoA�N����Ν&C\�Ez�݌Xʢ�ӳ(S�X���^�a.�	�a���h��4 �	�q.̊S�Q��2'�F��@��0]g­:��OhI��{���S�F֒r*�PP�� �����'	U�d,;$��.E�h6ݟ�O`�bM�8q.�8�Ek\�����tƣ>qe�YcR�
Q�Άs�P���E�X�'�����%	@@��aXa�����D.�?����(��Q���5%;�zT�ñlA������(o\QQ�k���O8���Y^�\�(������:K�
m��D�@�'~
l��4�`d"D;��[%&ߎ�* "�_"Q�AŎ=�O�ٳ��ח
̾AQHT*?D�f���g.�x���������ϡ���<�-O���A��>��a��|���ċ�	w�~�[TJ�8x�ȴ�h��)8�rS◚%䈁3�\�) 8���O�Y�,�'bm��k�7}D(�֘}�
�;,O�[�h��L(��8[t���	=@�]�F���T��bd��:0��'����F�<������E�;f{�}P�B�e^���[{�ĸa�/�A�,�X��dՆ_��)�w��#��X�Kzv��S*G�
kf���?��o����
WY���'�J�I�/�!�bݰ�A��[�+�xe����HOfA끇�.X�!��%��<��O��aʠ��OZq���T�va�-O2�v��L�|���+ϐ9�2+F^�H	e�Ⱦ"��z��Ŷ�M��ț5i!��SL��P��R�?˓�?)5#V'ɪ��DJ�!��6�� PQr�y���O� [*X�!�^-ǽ�uקI�'x�uA#F �l��e��M�4���/I��@��8���OЉ����O�NE�f��7o|ٸ`ɳV���e�D-f�}q��'O����U�y7ًM	�F	�y�
��LD	�?���a�	8��d�<���`��22ɫQ�N`4f2r�<�I7�;;��8��DR�Z�@�0�`�<$d�x��f���3� V	Y�lB�E�a��B���aW���'����%�*-�� �o�`��/{+��S��%|�$,��
mV޼#���r�8]��C�oxЩ�b��B�z�#ϟ�	����>�¥��AZ;7�1a�l��M�E�Ozٻ���$Cm��`x݅I+�T�'*� Q��S=j��!ṆI�\��J2e�8�ӷ�����O�����OJ���.If��bE
S"�Ԅ� /n�UcBGN	��O0�B�(������N��7kR?��� ��""��'3&��'��Ipy��.�y���NA^�*1'�&]�lAc�'U�k=� ��	�W�|��Qj^:�؀_� W�"�(��Ff�;ӌ�7f�37l�XJ�"[�<qǾ��d�
�2�M1�F̸���&R\Ñ�I�}�Ĕڂ��8?T�c&��\��%�B\�m�ڍa�K�[쓶?Q�Ovr�)sGۄ5�ZTb�'�#AN�P�'��M��FO�
L�q  �	PB�� W�(O�T��*
�$z�������"u��Z��O<��%���|b�'���MK�U�
�������5��pҠF�P�P������o����T�w��T��c����ǖ�2��p�A�'�|BS>��_�ڴΓ{��[孒fp�3&˿@��!@��c�'�x�c��KmL� o\�?h��O��j�@��d����pg�^o<`���'�bS��� )S�<��+��$�6ݛf��;O"$�R�#��c%O�G�0�3i�H���dF�&��ExP� ��f�A���d��.�8�S��L�JnD� ��F��F����'��5��N�. �j%�tg��nE8�Q��$P#%Ѣ��`��.a��/�"�۰.@eQ�O֢=��MJ�
0ʨ	gg�~��� �D1�N���<�ua�-�˟��y'&M&� w.�?Y�
I��ı�M���3�S�O���]<77�] �.1�8 �C�d6c��(	�q���s���,��Q�� �d�
EE���L>7$�4��Ü�3����$B����;R�A�eFչ:kT)(�KS�w�@�/,6��c闡f5��ÆCC�7t@�-06��gᇁ&�����t�#lP�bq>-��hB�
�jHP�]�9��	5��U:SK�
&h*�S� ^�x�⟌�af�{k����� �K�Tp��ܘ��'"���O����󉍿*~YIA,Y�e��Y�'��N�����臵TD�Xҧ!��?�[�/л/����f� P@���!1�_���jUg�i?���~��ÏAM��JT�V�_Zq�Q�	�4�Op�i%%q�4�#A��v}k��x2�����M���T�u��w��I�<�\��'_̥��������־�I�G� v��!7�Z�V�*B�)G�e�^yIX?2èk᥂Dr�ZB具��O��O���U�<W�Z@{���7g\t¦GZY=��	�'8�yw�U,������Z#<�ĩ@DX�WΥ ���CԦ�L>1"��56$@f_�]��¦��� "��c��50`*"?2eH&'P�7l8$�����T���6?r���	I�	�<�WE)?wT &�ج.F� ��F�'���T����F�dgL9��L�#P��1 VG����'4�0"ROѮA�ƕE�$EM6��ǢA�9�i5��%|R��e��1��O?�%���St��-o;*�+E��?baASV��Y��"�Q>�:aܑ�r�E�y��(rT�@;]����r�����̒I8|j�V:Df�ه�ONh���ו��#��9uNX�ȓG.��#��G����v�|�@؆���=0#�ʷ?q�๶l	�&nF���hX����G��<ٴ U�G`p����乐c�W>b��c��i�fe��tƨ0U�6kGȐ׏�)zBD��e�0��㎎�q*8m`��#(����]+���7	F�'
 ��ԉjY�H�ȓ�b���7y8���T�y��&�nh)e���j����5O�����oD 옦"ֈj����K	/ 
=��	��z�V�"*��k�)zޤ�ȓ�����[�,��F��j	���ȓ^8�C�NW�V)г��}5��ȓ&�<д��DT&�A3L�Qzd��l�z`iw��u�<ՋG��#��q��Z�����SH��k����=���%+Pݒ�l��W R�k�&^ 46}�ȓz��P&��+O9p��QUfDp�ȓ7�XM��FƜy�Vp�V�ڸy����ȓ��r�Xl�,�fǜ�a������Ԓqa�/
2y�I��b���_��<i��^Ѹ�挥AV���;pZ�Q� \2Z�N@c�B�� ��S�? \��DZ �P�rGLmi�r%"O4�+T�O=_e"��G�
�6`(��"O������?����i]�]�ƀ�R"O���ðjE�Ԡ�.[yN樠�"O2��#�Q%�pu��C�R]R`8�"O�ԐVj �A�̫����	]�U"O,�����f�FQC!���v9uCW"O\ cbң@C�ab2`I�o��8�e"OZ���.���T��) @V�0c"O"�Y�;Z���EH/6@z	�'���)�~5�����Å|k�<+�'��%T�ۑXJ�Q�
�z��p�'������,]@� ^&tO";�'@@,�f	��ib��W�␺	�'�����X'$(L��NJ�����'9���ƭ��PȂ������'���b��G p �1�1?��$	�'�
�Z@�<Q�����m����'���)`-��O�����i���
�'RV��w%Y�!_f�c��F6b:f��'��$�5�I�M�BT�q�ʱ^�4�Z�'�������u2�	sa�܀h}��b	�'�rcآQ��hqM,_M��P
�'մ�A�"�i��}*��>a����	�'�H����۽)˖Ļ#옠V責��'br]v�
�X�$I �V+�M"�'46�ʱ��&8���O_�\�Z���'�N��g�4K��xh����`(�'�����_0x BE��_�H��'D���'��o�D��D,�!XY�!��'�`�&o	�k�L��ÃN�Y;�'�"!ȧM�7i��$��&'I�  ��'��H��Ȗo�D@a4㙚1����'n$˦�U$^������� 4�h�'�Ř�G	wv��l��1�:U��'kH��/Д�H�2�A4"�����'�e��
�=rH��gͣC��q�'>��=�>H �+ �3��q!�0D��b�	L��$Au%މv�D`d�;D��	�Q�tX�@A�װb2aؕ*8D���!֜r�x���)W!|V��!	8D�L�� N	&mn\�`�S	cV�R�
9D��E�^|��\��H�H>ěb$D�| W�L�� �� r5PP��.D�<�Ek����`�AY*<&$�D�"D�Љ���D;QBb����}0��?D���r��4V<i�/Et��"�I?D�d8SmN�c��x0C�͂/ẕ��<T��q&�L�C�ʩSE;]t�}�"O�mh��R;M5��2��7&�bK�"O. �ukɺ�h0��k_�T��"O|Q�'N�2�|��!�*xȦ�"O��S�,J��X*s���I&"O�٦O�>,�3Kŏ�A"OXY�4hR?nsB����ٱ�S"O@�3�	�g�2��#�ֵb�D�81"O�[�C�#&�x:1*Ӷ5��IC�"O<���@O3(��HUH�kd.<��"O�`(C�δoN�Q`�� OR���OFݣ2�Y�s�)�!�0'zp0r# D� 9���I*� �ό}>J��G�>D�hy�i
 =Q>m+&㈹_,p��� D����.�["��*Co
�y�(X!%*�1�S�'C[��GS�"Ja�d�CU�`t��S�? P����ɝ3���0$�X���9T"OreA�A[�$41 ˏ�#��d@�"O�
�\6'�<��$�Fy��uR'"O|`��H*m�����`H�"O��k�M�~ǞE��l�\��%k�"O�eQ'O�|�b&�~�X��"O*�۵ ��M�p���7t`�dR��G{��i�03���0�.�9�0����<%!�$��N@
w���T�ʅ�S�� !�d��+Z����1+ذ�	u��!�DѤNyP٢����h[�����0J%!�_w��Y��<+S I(�j!�D)SX2աӍ�f�(�A'�ʪD�!��ُ}�$(u֛y�*�S��N�>�!�D��go��:3�Z�B�p@٢d�i�!�;]�Bi�4-Ɂ0o�����шd)!�d<	)�,a���X 庀ƛ=/���T��
���<@tL:*�\h��`$D���4#�$Y�h�Ǥ��3�FDB�E!D�,�w�6	I�Ȋ��-NLzg  D�0!7�,8�*��E��r�����>D��� �G�'��㥩[F��*+/D����䏽H ���@^EpȒs'"D�T��D�W�:�@��{�4��M2D�TyJȀX��ը_?�R��.D��u/PEbִ���/1�D	���,D������Ox�q�&ޑ��b�/6D�����A,�]ґn]�.��`Q�'D�|i�/�,�r����2	���֡&D�$3����a��t�1h��PF
�u�#D�Ȣu�+[s~���K�Q(@F� D�p�So���L�Ӑ*:P�S7�?D��Õ �s�ZB��=ja�?lO��xy6bŅ7Q�l[� W����;D���X�b��-���g:D�t�4�P��!��'�
Ɋ��:D�tJ$�H�R F�E�Tml��%D�̻`��I��(�! �;b`T�7D�ī��4%�Ȝ9���;L��A`�6D����:t�����8?��,�g4D���fG�wo2-�	�#����`�>D�:�'�1�
ur��ߓ:�d���<����S r4<��oG��A�A��mg�C�	�o�$��O�u���@5iB䉡7*��vH���T���{� B�	���帐�ˌu�.A��*O�K2�C䉑F�h�sPfW�A�j2����Z�C�I�\@��S�X{6�Sc�S�MONB�I,=>d:�Eɣs�ܩ�WA�b(6B�	g8�ђjX�-o��F��13�C䉯O� �]�DԱ֌UR�#<A�3/B	%�]"�£<Z��ȓ	��݊f�G�>z!����n�ȓ[^z����+0ʨ��@;�Ȱ�����E��1|R�`ѢO�<RC��+x�Yf��N�FSR�ZK�<A�MZf�0xe��pnТ���J�<����B�4�;���epP��l�<���e�
���H�nA����d�<Q'�M!����i��a��I`�<����/K��|�R�I�4�����c�<��o�^/N!cq,�,B	պeB�_�'�ў�{'��kt�P�R}v#���+L�X���g�������b�3? R׏	�lXQ'(D�� 8�+h�z$ɣ	��e�u��"O��A��y�,l2U��9 ��8��"O″�
��8�>!�6g�=�\�`"O"���l���Z���� %�$"ODt��:&���G��R�捙�"O�t�f�)=��q��'���!�"O�`"����H؜ӐeM�+��-�"OLѡG/�;���棅�X�ƍr�"O���Θ�L�R5�0BS�]���2"O0���U�H'Ԉr�N|�10"O�aK�A��&3كs�W�\�Z��"O�T:d�2�MߗK��i0�"O6�����W5��ؓk_�r���D"O*課��p�T8�F*9V��"O\�B��׶�{�)}�Z����Z8��j"��1ID�S���nF�`ʗ9D�h�&�P�6����].��p�e6D�Dr��#|�d�G�۵6瘝�Ua)D��H�m��{���b�c[N��R�+D�8�!mژy�!Jt��;*����-D�d���,R!h万��G����,D��8G���3hz�5AY�QܲI��)D���Qɛ<2��%���%
������(D��O��=6t�PN$k"��؁:D���" 	'5ʉ�A�̎q6�Y���9D������A_f��W��7ea*�(�!D�8a�Q�yNΘ��I�-i�(��"D��NJDm�w�ډ�#W$?D��bթ,��̂cm�82��'D��aA�
%ILh��1yqjdׄ2D��X�/`���E�-M����o�C����0Wm��PDx�*b�ǫ`��B�ɨb1P�Z�&�$�v�``�Et�B�	?q�{�M�l�B��0:�B�'M�<yc��j�x'(9b��C�i���M�G��|JS��
�L@�ȓW;���3�.5.����ȓu� ة�|y����
�r ��,B��S-� ��b-�'=�T���x��m�:@1t��v�2��>A����4!Y~Q�FI�y� �'��2�y�J%7�����B��+����y���Pkh���*\�xa��y�c��b��I�	{�̨�߳�yҁ?O�ȑ�-I.|Zĝ�bm ��yIC�}("��Eo�-n�@,rq��;�y��{(ι! ���e`&8{cH��y�������GQ�a}z��"���y2Y�c��I�GĚ�|���?�y��ާDDA֫��O̘�s����yªX�FJ|h��< �
\(@�'���Ƣ���`��"��e��
�'�� �3Mɵ^�*�k�
��m�tU��'���U�X�V�~��0e°2���'t�<8PBQ�7Oh|���V�(�:�#
�'�8��a�N:}봙ɀLJQY|	�'l����ONV��@
�N�*T`�'��)�D*J�c���nD"(��� "Om�0+�E��p���J�4a�"O����^�<礥� K��HGh��P"O�i��Kݞ0�A�̺Z4���"O��('��`톼��أh�p�s"Oxp;��6&��-���,�h�v"O$��AZ�e]�A��/��*��0j�"O� ��+T,�;D��E��0��<�w"O����ɤ.���R͟@hN�P�"O��`#@�qŖ@�򂈝Ve�0"O���P�lg(܊g�%/>���"Oj��� P%Q��%Reه%�Bs"O��炀�?�h���;��U"O,!"�̇d��d���=OFXa��"OBH�Eo��Q)�`򔬆�[6L�F"OZ��JX"W��h�l��g��h�"O��*�H�!���KR- |���"O��a�/Y;TI `�5l޼�`"O�eHPŇ�$I��H߳X���"O��"hI�b�,���=O����"O"K0&�,kzh�&�#�i�""Oȁ�c�UsBB�UA!J��"Ol5���^�t�� ر݈G�uj�"O��hf"����p�^�Rw�KB"O���1�Q�,��U���G�vp� [u"O��&�#Pt��q�_<mRjIy�"O0,렉K�L)���gȗX4�H�"O��G�O�j���-�7X`�u"O�����[����4�9.(�"O.@BD> +J1;��l���"O���!7]S�-:��4"���"O�E�a�^>MDӰ�P��X\C�"O��z���%K|��c�/. ����"O�8ѵgǽc�
��W�*:Dd�h&"O>ܙ֩�<pZa)!��K1ta"O̭��'�QxZ�BP�M;;��k�"O�i�EM�������]R,Q�0"O� %��#&TD��J�2|GvY��"OX��O�|u�ph%�Z
~EH��"O� r�A�v�EK�g:��`"O�iYT	.K.�y2�K�d�R "O��r�XXjz���j��E�:���"O�i�7�,�m���T%$�h�I�"O��!K�2G�Z��Q$#�Ɯ�'"O���ݛ~�J$+PC�����@2"O� x�C�x	bᘲ0XY��"Ob����|�x���E{R8�"O�Su�ѱ*���&�T�7Ԓ��C"OV��`"�:8�}p�πt���ӧ"OFxH����p�Q�ˡF���5"O@�1MK> ����p؟$6B���"OZ���	���#���68�H��"O:�C4�М	�A�8��2�"OQ��ĲzJD����D2�A"O�8��k��2��iC�&���#"Ol�[Q��t�DAX�(�[�ιke"O��CL�p�(Úx{ ���"O2hP�'��ck�M��I�,�"���"O�1�oW�+�� 5<Uw�D�s"O�������飗���V���C�"O��Xr��.�ܳ$��)�p�"O�����
y�,9s�L��|�2	�'� lP���G|��z�CϿ!�N��	�')��ȱӞ?"�1�ψ b����'�$��Ё`�j�S!O��K6�{�'��a$EAͻ�bD-{.���'p�(R�fF�cu.|� �7yΦ9
�'px�K��c%z\kS,��i��8a�'2�̂q�Gd���J8���'cbP`%ΏN��Ёe�O6K��8�'N6���+ߨU�h�����WF����� �03s圇C&�8RዯbRq8�"O�A�p�ۼB�C�/϶4q���"O<�!��n�z���+�XhP��"O�UCP�9%G� R�K�UGT�"�"O
Iw���DQ��Ɏ0OEX��"O<t��ÍM����VYOr���"O�-��
Ѫ"����qI�_�Q@"O`
a�ӡ-t|�;6��:�Ç"O��2���k��XKħΫ:Q��*p"O:@2d+S(M�9�dũVO�aY�"O����D1�����?�h� 0"O���o [�dɲ,6{h�
�"OĬX$ݿ<�
��EL*w*,+g"O��R*.9T9[�*ߘ/[Tͺf"O$(b�J�~|J��ygx�bS"O�a���9yp)2�I��yS��e"O�9�
CV1�� 筄:gM�$��"Oj5��(`M�$��![��A�"OPH耄�;}� �����D��1"O�)[�ˠkn�e�� R��4��"O��;��_�o�H|��W�l�t��"O��RuE
�e��pK�to��J�"ON�{����~�4"&o��%�F|:�"Ovx�b���F��1.X����"Obp9Ӌ��kf|�b�5_�H�"O4��ggb�`Yzt�?=���ұ"Ojt*�.	�Sa���ό���z�"O>��'hЀ�4yVfE�<���cR"O�uj��J�NpC1�Z;��E;�"O$�S��$O�@jī�⨰�"O� ���H���� +�3|�84"O(��"Cْ&�6�k7#�)M(J�"Oz]�d�*B'v%!��0{!�dY-��Cbl�>G��8ʓ7T��A�u���
�k>d�2�A)+D��fOɬnM�EÑ�Z�r�� �$D��rN�9&-�I���&�Q�V�"D�����##P�	ȗ�Xf0���&D�$�A!�ƺD�t"�K�Τ��2D��S�	��%E~��o��v��w	/D�ȸ۱�^�����?k^����h.D��zV�uVQ�D�
����.D�L#�	`�Jm�G��u�؁��g>D���A$�%FuX�*ؘ��(�B>D��� $3(�,��[$
�|�8��6D�D+�)ǌ��}�eģp%Vc��1D���vɝ)���A��O@mp�o1D��)#�r������{�k��/D��[�1���r�lW	�θj�e.D��8�d�v��s�o�0op-��!D���.6�NX6��#��U"�� D�A/͂;�$�83/G�EJq$�1D����U_�����#-z╂�*D�0H�V��W�W�,z���h*D��[s�طedF�I��U) l\��E*D��4�/`,�� A��tVd�"I,D�X�Bk��^k��bQ�ua,hc$!*D�Й1$�Ī�u�I8E�j�JE�I��y�OG�|�v�Ħh��E�%c�8�y��D(@4�B�1]��0p�/H�y"��-�^��f�B!YR�v)���y��K�ApV �lߊQ6��Ư��y�$C	:u����� �D�)W��y�n�@	�EXUkՁKkޜ�F��y
� ���D�P�FcX��<@�x��"O�`�2��2;�|m1$��o��:�"O���I�4>�V�Pv�@�J�� h�"O
�q�/�xDSW���`�`P��"O�t�u��)��4�W�!�}&"O&i�,�*4��7�uc�yq"O�`���� `���F��B�x`Q�"O����Q�9��e�S����"O~5�%Uk6 �ru�B�"��la�"ODY�U#�<���7�D�K�(��"O �j�l#.�
ř/#�BH�"OQ��_�r�R���Ĝ�6	x�yw"O>��FX�lhs�F�*���R""OXyj[#l��4U�/�܈y%"O��$GϿ'r�����gU���T"O|��$+�,ٺ�,
:B�#"O8�ta΅Al�0�Ùe��J�"Ov�' 
t�չ�
ĕ�Pu.�!�$ơj@��G�>� ��_�!�$�"ruN�2a��Qva�0��H�!�ĝ.n���qB���b�+@
t�!�D�3��[uč�X�GL�Xl!�d�y�;n�uƦ�{� �(�!�$�}W�<X �,Q�����E>Q�!���^8��@�<V���o�S�!��ů`����fظy��ia�	,�!�d׍'�|<��L`W���A��Th!�Ē�Pu��R'�OR0�����\H!�,Y8��¢��|X�S���!��8r�M:"],#��q��R$9�!�ā#zB�be/".�XjaE�{!�#E�jٲ���9���i�ܪAd!��Mt��Ĥ,��xY�*A�~E!�0]JX�����fn�KV��#+!�]�$� ��)�?ZDZ�i�`!�d�k��`��
N6��k2!�dȺY����@H�@7&�k�K�6!�̙fx��t�y!�4��Dd�!�د}{���a£A4�@v���!�հ9��5"Ӣ\�^�����L9�!��Mʰ:0 ��9�b�p�
ǵ#!�dj�� ��#�11�r��Bp"O���G�1T��zt+D�m6��J�"Oj�q`�Z(0<�����l��!"O��
eJ�>A� jA�
�]�"O�8㱥K�w7�58&IW}�y;�"O��ICl'8�(��"0�\��"OZ��+	�"�F8�����ˢ"O��2V@� ����?/�섡S"O~���X4=� B���q�X}��"OP��		�q�.M���	�FD"Oމ��ȗ=2diA�"M��"O�<�!��f�-�#���.¼T�E"O��6�V$ ]�t�!�p�d�r�"OB�����&@�j$��n�h�A�"O�0�B�/�Ĩ����W�Ÿ�"O~�U�V�y?\a��&�K�Ԥ7"OBiH���?z�\L���w��P"Oh�KҀ\��	�fk�4h���v"OLM*GdA?j֥Q��%Kd��
c"OҬC�kX*�,`#o�5�J!"O'з}3�mb�X�@��zf"Oh<���#�P%��Έ%�Lh�"O�p���5�l$�a�еN�d�Ò"O� �P�ԉ��C�:�b4�\�#��q�w"O��b֫�3��Ą�6�\�0�"O� a�Ş}�j�A�b +nHШ�"O&]�R�~& ��v��~@�Ȼ"O��C�"�#�0�9g/Ӧ52L��v"O��b�)7�D�z���uv�q�"O�$�A�{n2�rSc��fpx19�"O>0���WB�.Era�AUE��%"OJ����Q��K��4d3�Q�"OH���G�1
��8�͗�+u<��"O�-��!�[?L�p*W/"dBI�"O��"d�N�n~��ѬZGt*""O�TȐa��1]�H#�i�� A�D��"OPT��J/rJ�����	�F���+�"O��X6�"�I��Hխ%h\KG"O4��ԥ�wi����� �kr"O��S��J���3�$���M��"ORѣ�e��������ڷE��Msw"Oµ+c�E�W���p�_9�$��"O��W�>EY4��^��$�r�"O�I�CLCg�����ٗ霼"O�)���R�H�Փ�[�S�z��f"Op�;& �"SW�Y���E�~�n(Y�"O����Q7���!��̱I����4"O�-���<&� Y���$X�t�g"Ot@�r-�/��)ttH�"O*��� Q�B�p��4Of2Q:r"O*�Jc��n�z���C�:G}�ˢ"O���3OL��Y�"V�Cd�P"O��)��>�����o(cT$��"Oj���xŴ�j��!;�� "O�A��K]�Rq~xwP�p9�U+!"O~�x�lϏ1�������$"OVI���ã>�~=���`���ȕ"OH�X��>���4&�1��mA�"Oh�����CQ�0�TC��8�Sr"Oʩ;&�N�P:b<p�P�+�("O��z`-
�7������ܟuM`�y"O��N��qXFtHC��vl�%�"O8�[�Α=UJc��$\.P��"OBHaEW[��+��٫SP}x�"OX�rrG���(��׶p!`Љ�"O�2Pg=+@D+�o\+Q�6e��"OJ��rm�k�h��PN��y�01�"O����'^�)�$�R-V����"ON@���1�p5���k@�"O��&$,��IS
��/*��(�"O�-b�Y(i*��gI�zd�*q"O�ax���26�j�0�&	�T����W"O���SG��"g$��'g�1&DT}+�"O��r�+�"͆����k/h�;@"OvЄ]�=Ѵh�r#
7{*����"O�T�q�V�0��ϕ�{���0"O�`�5j�?��8�PA�Sz$qE"O�tRQ&˦Vm�� 	#M��  �"O�������b"+/�xH[W"O�p�tA5&��Hɦ�\(3"O������>��5�%HӕM׸`�$"O��G�81f�EA 	O�@�@�[�"O2�k��-.i��G9����"O�E�%N �����ѮN,��I�"OL]���_��J��%7���#�"Ohiqׁ�
 �P�9QKR�Z���"O�jw�� x����J��P"O� �(S��yx-2q	��.e�"O�ds�G
>�D]�i��6h2�(�"O��C�G�OS�;g��
=ZA�r"O�4��d��7��M3F��Ոd"O��`�C
�M\$�P�1@c��"c"OPl�4VYY8hj��Dp�2m��"O��HR6N:6���@#UZjtk"O`G
V�(����DJ��+Sȴ��"O�1p�ɕ?qi6��7���r6��3�"O�2S� D���! G�.@1&"OL<����>0��arga��a>P �"O���)�t�:������Y"Vh��"O��F���k)N��OF�)���"O&�YF�]=T�`|���7��M�q"O�x���B���wa�;S�zt�""O��á��6as�h�o��Ĵ �"O���Ȣa�1b��.|�Ւ�"O��� ��W.�'��Cfޑ0"OuKu	v)� �V&L�?F���"O%B�
�&b�%+a�g�X�:"O�<k"����jm(��0Q(� B�"O�{Dbx��cb�8"> �"O�("Jǳ9y *�k�d8��"O�=��EA�Њ��+��0m�"O�#�ԑ>�:�;�J�fɄ��"O��c�Ι?
��1�dۡ2����F"OB���HB�tCR5z$��'U7
�@�"O���EH*<� ��$��BJ=��"O�1��A�!Z�ZѨU"
>3P�#�"O�X!�f����pB�/ډ9Cّ "OH��2��K��1s�`�\7�-;s"O����ኗr?lС��N�1SU�"O�ثr�P�̅���̹fEA�7"Ov�sf��0���b��<:��"O�)bp�Z�Eۀ�C@#��"O<��AƠf}����\$�J�C�"O�uq�̗�(ߖ}�T��'��x�"O�L�c�6z2x@ږ�K�t�Bh*A"Ov�ۣ �?,0 �ӗK	y"��X"O��q���+V��"��ŵE�]�"O:(��&M�+�(������쪵"ONyz�儸B���Į͢��Q�"Ol��EĹC���`�mJ�m�d�!&"O� sp)ҭ1kh��a��,F���" "Oޤ���%��2&i�9�9q�"O�T����C�q	K�:8
"O��	����6��fg�*B��au"OZ���c8t&]��ܒ+!�(�"O���H&M�M����"O�-�i�
0	d�HGl"&�f���"OJ���`U�)��1˖�Óa�X$��"O�i��I�. 
Y���3KڑPu"O�)��!7x\x#��a2�-+%"Ov8�5��4w�b	@aKO��A�"O�k��
Q@���
�?v	�L"Oz�#���b(���S)� 8���"O�5�����vD�a�ɉOd��"O�ᘆJݶ�R �5.�70� ��"O.|H3&C�N���[�4�$ z "O�L��Y']���LG0@y"`��"O<X'*�}��%�3B�	i�03�"OF�QCB<�Fy31'I�[o4��"O�Mqm�<���G�Z�w"O�rW�ܧN���B#ƕ�:W ��"O� �%����pp��!6D��Km�XA�"O�љ2�U \��,t�ʔ	��E��"ONа4��(�0��W�߃zԞ�2�"O�����6�#�D�,�!"OX �E�OzB@VNֽ�Z���"O�T�aQ��U1�C "\����"OƙSP%D����(aM�S"n,Y�"ON0�Ţ�f���p�Js����y�r��+7톑��5j�σ��y2kT�[Xm)4%��z����n���y��=,��}rF�-%��8�/��y���#���)�.�
p�0IC`��ybj�:Rz,!�!޹b<r����7�y�A3M(� XG"�7)�|i`�ˍ��y"�%o��k��Pe�mCԩҝ�y�Ɨ�8�\X��<1���CŅ��yH� T���f��z���)݄�y2�L�0P�EĊ	$�8@����$�yr-��@?"!��!��`� 
��yB�A�!��ZPۚ�Xё �	��y"	�`��8	�� �p��hk�"�y"��&n�����i�`�I��y����i�8D8fZ�Ā��/��y�.4���PЫ�?#���gW'�y�nK��ց�ϑ"9$����y��ěq���0`��#�+�#Y�x�ȓh�{�g�v(wf��M�ȓKA���M�4���Ͱ{5�܅�/wP����f��"�c�����Y=r��䁀,\��@�v�Ï[^~х�'x�c�7b0Z��sc\�m�0���!N�!ch�wB���
h�݅ȓ]�T@��D�
Ht$�ɍ����ȓ\BVL��hݘl�b�I�,
�\O���[�����H5/���)�*�mJ��ȓ#aHR�N=I�HI�fn��y"��ȓ7<���D�w�M��R�'�<L��]�ȼ��%o�xL���@�j+v��ȓU�Q����8�zy"�=,u�T�ȓYNv��cB�0 �,�BM��5�A��EE4��#��8`��Y���
� %��[���L�<��d@)�0�~��ȓ0R�C���Jta���>&4ȇȓd��	Xs#JlU����$^�.܇ȓ3����FC]7\��S��@��ȓX!6�Z`ƽAC�Cӆڂ-�61�ȓjZ81�����2�O;@�����<|�� ��vVh���:G[�ɇ�t�$-���.]��U�7\:[���cp6��8=������[��Y��ߢ�p��Z�tT���"��=�ȓL
���!x
u��i�6Nߺ���G~~��t�;����h���e=L`��Ǉ��-\��d�4I���V�9+N�[O��S`� ֜��q	�Mi�Х0�ak&AM�A����ȓg?4�R��%U��r$��1U��ȓv�Q/H8a�kCc7�,�����b��D��x	��:L�ّ�'Q���J�g0���=d�Pq�'$�H�%.`}�d� ��e��M�'�b�����m�0"\3i�dt��'����p)�TRиjS$�&_��ݫ�'��}cEjL%@k��jBV�"�x�s��� l,�� ��r��`�����-bl"Ovt
U�ّ?lh�2�˗7n��U"OJ��+زh �h%�
Y_�A��"Od�y�m\({T�	�R=^�� "O�Rwm�I��Aa�%��=�`H "O��Ґₖ'dir6&3O( �d"O�Z����O�&ۇ�׷1/\sq"OZ�"�)b�dr���d���"O�m�tbԯCZ010[�G	���"O� IQ�UW`��J-a��"OL	
����,�S!)R�>k(�B�"O�9���W, "�g�
b��"O�U� �6�>��f�$\���W"O� ��=*�&�حiU�Bp"O��Q6핻V�E���0S���"O8qۗ얗cn|t!��R@@\��"O怛���=Ynd�4Ƙ3]UT���"Op-8B�E�-�e	��Թy\4$��"OduY����hZ�T��)B��p"OQ5���X	�c��oE���"O���h �<����&Ì�B�`�"O�HE��0b�i�s�M5T99"Ox5���{�-���7/*z`�4"O��
"I+V�m�0A��mx@��0"O�E�+�<)H"��[w��B"OJ(` �^�P�A"�8{�!B"O����O�����r`S�O�L���"O���wf�R.�%� �B,�`�Q"O><7���y
m4Q� /[2j�C�	�J��ף6F6�jr����C�	�V:D���R�@�gm�USC�I6�p�"�N^#� ���(K���C��1��ȳ�	�P��M���G*�B�2ZX*b�Ж9�(ᚁ�D�F6�B�I�]�ȩ@�#-="�c�j�!ONB�I�&cD�A-�&_�饪��
B�	�cU�+O��%��' �3JB��J���� '	�[�X�sR�{�NB��.h��붂M�`��0�g'*B�	�2j�Y�uk� 7�^QЄJJ B�$}f�-"f.�?�pE�0.$�C�	��1��/ֶch�p���ŵW��C�	7nUl(�תC)�İB��P�C��6H$:���S���Ff�*
��C�	�.����sfl9BA�z.�C䉁pJ�2 ES�$�f�(D�ϿH`�C�I,�.��r�˾v_>��f��0j�<C�	?\N�pC�덧*rH�d���C�ɀU�Г ����B89�/��k�B�	�L�洪q��:{��p��BN�8~�C��?��������MUƘ����z`"O�q���K�� X��D h��j�"OxD�Wё0���#ƦVV�X"O����&
�V���irI�t=��b�"Or=
�^�H�N9��F��^(��"OЁ����lV�ݢ��؍�x��"O�,���A���Z�@ܺ�X��#"O�E��"���\�"E/	�#�����"OD�ҕ��D-�E�2)��ˣ"O���d�]="x2��Q|F�� "OQ�Y)c��  b�v6�S��^�<�NT�-��C�eϬWV��� o�<F��V}�tP�&��m��4
n�<q�hƻJ�6DP���C���y� g�<� \� D5!�L��FL�Ϛ���"O(��_	\�x=iEB�k���J "O�Ô��'�zы���P��*�"O���%��'@�F���ba1|�"O�4ɥ)H*�tH�O�X��1�f"Od�'�УO�Fh�p�_E��qk!"Oje�s)ă< $�[��������"O�@0D��31��(��	�37❒T"On��F
�>C�)qwK� Pl��"O8e���m	ڰ'G�#uH�w"O�A���I�v�X�`��,rhPS�"O0��g#��^�R���)_�-�"Olu� �\�\'~50�͐�He���u"OjUҷFW%t�h�k�oΖpd�p��"O6�&�@e�J@��o�Z�\(�5"O"x�� 
�6*����K��[��,�S"O�A��ۡ3��8y1�D�<�����"Ob��k�2Yn�9"�M3uN�@��"OF�#�c�7��e��ť%��ZA"O����S�5�,qk���1\�th�"O^�qD� V(��3ۿ9B4=)r"O�m�r�C!��H���S�i!�5"O:u
�ΐ5���FS�?��"Or���5��;!�!j�Ѵ"O:s���Xaxh��!� P�|�C4"Oj�9A�Wu�	#3��+�0��"O������x�r�W-\2(�(m�`"O��9�d�Z�����B5`f(���"O��	�L�t�t�lPc��k3"O�  ɉ>����׋�%6�@ �r"O�Tಆ���H����Z��"O���U
�������n�<rC"O��ԭ����I�H�+w�V�f"O����Ђ$rXi���1�X��r"O�᫷��6���Bp�Ǒu�Xrc"O^�����s�ؒ�C�t��"O�m��� q@}K"
�!jl��v"O<�3H��;e$bE@��>��!�2"O��S�_�/���w��vܢ�["O$�k��]�^�4͊�#�.!Ҷ)�"O�HZqIU$o�|��dK�4�^���"O���T�A`J]
6��)�����"O�=8���hh!遂	����"O>1�D�^V�� ȝl>Jq"OL�*"-ͯ`G�T[#�ьY�B=Y�"OT�����D)r	¤&�8}�"O���IKaV�e�_;iδd�"On�h��,��)C(C2��P[�"O�Ĺ�;d�l,����8����e"OL��/7�����VJx�y�$"ON Z��"m�dd
��7Cr%��"O�|K�@LU���K!�*Gb&i��"O��Z'�(VYB���<�2���"O~ �'��b"��� �μ��"OB4��aP�e��M�I
N�R=�"O�=Pg��nf*!�����` �"O��`�+z�)���P�p��m�"O�(�a ƛIA�4s�*CO�Π[�"O��Ƃ�J�X�'4o	\И2"O�Xp�N�.����Q�͋i��"O�ͺ��Ŕ^t`G#A�2+�qp'"O��	f��|�d!Pńō1����6"O�*)P�+l�]�J�%�2!�6"O���cMJ�8P�	��\��%��"O� ���a�;0-�����%B�2%� "OT�AVNM&9KZ	�/D<O�t���"Oΰ��FA!u
` ��� �4��"O�	����@��,�����0�V �"OHQz��Lhhұ��/a�Z�R�"O΅Y�H!
Z(�#�b�H���	�'��5��@�HR*�k�!�x�D��',r�j&Y
j�v�#@�7l9����'5��[�O5`�D�G+�ex� j�'2����C�O`��b'B�c7��!�'���2ׇH�G�b��V@��V����' �X���94��[A�еI��(��'�2�S�@CF������n
�J�'�0���¾S`�K!��dD�\B�'�$�k'ЊBl$�'R#`3��P�'l�J�h�
=��9��g��)�$PX�'2�!XB	:ƎPA�	(5��C�'��U���:R�Н� k��0�@��''�5�tLۼ^������*�j��'�Z�7��{c9�0 qLK�'T�xK�!ʦ�t�h0 �9�ب��'�����_)�l�I�C�"RR�x��'����6
Հ`N������5NN��b�'�H\�P��>�b@��EД3���'��yaІȀ)��x�S.��,2"p��'�"���nߌc���S!�4�v=H	�'���B��% ���M̖/u��#	�'�����B�~�"I��8�ء	�'�53 	]�:�Õ�_�@r�]��'m0��RO1� :%�>�F���'������l�<��"U�Z2��'IčAsg��^xn��3��'�(h�'@��؆��"+n\���ڛ.�m��'��y�E
����ICE�@x(��'�
xڧ�ȩ_ ��Ə�H8��'� E(e��[~z�i"�Й|.�Z�'�p'\�>rL\��ӧ{�Is�'�ī�H�!lX�Nݱ]�b� �'��T�f�\�E���у��:[�����'���R��Êr)\82D�=L$���'c�}r�
�-r`����S�2P��'�Ũw�F�>�"�0��ف%�h�'��
F�� �A�3)�la�'rh�GAPd�`Vl�+l2��'A�lPp��.
����P�Ǟu��i	�'Pp:�ʤ[�f�S�~
����'�6ȁ��ŸS��*ө 4{A��c�'s�hygСQ�>L�%�T�g7|�'ݖ��@W?gh��)��؆d\�H0�'������vq5*�NO/M]�1��'�"���2���x*�Hj�i��'զ���KLu11P�̆CP8X�'7�)�C`FB�6D"��ȋk����'�)� �8@��G�]a��?���["=r�U�
j$ri��kQX�C�Sn��zf��� �ȓp��}�ևL�k�$�zE-VH�~�ȓ����M��R��c`ή'[
,�ȓ 6!롬�yc�PI�M(M<Z)��f��H��� h��� ��;��E�ȓC�= ��OY�����ڳ9�rT�ȓ_Q�c�	0Mo���éj�(u���9)Bn�4D�0���$P����p�l��@eH��y"k3F���S�? vqʄ����:�B =���[""O�@[�O5�~��ց��)�$q�r"O�S�����@� �"�0m�"O�}�EV�S<��1�\�z���"O�A�]�l(��LZ�o��4��"O�TYU��F�fU�0!�;V��A@�"Oΰ�GܽDK�h��@݀y�N�K�"O��,��@�~Q �	>O�0�)A"O,�AC��M�����>Zĥ�"O�Cu�I�\#֋=;>$�x�"O�������\����e��Jd�"O,�1�*�hKfğ>�<i�C"O$��p��c�Li6��;QylЂ"O��aq��C��ea��/pd��r"OJ��a�R0��	�&����@"O�!`����	���*A~T�"O��BK1/�����"�9"�x��"Or��f�S؂1�7�OB�~5"O$|H��>/�}Yw�ȶ\8R�"O.�{�]�$�0{2�ɖ/�6�µ"OH��v��%@�&�a��o�J���"Ol ����/�e����p����"O^[hݕr�<��X��D��"O�%����T�ب7S�z����"O��ui�_����"0�ZeHA"O�<�w샎D����ǡ��V$�u٠"O&A�ULQ&CO���SN4��e"O܅#�,�)��=��4�B�QF"OB1�͞�'?b,��KL=7��˒"O)�d�FZ&D�җ�"�>��"Oօ���C23���GR�Ӧ	)e"O��ö�[6tj��G��S��tC�"Or�3!�-V̜r��ȩdr.��Q"O�1JW��b▨�!d(Yɀaҕ"O�e�!�ӊw�\�'�E��\p�`"O`� g|�n;6�(c� �90"OR�9c�Q�4����j_@�@�k�"O���%)�*�.��t��P�Y�0"Or�� הv�ت��V�q���0"O��ԦX�jd�xU/ɗZ�P�R"O~�jԠt��,�3.ƍP��"O�q� �x�����_x�x"OH�a�ʄ���P�-*$i2�"O
Eց��y-�Z@}��"O��a��G���lĊ[�HqP"OnhHENR�JLEˆK N2ae"O��(L��bw��+c:���"O
�{���Cd��
�j�Ea�"O��S�C���Aç>E�5ʗ"O���2$_.d :�9|��h�"O�y�!ٿc�TI1�^� �̙Y�"Ox!  .ʸ�"� ���t��%A�"OF���g�#B8�s� 0w�d$�g"OF�t)݌�t0X�"��t�^h��"OX�y����/�j`�
ȵ1��䲕"Ob�:`�[5mM��(\{XD�ѣ"OhD�5�Q�Oe8��'ƞ�y��"O,�(Vl�3}�4I0'�мF��qi#"Oj��`�h�������_��ە"O�U"���	1�^EҐ.ѵT�j]�e"OT���F0Hp�Ui����"t �Z&"O��Ƞ����a�����b�K3D� *͜`x:��E܁Z �Q#�>D���b`��:��8/��%G�=D�� ����~\����\C�("O�9��ԲM=��sl��H�@!�U"O�iر
گ7������ q۬<ba"O|���X}H��Hȕ.��`:�"OK�jK��{�!4<�J	À�V0�yb�E, "����	�.��4k'�y�nC�Rf���/W*\�@ ��M��y���(H�,�Bt��V��X���?�yb 	 6|<��A�4`vX�����yB	T+B��%k���T���gі�yB��	VeD�aR���O~V<3���y򭁍p::�h1o1K�B}[e�3�y�"��N�
��t�7=�(E�%+Q
�y2L/�]�`��4;��m2���y"�<� #�ř3z�A�Bފ�y��7t���Tkѿ==�X�Ql��y"F�Ob�8�.�2H��!JP*͝�y"�̡W��J���9\@���	�y�B��=R��*p)3"Ƒ��y�iə�Q	ڇ e �RF���y��<9��A� �5e���ab��ydL��BdؠD�)h�9:bM@!�y2�Ĕ`���t��2��4�!m��ybOָAl�h��OA./s|K����yr��#�hx����(1�(2��[��y�e[�kxl1�C��v��=:S��y�J��?���򍙯i�켒E�F��y�^1�4 ��g�Tme-Ζ�y�g�(&iR��#c��e�j�#'Ț��y�o� 
�%33'a%��A�O�y2*�*H�8Q�t�Рc�DCgۄ�y����4���L�Zr|)j�h��y�-Xh���hB�IS�̈c@��y�&вzG��#���m�����gP��y[3�����*;d�<���U�yRnS;{0j!IՎ� 9&�LH�e\�yb
�2g?$|�M�8��=¡]��yb���+��� `J6�\� I���y��O�s�d��!�D�x��E`��"�y�+ג�������\!��)����yO��ZT�B�L.f}y	8�yRN�e�ܹ6荺HY5r�F$�yb$�0��Q��<̎\��Z��y��xCމI�ܝ R���S���y��5��\��	 Gq|	���"�y�O�)�҈�3�����Y�2��y2F�yv��p�Λ~0�s��P��y�V.Y�h��s���~��ؑ��1�y����<w�i#��C6vWm��cݜ�y�D��iI�izNg��=0@#ˏ�yE�H��8@CmQ��J}S2�� �y���5�ʌ����?�Ԍ��gF>�yң��b; �
'���ĭ(�+@-�y��dy���P�S������ݽ�yR�ڱ	�!�AF>z�zt:���	�y"��1c�/k�v�r��^��y�)�V�x�8 !� cZ�X���;�yn�����Z��@�g�y��޲�Zթ��[5|����"��yR�ˮO�\�P�B�����yRJ]�l��1Q #� ~�H����,�y�?x ¸X�BєU���JO��y��A?U,%#&��Jf�]����%�yB��7�4-
��M&0�E���y
� �����b��xX2GC8.� �&"O�a��D�]V�j5�ƝLN�91�"O�hr��Z,0�[�C�4' X�"O����EITK�IԠ��s1��� "Of`�P�F�+�*PYwBW=P��%2�"O��yg��?���cF��!䔅A"O�%b�A�j��Y��`��0���{*O� 8��[�RSJ� $�Z:��8�'% ���RJ�(�B��;H��5��'�ȅ�͋%�&]�2D��A��s�'u�%څM�-Yp���U�@��$��'�&T�r�_��R��`��&�L�S�'o:I �C-Z�9`Ƃ�#����'r�yz��K�<d�f*̵�BT"�'HR=b5a�;�|�v��"���'M���7i�� S��2� �'C5*�R�@�����а[�'�p��JE�3:�"B�ν�'.$��D'3�U��-y_6Ms�'T�ћ�j��7j4\{A��u��	�'�:�U/�3+�D��h�g���2�'� d�QJܧ]�l0�t��]��P�'m�=#a�5H���Y�N�B���'ILY��33���Sǝ3v�T`j�'��ySb�K�t]d�"�Ո"�q:�'�����e��Jb~�xA�N9f$�0�'��u����p��B�\���r�'o$m��� rܠ��_�kǔ��',qK���9(�1�E�4�T��'��h���~�n�[�Ʀ ��tS�'�<�w�\;s�ժ1āk�u��'���#�ңf���ڀ��j��M�
�'���Vė�J���/������.D�,�M�K�R�(`b�,m0~���o'D�,"#Α0��<�@$0�V��g�/D�h��'��W��uQe�[\.4[�k/D�0�0�4+�1��ـx�^,�p�,D��!7"����(�4e�2B�<�� +D��kU->�D�C�Э|���-+D�H�q�
M��ᒀ��%&���x7%D�X���t�R�"�o� 0�)�5D�<�G��}��t��*>\!�5�3D���L�hh7 �;@O4A�H<D��BwO9�"�V�B,H�a1*OȺ1�ܑ��s ��CMnI�g"O�r�A1j�ؽp��6EI��"O*@q"��
�<�"�-@M!Q"OdZ��P!)�r��J��Ma(-8r"Ocʄ�m�x r�,K�#\tP!�"O����OP'\��m���Ӕph�Ș�"O�P�΅�+������B� (�"O�,#�H
#���q7I1F@(g"O�M���$!� �xV̀I֪3Q"O)�áR�X9����!. HB�"O��2�!�_b�����>/>I+�"O`()�J� /�5�ՉA�3@�:�"O������4�p����D��"O�;����c��I	f.I�>�@u�`"O�*�g��}P����J�9���)�"O�)��)�\����4չw��ARv"O|��t�7P[T���a��}[ya"Od �#c�O�rL $F��0�9"O��o8���ia�T�^� m	u"OD)s�㑣k��T�aĐ>���`�"O� ���H��m0������E��PZF"O(l��ν��ɀ���"��e��"Oh�zD*�0v�AP �]nY���U"OVL��AD����P'��/n*��f"O| �a�Q�#�v�C1��3�Q�"OQ�b�$h�&�4v6Ry�G���yraB"<�C3��>m|pu#Fj��y�$��F�
i�P�T�x�,�buF��y���L1����D�q�UA�BQ�y����%&s�ƅ�8�¥��Ę�y*ɱ#�\Ń�욙4G@Y��a���y�V�Lw����'̼�*� ��y�J�29$�uh� ґ�vL�5M\��y�۷]Pf� �k�*2��烘��y���7l��E3�����^7���yB�46~�Q�k�?p�K��-�y�ሪv#N}P%˵uB�a�5��y2䕶p���zg+C�j>a�fL\��y«Q(��R�$ô����`�<I��E�>�����R- �L���\�<I��<G:T9!�&N���P�D�<YcN޲-
��W�B�� 'b�z�<�#]:	������G`s�<�¥Z���e �ߏ
I|�f�I�<��ߣF�m+�LA�@�$4���^�<�g�S,Z*��EVc��M�Z�<A�%ڗ�.Y;���k�P�C�*�X�<a�E�-3���o�cK�q�	�{�<�r��.�u�`�[�
�!B��M�<	`���d��L���C��(�#��d�<q��U��\d�J/�P
�]^�<ѷ+��%w*���L��_�:`zbN�X�<Q��]�T��蒲�U�ZH�#"	T�<)V*X$�
�����E#��EG�<�R�Se���u��;B��ݒf��J�<��/_(T��҂,O:������]k�<9�,�m���aٲuD�GFZN�<QӆտCҘ|�0/��@N��z	ER�<��GF��R� Q�Q63�r(���E�<��Ј|�PD��H�k���YP�I�<�q�y����֯Y�k��Á�@F�<9�S�A��	i"�ŷ$���3��JH�<q5���Z�RT�QH˗,�P��)G�<Q�<�xp���ɪ1�Z���c_w�<)gaїv*���,��k�"a�V}�<IM̳E|���Ç�&j<�u�Q�|�<�"M��WG,��0(C�r����A�]�<����Hi����=������W�<��*H��`v��)Q�� BpB�U�<!U#֌Ciny�V"_�ҊL{4f�\�<�JD-Q�x���y3���N�W�<�GI�<��I��������pbX^�<9�� �P��a�'X^$̲��W�<���&Z,���˦f/�5�U�<�#%���κLN��AT�@N�<!���,r���;$o��UC�U0�BT�<Q�ꟊP�M1�n��KW�`��]R�<�
���:%a^/\�h=p@K\R�<�b�K.d�аsb"Ҩy�$P��c�L�<���JNq8���b��-� �b���n�<�R��9�X� B�Џp����QUS�<��%\��)@�2_��K��J�<1���"����A�ñ1W�xS��H����U��U�r``�(����NJ3h�����S�? ��CM�
O,�P톢T�&�6"O>���hE�d�pe�h�z��1O*��ѡo����C�R�{@���2pQ�D���,���Bv�|�!�����B�"2w`E� 
�?W���2��
0=�B�ɹ3��KR�	Jj�ȃ��@-��o�����ٹ��JW[��.Վl��`c@"O�,ڷHʾ,�~� �&óT X�"O`�-Y�|80� �AgE�C4"O~p�Rkaj�(�A/}A����'�Q��yu>E)$�����*32t xrl,D�x02%K:N���G�ĎJ��p �%D�(KäY�sT��39XJ椻�l#D��R�Ƥ~�jd��
�j����Ƭ4D�8���C�uT�*�!�&xC:e��/D��Z#�������oqW 8�O*O.�`2�#9Lb�ƓE�n��U�'HQ�8�w�I
�*��qg(E�x�+2D�{�#ʹ�J�8Ceϡ3oD��s�/D����JG���cj/;b��1� �=�S�'U���K�ǆ�v�
�0{�L��ȓ������O)S�,�(4�Ċ�謇ē�n��K���Ժ�@ܕ,�I�"Ob�riב2��`�#�&4+m���i���P�$?�x��f����Bh���4D�l�u���c��Ds�[{m>��e6⓳��w��ju\�y�Mè5��-���@k��y��i�>Q��&d��AaQ��5R
��U�c�<�mO�g�nlBq��Z75ۀK�<�E�9�̱�
t��d��!�}�<�f�  � nZ�
����D
B�<�G�\�:��WLF�h]�̉D�<���Z�v�H��jؕRG�p���@�<��f�-sbx ���9|Fru`��{�<ɠG�=u��X�L%���a�I�t��p=!bh>D�F�Ô�4_8��t�@K�<)�dI5(X��B�G�G������o�<�q*3}�h�G� =��8�Dm�<a�aT�l�8г�M�8D�l0�$��f�<���-us�=��o�1$���j��Kb��D?�{��4��7#x4�;B��&^�|��զ���p?Q�O���%N3A�+E7L�	)�"O��jfM)C��	*'u:
���6�S��Gx�"��ӡp8M�$aZ�;��B�	�6gXYbǄ ���q�J�f�G{��9O�q"����q��z�+�<�
�"O&��sEH%}�<�p$�S
n)Bt�'$����IF��Ha$��7b�n�:A�*�ZB䉱_g�Y�D�'퀥�'>C��	7�ȍ1Ю�m/�H[�
�T� C�ɾr���ʜ33t��1 '�;b��B�I7A��iB�ן	6�-�4�O0���Ms�'�'��<!Ձ,X�h,�w��3?3�)@mJH<�+��"���"�&�J���+LzD��F�<q�"bZ��bE(J�" ���c�a��H�'qO���u "�s�V=)� 08�"O,���b�z�="m�'N��U9�"O2���T�.���:��0����Q"O~\���Sh>$a�	����;0"O&��uN�6�6�ɚ%��sp"O�D��˦ygv@���ZRɜ�� "O�u��o�O�.K�[�]�����'q�1�=AɎ>p3��BU,�8&�B5h�ۦI$������Q����~9^��teO�7�C�)� BU�� B/N� �A�=fiH�"O|�^�ڭ:�S�U�bL#��OI�'���Oz�t�D'@>iAƘ-�xq�'Fv�!���;Fr�<�!#� Vp��P��-�d�h?�O��јO$�@y��A� M�U$
J�����	{�����$w��)i���> M����Cg��Fx�����z�x������͐B!*D��s�H ����C�]˺1�)D�0b�iٯ4d�Q��&ڜ)�b��oyR�)�'.l�y��$zZ����Єȓe��m�Aa��s��M��V�1Ӯ�$��F{���bǺ{e
�� @E�6�ּ��ډ��=q-O4�I�`����8G*�@�B�"	k�C�I� ��RR��!S	>�r�L�p	�C�ɝ}�f��q��)b���@�֪P�hB�I�{d���Kפl���9C@A>�.B�	�T�Nij5?�ΰ�
�$�">�L>)K~JF��W��ٗ �
t뀮d�'�ax��
��;%�%(���Rf��y�D5�b�z���X�$-"�?Y�'��؈��ʰ��
�H�A�J�:	ߓm��'�:|�eE���؄�A=���B�'�$�1Q��r�Aa��7&��A�'���:�S�gybi��<'�1#�ΧR|�z�I��y��P�^�QZ�*؋,8p�� ��yb�ێ5K,t�%�7���'��x�r�|,H�Ĝ?f�Z�;r/��EB!�"ONdyP�
R��]��[�U���|��U������0�BK��J1]��ɗn31X
�'�Y��g8��H�Bd�� 
�'3X%&�J2%݀q����5���(
�'��	�,�3ZXB�j���<��U�J>	���)�5.�>QĀJ/(ցj�'�Q F{J?��=�UF�	=vI�큾w�����^U�<I"�	'jjl  (�d��j���N(<��4G^��hS�Q
��"en�!	(̄�X��4ʕ�7?}Hp��z�(��ȓQ�\<��%��h�5�V�/r(��ȓ�M��IӤ@��vJ	D$��i�'Sp`KU���>Q�zc

�3 �Ś�'�R�`5�-F�������	��җb9D���k�a�<�qQm
�Fy��E�7D�,���A���h�F�@�8�I�4D�КP�܍=��a�D��?A~�ap��3D���3a:h` 	Zե�=F��u��+&��hO��d�H��0+�L-5� ��f�r6=�S��M�F�יK�44��' �p@b�Mu�'ў�f?���􀊽4���шՈw���F-��R6<v���@l�����M��d�/>°cr�^tp$�3�b�<�%O�g�hx�M���!⡒^�<	0º ���!��-�	�sf@[�<� �V[�S̚�5�ĘF!GW�<i�)ݦ2!�x3���O<蔠��]~��)�'V}L(�`��H�: �v�	m��!̓�hO?j��ߴKC�H�D�'?�"��
?D��j���U*�z��b��!���0D�l�$��A�t����CU�z�r��2D��@qU.�8 �IB3rt�	�+D�X�U��ά%���޵)Ӥ]`��(D��s����y�b0�>)���!Vc%D��[�p�V�rV�T�Ry�4�Xr�<ᒯP�{�@��S�G�lK�L�n�<AկI^�|�ʑoV�`�!��ER�<� �5CF����� DgҾVR��q"O��S�oSܚ؂C�� Lp$��"OR��w
Št�&���&'�:E"O���&D\�R��q��;t��"O�qC$l�$h���AN�+��1"Ot���䝃�p5I,Бz��pk�"O�lS��hd1SR�
Zڤ��2"O���T'�|l ��!���)��"O�)�6=���ҡR(D��"O����G�Ov��v0*!��"O6�ʇ��H���r5��*1�	@p"O
A�č� Q����C�.9��@"O
y�pmW�}�E�6�F�uHQY�"O4�����5@��Ƭ߮:|Ő�"O��*d�دY���&�J�*h�A"OB� �gQ�A:�-�� Ad�$�"Oؼq��*A�0�������"O�;��БI�Z5��J4wh�
%"O6���Ǯ&�bH�#+��oL�q"O"��T�߷<wF�����&k!��W"O��Z��ґ�i�b-���"O�xj�F]F$T$���M�N:��!�"OTS��U�>��|a2��`�N�"O�q��jI�D�urm�~-��$"O�0���>#�p"��N;�fi�"O�9���N�y<����L���"Ox�:t 4������31 �9s�"O��Bf�&��J�\���K�"O��U(J�mXa ү�3ʔW"O
���I8  �4����z.D9�"O�XA�!�Y����í�^!��	"OD�9$F2p�>��$
T+Z��( "O�ر���	q&�ږ��M�r y�"O���E�f1~8�����Ұ"O��1 ��b� �Acяo��#�"Or�s�BV?:(,4�s?���;%"O�8���S{�	��B�D>F	�"O����q��2w/�&�Y0"O�P��بLV(	"��ȕ@ �4�	�'Π� �ֽw*�%@v
��zE���	�'U�ac�A�,U�`��}O�E�'����V!շP� �AE�.���'�+3�Ӏr����5��l����'�$�WGˏn.����`�l��'S��`eo��h�αhu�\�uz�5b�'#R��2��#t��A����<O�<q"/J�2��E._C��V/L�<��.B
Q�d�!nQ�3�����L�<A'�iU�����N,	q\\���DO�<Q!`��#����(�"��  &�n�<�
�h^��#���>B�Q�t��M�<�RMȚ<�PXk ��� ���BWF�<�F&H:
@-[�"�>4^X�JcL�C�<A�H�n��H��;�F�C �x�<�B#:^�VDK���MQ�����y�<a3�
p�C�B���Yès�<����s�,h�&ԕBfd0XR�<1��!�|�H��Z{���;�K�a�<���@�>���ހ!�D��'�X�<��m�]��*��INT�C I�a�<aZ�u����`.P	C� I��DCW�<����?c(�r� �=G��,Q�<i�@3k�8ecR���74�̀H�<��,6k�	�PԈy˵n�G�<� ����J�4(� �D�W��Ű�
O��{L�`�����9\p����,�`��'��P��=,ΐ�
7���������z��4[Fk\�ħU��=�q�݅������|A��e��-�7o�k�^�D�;>�\-�':�T3��^������j1�䵒∜'N�RI�P(�S$���"O5G
4&����ߟ$�ԑU�p���<E��<�pF-��3�I��$-;tӨzX�試f�5Y\��$�U;l�d��(���a���,9Ҽ`p����MU�������^����w�'�L���ͥ<g�">�+Ѱ�ܑ�@�� ����,���2a��$�~���'�h�j�d"O)�#�I�Z��h!������@C�=O����7SB����������Q�m@�LH'�/��|��MPp�<���\�(5��Y��C�\I�
7b��
�ٛ��T�4(�5Ā/v.���O��{�'˿t<���*K� s�Ic��'����:���@&B�C�.Ũ4��$M|=�E�	l,� 4�'Ĵ���Mҡ&��-y%��Ba�����X�6צab$�2 �t��eh�|B��4s�����M=ͪAC���B�<��˨ys lS%�ѺYJ��t���<��B7Q���D�E����)��'ix���aΪV�D��1�&�!�$	�
^z�󃮉�;����6�������O������h���1�?#<��ҝ5��&�� z����i����"�V?L���I-%:��l^#e�4���I��h�H�J��'��ia� �4;N q��Q��9���d��T���c�=)ȟ��2�_?���5�%$�,�p�"O�,���ֆ5t��ЋŞdǔ��Q������\)�0�����0|��'�5B�� ��o�/^�����X�<�gh��(����T�|���j£�{����q)����g�NVj��B�i�
 �5�Y_Շ+4���D��=pN�e��bނaS2��D�[:H��B��W�x�҂�]��-�R(%pC�Iv瘍XW�\�9#����L-i�XC� �dM�Lӎj��M�Ħ��p��B�I�vȲ�1���������e'3�B� u�
�a��Q�L�����ǫNLnB�(}��1'-�*	@�P�"�B�,��%[�%|w@P�l��%"�C�I-�n���'cM�0���ѧ@!zC�I$f���P��+��j%��%y�"C�ɀ���R \1P��\���
a{�C�I=ɚ� `HS�4�v�ye��)��C�	#X�*��&���\�y�`j��WP�C�ɟs��3�Ǯ	3p����Bm��B�C@����#�6YHe���5@tC�	�R�B���
�=-&�K0^�,C�I64t���K(s�vIHũ�#y�xC�����iB�m^ �S�"�t�VC��X�BD�$�_�����ܼ)�C�9	��0Ж*&a�)�D�*RDB�!1eŇI(.1��f(ÇW(B�ɀW�z�C�  �GJ�5�T�]vB�	�$
��#���T-��;c'ԁ@�C�I]�8��_Kz��AmR,TC�	��0]*�L���m�4�STC�C�I�S��`nV[��Q���K�`�xC䉜 -�� Rn&d�,�W ���2C�I�cc�A�vAX'�����Q�qsC�I<T)3�[t����J�1��B䉳r>�0@�R2�r)��E[�5�C�	�j~uB�:c��`���<a	�C�1g- g$τ37(�J	�a��C�	qwf)��ۉA8"�J�O�< C�ɳ05���g@�E�0�ޘE40B�I+~��ɗ�F
31uk��P B�)� ��(A��t��	WǞ�@ۄ(�p�'��O$a��[���e�͆a[4"Od���싥]���"J����CĚ����\�S�On����H�O��)�mۑO�B�'HX����бE����"5
B\��y��'�y�%_�+B@��Gn��,��,�B(׃�x��'\���'oO�#�L����Z�"�B���OXa�v燓,�=��BʦHG��@�'��OV< ��%��0���"b6��a�"Oz6/�	�|���3\M��"O���5�0 �9��]�x睊�C"O���ڧ[������P�g���`!�䕇k��l*1�@�D0ě �O�xm!�ő;�28� @;*!�իcKzJ!�@�x xԎȕx�+� /E!�L�-�;ũ>%��+f��+!��F0�<�@��&|x��#�!��Z��AC.�C�>ͳ�*L'
�!����������3Hz�<�P���!�X
Hx����Y����b��!�ʢ18�H Ǣ�{�`�3�P�*9!�ϧJͤ��G���ؤ��o>!��3T<�ʢ��NW��G��!��S$���8��>E��y��Ym�!��|���%NN�{� ��A�A�!��U�K\��A1(Y|��a�3H�6Cr!�d�`CtjKI���6�Qu!�_>$��IθCl�Fœ�]���°bY �B���D}�D�u��5u���E �ă�Kܖ@�R sn<m�<tA1�8,O8�8D��� q,���N�΀��Ã7*��ȓ/9
	PR��4�4�P�_FP8�&�Q��=	�qO���I'$�j
�f�7#+�eQ�"O��+�P�raz�:&&B b~�: �)2�p1���L<���D0`)F��d���"�aH<!a�a�jL[�MPh��R-P�Y�|@6�&�O&-3��ܪw�ĵ��ő�W��آ#�'�z�S�c�	�#����D���š�S� �C�	"R��$��4�lW(+�ޒO�8�$,7�)������gI�p@t��_�B�%J����D�,�́q���q�B�	^��5P�瀪L֌i�ì_1�B�	�J�T⁦��r�z�R�`!HHB�&g~��j��S �M�gm
��C�	3w"���%�r�ҥ���E�r��C��>>F��`H�R��C�	̞C�IH�Lt�@L.!]�չ�'4B�	<;�H�h��k}��1�ݬJ,B䉚�hɨ�nܒ:=ލʷ�
�B�	6Vb:ز�I	t1F��l=�C�	�RC�a9��Ȑq~���I%:BB䉝adP�SȀ:�,�3'G3[vLB�.����V�T�69h�*���C�I�EIR9Sq�ױ?.N�jd*&NB�	�eN|xsHW�$�L�b�B�	W�"�a�L�LL�iA���:�B�	0~５鶩��ą E!I�0�B��q��l��Jk��qyuB(l�B�I#�D@:��]!�����nC�H6�B��9 x�-���-p��/@�&�xB�	��"����dQ�Ҋ=�C䉈|���`��$�4m�C�	�e���L_�ո�(��C�	>�x���A�_e*�bv�=tڸB�)� ���f�d�-��7�l��"O~���f��bW�]ؗNܴ>���"O"h��E	1I�Ѳ�k�]�R��W"O |�e�5Lx�u��M,(�}��"O+�T�;��q2o�NKܬzC �y�'n�*��ӕzF(���<��I1$��d�BB�4p<U#7Mϑ'��4͌�l�^�I#�ӵ������݌v��B���>Np}�"d�!�y��)yȮ����S�3Jb��r��>��D�-$����dɳ��za�,m���q��
j�a~�JE5�y���8dw"�7�Κ{>�D+p ˀ�y"�ԇ7t�}P���?A !��`���yr�%iFZ<ِ��Bt��ㇲ�y�O&g�ҐPcd�
n�,e�����y�F��"��mcCB1`\y��)Ş�yk�7/���#7!�T~�"ÏK7�y���QDB]�#CZ$/l��ǡN�yr�FW���W9&g6�W��y���|���K�"C�wEӦeB2�yG�p����3�����!Fύ��y�N��L�f$�fˑ�z	��E�J0�yB#��c �� L�{Ob�+d%�y�iQ�U�D!���.t
�,!�+��y"H?>a�Q{�͏�k�6i�Ad%�y�[(�A��E�l�E�@���yOΰ]9����*ށnX�% ee�y���.0j������V����臬�y���P���%�?v9�$�_��ybO�,�6�p&�T��T4W��:�yrᕗH4�\Jv��W����ɔ�yb΅�I���Cr�+A`��:7��6�y^: ��<���<>�|��o�2�y2�J�]b�)R���4)�B=+F�Щ�y�!��^��qx�$�=��)�k�ybnݶ{Zx��T�=�~Z����'�v�����G"T!�l�sHXP��'u���` .�����r�t��'�Ѐ��#� �$4���B7at��x
�'��rUD��0Q2��vK꼹	�'a.cR�V�T�|Xɷd	�JaX
�'5X-;
��@�p2@�b����'��xEnY" �,as`k��Q	��'F`���צs�zd""*�1K=��9�'��k��Kj��vGD�S�8�'0bY��
:\�܀j�,)N���'��d�F�zf`�����S��A�	�'�x�3]���@�ΐ���{	�'������8
EV%���FIl�	�'?X��!-�W�2�;�N�2?2X�0	�'����{	�����#^@yY	�'�vѩ�C^(I6�xB�Q�		,8�'kRѩ(�/��A����7 ���'�.i# �~C*�)c�Z.<�Ū�'��93� c��A�2`�x��'���5��87�5!�!�z�.!;�'Da�aDA./�VhK�ɐq\"�Q
�'���ǩT/`&�%�s�� x��p	�'�ޤ��b�/u��D:�%�T=i�'��q��B�-7��-r��	��X:�'/i���R�A���!�$э|�����'<z� ���1���P�<y�>0:�'��j����w
h9��Ѽ	~�	�'��x8E#Z1Y%�%Z%B�9T��0B
�'�����:�<�
�eĽD���p	��� ���$%]�ɓ�:X�~�Q0"Of�!6�D� vM���n��Q"O��WV�O�$�z��5Y6���"Or��p+�$)��*�ȧZD0XZ�"Opa�!�]�Dq3m��
��0"O,�2�ͭu���%&{o��&"On� �2�F�gU�4�"|�P"O�2k�#Q,	����@㰘�#"O�86$�3�����z!&j�"O*�� ��y�I��̓�\��"O�XC�FD��j����1�J��6"O651c"0q�ꙈУi�6��"O\8��]Q��T�!v�~	��"O�A��Ma�2��*#u�dMӓ"On`� 	�!�*��(H�j""O��z��!+�Z� ��2�t��"O�	� Mx�<��'�)<�:�@a"O�Hv R����Q
�=�%5"Ox5�Â[8]����P���Er�̃"O�HR ���������� _u"�B6"OV���j�&!@1�woK�LR�)p"O<�W@�P�J���N��6�D�p3"O\؊�$*F��L�$+��s�\�"O�0�'�%f޲���Kɼs��9�T"O���W�@]��H�߹b	�xi�"O�1�"�:p<Y�ڝ�Z�#�'R�-�e�E;s���2s� �ti�@�'v�e��R�(:��2�7\�H��'�Z���Y8TB�aҠF�|��'�ش�p�Ͼn*1W�=Ѵa�'됥Ƞ�ZZibD
�	�4�:�'�XT���$.���f�������'�H\R�iB�&���0�����䅡�'�j�z̀�M�4� �%�-���'��PA)���aA�� ^Y�02�'Td��P�aА���.��QLj"�'�P�!'�9-��,��a�p��|��'#X�P�b*���WfzDJ���'F��j��� �΀*�%X=v���	�':���A	�������M�'�zh�n~NŊ���	�rX�
�'A��@"�]R,z�uc��<�c
�'�f�YN��Ӭ�Q%O�-T�*��� ���@i��*�b�-�8�t`��/��y��*��X�e2.F� �Q���TUa���n]J\��H��>���ȓi�F��nڳ��@ʗ/=�]��9��	�lə'~����xՇȓfp&����r.F ��[9Ad�@���P4u�
~�]j�
�5p��%��O=�����ȏU�p��e ��Z����0��Xrʍ�\m��*���%�.��ȓS�d0��!ӨX�4oE�hb�ȓ�0��I�. ь@B"`�J;Hp�ȓuJ���ֳs�&5z�`�$�ZU��	�!�p�#	��%�AdǢ?�" ��Bh�[�ɒ�zJ�Hq�G�L}b�ȓm'�I�A�¬;8��ъ�JY
���Wm4�Ra�)]��<HфY�d���7�bWLI� q��UNB�č�ȓl�zco<"| ��NF�FY�ȓi,�`��Dlv5�r��KM��jZč8%d���[�*�?)�Ɇ�(ք�j�Rp��#�b��%��S�? �I
3��8�yb����R0�T"O��G��~�@�pT�\�9��y"O"�ڳb��zpHE�ޣYxd�%"O���%��E]��1C�=J
��"O�0���!���	$��$HP"O�D�bċ�ͩ�*ݘP��A3"Ot��q/_�)g������3�0��"O �R�λM h�	V�B�)Ѵ��"O�U	�*F�̅R���ע ��"O��*b��JV���u�\46����1"O�uSW�]IK�`��#	m\2Y�"O�Œ�G�5,Ȩz����FT�c�"O~1
��"��D`wD2P�˰"O8���N%�f�@e�^ĺX�#"O8i�@M�=�>,�0靐T��H��"O `��
	K�(8B3�Z^�<��"O�	Ӳ�Б,�$���d��$��"O��x-��9�Ԣ.A9 A��"O��k5�̈_��a���=��ۗ"O��Z�+֪Ep��B��4Ft��"OL��"����ba�P��W��hD"O��r@�5�x�A0�	>�h7"O��!��9L6��iр�*dx�|�"O�D���^xe��Ц(,xdX�P"OD��Z$=v���d̺4�ey�"O&l���% �E�'m�B4@"O.4�� ]��@�b ��q�"O�%���B�`1�%L^��r�"OX�ەf��P����##�(�P"O�vG�?�>Q�Qc����H�"O�����������2�,�8�"Oة����
�p����=X�`�"OJ	�6� �S�6�(d)v��;�"OФ�l��
��=Ae�ۙ:�f�)3"O@����C�Z���ϑ=7i��i�"OB�$��}�o�u[^Q��"O��&o̦����t���W^��HE"O����޸%%��i�)F��h�"O|�KdA��]��H�q ��"O����CH�f����B1��"O�H�!Κ�B�$If#ÓR6 ) "OH\�J��(�h�RӃΤ$�H�"O��X�O@5��ٲ�i�Ը�Sf"O�[��[ rHa�e�?�U@f"O����MF�e(��8�kϓ��{%"O�X�h�.wV��@��M�"O:;��К% ��E@�^����"Oj���!C� X���H�h�&�+�"O:q��Kƛ::�H�ECA�z�\ 7"O ���+��9��|HcI�_�vق"O��)B(�>|����&�Me����b"O�0AޛmĠ�)�ݩ�JaYg"OZ��#$�-X�<93'Hˤe~r���"O@�x����Eɇ��B�L9R"O*ܚ"	�a�����B�g�l�'"OT���G-n$j����M-4R,1�"O^ىWg��G��yW$�v�|��"Of���hI$�#%L��XhP"Ofl��(,<�BT?�#�"OD�X�RI&x�7��H�e 5"OJ�¥J�]KxT*�G�$b;2�� "OԤXw�B�m�1�Ӆ��?t|�""O~@PTl%�� d�h'� ��"O�IH�53��|�F�! ��""O� �0��/��E<�;S$�a4E�6"O(���m�N�4��㙳��p�a"O��	t�T���VB�U��+t"O����L7�&�Bw�>|)7"O�-��>D�l��CX�
�-�A"O
آ�+)�4QR��,�N��"Oܡ��K*�-ʦ��-����"Of���W�[.��4FY\��D��"ON��'X/(�}����*U��Y2"O��#�Q�n(´E�����"O��ڐ�D�*���P[2=rjE"O�]*�� ��Њ�n��^rZ�J"O^�"�n^TR40��NA�9��҅"O����nX�e(�)�fb�hpʰ"O t1�E%	<݉�C� ��1�2"O�����!E���*ţX<w\uY�"O
��Vۋ/)Zhe�?g|Є 4"O� �nG=PD�����DiY̸
�"O(��(W+C�"qǅ��AeR�"O։� �Xy�tEb�枺-<n%س"O~p�%�K\׾)Y���!>��A"Ox���i�2Q�ܱW�R��)��"O�HB�JMV��Z�ğ-(ӂt"Ob�2g�O�v�LণD=t�aia"O<(5@ݮ1$yU����I�"O�T���D>Z�$���b��^.,�x`"ORt�-K�.��M9WA@�]���2e"O8�x�+�1L����e��:.�l��c"O�k� �-!�Ӈi�P��q;v"Ot��%݃SJX؆�O�l�v�(�"OT�9�k�'b���3�	��-��xS"O���pĜ7�����B�/z��K�"Ozx�9 ���ҋ�2x�����"O<E��ᘤ$U8X�5O�A0r"O"�b �ªo��#r�,mƘP"O����4X��Pr%#�;mVH,�Q"O�Tq�b&W	�	�a�e��Q{V"O��(b� <x��20��u1F"O��B�f˜�����-G�0��"O��"@��XctKͲ>_���$�/�0�'��(��x��'�Mk�O�7�O��G.pD>ŋ�f�ZY��2O�
/O��=%>�"Ed
� 9P�p�i_�;��� &�9D��2a��^�P�{t�ǥd�$��
�<I��Ez�)�43q"� Oh�����TCƄ�	��HO�>5`�K	�t�<�I�q�R!=E�Q��[�';CT���dC.�p����w�ҥ�>!5�=�S��j�x���"�"<�P1{��L��O֥j��)��%׊YP!+ϛJ:La{��d�D�Yx�"<Y��)�<OQ�e� bG;,ECԡ�*>���	Jy����p跮W�;�@hXv�="H�F�ɤh��"�nѩ:;p��	_0���!g�Xi�+u��?�O|��-��LȜ���΄��1p䦈h��݉!**�O�=����R��Ts�X�M9"������,��F��j>�=E�$Ï�|L�D�R�EƘ�J'�M��/�I'�0|��M̋p�. ���̠eK� �釂��'y�c���eJ�O(���Ȉ3�fU��^;g���"�Oɢ�v�D�O��>�Ɇ�v4��ϚRc�x�ǆ���D3�?!%F,���NFp܌A�X�闎�i����'�dFy�����l�dn=W_�L[ԁ 8��6��U��ȟ���$��7Z�S�F�G��գR�I�0|*P��2&�.��ժKl��*sMU�<�����4ؔ�V��8��,ˇ��P��hO1��[�B*yA K"�ˈ��IQ�d~Ӓ�O��S�B�7+ZvuJ�`Pw)�0�왫3.�x�>q���K���� D�����2Pv�סN�r��a"ObA#ԤH^�$1��P*7攥�`"O��2�<>��0hֱ���Rt"O !�dnJ�}"�YS��>�}K$"O,���o�Y͔m[c��n�	�"O>�+�gVk^�t�Waڧ`Ԫ�J�"OJ=��F�=e������Tg_R���'��2-F�<[H��Nܡ"LE�'�j�@qD����o5�a�ӆ�y2�1�Dk@���r�b�yqE��y2DN0	�!KcI��q�H��P�F�y��Q���c@��5�8-B `B1�yR�@�T&걑��
�,�LPЧҽ�y��O*<0����ą�)�5�G&� �yB��/��u�Q��`s��'�yBM[�tV��{Ci�E��TI����y"���`���!���	���8�E��y����fC��{��T�rD
�yr*P A�p�C+ٲl���iЦ�y���_��ő�!��aB�5i�gL�y�n�'�3Um��&rz����y"ýs�ĭ��`���p ����yrdS�x�R��r+ߕH�ґjK��y�C5J���8���v�C�y��A�I�	ӁӜT�,�5��y�!N�(�8�����;�\5�%���y�ŗ-p�h0f�G��%".e8E�� j"`�S��EY��I<T!���h=���'��4<E[��\�!��3G6��!�%��?�x�s΅2j�!�S-\kV�P����e�^-��,���!��0c�ш���W��S�+рg�!�X:,ÚHS�ÄM�6����W�!�$�N�đX�&�74�|�2�,-v!�D]&I��P�0k�*I��%��HV!��=dͬW�a�J�{�	�369x�ȓ=����pZV雴��Z�"9��3�
�tA�!�dpS��'^��ȓV* �ۖi.7B��AG�	P�����J�D��_��@Q ���2�yz&"O`�P5)+7H��7옲s�yb�"O*y���F�Lh��I%S7D���"O��T�\��v��dj�"O@eD�B��a�ȽV�� ��"O�A���$;B�[��]���#"Oe(񀉾W�z��hؿ?�5j1"O(�� ��*�)���
K�<�z6"O��j��7 J�0�'@�[j���"O�y��f.��H#��.P�$yv"O��9��K��27�ȷ/B��b�"O��Ӣ�9y�Yh��_!@�1ѓ"O�q���0q}�,R���,�Y�"O���u�O\�y5 6��i"O޵ш�9}l���Nލ�b�q"OZ��iM�r�vt�w�Ԑj��ɠ2"O���J�؍�F�ɠ{�x�"O*�b��*D��Q�@"N���w"O<�[F��<&�8�3Ø|�eQu"O:��a�S/`	��`/ �Oc�i��"Ov��BcU@�������?G�-�t"O�-{3ɍy���)#-�05�� A"O��o��p�,���͇�%��:�y�Eg1�z0�S�� X����yBF�1�$�u�����i�����y
� ��r�>-��P�q���h����"O��)��Ք^�`��f��<�ڸ�S"O8I��+�
K��m	�	�+lpѱ"O8�A�Y*C}�S)^&[g��2""O�I9Bɔ�X�� "ӨƾyV tQ�"O���޲b���DhG�B��I�"O�(�4H��8�H�BE��r3�%I�"O���fǓ�?@6�I�%6lSP�#D��r�E'N
m���H�@�+��5D�\"�"�fݤ5�7��gF>�{F�4D��Y�L�@�� �!�ەK"e��i3D�����))�x3���!��%0D�� Э� Tf`[��F�X�����#D����ϑ6$��p�r*48�HII5#?D�R��2w��<rt�M����I0D�t�$̟�b��g�~b�`��g)D��8�-_�|���*T㗳Rtvɸ�+D�dkT-A�
���ʐK+c �Q�/.D� �1MX�o6�1�N:J�&E	�?D�8b�	R�|���B��8;�DP8�E=D�8�2 ��x�#g��r1X�3�#<D����!֯
H��ڷ �[�P��@<D�ء���7�R����ج'ˌh�� .D�H �+��dw(H�"l-a�>��-D����Ok�aC�O�0�<x{�$,D�,����.�}	m]����f D��Sqf
bt@d��%@*1t�s�k9D��s��E�W�|��VA��pt�}Y��5D�����1�
�[F�B!yq �u�3D�P����t�T�����nU�Aa��/D��J�эhVL#�=�J����(D��B�͂6���'�?�� �-,D���r@��K����a�5�J���d.D�h��%�/�*��V#�\��2�&D�0��H��p��Q����"m��	���9D�p��B�@�LVHcN�2�N<D��q�g[���p� L�=�L;�9D��8#j"�t���VZ�~�@p�7D����x֤��!�T�!�h +1M4D���霺)U�-R�$�$`��1D�d"�<6��� �Qa-ȠcC/D��ʲ��(�:h�,��4��,y�.D�88�h��DzȈ�"�(:j0�F�&D�4��SM���+rfV�ND�#/D�(c�H*{��5�4/�#\�����+D�����.H�	�c�gaBE��(D�0�!d�Ve;J��e��`0D�P�䊝;KD�QE�P�]c&)D����ǘa|$��P2�!#wI+D���D��:�$Q�T'{z�i�4%+D�dP`��=f�uAV 7����,$D�,��N,9I��!�J�rY��z�>D��y5`:0	� 򶈉��xF�1D��a�ҹ8���	���Z��;D�ظP��-xљ��ݯrtԐrN9D�p���2_R����N�R�u�5D�S�ŝ1;��h6�̛"ۄpQ�O5D�T�w��:q�h2T�E�n�4��4D�<{�
�Pm#WD�K-��(��0D�Z̛3j�!�@.�� ��賦C/D��PdSR&j(��J���h,D��PfX�;+�;�I$�����/D�p����B��u��i	��� bg� D��A�%_��hj�x���a��!D�� ����m��S`�0�1"��0�Qb"Ofä��0,��X��+����T"O��Q�k�$E�(��' �?��=��"O�@E�7{[İ�d(ۯq�t}cD"O,����!6�(H1��G,�\}��*O��q�5�J���aV?8\��'[V�y�J�NxֱIe�X��2�
�'� E@�JX"#82!
M��_t�2
�'�L�`�'&�&��Kڑ�J)J	�'/ށ���^9&D	r+�p��p�'_� d��=^h�it�\7k�<�S�'PL@���=����^M(���'4���e*Ёm��|!�-�-�j�k�'��&`
oP.��(�l��'�V(�6��NnH��^90P(�'�ι1��4U�PD	wͳX
��A�'����@�*��qA��d�8�H�'*m��
����s�A�)�ƈ��'�`{![b��р�%mtV48�'ߐ�qR�21V�(�B!g���P�'VVK3h� '�A�$��-H��	�'��	�S튛RT�D�̓,zN��'��q�dF?*1$��)�$$d"Ej�'�dRvJ�>� �� ��3�X<��'���A��	
\��!�#aʏ@�r��'��%AQ��C����[(I�Di�'k�]�cG��V�x�WC@�DD���'���N�+�*]�0�L�t�T}��'�t���M:���`�hREI�'T̍���)G���a�O��| �'h��H�,/�P%0!O��v b	�'���H�]� d�=�1�	�Z����'����I���S�۴Pc�8q	�'�l�Q-5N@� 욧u���8
�'�����A�T�Ѐ�ףl�"D�	�'dxXR.��ځ:��;5V��ȓ|e�Lxvˀ�2x��k��5#�$<�ȓV�����\�mSP��/sƀ�ȓ0�d��
�6 ���3)�ȓ?�@��
Y��.­Ƞ�B�<9�M�#_"̸!�̒m��(�ac�<� #U�����T�Cu����D]�<q4.� g��Svi�&ل�Q�m�n�<q�CG� S5;j�\�/�m�<�7#K�b��S5m��-�*�m�<�5욒r�BP/Q�&� �%�Kh�<	PI�5��{�-H���Y��Ta�<�tA4j���mI=t����i�[�<�3&C6P��˰��1D�+���S�<��(SZ��p�֯ͧ~��
Z�<�%ER���Sɕ�{�2M3�@WT�<aV��
(
y�$%�(rΨ �O�O�<���OLƴ	�f�Z��T�O�I�<�R�L�i��:�I� F	�q�f��E�<Y�ךY����M�sD�Aׅ�z�<��޴�~�"�B_ �Z��}�<�1e�2��A��K�I�zDB�/�Q�<AH�Wt�Q���3	��e��aJM�<	t�]���a�Q L��v`jI�<�!H��)��_`��
WA~�<	��ݪQ�&d�u�֝M���T��}�<Q!�2s���҈�//\HRÌ�w�<�#IVM�"��`�,���r�<�a	¥U1P�6�D�P�Hyr��q�<� x�re�H?��c $UD�Af"O.�2��N.����� `���V"OVtzVH�]�y[�E�,n�\DH7"O`��4�Q�0����+��"O����   ��   U  "  �  /   �+  �7  �B  �M  X  a  6m  �u  Q|  ��  �  Q�  ��  ֛  �  \�  ��  ޴  "�  d�  ��  ��  /�  ��  m�  X�   �  ��   � �   # X) �/ �5  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,�DP���|�I	$G#\����Of�Q����<Q䔜Z�,`:�'MqONˡ�̳(����A
D�~����5�S�	��������=w������Ui��8E{��n�)Ϝq�c�ߖd��"O�81C D�I�dl����5jyR�i���jӮ�O̢>Ir��v]dvB^�Wkʄ3%A��$`a}"T�<�% :�@��g	U�f�=[�<����i��&&N�S�����哿4cV�=i�'��>qz'�k���SbӰEW-*3@�ϟ��'x��Gy�g�{�I�j�:I�w�2Y���c��ʭE4��<aJ<Y�rL�s89���7A��)7c���yB(�$<�(7��?�XeI�h���:��?�&��ome�H�c�j��cP�ώ
�R=lZz<��	�K.��A�ƋZ]8�FE^b�IF}"�x��O��O*�kP��k����RMܘ{�����'�<5�7��}���)��{K$p��'�	C�)�L<�q�0.�b%ڢ�f��E�2��Z�'��<���7[th��"��DO�E0��Y�;D��&�H��8�J��NC"jh�j`M{���d,�S������j`|0&X��e�5H��32!�d#g���"!�*ܓuB�"�IU���'9�l��y�#�,K��2�ȓj`�Sb�����**>N8}�ȓ>�-C։ӫ	m�ҡ'O"1s���S�? �g�Q=����i�0z��(�"O&ts�!g
���*�:io\����~>U�Df^���1g��Ҹk�m&D���am	6��G�3G,���s)2�O�˓��3��ؿ!^D�����+	�6��ȓp<�(h6H�Նe����%{����q�k�ެF�(�bd���2�ȓ`��`�A�(5�z���V��<(�Ɖ8����$GF�r���?i
ӓ7�@�y�@ϭ!� d8���p�t���5.LI�0�A$4��d����Y,>��QĄ����]ʵ���	7�Gy"��4lZK}�U>EX��Ñy�|ġ5O �/t��C[�hO?�
�+�:KA:<��p���7&��'xў�>��C"8��4��윊@
�[��9D� #7L��@R�q��f#�q��YQ�'u���Y���s�?�a)b�V�FX�KE�$D����(�3��Q��R���q��@.��M���iO!�Xa ,Ղe��ԃ �RW�z�i�O���Y�yFh��6i�#TQ�xC�i�'��>�	{����Ҋ�"Fj5 �6k<6a�����O����.22��h��0:� H"O��[�/�4�zqAA���۰�'2@�O��[ը�	w�4kd��9���"O��@Ώ�Hp�rW@43EV�c��x��'�2��.U�t�fT���!&��	�'���l�6�)&�T�d���'�"ϊLS�Q%O���qQ�'.&�Eʺ}���q�éJn<��'F4 �L4��X�e&X�9�8Y㓂�ta�G�7�< k�C�i�x.�2�����U���"u�ȓpm���� QH��r�'Qn;t�D|"�'Y�>�ɲKD [�l�`)ԫ>�ũ����hO?�d��{�̚ �N��uF�

!�$�Y�����j�4u����%�!�$M�Y}E�5 ����͝�c1Of��d��T�5Q5	=\�^���O%SR!�3W��pJ�N��Q���e�$E�ў �����ف��7�!��I�Um�<a��T>m{@���@��+6��PΤ�Âb��=E�ܴ71�:���^��Ygl�,	��p��n���B�*�z8�q�$��pr�\�'�a~��$7xM�n &"(@Wh�yR�г6��Zb�<m�X�`�JY#�yRG�-��A)��e�L�IAf�>�y��߮F�)��f^��:tD.��O4�B��	��uڕ��Ԇ)��,�ҥ�|�!��8s1$4KAC��Y�^�O�7r��	��HO�>�Z��c�M��%�
h�c.}��'\h��w�F�&"T���)�B����
�j��I�G�x-�eV�6D�e�N�P�VC䉯ߎ�yg)S!�*XF	�+tFC�Ɋ �8a��3e�9���
L�\B䉴wM�&S�L�u+2k�N߄IC��)���9�*бge�\�[,L��!Yu"���E{���8	9���%F�(���4�7�!�dr6��6O&!rm��+��b�'�a|��Y�h� Pf��!hNT=��J��y��@�"�v��r��*5��ҷ*ׯ�ē�p>9Шǁr3��ɷ
�4�yۃ��_�<ac-�2
I2Y�SN��L�B� ggAu�<	CB�(���T�ڤs<��j�MX�'?���D��0�5�C��||�9��f(D�� ����l�C��4���ϤVz���xb�'2�QQ��t��:�g�!3t�(	�'��e����*����C��&č0�O�e�TC<�,�З��\6���'��	>�@)�Tiӧy����Y
Ad�������OH��nU�D�vM�&+�#<"���� �ȟ�̸� 	�0���A	ڧC��"O�A���-><�	W��_��Ͱ@?O��Ȣ�'=j�@�3f��L�<�^6B\���ȓ8t�;@$U�0��d!͛M��C�I�_pdI���0����@�g�xC�	�<]I��0YI❋�%� �F!��q���Q$(�����
T�8�LF~��	�?��
O�-ڂ�: ��x��#�/D��3����}��0COV�b.v��m� B/OF6�<�O�q��=uE�:t�D@Zfi��vZ��c"O��K���/3P|y҃�S�{j����o8��<E��'6���BCm��c�CQ5&@���Ib~��R:w��M�Q�ܔ|ZX{r���hO
��d�"�4U2���t�rF���{󄊑�>C�o�/f*}z��־C�!���25r�v0����M؇e��O8ӈ�~����o��2��	Q�Ę�A�b�<Q�ƺ^<�V�^�J�
�
�A�V�<�
Jh�z%�DD��sJ��:�	�Wh<���Q�`vR�I��36d$s���$L�����	�Y-��!�C�'$�̠H�-КEV���3?y+O0�a�:�b4����J[l��=O����)+P�`�**>n�0���4b1O*� ���ɉ�x�r��ԥԾ,F��嗕b!��=V<���Z4���0�����D`��"<E�����0�Jե�A|&��P�[��y���B��eP�/��:%�HP)��y��0>�
ej�Ғ]f��x��ҟ�yR�Ȇ�V�#�MGX��kR��y�W{�0��K�A\҅:@T��y"O��2��k���o�Bū�d	��yb�	8^�~����Hg��0�����y2	^�5WL�����6-g" �GAJ,�y2��j���M���0�;��V��ybW<�
��e��8r�i��%ق�y�ƄV�ĕ{@o,��AfB���y���/�j�h�-G =�x�q�KJ�ykW�6�n���4�m�UaB�y2��jz젫Ƙ))  Q�D��ybO�	mL@)b�e��
q����/�yb+M+@(�Yef�[�J�@�N	��yr`���Θ1v�P@�+`NL3�y��]��a)��s7=�wa��y�&O6;��2���V:��T+�!�y����*UR�@g�ȩK�TY���@��yNщp�������*9��aKed(�y"&��V6��A�n�1b ���ͯ�y��W�J�h�`m%H�<q�� �yr֧=�F���+�m��Rg([�yҍs��p���uZ����y�M���&�"'��ؗ[�w,�Ňȓ&���@��սW�l��4��Ԏ%�ȓ��<Sp`ͺl�^IZ���~��$�ȓeH4ٳ o��V�6���c�ø��� �|�*S��VE��@# ����ȓp��a�Ҫ�S�n!��2[a��C���VJ�#fzYuרek���;|D�P�!Ա6Q�������J��S�? H�nF&#�t-�q@P�d�xP�G"O���僟�4����H=�x�i�"O��ڣlXj�"�P��#�D��"O����O�Sy��d��!_@N��3"O����#��
e�آ	>؜���'�B�'
��'�'�r�'���'���3��o|�#!���"`� %�'��'%�'d��'��'I��'�>�ѣIM�xP��1!ڃn~���v�'��'#b�'A2�'B�'��'q���3D�(�`	]Ƽ���'���'b�'YR�'���'a"�'��jR�R�IZ�8��6 Ur����'�B�'C��'�B�'y��'�'�`A�D���~-�QCk�20(���'m��'���'"R�'o�'5��'.j��V��=!ۋ��}����#�[6�?����?��?���?��?���?q���=�������a�H��R�T!�?	���?����?!��?����?����?�3�+ma0a�b�M�~9F8����7�?����?���?����?����?��?�s��QB����>�It(�(�?���?���?����?I���?��?��F��� 9I#F�9dfr�0 Ϟ�?���?���?a���?���?����?��n6qWR3A��|F�=�@fΓ�?����?���?���?����?����?����8;�8@ǤY5~|����1�?I���?9��?	��?���!}���'G��&X{(�"�EE�u�U{U��� �<ʓ�?q/O1����MC��)3��QaH�c�`��-<�ޕ�O�6m8��������A	RCV��^�|"V��$l	��M���z�vn`���+�ƑІ��!���Oh�ZA�6t��@W�ڗ�у�yB�'��I}�O7}�N��h�����A�H�c�wӶ	����&�'�MϻGH 1T�޺x�P���Oԟ���z��iF�6�|��ק�O��9y@�iq�#րh�h�;iK�9��ҜU�D�]���6�@;^.�=ͧ�?%�ĵ:*ZH�b/X1휁+B�<�+OR�O�Pl{��c�Ё �w�dԂ��׾p���x�JH]�'��	��M��i��>9N�d:�᢮�.Z��<z4��`~bG]1Z�i0�-��O�
A�v���V��VL~�:��ď �iòQ�x�'���9OF� �B<O�Ⱥf�83�-��3OL<oZY���'a�v�韪�"�\�_]�	r��ǌ��S<OJ oڌ�MS��F���ش����/���B�kʁ��|I�B�4{�p{�B��jhJ'�.��<�|�<9Z">̳B��S��)�GX�eՠ������	cu�������X�M�ڬ�3�H�[��u�aJ˸m�	��M�C�i:ɧ�O��}��H�Z��#Q��	��s��ފS�l�3Z��c |	�E�;=��'�	
G(tx�pN�����qb����'}Z6-��>X���4BT�`�ֽH�������!�Eզ�FxRQ�([ٴ+p���'jL���Tg�ډ۳��<��E�Cf܁@b�����e�9T�X!3u�e�l�P%a�A>�
h[q-3i� ���L8�(���,���z�3'�TEs��!b	D0�z���.9}�p��t�I���idK_�C��1+t�͍x��,�j��H��5����T��(��˭O�>8)�IZ�_���e��o�JTH �Z��!b���?z�)��+gB����%h�����"�t܂i���B��"��
0釬�!s,�a�3D�uR��� "���X��8/�$�0�P K�\�b�ۄC�PS���m�`�u��>���t�	2;�t}pv�6f��Hi+Y�5/���%� /<�%ȴ�o���d�O��/7����?���?A�'�D1�G5Hh�EKQ���U�ʡ�}R�Y Fm�'���'7҈O8�H�2fJC�L�à)��.��7��O$Ցe�<���?������2B�4C�ȵ��+_��̬"�%�n}�� ��RP����Ꟁ�	Ayb�׌9N�p�w�Y-2��1��=)�6Q��V� ��ϟ �IS�ϟ�	�p�Ajc�çB��+�O�&;����0OQe��ꟸ���x�'/2�3W۟vy��B[�-��"RK�1R���w�iS��'�B�|��'��N�,^����K�LE��O[��X��� ��ğL�I��'��e�S[>�ɤL� z�J1`��гA� �i۴�?!O>	��?���@�8'�QЃ�B�9^ԡ�c��?�pm���Kybo���ʟ���?I�P��:<�H$�d�R�)�
����?��"܄����nIsr�3\<-z�`�F��4"�iO�Ɋ1D��	؟,�I�|�SbyZc-x! �BAJ �#�d�9����ش�?a��s��UGx��� �"��	)#�G��ɑƏ��M{����?����?�����*O����Ot87J�eN�9�d��6�\��j֦�@sÎ~�S�O�	#b��&�;m�|QRV��;��6��OL���O��	�ǰ<���?���~�e
z.�$�GLG�Y7vt����'�xٚ��|��'���'e�1�	�(P�q��O%#�4��kg�6��̇A���?����?�J>�1s��$��G�6t����aM�@�ֽ�'qxpƟ|��'M��'j�73�~��BNH+H?`,�����F��
�ay��'b��'��'c��'����c�7}>���Ȕ4#��#���'R�'��W�\jsLOx:6�t�p���Q:��Kt(����Iß���V�	ß��I^~Q��z��q��U�8,�����GA�'�B�'|R\�l�ca�_��'ӆ� �����9*�\��eW�I��u�3�i�B�|��'�R΋�qO.ɒ���7�t�	p��i���'�割S�zE�O���'��$\:x1�hy`c3Bv��H�O����O��@2�O�ӳ^��QK�2d��n�#r>p7�<�RJC*�f�~���ⵞ�����£2(%ٓ�{�Er$-g�<�d�O����O��$>�^��4�fX�1a���,�E�5�.�l��`^8��4�?���?���"���\c�xM��R�{��8 �L�WA4Aٴ�?��?�����|�'������l�� � ��$�x�����O��Dۦ�'���� �ɺ
0LA�0�\���aͱ>h`�:������˟��'2h��<I���?����@)J��iQd��=��j!�i���Q�*bjO�	�O��d�<!-��Lr��b2o[+K�*U��z��Y����Dy��'	B�'�I�rݺ�ѥ-F7�\ ��^�!�F���Kʧ�ē�?!���?�+O����?m p��*Y�AÃ�7��i)�By�����<��3��s���	�K<��'Q���RGJ�U?Ҹ��@װ-Mp�n�ޟ�	J��?I)O�%颰i�4�P$���f�X�p &	�# �� L<�����O�|j5��|�����C��ݮ��D
��ɚj����i��O���<�VIe��9jܢ5���6�U�J�Hy@�k�@���<��t%�(�����O���ƨ �d���K���k�&j�&T'�x"�'��	�D*�#<��3+Z��T��?8# 4�Ά(U�<��'��sw��'���'@�dW�֝1m�x����%g��!�)�"lT6��Oxʓ2v�4GxJ|
�FD+j�`!Q��@ڦI��!]�1�!�C��M���?i��J��x�O!Za;�f@>@��)Ϝ^�����'o����Of�d�O�����0P�)!\�`�fV�`=�Ɂç�$�M{���?I�/�4h�Ӗx�O��'��3K(����hT4Ʋas�}�<�$�O˓?��3?q��?�ݴI	�� 5m�u�~s��7M�O��JP.o�i>���Ɵ��'Ќ�gA��3>����qe�x��v�(��?qJ>���?y*O��gh�a]D�0�3>��	a��*B�6-$����ßd��Cy��'���,+(y�rh@� ��D��c�8 ��f�'}�'\2�'|�W�ء*�O��đ��]�.������ )Rf%��Ot�$�O��<�����O�H*����B<�����r*�SE�UG}�'��]���	�.Z̵�O��狉! ��f[2�HX1p��,�:7-,�I����'
���O<����j���a�E�M���F����	Ry��'�E�\>���ܟ(�s�������p���a'VL�/���OLʓa��GxZw9�h�"�m����&#ҏ	}DlB�O���#*����O ʓ�(O�n܈xyt1���Ri��J�8ED��' ��/�8"<%>Y��J/x��0�aɇN�vu��eӺ�V��O��D�O:�$�S��J�|��<3��X&�I#W���h�p�A��=Ex����'��Q���88���P��Q(��d�����O"���'Vj�$��ϟ��I>Jllc���,�r�pÉ��wA����4�?y����d�m��'2�'N���I��qұX�|ڣ�۴C,�6�Of�z�٦-���������"��J��*z[}�JZ&|P�p��Z�>>��>�x}̓�?����?9��?�)���SA��	��1��ڰ{r$��p.!{ �lӟ��	Ɵ��	���ɻ<���+_��{$��?H�h���j��9��V��c~�'J��'�Y>����Ms$��njzX�2��q���A�F*�?Y���?��?9���d�O���?�k�C$C=nX�p���;�6�jG�����4�?1���?���?)�pJh���i���'�+���M/�4�oI�f2n���3�M;���?�������O�p�.�ɪ
L�y�-n� �iBh��U�Z6-�O����O
����aH�o���I�D��tr�L��&֭z�-Q ���B��9a�4�?A*O�䉹c�)�O��D�|n�zf�L��-�3!��(0��Y�~6��O��է-
��m�䟰����P���?M�I&!wB� "��Q{�["!̂5x�Ρ>����9��G��IOy�O��'T�VQ��*�"hµA��� �*�lZ��D�ܴ�?���?��������?��HT(�z���1*�!pdL[/H�ʍI��i0,l�W�'�"Y��SU�����b6N"}y�[���I@�!���	�M#��?Y�Z����v�i���'�R�'�Zw5����@N�a����U,*e:ش�?!(O��`f>O�������t�@��8<����|3��"���������4ZhTa�4�?����?��"L��y?�v�ҏ�|�"k�%`�l��R�F����	��6�����I�t�	֟��I͟ ��'q@�4�"��>Ex��ԙ��
�4�?i��?1�Z���|yr�'G��i�!��h�$݋£M!-��Q���C
�y��'=��'��'��S�t�pH�ش�hD�P)T�}T�#!�ɼo�))��i�"�'E��'��Q����w�&擇J����,H;R�|V�(&����>���?��?	��<�f�`�i)b�'���cTOZ\���9r�ʞ9�L���~�(���O��$�<��e�:�̧�?i�'��u�B͒��D��ß԰��޴�?��?����u�#�i��'xB�O����o��-�~���j�0�Ӧmx���$�<Q��P���'���|n!�l��%�ƴZz��)u��;Z��7��O������&9l���	������?���ۀ V��UOP	� ��E (<�"\���	�*0f�'��i>�ӺSl�+t�(B�SC��bh���H�c�M����?�������?���?Ed۠fLnpʃ��)�� �pi�Q̛����bx�'�i>�%?m��!&�J�i�%��� O�<zV !�4�?����?1pB	\g���'�b�'g���uW�ē$����l��m2(\��yu7��O�ʓv����S���'�B�'N��
��"OD��#oZ�F$�I+�$u�n�:F�@oZɟ����D�I���>yԭ�9&e[e��<JŲ��>"H�<����?!���?)����)�<mZ�l��Iˀ~p��
��P�sؤ��Ue�m���<���L¬����?A���O�P�I@��N�Ȥ��!S�*аϓ�?���?	��?(��܈g����y��jۥir�iT�R�ACd�������M��?���?���$�O��<�:MӐ��"���PҎǞ=��S'����Iݟ$�I⟠ۭ��}!�ަm�	���a�n�c��I�HE)@y��HY�M����?a�����Of��4���':8��A9(���1�RO���rش�?���?��
!kܦ��	����	�?ً���G�Br�?����CD�)�M����d�O��x�<���$�<��5��ʪ2U$�'�Y�C.�x���k�`���O�K�Hܦ��	Οp���?)��˟8�©F�X}~�I�o�g5j�t����O�)E	�O�ʓ��	'�t
����c��	,Z$((�(�Mk���O���'�'���O���'9��E� Q��,E�(��E�_��6M��wf>���O^��|�H~B��v� ���Eb����ՓQ�ݡ�i+R�'��P9<��7M�O����O|���O뮊�T{6zG�Ӏn��M�E�[��'�r�'�������O���OP���`�06���u�ԭ[��Q�ভ�Ɋ �0t�ݴ�?���?Q��&��SB?y5C�5"B�<����(>:�Z�E g}�-��y�' 2�'��'q�'N�}8F�nU�q���$�pT	U)�D�b6��O>�D�O��$QL�V����mL܌�FT-�<�����"~���ѡh�P����������IU�E�a�`6ML�#�l�H���[��U����u�0m��	�x�I���'�2ș����4B<���a��1ǆј���Vi*�lZџ<������	���)�*0�V�l��|�ɓ]����炮.4��0�܌f�v��ٴ�?Q���?a.O��� *<.�)�OF�ɯ/�"�I2W��,����FAa�b��Or���Or�����I쟔�I�?xf
G��$���IC'1����e���M����$�O:k�7�8��<��eR��[Ԥ�cQ���'�p��!c�h���O,������	ϟt�	�?=�S̟(��g��\C.����ep�uy�����$�Oքz��O����<�'���!c��i��u��Wf�Z�&6-����o�ן��	���S�?y���d�	�A���n�`�s@ݦ�
�ߴ(T��������}����'"��xӇ�ю�H�C�9�2��qӬ�D�Oj�D�T�1n�՟���ϟl�I���p��-�T
B��	#�L2G�0���_	��i>Y�	����	�~�X�1c��$�v��F��ck�Z�4�?�t&Jכ��'q��'�B�~r�'��uQ��G�ql�٢͎+/z�$��O�I!5OX�d�O��$�O����O�$Y�(;��A�,�5�\3h|�A#S����I��D�I՟$
����?���Q?MXщƇ�^H@��&��"I�d�<��?)��?���"o�҃�i/�\�ת�5trBu�r�̷A]�a*Ӱ��O����OB��<���I�9ͧQu|P�.��JYh�4�ͺA�VE!fQ����ퟸ�I��I ;n���4�?i��q�d[�&H�i���U�L���9v�i
2�'�"]�,�	�[J�����ap��2Ȫ�p��hl��X�	uyR��#6�&�$ꟶa P���a$��*I��b�K�>1$�(�I֟0[�D�\�S��(Vh�f���D�c�N���_>�M�(O"�1�����=���V������'u0E�V�K�u���+V(�����4�?a��I�Fq���S�' @D��(Q!�޸c�f��$&�oZ$UE�4�?Q��?)��Ta�'�B"� �x��7ゖ��t�wǀc��7��e�d�D5�����5�^�My��8��'L��M���?y��(YH���x��'02�O��XR[YP̈�FT4iW�]��iI�'��Þ����Op���O���$�.�ы�I�/I���i�AC֦5�I�'�(	�M<A��?�J>��]jmz7$ЂOJ�Q��剃l3H��'�.���'K�I⟨�I��(�'8@{a�7%������g��O���  F�쟘�I~��쟜���v)��l�D���:b�ȐI��(:qCx���'FB�'�V��C	���ĤغH">�X2�E ���b�V����O@��5�$�OB�$U�0���	�-d|cV���>F�
���.�4��?I��?�/O�9���H��#V�ҥ�̇{�F�)��Ъi��q�4�?qH>����?q��L�?IM�8����w��śE� 	���5�kӢ���O��A�Pt�Ğ���'V���
B��%BM���IS�2�O����O0��8ON�Of��yv��d��:�4]�1�Èc�6�<��$������~��
瑟����	V,�;N�}Vf����eӺ���Ort�E��O��O��D%xe�Im�h��H�,V��6�i팠�`�c�z��O��$���u$�x�	*Km|�����0c�8��󅃾�9��4 #�����	�O���ujK.R��|S�.Z#�葤��覙�Iߟ\��U�*�M<���?q燎 �D0���s+ ��!��u Ԑ��i�'9H ���I�O���O � U#8F�,;�:2��Ö�Lݦ��������I<I���?�K>��j��UhWnF84�d`T�d�^��'�8ِ��'��	��t����'���yjɻ,x�E����	i��Kq�G`Y�O~���O��O|���Obգ��ʞ5p�]Hpd׶Z��|K�▊XL���<)���?�����Ě9G"���'TEAX�ʅ#+H b�������')R�'�'(B�';��J�'� �	��<D����Y$& (e�E��>���?�������o֪-'>�!�&B��S��@8j���,P��M�����?���D��!�{�#���Z����Z��q ��Ε�Ms��?�,O���1��K�Sǟ��s�)zƈ�-pqR%n	�\�v�RS�#��jyB�'lQ>Y��N��<�b�sDC�CP�A˱�a���[�$ꧼi���?��
��	�2|j�!R3@��4C��Q(:O���D�O�ᓽ$D�ST!�;�j]�ÏQ�Z6�6-_+P���d�O�˓����?�/O �p��e�` 8���6�����|}����O1����~ġ(�Ē4�H)�QR�ƈo���\����'&����|"��?��⛉]������Q�Ҡ�Ǳc��Oք����O~�D�Ot!�'H��Хǂ�i�2�Ck��'t��S�x1��*��%�d�)����FK[#���Bs�B�i�'�0*r	9?����?)���?q��)��e��Z-���s �`�F���m�5|����'���'~��~B+O���U�7U��G�^%�����V�)澱�2O��$�O�D�O��'�?a�iG�F1�hh�&�΂h��,���֣f�\7-�O����O��$�O���?IbM�|F��a�8����ՠE�7+��6�'���'�rŲ~Z��y�V�'_���[�$�y�R�#4Yy��ҨK@�7-�O��D�O���?!�d�|���~B�=f0pM`5jH�-��AXD���M����?a���?�ֈ�ϛ&�'���'-�D������f�@��}rׅ�P;�7��O2��?��̙��ģ<��ŊCJ�/VT�e�]2�޴�0*y�J���O`	

ۦ%���|�	�?���lQ�@Ք1P��{VV>w���%����O���T��O��D�<�'���-]�$t��P$��Q�b�ْ$�iGzԺ�pӶ���O��d����I�O����O�I(6�X�I��Cɔ�D̲ �����Y�d+�����Vy�O��O���	NN�!�
W�?�� ��R=q�6M�OL��O~Y�Ԏ�O撟������phW�z��voCwHT��Ǣ��O�i%>��	ß��	�]�zhhR�p�����D� �h�4�?��պ#��'"�'Wɧ5vE$+ $�t鄴�h5X�����O����O����<�Qjݷѥ�	s~DX�����vSd�b���ē�?i�����?a�']l@Y�:h�Z���I��i�@EH�}2�'T��'�剰z�^�S�O{.e�k��M7މ�A�Z#k1��S�O�d�O:�O �D�OH��0T�@�K�x�ض-��C�Șrj�>���?�-O~��  'Բ�'�?���[.6����S×�^L�csĐ�:D���'b�'t�P�9��!�D�#fZ�%� .C��q2#҂0�f�'!rX�p�� ���'�?��'nZ��g �:_؅�&+řU�:eHg�x��'��z2�J�&��r�T��W���M�.O����������D�p��'���q���E�dӱLY����4�?�
�$�=��_�`��x�� ��j�pxn���^uQ�4�?���?���R��'9��%Ob�X5�"��XV�^�?��6̈́�I��"|��1]x��Y��t�ڀ�<<�F�a�i��'B=T�O4���O��	��@A�$��X�h����3s�c�<Y��,���\�	ӟ4@3)�:0zQ�u =��H��;�MK����By��~J���u`�:K�VN�%cK�dт��$�xҥ)��d�Oh�D�O�˓	jl�c�b�d�R��JG�]� h p��<b,�	ݟ��	����Ir�r,�\��� H���>^�{��i��'1R�'���'�Bl�u�	�(�z\!4Jƶ1aX`)����VU��Iu�I��'� \�ݴS��,Q�G�5..P5y�ʙ ���'R�'�R�'Jbj֎����$Y��%e�xzBf��&�p�4�R!�M�����?�/O��w�x⥑�!�8��c\-RQ����M����?�)O`q�!HP�S՟����!�pY�#h	�!ܐ�B�5X1ܴ͒��'�,-"���i(]�7��G	�Yb��  ^
���4�?����:\���?����?��'����1SC*؝]��d�5W�T��x��ik�[�X���8�S��S�4z��.h�B}���%��7�u�x���O����O��ɥ<�/�z-�aD�1�����/��*��Kz}baH"�O1���L�-���鑋�8=ń�RBW,'��Mo�̟4���ؒ���|r��?�a�R!XiT�:%i�0�ޠz��jɱO��2��O
���Ob��C��S��!��Y'4����s}rĘC�r�'��4'�0�KV�tK QH������IK��ēZ����'��'�"R�y��#}sf��Ud>y�`ે(��O|���O<���?1K>����?i%� p�e���aX�C,{�- �W^��?	��?y(O��D���|r�Ԯ"��A���#u�0�ۖ��C}"�'���|2�'��R ��$W�R��@Xg�ݖ��j�$V�A������I��' !�r�/�ɔ/yY�����0=[:ٙ�a���|oZ�t&� �	៰م�!��8J&��5B��)[��#1oю&|�7�O��D�<Ư�&gm�O���O6���R��r'p* Jͬ7�Nm�&�&�$�O��B�5h��'C�Ќ� �e��y#K_���Pi�*�z��@ʥg
:����́L�ӈ;��OFP��g_�<뺈�$߯�b`��"OXC��!S_��2�����ҵ�D��X��D\�"G���L,Wf�K�c��Ay�uʳ��k��t4�C�/(��F��5bd�N�/�J<�T�@��T&L��42,�&Z�� ��>X2��E�H94�0�4�H�`��V�C�1�85�A�b���zփφW�T� O��a�T��T��O����O�������?W��:@��U�'"�0@����iL��	3T�:	����.t���j	Ǔz�5A�b�;<���d&ã(�:���1� }8��839��`��'��z�������0��ęl߈T�⇔�?b�';�����O0ʓ6_�)���UPX�	!�Y�x�&чȓP 4�բ�J�h`��V~4���	.��<�P�O�Q��?vR~L[w脢~��µbƣu����O����On�9� �O ��g>�ۖˀu(`b&��5G�<�R���	��4̍�Q�*���	.�xK^� R���۶Z�����Tx�̳#/3F��`Iu+7'.��i���<�8���遍n��'�>�����?����(G��9 ��H�R���ā��?!��s�<���+K*$�3g�~�,9��'�ў��u E$<�N��
Y	8`q3��r����4�?)*O��� ��A���'���(Q"����\�7)j5�C�Y���׀S���I۟�n_0Ocx���)E��@#�A�4J���J̋�C5Y MIG���(O��٠����L�@�O�mt�MAD	�:���r�]Xc���J��MQk��fo��Q�F4��L�fO��'4���B���u t�����,��!�>O��$\�3���r$�8X�p����|��g���t�(�A]��fg˵-�N<I�$��Qg�R|~�\m�ɟ �IO�t�΁p6��'m�A�3Shl�)Cf���Z�m�z䅒 ��1��T!�i�4���T>A�|�ɗ<;���*P= �IG� ��}IAEҋ}�Bi���	Dxx9�S��?�P+�L���k�	�1�tQ��������?��O�O`�'�Â�� \+@��0=)n���'��ٸ��H+FJ��;`ŕa�lU"��dBR���i�=v�x�C$��`�iԬЭ'�4���O�5{#�K�h�*�d�O|���Obԯ;�?�F���m�$Jh-��~nZ���'�H�[SBۺ9�n9�� PF{���{
��Oޛ|��t�3��./d��0;�:�6@/\���hO�D��@%?}�=c�I�&(�A�2�O$���' 2�	|yb,�� �2TG�E0�!��y�A� 7Ҿ��䙲S�=�"�!}�"=�OV��9~Ίq�ߴY@1���e����P�Q���?i���?Q�œ�?i������ #��� �!�?t��,9A.Ռ��[�f���h�É�0=Y�̋]c��:E�J�*z�)r��ˢ0��8��Qewq�QA��� ����O|��W
;z<���!��~�D�y%���a�!�d�22Ꙃ���-oᶡHt�F�e�!��K���*3�L�c�[�$"��t�5��9�#]����|�$e�\t}��+��P'8\��H\�Vf�#�'�r�'�bIx�� >���٧gg���%��*8���+�������<�v�	���/��<�����!��d�9��i!h�5,�Τ�Yw�p��O@(J�8T�$K��?�b���֑�r`�.x�~b����`l�,�2��/S�ri4���<�����>�G�%Lr��+b0@	�H !
�v���O<r�Ȧ��Hu�ɣ�x�S��<!ׅ�Uu���'["V>�B���t��ȟ�@��"z6Ll�RG#c���Zr*\%#�ڜ�$�j�S�����Z'���I�V�锃�8."�}��Ĝ�a��c�"~��)/��T\�ey�9�r'�P	:��R���d����Ih��?顣�3{��4���2*�T�.��<����>YqFU�.��d���6l��O�}�'�"=QЯ��t�0.�Hl��M�#l���'˟��I�(��AXV�[ݟ��	ٟ��	��u��'i� �5<��|�NQ�#��p�����~���
��>�+Ҡt?4�1��48Q���N?��Tx��s��ʇK=�p۶���;yR�{&���,��#��x��4=����$�O��g�|3�E��F����`ψ ܶ̅ȓI�p��"fȪ.mN�@E�LH��`��	i�D]�������M+���((�n�arcͅF8|����>�?���?��LJ��#��?A�Ok�l�g5u.L�;ƪ<�NEPSZ?wopT wL:Wޠ�yAjY_8���r��*;Ȃ�c� vQ١��9�~�����K44D�L�	/ʖ%��'�(���!'���@�r�&�X���+r������a�6M<�I?�H��i��ıFL�4Z�z�"�%۽,K!��*QiJ�I�l�?x������"�DKb}�Q�4��  ����O\ʧT��k��${���A��B�!&�h� W��?���?�R�Eaf�E{�5J�2d�S�dB�̪��!�\�$�,�yҗ�(O�����fP��B��O]�\�o�]j���A���od(��F�\��t�Ll�~�WT8Bu�c�EZ�d��,�<�����>��n\��D�R�5x�BD,�v�TBO<Q�LX�n]���� ��r��<As�\O��F�'"P>X�H˟���П8c�H���8�B ȋv�Fq����zf<��l�$8�jT�/<L�O�1�ߥWX��4"V�!��Ib�~�Ӧ#̊YLΑiS��}@�9�ʑ�W*��%P	'`����嘀e˜]��$(�� �`@�2eW	Y���Iǟ��I��D���䨵�B��q�6u�é>G���Γ�?���<����`��֣M�
_`�<��u����Sʟ���i2�>T@����H��k3��ܟX��8ݔ�3�(\��	ן��	�u��'n��Z��4hƭ�@��E �
'@�$[�x�\��
@	mv�e���hO�
sB��'r�1:TB�W\��������1!����n�$�z��hO�ԃ2Ò�2���s�%G�Yњu����O� ���O�l������꟬��ϟ�iޅ��̌@�n�{0�IYX<�<D�9g)ǀ{kX��,Nl"P�/�HO���'c�I~ʄ1�4�h)p0N-\T�5i��N�p0�]��?����?iɖ��?������$Cr������mM��3�5f�\� �Q��  ��b��yo\60�����d	zS&a0Pb |����u��(~D�$�_4B��@MFa���LаEJ�l��b4��=0
�r-�H�'!џL�SA��]��uYs'0/�uO3D�xؠJL�R1%ppj@�6{���.e��ӪO�ʓa[��8��i2�'�哳t)xXRD�6oT�<R�B!U�(�V$��\������ K$��{TB�T;V,�S�T(ۉt��(27ٞu�Ģ/� �(O��9�*��C��3��L��O��ѐ%)L$@pJV�_2���d�*���r�Xl� �O�R)�a�(���怕8X��z�'Z�O?�I�M/ڄ�Bеu�n:��C1���DF�	%ttC�j�d����8Z,b�-��8�޴�?���i��w�^���O��D5]Yt�����H�s�b�]ĄYB�c[2E��Q�.H<!��V,j8�M��%3���`qH`I�;8U+vFǲ�j�*&��=��y��Y.R�,+��̵Wǌ�9s�L*Uq�EӮ��<ꇉ��w�R@staN�^Q2�
��'h7��Hy������E?u�0�y3i��k7J�g	�y��'��}B��$N����%��x�H���o�O
�Ez"]>A�#&�6C\I�T�[�x�$�V�T�I�>��1�r��p��˟��	�ug�'��bZ�:� �3K�s*�� �zl} �H 7o�$J5$76��@0�O��=���q�|j��#£�a2*%���W�l�0!S��$�d�&#ӱE�E���z�#Ϫ-�Rc����9k��A���-m���d��T�e��O�o����?����d_E�M�X )�b,�V
�!� ��ZH� �QFb��Xrnŧ8��MGzU>!�'@`�J%�e�&T��i�;:���D�ծ��u��O���O��dZ7m���O@�$�B�җ����4E S@ҖZ^�����`��(y�El����T�>�x���=�X����;).)#ʖ�X�fk̭*� �����d�O�pm	D ^���T� t2s��O"�$�<q�����I7�(i���Ӂ**��]8fI!�S�4��ᮉ�Z�Ƭ�FT!1��_}Q�̸ώ��Ms��?�/�=b��4`�@��C����Q�TQ ���OX��͝*��5�1�͔����JƟʧ>�h *3�H?m���B�D��a��Gy"@��((S@�H�_�a3ђ�d픑N$�E1��'N����wIE��(OP�� �'@R�'�2Y>-i���I"��+�L,X������֟p�?E��'T��;q�P�X���6�;f��u��N��'h��
@H�#^<�d_�Z�t�Z�'��E1��cӎ�d�OD�'a�<4c��?A�_ޖ�䅐2 ��-bף��Ts�臬}:¹
c��:LU`����`��SP���}���S�h*�r���t�`B#Eއg(�%�� ^'d�i	DOX� >�q���w� �J;%16�s�l��Z���J��	��(s��d�����'��q��,!ru0Eo�Q2N(!�'���'~j���� �Fܻ��O0���ˎ� K�'�哏	��B75ROt����@P��Ɠ6��y9ł�Ѕ�B#�5`F�Ćȓwp� ��5F!r��K�z��t��S�? h4�W�.}����ڹH����"O���V`Q���͛�e ����3u"Or��!�Ne��eHW#��|"����"O)���U%T ��қ)�P�"Of�������قcڥo�dis�'�R4{�C�6!\rt��r�0,�
�'� �x�Ϟ�d����P�nF:�a
�'c�E1a�|j�K���f���'�2��ve���"P�+TvG�l��'��t��1GyV�JS���h �C�'��ڡN܇}o��Q2
R�]�tr�'x�M:�� T���
Ճ�1���8�'����&�z,���1}B,z�'����h=l�1�P$�\��'',�I �@&!�"��$��L��P�'��mB 	��$�p�iA����'?��ȁȞ9��I��j�*0Ͳ\��'餉��%M{�^%��-�4(~��Q�'D�ar`�-7��������'j%�2j[�)l��j��;���
�'���pb�$ ����n�*y�y
�'N�P9#�*��L��d��D�
�'!�+�/� ) ��������*�'K
-8���+������rG.�#�'cƹY���H�ZI���G1raF@��';H�G`S�0�hB���"��{B�ê�O�O�p�w�9(b�!�R�f�T��'��(W��Tht�듮� {�: ��"�`�� EF��O>\��a\�{#���U�"O�5 E+O>����e�	�]���S��H#4�5��]�V��ر��ekax�K�E$*(لM
�U�� 3s蚝�0=�"�
:���;p�^�h�B,@��N�\v��R͛��)���:h���	����%�M>�$x� ��8Ab�%�x���Q�b��Ë*2���eB2}�O��pui]�G�:uxD���7����'k�=����ӽ>�(�p�G�9�܀�A�v�����-��8�G���S�I�m��;r�%���X9tTâ�Y�^Vl��'�b��M@Qx�4H��u�r2��uQ�b)��I9Mj�9r�B&f`� ��B.& �H��#t���5"�諣G�ZX�%I}*t,9��'J(W�*l���Q�k١~�Du�S�U$m �-���g��q�p�/�ZD�j˂x�x�S�T(�I�i�&b��Ӟ"�,����Dr��5��ɟ�D%8��Ĉ]�p�s�l_1Nؖ�=Ѷ��fV⹑�$�?�T+I\�<a�%�}F���I���в��(&�⸓�ܟ���X��A4c���pD/QSص�tA��Z�$@��I�oڑh��CjΌ'�0����'���"%A~$��zFC�Y�:">�����v'\�RF���c�ɤn\�iZ��Yw�'	JGz2 .D�RQ�J�%:MPW`]9��O��� L
jc\H ��T�Ij
�)�<O���&�E
f�҅g�#w��fQ�(���|���� �K���
G%[�<v��dm�-@4P��&�ױ�y�kG9V6� @	/�x�G-K���Ov�Q&�2�؍��o�P�d�p��d�zd�r�fG�_��-�U��8_|1O���qǝ�}�����Ȟ�����ة�?����HO� ���,C͠���8 �r)�!2{���0��(:^��d '�e��李J���"�޳���Sv#�)���	v�����vQ�H �jɅ3�L{TD7m�݆���#7�D��(��Xl�]�\
�4�!I<��'��OЄˡ�L���� �>U����Ʈ.<��*�/�B����U6�q�U�F)u�0y�� <M�&�Gw�8IC�Q�5������͸'��iiuo��r�13�Y:��kI>Q���7��P(��ؚx5�<�SM}��R�/F�ũ��mj��D���HOڴ����3.��*�, }��X�b�]�Jx�=��� �bMB�#8<OP��/&SV�@K�9l��aE<0�`0�h�aX�� &�{�6�+,K�Zt33g��A�Y��y���C�D8��U�">��AhE<_p�$�����EM?!�*�x�8�S�ɰLL�1x \6=���	��O�d`�ѓH�(�.O�0oڨH2�@ꕫ��B��C2c_D�O�@�'"FD�UB���)��'u����'�t����8Z�D@#G��H����O��#

x��D�)O&�8[��#�*������(�(�L�2t�|�1��'�x(�d�R�H�)A��W:c�*����  ����7w��Gد%�2�B�W�<AH>i��s�f$�G�=�F����7"��� G�{� �Gb4<O���O���SB-B�1;�y�W�]�du�M�`��eT"�/O��#2-�R�iOw갉�S�I��)'�@)g�Ek���1.C�(J剑V��p��CԘL]�)S&j�)j���S�3���
S**��PFL?)��9���p�|٣�Z��*J~BvJ	m|�or T�0HWT�V���L�r�H�y��l�����$��ħU�b,(�t<�pE�.��I�f�ʸA`u�pC�8���j$A��*֮��	F�H��LF"����uc��\�b4b4A4���D���+r�]7V]�d*B+V3�-	���bw�ta��]�f<r�OX��˺���� ЀA򇄕�X�-��o}�'߾��d,��x�f�5<#�Xx޴Bk�<��:Px�\�	הqhQi�٣p:؁A��7;pL[C���~J|ZG����p��O�Hq�e:#��Q�~h����>��&�9Yv ���K˜'�z9��/^D�'�����.*L���z6� I�PpY�L�xd��`#�#+(�p�EI䀋��đ�+6h��bX��$����x�vi�&z���Gz���v�'f�6�Ɛ3�dm4�S�V�ҝ��iF�*3j;W�'����&c��$*Ǵ!Zƹ�˕�Kרb��Zc˔_�S�p��!f�����C/M���X�.�1V���j3�$�(�zh R/ע7���@�NG��fao�[ю��򨁘U�`�A�'[�~��>��Ho�[�F8��d��%��"V�ؾ�S�Ǝ9Fv���>��e�*�v�3�kW$7 ��h#]c�'f�Qx�1T�n��t�@�YF�}x�'��8pc�k�*�0���#sN(���d�8+RT�t�\+�@�s%�F�l�ր��*U��ȴ��IZ݂٘�LD�|������ e4�D��%��iHD��	��S�䄈^8�:�-�~�P���O��Ԁ@ŗg�D%sD��)����d�Y�.T�׮(O�M#aL�{M�t�v�H�6Œ8�A�i�R`�#�3DL�`i�G�r�qO�5���HxL��
��X� `�|c[�]��|� B N3��I�����D�@fK��ϱW�`mɳ��O���C�������du�p�1p�ę{��ΪA9X��CDFȰ<����5*V��@�1<j�U"�
9X�\�f��T��_*�<)2Fڍ\����-��P�����wo������7��-B!�[	�?�$H�����I�#PI�R�ęon��[�BQ�C|P!���|AF�r�F#O���b(A��	6"�;v��,j�@�p����l�fe����	*w1�ɷF��0*��i���pK�0p����`�4�X�K�p�`�Ɨ$B�zi ��(�"r�0?�� P�P�A��N�����LX�<7l	:�.���D-Tè�����*`�4��#nيg���B1�Z�*� 2GS�}b��z��)O�d��h��$�.1z�K�'���s�X�8YI���W��dѺ7
e��d��D�)r�͢8���T��Jy\�Y�7�����wxT��Gı-�\kA�$3����w�O�=�ڠύ�6D�)��&�1���^���+�h�%s�na@�,"��$���MK���r2&Y�z��>q�)چWʶ 2w�u�VD��#�'�lz�h2W�*!�f]4H��}̧7
61q� ��5��Ir�!�,�����Ǐ.]5�'��L�+�?:j)�O�)^._r���l��RK"&�>�*�*P�
����fIᦅ�#�I��:uCw�Q1�-+�L<���}���fV��WkۈF�r�Ӵ�,}�ƖQ�H�%m��kub4r��Ԋ�򉞤)n.ek���w�܍J�&��:(*�r�N�bw��;���J���n�7l�T�5C@�An�苣a/`�yA�G'9����ꕎx�6�P�Od�t��KQ�����'i����N% BᏟH�]!p�������?{��Ƙ|��%-̤ZƬ�.Bޙ#�.�:vM��R��D�E�*�#��+F���#Wkݵ3�f �s�{a�@�,k��ݣ{7~LA��$��iqd�ݤ~�xO@X�f���}��zt�֯i���&'�Ll��ޓ��1J$`F�%_V���(6֐�%!�`
v��mU*)plQ��k;�21I"hV��HOX`��D�"-q��j冕{�@�'��B'�2�?��fQ�sG�Yc��	<$1�6-O��-kwڟ`y���yU�%�BcNPzU��ײ3�Z���MJ@��{3�M!i�ށ�� ��&�����mK�1+L4Ӵ�
(Dbhi�I_���Lc��GB�[Q�i�6�O�h�rJ�L;�!�G$oDڝ $�?<O� ��O+�ʼB ��6lw���`��1���f���bM�=��L� ���eN~�k�(�*s�A��T?1v�N�F)p�k��e@ɀNU&D�cK;R�� QF3�d״2,,����{ )ԡڤh�vm�'_�Ji�Ƙ�,��={�F�)�D���`	5X����͓W�h�DęL��q�q�'��XR��1���yҨ�6cK,�$`�a�����gJls6�Î
��[T�x�d����/��P���MM<u)b(_�yy�C�	�^��L��%��i�1�`�;\���FH�+B�ٴ�x"�`��i�l�{�c���yb_!|K�]Z�虤vS�%9$"P�Say�L�e�aI�HE� ���)�gY�d|6�84�H!#�N�;R�����'�\����5/|�#qcP�,?b$��'��9YƉ'�����}~���PnۈT��K<Aө͔U�6����C�p�y@��_4��l�j���~��[Gsj��C�ń+Yvp��L��>���s0��	x�\M��m��0=��E;�{E��.. .,٠o��9XX��������	�����O{���g���_���H�,�/�����m����Ì��5��10p��t�sV��
?D(�?����9x�Tq���I�'��� �m��E�=}$��؇-&v�`���'�J̃�:�\�ed��nf Yr5�v	"�'�!2fAI�{� �A3�%1���1m��I�O��Ilp� OF$f07�ɷeT�EzBo�v�tT�#+C��������d٦dݠ��eZ�Z���.�lH�-^ۦTk�-Z�n`r�󄄛9b�)V�W�~\�P
�J�a��6O��aEJ��ԇ3
�\��$)��O�d'l�t�YPb��=��Y�B*>4��XR����e�[^�Z�G_ax-��IY���Oz���`�|zZ	��w�Ƅ����=F��<)g��}A�]�'�p�"KR�z�A�2��z��`��-�I�7��U����0Rԡ��9�l�Oly��M �q`ܥ00.��F�R��'�ƀs��pYq�@@�8�����M���k�h�|�+7$ �l0!��j�((|�)3,(@
m�ub���4N�`�@e��_}�,P�'A����%ڟtzX��FV�h@���X�%y��� �<"�Μ(6�K*	��[�'ll99�E�OP~d��8R t��Ά�3a^�� �W��hOB u�4H]�� n��\�R��{5(��.�8rVC�	 ..�ժ$����ai�-�� ��#$�	9~��QA p�6X����&]��'%����S�E{D�H4�J�c�.�	��,�'�U�	��r��RA@��u#DRD�0ĕ�E�n9����B�5(U$K�\�Y�冓Pi��$�w�HH���Qjȁpg�Z |��Ƀ~�ԑ��ؕ@xԄ��F)i�"<1�
&Z��� S��w�`Q*�d#�C��2i"$@SW�'!o�H��ʚ9u�-�"J50y�ΛD����-y���ݥTx"�#FB�<�<T�����B�	
%����b���P�Dј�$���R���OIJ�I�	�� ��gn>��f���D�&��`�c��I薐��K��\�(�g�(�O�rH�k�J�ⵥ� Q�X��'Z4o�ֽ��H�ZFJц�%��D�b`�	t0��	�C"��(��Ĵg����[�9�"<i6*W0lD��UJ�)ON�y͟ן$��@�)��8ak�#WNμSP�7J����6O���,P��Lh�C9$w�!p�!0^� �Bܤ&`8�Av�"A����%�m$>�:PZ9�k��L��}��bK(B�C䉖v�"xK�*�	�0H��Z�on hk�&�O���
�0ͬ���p>yI�"	�_��1JK<Y�&�w��K�H�2_J����&�u��P�L�wQ��Q���1*����M��U����U�d�����{ZY�AˎFH�z	˓n����@1f,�it�`�DxbKW���J��ǡ"L*Y`���3�?1��ޯp��ɒ1�	S �I��a�-v�%r�D<$�,�"��#eL�,�J�&�uq4��"j"�<P��܂p�eif&K7�-�&��!��ZM~���l�U�@�8It�!�F�5��C䉳g.�0O׆+�����ɯ��	_
d���ӀG�e3 ������nțS��B�I�(�����nα#�E�:�B�	�y$V�G��;Ȧ�r2$7*bB�I�o{�{T(�`��	�!%P_�`B��
[�0�[q�NKt�\@D͐!Z(B�������$�@��%x���"O6�z!c��UJ����Ti�i1"OB\PS��IMx!�1��ZZrm!�"Op�q�B�ƽ#rjYVTΕ�"O���"�`~��R��:ڠ�F"O0�z�_�{�z�J�6 �3�"O��X@KD�{b��d�$�!I�"O��#獀dp��χs.�Xҳ"OF �l�'+��"�"OV���jO�U]��*�oN�9R)�"O����%6J��t� ��I��"O� J/}��2/\'EY�"O�P�ۼ|�u1���=Y&a�e"O\���IY%�"�RS��c�Pq�"OX��CE��7�,;h �i�D���"O m`�G��n��H blD��x@ �"O�5(gΖ0|���⊔
#'��R�"O�C �;<��Ѓ�&Ұ�$"Op ��O��16�%���T%]��q@d"OD,�姖8h�h��T
�"}e�� "OK�s^���L�F��a��EV��y�.�W�1��P���S�!U��y
� ��ఎ�"< ��
N�]����5"O"	P0��@xEJ�Ր&���K�"Oj�Q�3��	s�N�=(����"O�����Es���+x%n�a�"O�zv޻E ����v9�� T"OD��K�*x��IE��hX	�"O|yz�'ȆF	΀�d�R-�p�!�"O8i2%O�X���P��`h�`*4"O��P��$)Vz� `�GTb5�Q"O��9�ɚ6x���ԅ��[o����"O`��@h��г�E��i|y��"O�Qx��ȴS����@R2�(S"O.�I\����S##Y�@�2Q�"O2!`�͚���֢ 12�HC�"O �" n�6N���B��\L:�"Ol�b2�÷�P`��H�
�
Y!t"OT��S!�tY���s���"O��2	�E��H���#!��i�"O��@E ض,�ӂG�P��"O��+0��;l�(󗆑�MB�C"Of(�m�x��|��f	�mX�cp"OȀ�@��"�(�@��ŉy�
�
C"O��1ʆh��Ik�?<����e"O�KG�R �h�r�
&jf��"O$�RĊZ�xo&��i�$ef��"O@�:�ċdO�AP�(D�/��MXP"O�A��}�@12�HE�\�"O��  X�̈@���=py�"O�Z�'�o�ժ�
�.�v�(�"O04x����z�(\%2LΜ{�"Ol(!"��8t.:§Q �¦"O�0���SL��)1f�h�����"O�;FD�y4>��3%J+��}B�"O��F�-���ǆ�p��"O���
6a$%���Ā���pc"Or����?�X�iR�7<T(%"O<$���݋@;`1� ��My^�;�"O��r��X)u�F)t�0\,�W"O��cb��i��8��*�M��Ԉ"O�iqf�,{pQ�� �x	��"OX�!�	�����O [� �"O�a�a,�{W�Q�O	+H����""O&1�rEȃ:�̱3���:X���"O2����.y��iէ�-9�`�U"Oع%��)o�ꍪv��$���aU"O*���NC��d�A�5V����'z1O��"L��h��܊��K���a"OvQ+1��c5�9	'���n��
 �'����)�|r˝�=���p�D+U~�`��͒�y"oԗ'G�q
O18vL�:�.�yD�.x�"8��D�3y�0��ʜ�yblY�sc�tP%��L�X���,�y��4�~�!
���ҥ�V9�y�䑕>�RLA6�P�LC�(��O��y�K�(U��[q�X�E�8���F���y�ʯT�P%�Ӯ�<�,ْ�T��yү"o}��K���5ݖ�� �ylĭpt��­+�\E�ؗ�yiXY�1�t-�!�nQ5�J��y��K�I�t��fGHA@Uk���$��'�ў�O梉�3�ܳ/l��S�o�v�����x�bͮ^[��!�ʃ�H�v$��N��yR.F&vЬ`�-�N��	sU)0�y"a�
(��ܻ��іB5x�jpn"O� vp���D�#nj92'�Q$ 3���U"O�@9V"�M)��
�E�i��,��"O�,3B�X��y�e�	�x����3�'��OޤI�B�6wٲ	[тV;H��`�"O,�)cD�5�x!�AD�e�����"O�Ћ�����дb\��x<�"O��$ֻJd4�&�W|Z5"OX����<C^>�k3�ʁZ�~��"Ol�BY-Q��� �	A���"O�d��H�cM�,��B�|���K3"Ov�C��5����D%-?(�y$"O��Z�͒��V��c#�3�xH���O�����q�T�B��*0��_�|&!��_0y���3HߞB(Z!y�'�^s!��P�Ұ=�W��@M�l Y]!�142�rT��/ ��J0�*=\!�$%D���׊�;5��2Ո^d�6�)�������S��quK��bt�����6D����'MT��UR��2Eƺ=[��3D�Z��?6J,�G_���A��4D�<� @PCd�B�j۸G��HBw�&�d5�Sܧ9�d�@�׷;lhS��`�6`��	t}bfܜ_\��f���hR�4B����'a{��"	.q��[_:���O��y�ٻugt�@v��;S�(�!�[<�y��ȄN�*0SCoSR�Z�B`+'�y�D�Gd���J�L�4Ċ���(�yb�F!U��0�J��W�� �ρ=�y®�,߬�c0�L'UL��y�`��y2�їf���g��M�"��B���$$�O�
p+�z����H h~r	"6"O�t�v�[�	q��fI�Eo4I��"OJ���qp
����iSR���"O~�Qa¨]����c�6I�x�@"O�A��ڡQ���х��e�0s"OxDi3N�:^\�r�}�R
�E�ȓ)��е+1C�D�EW=^��i��Xa ����B�>Ӛm��(ͱ<���4B�d8q$M>8�j�xAG�S��Ԅȓ�ڬXCD�x�� �c�-\q���+������'1�@����Q�w��P��!��M�sl�X�r�&Q���Q�ȓF���J�*1	l���N�Z��0��MQ&I��0�Q�I�R��фȓ
��l����D�~p��f�]<��`.�D
�/���ɒ�8f�\E��3͔q�"bK�B�)��^�����E�İ) �e��-YÜry�h�ȓU����MY� �z�W(Ε/���ȓL�U�E���
o
�ز���E���>����Ԁ*b�5��-�Hы�	�y�@ҥ�,�T��$;��E�=�y���PC�|bE�ͱ_������
�y�f[(Փ��F_�� ��6�yr�"� ���F$\hD��:�y�"��g��!�l �T�+uA��y�j���1�X�x�Ѝa�a�&��'ў�$�)���=!l\����x��Ps��-\O����H�7<�ބ���1p �0��"OB��D(_}.ȩ�Oҳ*��-��"OF ���dU���e��e�9pb"OL=��*�^�0��y�XD�"ODTK'��G��\Fa߀X�4�e"O�d�E���<e�b�o[�P�Q�%"O� |eCDおl��Zq��r�V�X�"O8%*%�f���V-��&� (;�"O��K�Y�J�h�WŊ�r�z�7"O:�� V�*�T����ԩ�K�0<)��č�m��=JEd�K��ي�It!��#��雩r�f��e�H��!�D:My �� ꀢ4+X�kʧ5��y��3s�����MFO�t���Q��B�ɑ��r�%t �B�o��g�B�ɛ~��y��>��y���X$�C�Q��́����i��CYv2B��:��P0'�0�"���n�SDC�	�-+��r�Ǝ�+F�`	%.�$H�C�I�s�>�0���'���
2g�C�n6(��<#�\e��iƔ(�C�	�_d��A��M�`H���C'�^�C�;$4(P9���XHZ1���.�$B�	�Z���H1�]!~�f���	y,�$F{J~��!r��xbu�Y�S� !1E�TA�<)T�f�*�H����a�
H��gz�<��A��E��h��ƛR��P-PZ�<!`�̔@���S��&� ���Y�<a$�3-�L����Ѳ>�H���X�<IӊԜ>�H����`��2��UQ�<�wbC��m�S,5�`�F-Ig�<сf�5	����goZhK�hqք	]�<�G�<u'*4"G�2my�S�<�5�ݟB9�){��3�B5iPOx�<�Q/�>|u���c�$ANl��
|�<�ҋa�|()�ɫq�N,{@w(<��4��͡��_�A���h!�����E�iO�+t�U�a��h,p���l96����>n�I�uN��9�xQ�ȓ>��a+j�
V$ɔ�;rv`1���s�pS҂QLD���F�v��iSRA)D�H{!A��#�$��`o�9֭�3�'D����j[��6IK�����f(D����D�B�`١B�'� �9 !#D�܊bk2 MҔJ%E�=[�X�Qh D���3HP�l2�HR�==�*h��C?D�p�äE���$q5ℙW���;D�tJ����%@'l�!x��,D��I%��>t&D	XC6h��@i5D��ؒG�z��]��iZ2=
z�Å�3D����C%E��(�P�V<�\<z�3D���݂/	�p�W�V�}��z�
0D�\���\�c6�S�<�Ƹ9�+D�d�'��kL��Y5���{ż��B'D�H�ul�,0t��f�)1�t��%D��k�烷{``���Yt�t�$""D�h���D)[�
	 ˘8��k�,$D�r夎352���Տӯ;�܈9,!D�� e47u�'��x�1�?D��)�锗/�` ��M�d{ת*D���2�<��;���:!�W�'D���7�H�tHa�\�,7Θ�j'D� !�N�*��Ո�.��D��8���9D�x���d������b'��2�	9D��f�P�J")�%߇^Br��(7D��)��3gO�H`��ݝ]/5(V�4D�`1��:��(S��7�4=Bd�0D�����R�5F��&4���4D�x����"����u�![J�aU'D��y$�F�LUء�E�P< �be�Sm1D�� V	�@Az� �������)��"O0�G�<Q���A��^�W���Q"O��hP�G�"�$� �IǶ*p�;�"O�\!�/J3:��j����i��@g"On�ٷ��1\=���T>Gg��� *OH0���H�w��|iAZ�V���#�'��mɠ��bAIS��-\�=��'��x�� Ts2^�8��[�P*F�B	�'n��*�G��PB��I�(	�'��)��P
����aЈct��B�'�B��c]&>�ht)A���[L�;�'��4�o�@BĞ�b6����'���E�هG4X��U�O��M�
�'�n��V�j�d��"�ߌNKX�s	�'I�l��gJ�t{�=CE9	\��'�Ц��Dk�h��\������'����ϗ��F��gؐH����'1��r��H=L�ɕ@��
2���'Ғ��d��ڶ�H��

3/�x��'Fh!p���9�I��-&����'���B�ڱP�f(��,M�P<�l[�'/��p��(6>���Щ^�Vq�'9<\���ޖ3�|����59�Ĭ�	�'z�� BP<6κ��.�1>��y
�' ~���/F�g8�Z�h�'�x"�'�@}�aNK�vl!"Q��/J��9�'�^��d2 �j���9A<<��'��4J5H"wZj���[�2�`=`�'��iZ�c"=�B@�A>|M����'�a��A�4���Cԯp����'�ʔQ"(�<=9Z��U/�e�@,��'�:�dFS�����3^���H�'�V8R�5����D����Uj�<�I�b��I�뗠8�8�XL�<��+�ymJ�Y��Y
���mS�<��Ɲ	h�� �l��h(iCp-O�<�7��CJ��xňB�&GD#��N�<�G��.�l�
��t����FI�<ys+>�����_������y�<)c�,E��Zp@�'�Ԁ*%�_t�<��C WM����� 	o0P�U��n�<�c :T��9M�������i�<Q��`l�ix�l"��9�qP�<��X-R]�!X��$ը�rt�I�<Y�#�6Q[$�D޼exVT�RE�H�<�*��,ڜ�A�93vH�(e@�G�<�&�fx��D9b�,]8�)�}�<�r��Lk*�!���>�����Ic�<�&T�}��DIв@J�#@�S�<����8A|�P�A-��i0d�(�N�<iG#�!:�9��ѧ?H��s`�F�<If�Y�8-4��0ş�f&(�(�ERH�<Y6�K��a���%M�Yh2�M�<%�% d��ڥ���d%��k�@�<�m�f�x6��8L�CvF�y�<�%��r�4�l-%���cFa�x�<yA`^.A���8%n�D��̣�Cn�<�Ň-�]�`ULE�P+��Q~�<ɔ���(BA��C9� �
b�|�<�w,*9���PѨβW���0B�v�<�Cj%L�X9F�ϳx`y�7�l�<��J�bp�(���_�R���#�j�<q���2)�  ��;XX�H�O[q�<��M�I���ʐ� �s��8�W��T�<� �(B�g��]��6��D�Q"O
aY�T 4@�z�l�Y�t"O���`ݰT#�4�����[���%"O��P���%��l�sM��}OD@u"O��
G��"��i �KԪ9+f*R"OֈSS���DM&aӱO�
����"O(U%�R�*�p����>(�F��"O� "Ү�!\�N9���Ԝ��"O��w�)�4��+R:8x�u��"O��1E�RT:��䠛�,DV�z$"O���b���Hp��Y[�  "O�0����*#���oK��Y�6"O�����F��4�$.�3��p2"O1Сn��J�8�c�G�2ըh#�"O�h�%aO�;X���Ũ�"�lp1�"O�CU��	��� �r��P;"O�)6�J�!�.�rmE�C�@L�"OV��L��I�,��*ˮ�z4h�"O����l�����&
�3NфYRc"O����M���yDn�HȀ��r"Od��G5��Y�`cY�+�𩘅"O�Hh�`߹`̠����9#�z�+�"O�]��/.a��0c�ˣ,��(#"O~`C�,�$6V` ���B�oB��"O���S� Z�t
X'Q��Ӵ"O��[�Vî���T<8i����"O��g�V���i��#۔�����"O��� l+���w� �>N(�C"O9I@M��0K��c� ~-�l�2"Oс�K c�ʁ�ކLn�ht"O�Ī@�V9$�"̩D�UlR�y�"O���H�ࣆ��<)B̔	g"OJT˳kR�%/6@АF�X�""O2-*�c��T��a�ѢԴy�>��1"O��Z��c�&�Xp�Y�A���'V:�'�ˎw�^�yt��0&�y���.�z��� 8�����Ŵ�yr j螽�gA�F��&�H5�y2�+M�40�䆁<2���&ʟ��y��S*rb�s���"���z�̍:�yR@]yi<p�Կ���j���y�c�Q��P�g$â�Y�솱�y�l{=V�Zc/�d��Q��I��yrܕ%~}q#(�qXB���Z�yEX�`��P��Ӹkx�2B���y2J�T�q&	��i�Q���0�y�%C�HS��`+��.�e����yr���M
�h�7AJ=2��H�����y�C^,@:�X����$$u�H�tGC��y�!�(0~�)�lO���$����(�y2@�xS�����D~>x�U架�yE�r"��6����h�5�y�.���c�Ŗ1��H3���y�*M�d��̙b!շ2�@����'�yb��?;��%{wJA00):�{ ��,�y�%�6g!�1��TF:h��l��y�b��a�ą��C�:{�Fԡ���0�y�ቭR]"}�s�P`n��d%A��yI�w509��X	=J�͜ �y���7O�&řV�-*N�P�����y���)E6l��%���h��K���y�'!OU����%Gm` �d�X�y��1F6��%��9�(�����y 9w���'De������y
� T��p,��bܐ@qLW:x|5!C"O����
Nkq����3#m豚"O�J��ְ'�2��Ӿ�B��G"O��Q���"@��D	��Ȟ,���"O|�*F� `9J�h�6 ���"O΍�ta��n�@�B)0b,bA"O�5YWEJ�:L��qo�<��a"O��p�F1x�<�s�	�w�Z=K�"O�<#�'��rt�I���dx��1"OA�_�������*�M��"OP	Ke��l*D8��*�34"O�aAtc�8�6�h5Ɍ���8T"O�u���.i)l|���C�[�Di�6"O&����XKb��E)��0r"O"��E�G��PJ�F)�>�)7"Or�[�)_1d9J0�Y{�J�B"O\�rb� sԠ�Ca�&$��8�"OJ}��E�*q^Y��,dDH�s"O�Pib\�=3S�̩@[���"O�\KUKO*x��YW��'�E�"O
�����F���р�)ǌ�"�"OL��LωH��@�S-��v��!��"Ol���<=�cWK^�o�NDQF"O\q:��G�M��4��)��S���E"O1�3�	������F�K�"O�]C ��`��I+��)"c"Op����XDy����S�����"O� ��ɉ=~0��'#� ��"Or�Fa��
��Uz�F��V���+1"O����H�-jC
��$x��"O�j �J6?���0�$%x �J�"O\ԀDbǊ]��0�� �d��٘�"O�ZVYJ��Թ G��6H�#"OZ�jPE Yj=ip�	�����"Ox�U*^L�lDnO�p߰�t"O��#N�) ��a#mPt�}��"O\�*֣9	̄ۄ�!D]����"O�9�',�e�-K�'[ /L �
�"Oh�9��?rwV9Y�,����:D�<�¡	+~�&�F�8"�`�#�$D��CW�"wQ��x��<.j-'� D���B��=�1�C�`��=��>D���Q`Տ�P)i��Y���2�*D��C���
&�:aŜ9K�^����'D�HD��+Qc��4gZ CAD�3R)D����ˌ�/4�1�IƇ#"��3�&D�lB�G�H�v$9&C�H�	�F#D�dȔF �8�Ƚ{5�A+ �v�D�-D���O��z}Fx��Ğ�F�0�s�*D��BCDl쮸�`霑e6D�$D���G���
i�)�U�_C�pSF D���E�jU�e�v��9?H8a D�P N��X����]���p�G D�T
CK�o���M��j�Q$M=D�(�������S�Icp1d:D��LpCA�_�j,Z��Zu��'0\9���F�G��A�шͶ[e̥S�'���b�Hܥ ��T�qf�?)?*a��'�^��s"�"g����I�6!�v`��'�:yr(smRjA�,Gbx�'c@!jӧQ�F�*U���6R�#
�'�"����	�k'�)�'�{pv�(�'�t<�����ͨt��;c6��'zV`16nN
(���Hi�_aH��� ���dO�i�� �!&>p�h A"O&H�mN2~������ݤm�ha"O$��Wخn�|9#+:l8J""O>��֤]��L���ׂPavH@G"O���c��+٠��e⋞}/����"Op�y�#�0��P���%���H�"OV����e#w��uV�	�$"O�L���>_�t;3ŀ;4rZ�J�"O�gW:�J�� ��Wꤱ�"O��Ác��`�=���H�%��0�v"O� ��(߸��g��.l����"O�   �#t<L�b��%�ҭ��"O� ���|ɾMz%�A	J�怱W"O�MA�"ԁD�x-3�R�!�F1P"O0Lk�A>y
쑗
^�/��d��"O���p�85byp b{x�r"O�u��
M�AN|�2�;�*��"OX��K�[�lҐ��o���+�"O̭�!铵xAtcp@�[!�Y�q"O�*'��/bƂ�,°"O�����#�6!���<I�R�S�"O�i��%S
WN~ёb�m�R�8G"O���� D'FlB��Q>?B��i"O�%i����%�bE�!@K>	�"Of� �b��A�("�A2�K�ybF�F�|�ƅ; �R�&ˡ�y�g�6�a�	1����v���y"�͞�"��sbݥJ"�a&��7�y�F	�]	�8���9<L������yb��=#�!B�J��$H(�N�y�(ǵ,q��k7l��"Yk2��(�yB��D5�p�)�'-dݩ����y��!$�@��"]�=�@�u���yҡ�?5C`�/ �Ԡ��jک�yB�U5D5�M��A���D�D�W��y�j\++ȴ��靌�^T0À��y���>Ƙ���D V4�+��V��yRo!=��r�/@<z��ʲ-�y�C�-�̘��sg"9L���yf(tu����,s^L%b6�y��J?�TrV�L7l�H(�eN��yr P�pNH�@E	6j�m�Q�T	�y�
�.j�v��EȔ1(���q	��yb�ȵfNF�z�V�9��aG��yҎ�q�����0Z���p����y�H��X��%Ʊ^WH@�`���yB�ër6I���Y��M���^��yC�^��i&#��ݢIE��y�딏Q��iA����i	U�V��y 3dޠX0V!�����IS>�y2F�"��tPV*�#��0&���y���9<>���&Jb1�� ���y�k�U�|01�T�a\��o�;�y�Ԉu!t@�� �K�2��I��y���L��!��S�B���*5�L#�y��Kvyp���N.6z*�{SEJ�yR�X�&�L����?)Xn96 ̯�yJ��R��5�Ӭ��P�k6ϒ�yb��l��q�O�	��`ZV��y������%�Ā	����u�*�yJŉO��S�/�N �%�R�yk��'$��u���s��D�E�[��yB�8��KS��}s��8dψ�y�k@;?2��+�M�B�� ����y
� &�)B
ݔo�zle8�fT��"O�X DcT|b|�97��gI`�"E"Oh�j� ƻzN@���۠S;��g"Ov��g�÷+�ձ0�Y;I;r�IR"O�ԡf�7�@D���ߵ`9"��"Oz�ZF+�~!�b��4&� :�"O��b�/]�V0X�i��R��)�"O�kê�!ed%�sǁ//��0a"O������(0!��Y��'`��@�"O8��6� ]�R���f�.���"Od���@c��Kv�_.�ތ
6"O�T�p���{X!`�ƃm4IpR"OЕ�IW�c��(2�Ӡk�|��"O:EXT��l d�yĉڔ��R"O4�Aԩ%%j���Z�Xb|���"O���Te.'�"�*���##kz��"OX)&����!�Ve��)ix�*�"O:t��@?J⼘��Hc��|3"O�T��fO{n�8a�W�L�<��"O$�[�X��ЭR�d ���P"O��� L�m��X�"%���"Odͫ��S��6-RW/
�?��"O�) 1l&b��}(�N��죆"O��B�	ֵ7"�ۤ�ѯ��YZ�"O�IyGl��Bl��R7�l� �"O"�z���m��8��	�3~t�{�"O\��ᮓ�<�h��\��3�"O8��C���Q�B��0�@u"O�<Т�ҽ�H	׌� �D:�"O5��N�lm�%�qL��c�:�r�"Onŉ�E� ���;�m,'P�m��"ON�#1*F -2��@�3l2�dZ#"O�\;��D�"�i�(�;ڠ"O����_0W.��T�� |��(�"O|Ix��{�t
����F�|�<)*�.U>���\ȐI�
�l,���V�TXd(�8�R��G��:8�zE��Ab��g�$,��(���<Ivt��Q��h�:�Z�[eO3}��%��Z���{֥�����K�$y��M��g5d����9x���&�M#|�,���'����J��Z�Z��s�ZqVq�ȓ<p�A�ua�,�nM+S��{��u��5��]S�BL�$\0a8p@8'M�نȓ���lϠ,ٖ��'�
5?\2�ȓs�F8�c$#3�tP�O��L+����I6ɫ��،'��AY%! (��h��q8ЭT�]�Y��F'l漄ȓT<,��щ]��c�*��R�<��ȓ/db���ʙ��.=���'K l��y��̘�&�r�͟kZh �ȓ{��	�䫜�g���d�Jp��<�@L��E�.V��H@��D��e��r� �#�.� V��g#Z�4u��Z;��֘���Â�� 4�ȓ5�: �pG�~��)��� 7^��"�^�@u��w�ĸ���9��T�ȓV%��/E�@��E�w�T�g�j-���f��,�3�M����}؆ȓ,�~U��y�	;���1h� +�"O��ig��(',hqRs�E*X�h�+"O>���� N�l�X��ɀ	׬���"O�$C"+u�V�`V��j�`!"O���nѠ?������2C���"O� �r�Ťr��(��ڇ�fc�"Oz�Z�"R 2�h�*T�5�S�"Oj�i�#%��W�I��Eg�}�<yA�8Gf:eI���"BuЕ0�@�U�<�6GЛb�@K⍙0�(��t�SY�<�ɜ=r;0���K9���"-�T�<4�R5@ @`�����TnO�<1�f�;XD�q["�-�jwC�c�<� (�2=~�qA�ʇq
�9�&�^�<�"iV;_ֈ��6�K�V8iu`q�<q�)�X��I�C�Ub��)�b�<yw�;(��"������Z�<� J$�]��Ě<���
�W�<Itg� 2��Ġ�6WF��{5LDT�<1ǃ�o�Rp�G��k~ ��i)D�8�p/�"�(�)���p��ע$D�<`�
�dֺ�)ԧ��8�t��!D�zRI�g#(�0lݙC���,D�胂��1v�rq�l�3;�
�+��5D������� �rX�qhǘ�<�b�4D��*��?o��A�Ɇ�UP6��3D��QQfA�Y)�t%�+-�5#j1D��@�]�N�A:6	�\Zԍ-D�\�g��xԌu� ���4���?D���Z�)�~`0dr����>D��0�*��D�F�.M����2D�dÓ�U��4��O%2��]�'�.D��(�AV�	�䬲�*@2�����K)D�d`���2�~q�L�3X0��Dg'D��pJݮր)�( "����Ǯ D� ���)` 8����M��{p�3D���&�#<P&@!�¿0��$R��/D���A

�_���b��@��6��`-D���V�ӓs�J$�R�ӭ*k̩�?D���um�Ц,e�ѧ*v���=D��a��q�JT;!�ӫ�}���(D���F/T�m��� �<%� �p�N;D�X`d'�}���Q�*�!��@��$D�Zv&�$���Z1��%�h�"e�$D�����W�
K��襬��0Xc#D�Ī��ʞI(EB+�
#0�	�'L ܹ�G�=@��1��K��@�	�'��p�%vIXפ[J1�}!a��K�<ّ��:�f����7~!�q�ZD�<��O�C�xE������qSjPA�<y��Z���r"L
6=Hh;G-�@�<!'�Dj����Re�\���x�<��R���l)��N�pB��Zv�<�3	K�x\�w)� �t]�4�n�<�$JD�cS����J��U7��ӓ�n�<��aN�2���{a3V
�-��Ùg�<9�4�0A4f,u�6a�K]b�<�w��L���T�@)�|2��C�<AƎ�wYTh�U�D�w� ����<a�ڙ)�p��īŸ>� @B���C�<9a��]�(|���	1��@�Ëf�<�$HM|3K�3n?؜,i�B�ɒ"�vx'IN�W�Ɖ:��!��B䉬H�P�-Ԝ�ڰ��h��(��*D��8@029 h���0�\��a;D�r�ZV����`��*lWX�H%C;D�L9��A�x^<��A� �~)v�,D����a��l�[�ϟ�i3:K��+D��rt�W"��5�ܠ6� A�#)D�� �t� !>qY!��?e��S "O��6gٖb���3�����q�6"O���B��0~!s��.4ɒ�0b"O*�i���&$ŢH٧��,/$r48@"O޴���SIk|T���<�Ȕ"O����ቅ[�����W��!�3"O�`�c��f�t�x7��6�N���"OE�?�F��b��׮��""O�ɉ���\RTH�s�HH9�"O<����S�hE�0xf�Ы'����"O
m�&I˃1�M�˹i��T`"OZ���V�
�R0x�X9TD&)�"O�����Nwڠ�Z�'T]�m�E"O�qȶ+̗5���k����LF2���"OD��� 
E+���9�x�"O�t�a�!�Թ!��
= X�!"O��Je+·����G��.��I�"O��r�Gq��y����H����"OȵXt#8l��հ�"�2�0a"O��cC�g@�VBL�a�|0�"OP�A�� `���#LY2٢�k"O�d�� q��1�ӛX�ƽ��"O�P9�#҈�ٲ�˸q�H�p�"O, �q���n��E�KQ�@���"O\�iQ�^�&e���"n<��K�"O0����^<W��l��'�),^�r�"O����j2&Tq�G��o`��"O��X���z�4勵���'	���D"O\y� �=`l���f�=8���r7"O65c�E5=Fݢ�
\�ٜjb"Ol��fJ �ZёS*�5�(�"T"O�IQS���gc�YR�\�_猘��"O�ɘ�d��Dj�Ԙ�@�N ��r"O�0�N�IQ�C0C�1�"O�eqSL2�2�l�(6���E"Oȼ��	��[��0��� 5c�ׂ"Ox���Ϛ
�9����\$��)$"O�(W�O��J�9�eǕg���R"O\����\�K�Nd냆�Z��2T"O~�:���K� �%�!�&��t"O���ɍ3ː��
@gb-�7"O�]q�� P<��)�㚁2HN�x�"O��B/5 ����Y�P<���"O8�˴�Axڎy�4b3E:b"O���g��Hl 鰧�D)
�3"O:��B�U�a>���CJ;��`p"O@�bamA�,w�Ȓak�=�tк�"O�㤩��f�t���,A׆c�"O<�+�H�G�n�2[3���u"O \��§n	@��a�	q  cd"O¼9U>*G"���Y=h���#"Ov����ܝ��yV@��F��8�"OmAU�R�ZƜ=�g���L�%"O��h�#B�����plŅWM����"O2�jM[F���f��3;��@�"OAf��7},,c�N@�LMB�jd"O0�9�G
B،�8���93%DU"ON%4W)nK���g�#D �2"OKC�U�T���͝�1)��1����y�I�Z)��W�W�~U��(����yb	�7Z�P�SGΐ@��ŚW���y"`�E^��ڣ6��iI��ը�y2�I�5X��R"˵(W�"0g�
�ybEu��s@њv D9%-M5<�|��S�? ��H �W4�*�i�<6�`�"O���O�����Mq�4�"Of��6 \:N�T4"�m�V��@�"O:-�r(ӽ*�<���\�`�n��Q"O΀ >t����4'��eN��"OY�DN�x2���R��2�&DpV"O��JR��%_�$���.�,c"O�'l�&�L�CW����Αq�"O��{��J�	�,�I��� ""Oh���o��n�R�BDEFb��Rg"O���4^-�Y"O��oK�4R"O���1杏�803eN��>���"O�!
�M�wڊ<���ށ0)�P�"O�`�gN&	��C, �R"O�������z�VA����Z�@���"O���NO�K��Mj��1Xƪ���"O�0� c� 2ؑj�	 -�̹��"O���w�^�%��TZ�K�t�L%
�"O��Z�Ll�TXb�lپzDU��"O�\����tV�v��KY�Ѡ"OBat�Z#f�&�SF��_��в"OT�I�O��x�S���!��ؖ"O����s,P�R�T�a��@�"OB�y��-f�#�@-_N����"O��VB��~L�	��_��~��"O
P1�o�*}�hqo�9��8�"O�@z�i��"�r���C?qoj�b"O�-�5��ژ#�,�G�ّ�"O|� iD$1�"`�U�܁����"O2r�I͒B�|�wꋟt�>���"O���4#�-JE}:���k��PQ"OPP���FW�԰AaȖ�p�<"O�S%(ɕIL^i+Fa�.F�0�E"O<\�� ��J���o� $�&"O ))�NP a�8ԑ��ѽ.¼�Hg"O��ڴ���6@�I0��U��Z"Or��'ؿ>eDq1��vGZȊ"O*l3eĎ�
&��8�+��@���u"O�����1j���r��ɹ���ѳ"O\)��ҹ2�z98�I"Qn�q�"O�h�R7J1���DH�p�͚�"O���^�SА�
���q�L��"OT���*uQ��A0OF�� ��"O���/7��9�ç��z���"OQS��N+H)'ʝU��i��"O~Ԓ�@ˎ_�e��&Z�I8T"O&}�#�e�
��q]�H���"O�u�5��b�iQe�/�*HR"O 59�gΣ8�2�Hڈ�=bc"O6��(^=2`��h�2@$26"Ode�ä_, ,�d a)N�z	�ɐ%"O��R��y���*7��M�N�K�"O�"���� LPԐ�aD�xǖ�"O��a�o�vDi`��T�;�vmh�"O�`Ք?6��T��,sb8\bD"O��4�L�Eڒ�5��-	����"O���@I��RH��	��Su"O�(p`��	UҴ�C���$6ܤ|a�"Ol�,�*3Y�}2�V[���w"O<�VŒs�Z�k�ȗ<�JX��"O�Ir��*�ӂaL.�2��'"O�!�'��*tv�ȸ���7,��X�"OP�`ӄAoB���!L4;��pk'"O���͉u�z���Ȫu�Vd�d"O� ��+�#{���S�
?XW�)J�"O(3�
C9I�jxh�d�^��"O$�1��ڡL)�ъ䒩R��Ybt"OH݃4A@�?�<A1���#�"O$�	�$�� �TD ��	�*̙"O����D&n�v�B#	����"O��)�`�-_�D�F�� n��"O�a���^�o�J<�����}�����"O
�2f_`����+�	�nًE"O��r�͜
-:E�F�F��$EX "O�=A�&��XR1�U%ޥ}�\��!"O�}Y D����"��J�~4�"O�D�`-/(�b<`"CM��H�v"O�HRa
�>@n-�4��	���B�"O� 1ro�(f�<R�ȴ&��Б&"O���� �� 8$�&A�iH"O��ɸ[��mCb,�m/hk�"O��c/� ��K<k(��f"OJ�RwN�>f���R�ȥuH�:�"O.LQ�K̄N�h9���2D��C"O��JIWL�J@K�
D�P*�h""OTy���X�Ъ�iY���$rp"O<8�#k��D�a
�(�����f"Oؘ�Hˠt��q���ǒ=�H��"OM�AN�-3�*B/K)��l�"O���T�C'�\�|�|�A"O�A���I2b4�",T$����3"O�I�%��@֦d�"뚩�Z|B�"O�5�l�1 !KņQOܑR"Ø��yҠ[�1�~)��IP��q�N�y�f/$�sQN_�Uľ)z(���yV�z!k�i�Z|`��/�yb�=���GG�~�P�Hԉ�y��q��)=��8���\��y.�ac�B�55�Ũ�f[�yR��$R1��k�c�&1���h��S8�y",1e��%>��X�F�O��y"���X(ܥbSFU�;&x�S�����y��I�/��)�%	$��tH���ybGD/J�p�Y���o����N�yB� '�X�Y3��)|�XT#�!��y�S^��9��,T�n�}���I��yro>0�A�/gd����@:�y�g5_�f����^�x$cV,Й�y�o�m���
�(�N�(}���&�y").�ph+��I !R�&��yr�_mZ�*��m���/��yr*R;29����l��d����d���y�慳O�"���(9Z�N�(4���yI�e��ɋ�,�(����sFʧ�yR�gP���l�����у �yRG�x4(0`����`d��y"�#`Z�X��^�q �R��yR�K�	dZmAb��D�2�-�yrL� [Ejءq�ڡA%Š����y�h�g�4��N͟<���0�A�y�D�p��f~��&�SC�<��L< �� ��\�j!r3�E�r�<���]94 T��'�I|ɛ�!D�� �LҨl>�ū�3*U@��$�+D���7bK��$A�̎#i��&�/D�|I�n�pf!�����jAAR�,D����{"B���&�9�n� e)D���7�%b$&  Ÿ<�(ݒ��&D�� B}A�M=+�r)H4HԎ(�X!{"O���!PK�9S��L!�	�%"O���-T�i�X`A��q�"O��J�~������%�=�"O�ܫ3[�K�@�ZjM�,��a�1"O:���	i@���+�p�e�"O>�H�$ {��$�����X"OJP�q��p�����d�06�Ș��"O�L���ſJ�y�"
���Y7"O��Y�ۥp�~`�����7�:�#"OB5J@J\�&s̽B�N�ux�Ka"O� �Ś3xVPS� �����"O��7�J/\ ̹��ߧ �r|´"O��F*��晫sO��Vs�A�"O���@D�]�h}(R�?�(p�"OR��w���E�0�e�D�y���"O�e��G��D�e�ċ��1�"O����9a� 0��C�R�d��"O�D��'��Zt��5�R�R�b,��"O�,s��K��N�
�F�4�8V"O�<ڡ��� �&M��:|�"O� ����*o��#�+��a�"O�H��
�~D��)h�|��"Oxe�r=L|���P#�x���"O�4#�M��-����bB��%�!�yRn\�bGI
��F�a�t�d���y��^�gX��X4N�?Ut�Iz�����yr��?��rF�Q )[��	�y"�#^
͈�*�=`��`A��y�܏(�xPm@V�tu+ql&�y%& �f(�U�}�"���!�$�y�h�'$�=�4�I+R  {3I�y2e��h��T�Q��8'�~U���y��5>T�������~��k���y")؁Bt���舔g��A�B���yb�W�~*�Tz���D$��D�.�yroίD�ƨˑ��@�6q@e���y����� I;��ٟ<B<��&`��yB���;"��O�6t�2'��	�y�DI���%��y8 hB%Iݹ�y�jޗo��H�t�e)�F��y�F��+C��h��:�,ئ�y�H�:�t��Vh=c:���0b�y)[y�!y感WK��
��W��yR섖CW|�*�eD�f�!��@��y¤O,Q��pP�ؘ[E�rg-M<�yB���kY`t���(��`�'!$�y��S�\��i�!�4
D�e�化�y�#TF|@�bF*A�*0K�&�y��C'����ĭh񒅹�*%�y �'i+�aʳLɩaa��y6Ç��y�X�Y&  �� �o���]�$�ȓX���@���6��m9�J�*[�E��1d����GF�kP��p�ĝ�P���~� h����;~nL�*ւ.��͇� �����MB���U���pOJ(�ȓ �̊ÁQ�r�
p��!�8�L9�ȓZ0�p�ᜆ������-�2��
0���=m*3#��h�2q�ȓ|$>0��i-v*Q�%I��2���ȓv��9��!V�Hk,�4��e���ȓV��d.
%w��8��E��b����ȓ 1�%�OҿO�f�7̔R>�ȓL�@�3aA�=%k�(�B�E>S�(���S�? �����rsQ��V٤-Y0"OvQ�.\��!�,U�La8�"O���w�	1��s�J�Q�����"O��°��2`�T��$J��@���!"O�a��L����(�c��*��M��"O�)A1�$����AD$�K�"O�A3!���-"�OP�.��C"O�,��+�L�y .لEp�d{1"O�d V!L"L8�R�lY C�) �"OfE��֍Z`�5B����I���)f"O�er�ڋC>XĀ��'7��a7"Of�Y�@�>Ni��T�`���` "O�
��ǵu6�X����%V�䀂�"O�@�%�<W��Z�H��P��w"ORM`����Z�E�E�? �&=D"OX�c @�F�cF�V�n�PeZ"O�(�	��** ��( B��̐2"O6���c�L���'�рq�^��"O@ݻ��I��Y�����v}*�"O1��('?�Ѳe�Wl�8%�1"Ob�k�D�qpP����Y�,Qp�"OJ�B��ۯ�X}!ab++ͼ�c�"O����"��p��B� �v)y"O�e�Wi� `����ᕠ'�j,BP"O(��(�&w�����F�?�J�(�"O�r�� j��鰠��C��U��"O8͠[�0*�N'E��2���J!��*;���q�P2��sb�h�!�D݆~`l����9��8���<�!�d�d��,�K��My�#P��h�!�d��8��I�:e8؊3���!�ă(V8�����3q+.�`Z�d0!��_�`�5Y )�<�K�1#!�Ē*=QLHk��K�T$F,8TjF�!���16Ն�h$�p$(�R��!�d�x�2ݫ���i#��(`.Me!�A�O>4j&��"o{��I��Z/�!��ۥ&�5�c��

0��ǅ=k�!�$Ԡ�
Is��w�-�sd�-�!��AH9b�!Ҥ5��Q�#��!�35$u�����8�WM֒7�!���)�$�kC�_�W�<�P�&qo!�D�1� �0!��`�0�dgF�I�!�$�L�l��$̗H�����&[�@�!�ٍ�N��!��f��8j!򄕞w��pK��񺕱V��"}!��&~��0�0Ώ�e�ĸ��/J�.c!�$ �"A�@��X6d�ĉ@�WZ!��9�ċ࢑�F���5o��f!�E(_T8�R��P�A�����N<b_!�O�vJ�%PFC� �5RL�TB!�ԗ5����ֈJ�q���:#.!�	1�iI�cJ`�Vy�� �5!�� �p�N�I�ǒ5:��l�� ��V!�ḏ��M:���"%Ɇ�(�NÒF!�&K�����\�Z'�$a7G�td!�Ҹ;��  u��	I��i���.D_!��n�l�QE9~�����<US!������{��o��lJ�i��&�!�4ecLy�H!{д�R�Q�R�!���4u�t��3�&I3���%�!�dKQ��L[��]�O�:U��퀮n>!��7!l���"B�$��"�c#!�$�$l!*�Q�h�t��!��ɋ3!�� d� $O�� l�@�ULق��@"O������~}p�(�
Ʌ)�~q;�"O��������zi��*#��q�b"O�Py��c;���%0b�P�"Ox���F8,��$��|����"OTy'� �EӺ�JCߥ{�X��B"OF�;�B̭H�(A)wa��tb �"O&��G'y�rq����>�,��"OH�R��_�
H�tI�d�а�"O廁Ú�B(��Ԕ��	��"O�h�!�V�7�a�P��
Fwd%��"O�4�n�[<8���fܢB���Z�"O�a�$�R�C3��!Sf	�XN���"O����gʃ�|�aGl���%��"OV��`����h�{�`��#�@��C"O�c� �v�tH
@�A3f��ea�"O<�!2Oʔ6�f��b��#�� 8F"O�I0��.�Vg w�	�"O~��b`�D�b��QR;
��"O�<�$�F	6����gI�w�b��"OPP[c�$-֬��oH�&':y�"Of�$�A�h��i��'"Oʴ��R=a����̛k���1"O�sK
v�~yJ ̌�)�h��5"O0suOX�^O|�b���**����3"O���h�@��0����	,0$�h�"O�\�sBP�(N��FgM� ��$��"O�eQvA�;P���`r�՗)EZ�ۣ"O���"#ކl�X$����w���a"O!��)�C�e#��۞2��v"OF�(��<�P�3J�TߐUB�"O���3+�j��lڕ�
���B"Of�1��K�r_����l� �H�""O�}�r�^=^,p���©1yd"O��[%%ʼi�e.	C�y�D���yB끃<��8�e!�v��c��y2H�\v1���i�(�@b��y�l�9{�qk�'��q���y-=]�(��g���̼
a]��yrT�=&��p��ٍ��1����y�	�X���R��5����R��!�yOV
d�ճ��ڦ�&���g�y��A�W4(y���~٦�����y+ĂG��!d�<~#~��1���y�`խP3����o�R�8�B��yN� F�@�բϤ_�x����,�y¢��f�dp��g�j����/L>�y���9"|�Y���#g�F`83F�,�y2&'K[$eh�l�co�ᅤJ��y"(�kZ�!#C`N�^�2��0a���y�!�6�4[��=e�B�S`	�4�yR��z�ʄI6�>^�ME�˕�y�
��!�L-�b�Q�]�*�(dkP��yr�D�(t60p��O�-WB�ɢ���y↞I0��!V�<��Ba��y"'W�P>����̙73 �"�F!�y��ب^���k��J�0�ybf�&�y
�dj��e���}!�y��D6����lb�ɞ��yb�U\ݰ$�q�@�#t|[����y�.Ά6K�����?�:����y��a��ǍI4J#��Ye�9�y��9z��qc�w[B�'�	��yr��HX�1S�mդ  �m��nN��y
� �9�J)�l ���أJ}"�"O��[u�H�;�^ A�aG(?����"O2�J�"���!F���Ȃ"O8��	�{jJa��%��T��"O�j�.MZY�P��C�Ԥ�R"O"H��ܪw� ���V�s	�d��"O05�bɌ;(�8�DAJ4p�!�C"OĠ��7�I��`�`宥J�"Ol�k���I���,�	^ߒ�4"O����ώ�'A����b��5@�"O���O� cH-���3 �@�Hs"O�rB���#C��sɈ=a@"O��B�l�:6%�`Z�E�91�Xiv"O�=�(�`�C�C֔�(�	�'�bz�m�}|���m�(���
�'�B�� ��D�
��S�E��
�'Y�-�D�� -cN�؃��-���
�'�$`���-Ce�@
�����I�'��9QV�T�<.��)L):fك�'�r� q�J�&���֬I�<��3�'D`,N��4����0��@3
�'�Hu���3g�)B�i�/]`.(��'�x�Cj�A�J�µ�$P+Thk�<!��G�-����_����@�h�<Q�a&P��ȱ���$�`��ʅ}�<�sj�n�����pA�蠴�}�<�!M�3Y��x�򅗃,�L��Yu�<9�o�(S�^q����n&X��s�<A�-�1�h����K��}��z�<�^�%�N��7M�'>����q�<ɕJY�9�BQ�E��K���� ��c�<���ar����H�;Ϥ� Ch\�<�F-ʠ4�䉐$�qHHp���Z�<���5�&sT��\�d`��Y�<��� �`��鉓hۑE�!`��(T�k %��O� �ؑ�ǕI�F�3TD6D�$1fh�9Y6����
���1�`3D�|K* &ݦt���9R�PP�2D��ْl�'-�J����C� RD��p�1D�����2���Ċ� 7"*PhU�*D���@
E���i<6��Ek(D��[dS�>���6��j�±r''D�p��<}�i��=e��(��2D��8�Ýx�BѢ.�O�(p��D<D�\��92��x�@��  8F*=D�8+u� j���o�A'�AD�>D�8+!		<8
tXw�-_�H�6E=D�\�r��,���ȳ'����A�a.D�p���U�Uu����^r�!��*D������O-����T���H	fn5D�4�pkP�,� "�c]M��qU!!D�z���5� ��]	e�,���B"D�Л��;HR���Z�"�����:D�tCD�5K2�M{�ė)N����:D��ZsHG<G(N�� IV_�.���;D�p9#%V*tpd6eη��Lz�k$D�|��,�?���� W�Qs��P�F#�IW���'�*ё��@,p�Q��(5�ȓ.b-��[3Z����D�B-T��'�f�)�'_T�PаG��Zk�͠��T�K#&&���0�'T�Xv�[%>�D�;�M�A!d�8�{B�'ߤ�Z�&�-q��E���A�T���'�ְ�7mB�FJ�HH%K��IŲq��'lTX@
�;I�,���H��P����g�� �Q��AɅ`a���Γ%hw�	�_�LD{����13 �{��	zނ� #���@���S
S����`�
Y��ႏ�UC�1�>���3$s\�٥L(s��B�I�e$�h'2s��d�]�+A�B�ɢ1,���J� ���gܱ<�\�K<a�O�b>c�|!�j�	(upb@�Z$D�ФᲦ2D���2Y��}�r�EJ��,"�{��7=�O�q��̛
|p�p��Le8����'��$8}"-f*�)`��WV�jB鋄�yB)�8^t�v�B��rF��y�G[�Jt���'6���@2g[��Px�it��9��̱X/l9��(��pڄE��)��<�����
��Y
��0S��A�hz8��Gz2��\�I���J
��-�B���yr�$e�����.6@��R�@��p=�}��L-�n�+@�
zt�'"��yb�ҟou�@"�n�q��P@n҈�PxR�ixԴG��^��T[�L�l28��'6p���@N�k>@�v��]�r���'~D�b)W�s]��u( 
�@��
�'v���gҴ|�<59q+ɡFYt�"O���Í)z�T$�D���I�$��"O�ِ��:209Q*�|.�� �"Or)�$M�.P�����j[�p�=z��'*�'�vԓ�Ѹy��D1Ǒ�
g�P�'-`B "�4�̭qDo^�~y���'������7&���#V>nXTm�
ӓ��'>t���#@�Hz[b�9m߬�p�'�:%�C W)j�~0B+O�c~����'�� �)�Ӟv��ւ�\|VE)Ǯ�.1��!Z� T�y"���P�NpIF��.vJ=ɖ���(����0L���f~2�iq���Ə�D!T튱$ʺ�s�'LO��'���..����Jc���Ǆ��?S��z�'=�V�)ʧ/l2�p���B��aBፉst)�ȓm�渁q�¸+�*萒��/����=�ۓo6*�R��]*��ؒ!O�&�:����d,��?c����\�V��5�v.�H�`���e�,��I`�i�B�3ENe�gɓ ���<y��D�K�oǞ��$e��J�De�`�I�����?�l��(X�K�R�J��&���r�0m�~����sӺ�����!8hP�k��@�1���'^z���3A�ݨQLV!&
��1G� І�ߘ'�axB蝺ysTt�@�M��X�H�?�ycQ+yL�%�g�،D$��2b��-�y�B+}@vl+��<&@m�����y�`A�{�"���M@K����H��y�(_?h�г��S�I�����)��'r�z���4�"N�H�h� ��!��x�G2�8�a�����7��	W��C�	+{�����ŵD�lZ��L$>B䉗#�r�QQ�Z�C��#���(��B�M����K+\���'�I/����'x���S���	��H�i}����oU$�*B�I^�b�[��0���� �$:�B�I�`d������{�F^�=c�C�	�Lg��PbC
 Ֆ���@��o��C�I�4�� ��;B�� �؛H��C�I/r��N֠N���h̄3I�C�I�c7��£��72�0�X� �����D��O�9�U,A�o7$�20Ↄ
�u�p"Oz@���F�8�P�X�_bEZv"O��i#F�9\e�=a�Q������"O�t+�bE+t��PC.�]w�����7|O� p]�#�hv�;���l@`�'S���隖 Y��Zh�X�L���C��O�C�	�g���`\�%YmQ�׌:�0��"�?�{��JSL޹#���i"�y�`nH��0=�,=�	-n��,ІWz�7�[�� �������a#�)�SNy��O%�:�q���]{����A^��yR�?n"�i��*�ѩ�c� ��2Yo:�h�A�̴��"��OaB�O0�:�Ŗ��fN� #Z��F�oӀB�I&u�L�H�g��@��ʁ�x���}�'���4C��#�H���;v��A�a�+�O�O�}c�5�F��𬓄Y��4��"OИ���)q|4Uj�+LH"����	L���iB1{�� �L�i�L�S%��<v!�d�M��
B��#=ql���G�zz�=�O��O��{'@�6w�����gۙM\z���"ODeᱩ\7P���	�+N>�T"��$)�S�'+�McB���z��M;� �M�F<�ȓ@�B��M���ZPED-7R���ȓ-<p��e�j��J'jG��\a�����M$-�'Wń��ȓM�DY�)��&D�!E�ŽO��ȓUN�A�� ��H��ثF�.��a��LB`�rGJ=> �x;Q�][���'��d(�H�OF��2� �dF>i�Q�-s8��'3d�cV��t� %�0m�>a�)�ObY#������pQ��o��������Y���VO&�O0�NuNU�ń�+ŜM8e@�+H<̓]&��?�z��D�ØT
r�Z8�2=(S⑦�y"g��ZS�P��	A&���� �yB���q�N�ZelÕ�4�!o\��y��)�`�I�A�\H:^�t�Cq�R��ȓ�D�[i o�ꉜj�N�'E���ɥz[b�ن��;>�P�$m��0k ��ı>��E�!��x�$��+��C6��~!��	��)�))�4��eɕ2&may��	�n�[g.CA���C�� ��C�	�8X4�
p��tjU�fc�<|���hO>MP �A�:��Y�Fߎ\b���:D��j5����fH`)����Eh�w�|�'Jf%�XE{2�г���oΈ ��
vo��?��'�v0�S�^�G7��y�ȍ$RBliʝ'D�'yJ�ƃ�h�D* o�G��<��'��Q�ɩ~��-���P�>=��a�'Hz�(��,���js H�* ��1��D5�$'�'e*Q!����d�6T�WL ��?BX���*�<X��Ў"��iA���s���S�P1{"t'L
��`X{wk&D��Cҧ��a�A0�F�f�:��$�d��=��#�;Үb#�*�%E*�D��4$���<Tb�'^�	�2�c:y4�ȓ2c�� HU�=D�ɴ�9uPt��<1O<YG�1ҧZ$|��F�.5J��I��ĭ����P�8�1B��*x���-P��ȓwl�0 �)�Jq��&"|��ȓN: ���� #���0�՛>����<q0�4\OhU`�np�q�qC�Pey��"O�%��32�4��V">{Iv�"O�Tqs D</�f}2�!F>L��"O�a"��A}2�
RA�$X4�ʡ"O����Ü��1�6����6�!�;D� (��	b�5g�Ol�hH2F=D�8�JB:����r���v��@/(D����s��bB��q���Ӯ$D�� �����JR4�U��ɚ q�"O��+�c�R�vԫd@��7
B9� "O�m��X>
�ro�MBtv"OP5J���xb��3z��"O��6mԣ (r͂(G�FybD"O(�I,fq����M��T��"O\�Z��Z��Pp���h]��"Of���AI/U�r�B��94R��"O����-�0!�s�.]a8E #*O�Q�Uo�28�C��6��T��'�� �%�ݪl,��(3F�Q�''�x�)N�;o�!@�	,�Ɋ�'P��צ�`�����ܛE,t��'IکH�k��t����@�9�,�j�'�����3m����g/	���`�'�^EhA]�[F0T��iƴ"�ұ"�'���Z��QS�HApdI��KB��'�\t��*��a{������$��'����@8���$���j�œ�'��	3aN�M�$Y��KR�y"`X�'#�ґ�P+�tA�h�(�����'�t�Zu�n�BP����(/0D� �Z{ �c��p���ڧ�#D���C�&B�P���o��MRG!D��a�K]p��2�S�,�dH3�� D���u��bLxs��)v)R��G�-^�dY��'�O29��A�	kxl�t�;"昱�"Oh�JP�h�(l!jZ�c��9@"O&|)u�_�V���'^�N�m�g"O��M��0���BfE� �`�E"O�l�M_'���e�G5g(�3p"Oz0�bE{.���ɓ�fJH��"OH�[�GZ�E֘�kS�?x(}*�"O�hK�j�
��\I���
q��+"O��$��Z�"/r�\#�"OlHp���q���	Η>V��a&"O�,p��l��S'@Τ�B�"O�`�/�%A.���F��ށ��"O������r��(�2Tdc&"O�A���^F�RѥgX�5@��"O��Ya�Ƶ��,��̭H ��"O:��E�V�U�;��	��X�t"O�qDнg���80mؕ��#0"O�@����V<���@L�#jw&��G"O��
4O�A��a�ȿNad�h�"O8b��ǰ3��-�WkA�|b𙫠"O�` ��9Y4�pcԄ;��:�"O���,
)�hX�j_���@�D"O�pB�]�m<J��i���xY�"O���J)*��)�D�s�� 4"O����ߘp&(a���)#��`�D"OL`��ѽ>ꊄ)���z��Ia�"O�u� 퇣*�j �	
�>Y	W"O���l�4�Z�"@��F����"ON! `^����k�@�f�؈���'���(��^�Wɧ���E�ƚ�[��L����m]�����>D����!��&J4)��	d�l{s�>9q"	*%�X CF;<O���t%��=�z��F��%>����'�� 
L�o�,I�� ɛY��ek�\<hiI��]!��� N��6�@0H���ⰃVy�Q�̱g̀�*Z��Vb�p�j��1/�M�`��)�i�ȓ|4���$� 'є��u$� f����_y ���HH7`�l����2'��`��ӕH��2Wm؝�yr��;`��F�dar�aGb��~��Î3f�sSͺ�ay
� P�+�LܤNK���KY�i4y�w�'�p��$�"R�4�Y&p������+PF��t&�R2!�Ď2d�(�x� P�V�>�Y��C�6bQ��IC�0a�<�8ŀ�I�(;��k7���v�������=B��d�ȓ
��9rS�L�>=.�3��>8e05�`��"4R�8ң#?��)�矼��"�<
%�114`�`D�bH2D�1P�xS�mR4
աy 0���ʰ>����#S��#��<<O�9��J/&���p��
!#Q�'�)3q'�=�jib`���_���'e~B�8�"O
p�	Ѻmޠ��K;z�n�;1"Oi�l� X�����G�3NL���6"O�Ȓ��˧ � q��Ї �fa�"O�S�B�1�ip����$��y�"O��#��!_ b���N<��\�"O���T�A*t��Ty��<d#%#0"O��1U�S�E��Q�ƺd'�|JC"O�<�%AP9{�.ēE�=^JG"OB�QUFF3`gVHb�'Кv�x��p"Oh�����F]��]�\��"O̼�6�]�O����΂
�P�"O�!�$@�͐b�
+a5F�9�"O�H�GF�Z�b����^+d�(�"O~\�e'�W0T59`o
�d)�}"O��	��ꍨu)�<ɀ"Op�Z�D�l����3�L<:� yҡ"O����Nת�^lZR��/{f\Ab�"O� {���7h������k{~!C�"O�mz�@Z=�^�P.�0xW@U(!"Oи ��;3��\`��+a��}�"Oz9�D!�&G�lP;�B'�.�q"Of�t,��l�><���u�0���"OL��c�޹z��4��"҆Q	$�	�"OT��g�Ӻ\a*-��*
�J��E"O��IŔ�}�`�3�*�52e\E�u"O��)��6H#��x�,�+_��Q�ߜC�,h�$�'�@t�J1�|c���._&�ӓo��%ӑh���$*���!)&>�QKC�k�!�<E��͉Ы=��؃u��H��	�c�H��"��mo.���>�>�Iʙf����&+�'��ڤϊ~ a}�	�JX)�,���Q��@�<=1x�bSjA�;<`��$��I�xqh���O��2��6.U�Z5�E$,����	�=$��
���7/T��Z�Gᖴi���	f tB#Q/vfۨ���'��>�1��z��p�B�Λ]_�ݓ����5�7��5.�䴥O���(����5����5\z�ꠂ�';ʀ̸��r/tB�I<\���iC"b�� ����-@��ɛF� �U�X�/��]Q⏞n��0iUn�'(u�t�D+��o���%h��8��=��	 +Y�Z7D��?��IыJ��u���^=2��9r#(ٚ���OL�Cd1�3}�Z#p�n��p*X8RiqtCD��(O@``�[ v�`���'��0���?�C���=�p4KqH��Iu��2��5=va����a}��K68��(�3�_/%�xD�Ł�!ʺt�#� ?���B�'P�1�LK79��$�_�'�rT�5��h^�?l�Q������.�y���R�X1���	�,����6vt(�Nzj���L���Jic�O��C��'����S�<�'�)�����ɝ�"�t�G}8����nQ���٩@��cc��"abE<���`pL�9&��+,B́�	ZK؞���Twč#�`Ҧ:���3��+�^���d���Wr��$�'9���S%˻�uMHg��y�q&�%~F�-���yr�=K]�r���m�d�h&c	�JD�d-�D<���g7�8)�`��>N�?��ã;���A�I��0�ҷ�ךZ!��TSB���U#� ���"
8CD�a�d��_50B		�0�4����%c�c���pWER,xJi�g�[�zbN8��ɦy��臦��x�Fɕ������۝*@ʁ;@��ҟTQ��}��ŉ"�8��<��"�1�є�S�)nPY;anO�T�H����N
gQ�,�wds��DY�*�pur�Y�L
��tUP�b
 v�Xˇo�� 2��	���pyJA�+V[bmy�� �!g-�F@�*5%�D�>)�Is��drt��*U\nyi�ϓ!��DM�EP� ����-ѝ2�{P��*-��\��'�ꄩ /�@�Rm�O���HP���q�H/2��[t�'�
)8 �'�(�"���D6����萃 ��Y�HҮ0����O�i4��/�RA1Gۮv����'R�lZU��n��9r��H�)�;�f�4_=��2@
P��8S��b���ee܋x��u��'�&�!���TQʡ�w*�~Fx��r�$�ׁ@�H5T�rs/¯w�Tq8�Q�L��T}~�����Z���`�',N���Aֻn�(��UMD'���^�d�e�'�O�[���"
��=9$K�'��J��H�]���Jɼi��m���.�@4>����[�,��z�R O�m����H��m�=��" K��}2�)3"��[`���ቁZݠ��!��T���*3�?):���-xN�SD�e�(=hvC��r�@�����2Br�@��b0 �I,|X�z�$F	a�"1x����@�DUo��Pwc�����_��Y7܎4
�+��S=Ac<��dԀ �5��5z�!ĥ:����J�5���A���J��`�c@X�0HC�N�W-�\��h����?z�,e��'
��m����&D@��G��/~�dއXРP*DaD=�>Eᒧ���?�%�J�A\��H�|$������J`�`B�ˢ/�&X����.6U��j�P�bL��B��w�Tz@� 7ᛎ!*�Lh��D�t��Q�'�raQ&�X/����l�+>%p��2��id�l�f�!Wm�Mq.�ؖ�'�,p�d�͸o�]��Fv?Uo u�Ph���"4M2E[��	p��PN�vjS@'*D�`cO>as�D�(A��c��T�����U� ���bF��'�<D�U-.˔�!23�"̞+]U��s�&5�x��. *`>|��F�N�>[S�qܓQ��E��O����J>@	MQ�Ę�Mv�h�Re
{���L�0�T����]�'hA�(Ȗ�I�OW�杽xi����4��q�C�L4�lB�	/[���nE��eC�h��6�P��En#M�D��1��&�����rBa:7�D����]q��W�F~�P LW=.�$"^^azR	@1^n�����F?Q�o�*�V)A*�5\{dj�'�r�,E��fi@ �1D�:l�g�'H��J����a�2n�a����{�Kʱ@��R��x".�M��	3T� ��I }��\����`m�i�Gߒ��>	É��Vy�mi�o�K7�D�'��1�� aM<�$�Πf6�y��O�+��	�J����wb�Y(qbT�_�̩��%L�R'�`��'9�Y��h��[�L�K�Y㦑1�Û�by
�%Kv⨌ɕ.Q=��|"�w��c%F��!��b:gۼQ��'�$�i6Fе.Efl�7*�D���ȃdcu���Gy���:0�E��zf�0ғ��4��ӹv\�� ?�^9��I�_v`�3�T"	���uH�4D<Ba2�]�y��%�Y��};cՐ$!a}��ŤF�x����?X�t`3�ʹ��'`�Di ؈L�����̚z��ِT�U�4F�BA�5�4Ȁ�m���	r.��y�j9HX�)����Z4u�!���k���$圀y��\�U�Sx|��*1ʧ�y��
;�7M)tC̑��(l�!�$����E��,_7;Z�P�!j��%i�
]
��iS��D��6�O��QEzbmOFaq �Z�y2�j��ߒ�0>���?��l��.�*�m�&Y��TK�\!~^$�B)R�=Վe��{���㗅�oH�E��'ޡJ!&�Dy"B
z�����nM�Y³瞠K �3\�$�#+�R�<EJt��&E�B䉖��!"�.Ua��8��c��T�O�(�Q#���XxY��I��3� �QM9:a��S��
�!�D�w�(������z.��g��A���!_@�����y��E�D���#��,�A��C�V�@%ˍ�r�t�ƓD�l��J��zl�`�İ+�$h�*֣o�L�.���D�
�ET�9��X��|	����y#�|���/�h9�d��{%�`j$Eޑ%���E��3 N�[4Æ5!X�R
�'g�eq�䝹S�^Q�����o�pqL>��O��j�PA&�E΁%�)��i�:�+wFˈ-��DA�M J!򄐷F�^��䞥� H��FP27(ۢx(��c���I���	I���e���ȅ�)\�PW�D6!�[�3��u��
�)v����ܿ$���o�+����Ɏ�r���D�Z��Xw/W�2�:�ܫ	��z�C��M��,W��,S|f��U��+h�F|8�X'i�r�c��J���xHV	�*Uc��&0��U��Ć�HO2(2�+E�`�$�!����A��]Z0@�(���(Uk�#�y"``pJ�`"U-z��R�`l��bw^4��bцW/�S��M#2J�hS��A�?_���q��A�<��M��xh:�e�#%PIG�x}��S�*�4i� �zx����F�B��,�����1��]��;�O8����6[|����!n���SNT�	��)��+^���x�B.�p�H�-W�.y� �����hO�H�� K!^4"|Z'ꀚ+%�`��B�v��YG��R�<� v1p��a .�q���8��u"!3O:�&��Ǹ������2	�i~t���L��1w�q��"Oz�S�iI"X�2�y�� +��H "O�ӊFW�+M[iMri�
r�<�r�M,#9�0�N�~/L	�/^m�<1��F����ǎd���q� �h�<����'-����ţ�3�@D�ÅH�<�2ȉ]d.i!Ȗ��&��r�<�)��r��=c�^��A�n�<Q�I�9D(ysĕ6�\��/�}�<Q6�H;)ֈ4��ݬ7#����ePg�<Q���	�⵸���c
�KR�CO�<�d_�6���	w�[�4�|�W�C�<�P
\�n��L����C�Mz�<y����, $ ��ꋠt누�0`:D���� �Yuؼ)���?h�R�4D�8ӷ��6?60XH�*?	���T-5D����J�!�:XQ�"E�>���?D���F�#@��������,���0D�cF�dֈ��&�٩R"���U�1D�d:smX[j��P�+��	R4�8D�h� 哄kƄ@���[�%D�*$�� dK0�#���kK�Ah�� D���Gg6}2���G`��=��b�N5D���Ga���r�Μ�ȁS�K,D��BFD�>��xYTm�� U�� c-D��2��I�$�8��Y7{��J&*(D�d�ao�'[r,;7b9,H��*&D�Xa���3�T���I�`�$�"D��ㆧ��*\����9 d�y�6`#D�pq���:e�a�h��Dl�hC�* D�����-�����>n�T��%D�`KP,�+�f��1N�+2�)T	5D��Ad ��%/ȵ"���hm�Y5!�@�h2����	,pRiSW*'"�!���C�(1�DN0xX�!C�)���!�$�<�L`s#AÞ/k�2FCm:!�d�1*�p��GV�2��6�MC!���&����Ά�V�l�HU�EIO!�Dԗ	��#!e�a��`j5!.	&!��H���GJ%yz�<IR��	5J!�$%�JQ"S6A�0AF!�d��FC0���ŝ�a$,TA�! o�!򤟩X��EM( ��c�Ax�!�D�&.TX�׬��j~���eW�1�!�D��6�HY�.�3f�R�!�0�!�$_( B�BvlGl2�z�aH��Py�,��#��đ�Ѝ���:�߾�y�� wTdpv	�
+DÇ�	�yE.˨�f�)bQ�EDJ��y�@ʞ1h����I$+�0�X5jR��y"��Y�*%@wL��$����'1�yr�N��E��D�.Y0YJ�NC4�yR�Cwb	�ŗ�h�đU���y�,�'ō}�O�~���e����y��*@��Ռ�w�AIEEU.�yi��U0���h� )jE�7�y�/ϒGQh8��ĉe u��H��yr띧?_2)	�mƟYk e����?��e��b��M>E���ʺF��M�.�2)���(ԇ$A!򤔢��)r%j��`ـQ�B�t���+PϞ�V,��!�y�J�>-�M��
�ݾ�����p>�"`ƭ*�$�dgZ2�ۅW@ ���
�v�C�'$-(���  �6��$[b�v�@��$�W0xv��"�2c?� H�P�-L�D>n ����1@�hȋ'"OC��D8J�r�x`-�\-r,��$ܹF;Z�Ä�ƈ�e�����@��av93�������@��y���L��q��M�-��q�ǟ>�~b-�j�rip`�L<�ayr%�jx0��djڔ��C"f̌�p>�W�	�7?Flifځ&8���%�k�&F�	�'��qb�04�؝�kG)�4y��N�D��YX�"�27��c?��I_�)�"��fQM��@i-D�`1`㐼D=\�9��C�|H ��ih��HG
?�z,3rX�"~�Ƀ-��V*�&%@�9�1�' �ҥH�$)�L �A�� ���O�-i!�B(_��	ϓ�􁣀@юh��x*��	�`�ɇ�I�b��� _8��:S���E�(�g"��/sT�ȓ~'����D�J����P$�
��ф�7��c�׺g?����\�>vp=��t�yF��Z� ��W��But��ȓ1A~1���ҟ{��P�ud 7�X�ȓC�Q�C�	3>&l�E��.6��$�����+���y�l ����,v����ȓ��Y���I��K��ؤ77�Їȓ�n���hQ�#&R��Q��[�5�ȓh��л��@S�$:�d�]�(��ȓ3��l�jF��G�]�� ,�ȓ9��h5�'#�yJe ��R }�ȓ^��3�{c"��a'�&t�ȓr((�:��	-6t�\h�oF =�L,��v�ȍ!"DS��kW��C�.�fl� Z��pC��^�u�P��0�.��bGƔ/��,�5@@����ȓ;
p���+G=�$�7t�l��ȓL�<8���P�k�2}��1H����ȓG�bH��Ú@�x`0M^�[�b4��i�<���!��*2%`�
�3*��Շȓ��-+5s��(���IG(L��.�u�
�=" �JBMV�#�����hD\Y�I(a��Y��
ĄȓY֌�W(�Km´	�%M�մ����!�$)UBF�C)�9I��#D���*V+C�vh�B�9/�m�p�՛k�f�"L'�O�$	���x��)RbE�x�&�3��'�9�ЂB�d��	:h!޵��hN|�HX���S�NC�I������	D.��D�y)EY�DӢ�E"zw%h�eT�y�D������r+�p؎(a Ɔ8cƘH	��'ǈ!�BH��uUn��!\�ƅs�ʐ#��ȩ�P�k��`I���3-�c�g�d��?�	)G
�� H��80F̓ixQ�8�֧[ 8�9W�������E�r�F�D`���#�*�����P(��>�U�@�^|�x� ��X.�׉Q^�̪e�5耤O�����%��y���M38Ѳ����s���k~B䉟�t�p�ȝ���8�+TV|$�	�G��8%$�[�z��Sa�K� �F�����둇;̜$�A)
�`^
��%*ÖIQ�� �>���c�G"H�HA�.;^��4���ߨ9�p,�O��Yց<�3}��F<��褎�8c?<���E��(OX`g`G:�
���'�L{���?�@�~&�q��Ύ'qz�얌<���Y��a}MH.B)�	�����N4	�T�޷Gр�B�6����'d�mSD�H/C(��ÊL>�D6��P�8l!#Aٰ9�,�S���=�y���H"AS#
R�'HF8;���g}�0�T�55�,9C��32�@x�O���!u�'&�����<y��Y9�l�6	�p�\��hj8��S�^�4�� �$"�<*���s@+��}z��p���>���h��Qg؞�9�l�� �X��i�&a�tJ1�=ʓ���YP�.%��$çb�l=*�hݞ�uG���o���íS4x�:%��?�y�KGʬ�#�#ۼ}%��˴��>��$IL=d7�����M�$(�ˏ�DϨ�?�|Ȧ(���E�D���J��]�!��ҠTΈ�rn!5�Z�
�3$�$5g�*�)2�� /��؟�|�1�������H�;v��(��Q�$���WrP� �E�ǀ �1��>�E�tK�� ������' ɫ�@�N�l��j(<O���ĭ��$�!�,�� ���s��;v����m҉%~�lԙ���C��N�Qe�ĔId��l-d)̐P"�PP�� AE��[�fB���%�(�b����<��@��V�v��S�'TH����B�j��s�\�[`��O���jCNf^e��nR:\���=Op���Ӽv���H���p!?[�$��f��%��y:R�X����Eh��i�D�qrJݦ!w�˧	$��R�G�|���st�A$�҂w=dDـIY,��ʓJ	��a�çf���
ç\�m�bM�'{����cJ �$l�a^��?���X�<�|H8@�W���d�0]�ͳ���!�bA+e��$o0�Y(��>)U�Z+~�2Q�I~�C������͕;i0)�Q��8�0L"慿>�8ŀF�m��ۓu�`b�"��}2����MV*d_X����i׉)�D�$����N�]��|�@��|� e�m}��B `�9���
D�'�	4��:������K����e�,pdHȖ
B�+s#���y"��%�x�`���25;�$��S�t���Z���,�Խ�d��i��Jj�27ƒ]6���r��e�OV^�!U�K�V�B'��Qeࠥ��Pg�)/wņ])%f���቙|82A��b��:�p��1��~L��GcҥI*�Dǫ������5�Y���j��bHp��ɐg�\%R��&9;�q�b��,I��5lO��� ��1"l4��թY�"�tx@�Ʉ6���9Y���B�|�F�9X���12�����H�Obİ��S4CTn���L&(a��
�}���"��>cl*i1� ���Ir�GRZ� �?����(�Y=��1�.(�~Y)�A;"pьܢ{��U)@�>��9G��Ӓ��)�Q?��s�͜k���u�ڠ���cgc�?�qO����3?91�M�
{�}v+�(%��Bo؆?����g8}������gX`����<��Iå
Ҍ�U(ܦQ���㬓@�<))$@���:��ǝ3TN��q�K��~`Rd�^(`Ir�e9��`Kz�>�A��վH�8T��)h�`հaJ&LO(p{�fԵ}�`�8�'b<���\0�k�O� �t� ��P;H���ES<���0b ʦ����$&d�r}����	=.�l�����DrqO���h#;�2O�d���i���)zu@��&�N�&���67������k�����>A�(!�oѮ6@d�¦V�Pf��7d�R�	������'���&�	/Z��� �A̼s$Đ�M*5�JpzP�ᦅK�<#��5d-ށPӅL�zL��{���,3d�pv✉7Z�t��]��(�2�S����^���z�Fd�Gg��[�bC�	�E�ع�@�D9E��-@��A(	��;d,���R�3�-��w! �� ���ܭو�$
"N T���aa�
�y�O���{�P�R�*����#J
R�P#PK��ô��Yݞ�I�d�-9����X�ĩ���?�̭б���4���g�+�I!��L�eB�"z�c�#N<Oe��_?a)�Cǥ�:��&�[]��i4�&D�T� �S��L�c� V�*��ip2.S4

(	0�:
h��"�:E���is�Œ#K[g����e̴�[�2D��!��u�=X�R�"jjBvf+�x�zg�V�*�"��֡faH�).�HO6���+�������&�����F}�D����?��CD�<; 		�x>"���A#??L��ヒ��>AS�5"aZy˳�_�C/:��	�f�'�taRs�F��|��'�@(6��Y?u� ��R����2��v?�ց0D�@�1lΑU��Ih��/���g�3���.�
�����ȟm��7	�`%�'+�	E�t٪�"ON9��&ބ�Rc�V��>A�o��v�{�ȩ�yH�q���M�Rh�#oź;�@'l�E��N>	Ђ�,��!XwI?G^��ٶ"��¨^w�\�{ӓ$���F5N��Q�Ǉ'>>��牵I��1&�%80�p�.<l,B��T _��l�H���b���'��PQ�nU�/fD�ѩ�'<®�"H>��i�%9Ⱥ���� �F=٢�)�'5Y���W9r����P!�d�6B����QlP#��C%L91�To�@I!�`��[ H$�3}嚐r�P���$^+��Z���y�P�G���8Oہ�)��"��p��P�la��- Q�_#H,�y��\�<����N;�
p4�\-�p=�3�N��b�Zw��@	��W�a;<�xW���>�(O�Th<���W�|�Xā[
~���TkS~�'���ڂ���b9~$�J3D�vְ��6�YcK<\)�u�<Y�F�+T��3dܛb$���j��[�
�w�x�Ss�>E�ܴG(��b��`�P�韒n�ȓr~b8r� Cl��0{��>nhȇY�l�㍓c�$H�Q��� ���O�8)�b�@�+ƣG^r��R�'���E�=C���낉����Q�D���J��)��zh<�a����L�R�J�hj4�hեTf�'�f�s��>m+3L5jF�9D�{�D8��D%D��h���) �U�7��	�b���kb����ޅ{"qO?%S5�E?IZ�kV����>���
>D��DͭL�N�uJ�B<$�q�1D�TQAJ*<��C�	h��P2m.D����'>O��c	��t��iQ��*D�l��$�/׺@�a$�V4�Ix��(D��#rɋg1�H��.���I��;D�A��6h���c��:�da��3D��JQl��]�1a��)8r�z@"D�YRR�s}�eĥ%JE+B'5D��#c�V�.����(N�P�D1D�|˔H� c&���ALƂq�@���,D�tJ��U!��ҡDƖH�F�i"�)D�ȡp�ۙv����pnF,PA,�t�'D���RlԂi��3�3GS�H: 6D�L���*�8���O�h���*D�HA�0nY�cI�E5zR�(D��BЍ�	L8QJşc�܀�`)D��xr�ܟlä���E�fp�<sdo0D���,x������5	Rb�$�/D�H���R9H�ՠSG�2xG0QЕ�6D�$�휢�jHą�a@
ՙQJ+D��j��H�Ҙb��R�ML���.'D��ǦؾB����%O���${�j$D������/�R\�eK�b��TY��$D���D$��8~�D�b�z�D�8D����� L��{�j�)�n1˥,5D�$â�� 9��+1�O��z�Cg�2D����!ܖ�ՐӣF+b%��L.D�R"��%)��#Q�;Jƒe��`#"�4�)b��Oڴ�t��4*�Y�P�|ڴ�®�.|��,�(�T�'˒�[�.����:�u��jm?�� E[8�;'�A�Q�B�C�C�,�J#<I�%i>�x�@ZX�TSD$�oo�����3�I4on��<%?�!��qR��Xt�ޔQ�x�Q1K1}���}���O�H�i�$�~\�p{7!YoL��'h
��r��;	Ȑ��<E�t�TH�l�B�c�v��m�*�y�d�6,�'7��B���5��@�5}����ŦQ�����]fE�V��b]8с�+}iL�[t�f����D�"s	�ɦO�<� ����9<�a�L�^7n�I �&�� ��Ӈ<�����HVX�Ms�DƎ4.|�3�O9�f㞢�AE�Un���/��*�*��a.;UV�X�yrN{�'
.r�'4�<���_�.��y���I�6(KK�@���?��iXçm��I��͉i�E�Ӯ��S�&��'iLH��
v|6��<��!�4�D+�}V �"2���S�E;QiP�A����O>E�$BĿU7�i����S��s�	�0#F���lȔ�(���?ͪ�MR5AQ ��Ǆ��.�j=�v�,Z�&QL>�f/+��Y��ʧ>�$8Y�E�h�~�!��\)*��]�sZ�󑦜�s��@�f�Ok�\���V+t��9��G��Dx�'�X��YX��9�T��>Ap�i��s���.r�H�E\:.�z�BdѺW:�*�� D_ơ��G��"~R_wǺ�*D��Sb�Ȣc	Z\�a�/Be��� �,;T�(��U0�0|���X�J{���Ł���aF�$;?�Q��gρ8Z\� ��f�<M���f�R����3Ͳ�����0Pub���o8~:�[�8��tc#5�d���a��4�p|�ԢT��P�2|6)��yҧ�J�t%�g>�r�̕�/Yz���G�+S�@#K��<񂅇>-}V�: K$1�����6�"M��I�4$��)��Yd!�ǪX<P9���Px�P	!�N�R^!��8b�D����C'���	g͋<8T!��\/^9yb,9R��l�$kS?x@!�$��)[�ȧ�ݮA�����C�-!�d�c�Bբ�e�]h�i�7ʚ	�!�� ZؚG}p�ӣ/ߪ��YA"O$Zӂ�%F� y�ԩc}� ��"O�4��%�|Oh�&Nrv�"O<PF�3_2�y�,)�`�F"O�="Tn�"�>���lW+X�Nd�&"O��ơcR���$"ؘ9��"O�dR�Ǖ:Nԁ�d́v΢a��"O*L�K�:��x ����B���C%"O����X;;ID-�V"��q�@���"O������WD�Kg�ī-�܄ "O�D�V�T`6D�%1� �f"O���G_B	�uEI�8����"O��Õ#S�g�D���B��BL��(�"O��#N���iՠX�8[�"O�t����?˾�yw���J�r�3�"OZTh�h%T�i�G$��1���r"O���d+RN�p�T+j�
�ps"O&|ȳAċQ����� 1h�D\c5"Onae."�\Pe�$yhH�G"O�q�!aڵd���P$Y�Y4��"Ob��QÃ	�ȥ"K�>�t5�"O�����!�<�1B-���j4�"O���
 �s��k��_�L��$"O�<g�(@05�qʟ�7�]J"O0���� �KG�� ۰���"O���@Ɯ@�Z��ȑ"zY��"OF�;�*T�xF6E����+�0	i�"O�5
�^h��(+"���S��ID"O�b7�#]�ʄ�I[2�� �C"O�}�#�@�8Q2x S(�.� �j�"O������T����Y�:�{e"O��z���+
�Ps�N�+=Y$���"O&i@�LH!+)����LƉrGZ<�2"O,;#��"�m����R�(�"O�Y�6��#2�0��jθ-����"OV-��(�?$��:���8��\��"OY����^V4��#:pV�0�"O��uOVON�$��D_�YR"O6�xe��;l��̰���Up�Ő�"OH0���:z >X�#�n��|H7"OD�׏�:�ԕ�֥Q�z��A�t"O����˄?3 �@�C��R��2�"O�j��!g��%�S�R���J"O.h�)�'Kc�$���S�!�Լ��"OLH�4(Ĵ+{tP�B�t�J�a"O�y�����
v�!R�H:o�ԋR"O, �
W�3��P��%q�D���"O^��4���w�8�#��^Ɋ{R"OD)������!��J�k�T$��"O潒g
,�Z��2��^E�HX�"O�X[�k® ' �PB:K?��D"O~,�aU8\]n��'�Q#H�s�"O6��S���g���v��"Qx�"O�ЀҠݲ$I���℣^b1��"O^�Y��J20��0���kRd�"G"O2u(uA36S��H֧K�6(��(C"Oy�p���@b�%�(a����"O�JŦG'/s&�j�4Q��j�"OTH�Q���o������M�d}�R"O
,ʐ�Ղ��R�<FT���"OD���܉c�d�i2�OJtIiU"O>��b@J�g�MR�������"ODx'� -��H���2�H���"O��[� 5C�F�Wg)o��P�"O� had�K�<hJǆړ��Y�"O$ݐP��*�! ��$���"O��c�N�N<Re
��/���S"O�mp'��J��P ���eɔ"OD򧎏�3�xӀ��
z�^]Y�"O�D9����N�x���0c���:�"O�� ��8DvDqs�U�2�4\��"O�����^�bK��M3X��ى�"O�(�"J��x��c�y��S"O��@h 5���XPL�/)�h��"O���CG^?5u�)J2,�z&\��"O����IP< &ȥ���M�d9J�j�"O����&�(!��M
C�W�L�C"O�]!׮͉ Sd};b
�&�T|��"O����
�	On@�$gN1E��I�6"O�	K�Lоs��"#�K����8C"O�0��^4^�ĥ9�.�X��"OZ=��!S|F�)��"di�c�P�<1t�
�J�8\;���J����VD�<)�E+Q�� ED�1p��y�FHz�<!��~xV���nN�z�QA��s�<!@/ޯht���Ū^f�9�EK�<aWD �C~N��㘪KPN���*�O�<�1G��S�,9# V)Z��$�F_v�<єXo�0@*R��$u���9��l�<��X2ShQ�Cg_(cr�9	�e`�<���Q����zVd��M��(���[�<�+P�t�<��(�#aȵ8l]P�<	0)N�"4�M`lZ<D�i`��_O�<�`l��(l	p����;;�H��H�<у�%v�f���Ċ��X��Lj�<)��$o[�	�@�J�T(@�H4�JO�<I��]j<8�eT7,�dUg�J�<�#�#1��E��*SF����a�<)dɝ(cVaȀ����IX�'�B�<� %A.J�<Y��Τ@RJ]�+MW�<	��S��`8��j�.U� �`��V�<1fFJ�NV*iJW ��}�R�&MMY�<�a @���=[#Z�lG�mpG��~�<f�JT�<��7J�4tBp���~�<5h�x�r�Y��R3[�x���|�<�# �6��)���[a�p|+�N�u�<�֮ܶU�P� oL�`�cR��H�<���y$�mR���A���b&�n�<I�==C myr���v��@���i�<�D͉�n0�T+e�ڎ\�޵�-Ja�<�GӤ{&���(��:$��`��d�<	P��.$�� REb)�t�cCy�<�Č �H��	�&/��ŗr�<y!��?��ݩ����,�Nq�Nm�<�TP�$���87F
 _P�"&k@_�<Y���6Uˌ�Y�kX�U%زt�f�<�5H��I���u�ŗc"4<� �e�<�&�ޯE\��(�L��j��4hW�f�<�T�W��X�F��%L�[�h�<y�J[�@� ��N�-'~\�k��d�<�4�;]��C%�Д�&�i�<����BY0�@(����2��J�<�����$"�K�=X�z�^�<�����a�����
6Ȍ��g�c�<��@�S�"�����
�aڤ��[�<iHU�Z?��C�C&��2�m�<I�ECj�����>c��\��ˊc�<���v�h�`���+pR|H0$\j�<� ڄ	a�کx�ֹ�����T��"O�9�cÖ6�d�D��l0���"O�Q�����S��S�K�3t^ؙ�"O*�v�9%
.H��Y$\��qX�"O��۴��	iKZ]
4lQ/� �3"O> ����iD��0��5n��a�"Ox$��搈[h�!��)gc���"O��I�J�0��L��C�5R�xa�"O��{r�����g�΃UV�"Ol���N^'l��aA8_*ؠ��"O:����Ҍ��]x���<!PA�#"OL%k��8�H�IW�
u�u�%"ORd��PVdF��@N�f��*�"O\� ���;H�MP&M^.`�3p"O��t+�^��p􁍏B ���"O��R7�������\^�!�"O�M�	DƆq��L�),^)"E"O���L@-k2��)Bg�;c$�0`"OfM�!�ʿ�L��v�Wm�Me"O8�1wGC�	>B� &˛%�	�#"O8�94� �MZ^ѣd��(kU"O>ab�K3���K�c�r�Z�bp"O��J��&�2h�3#@�=�.�)%"O<	Ҕ�_�e��Q��ݥ~�^�h"O��4/��c�ͬ�2�H"O6͛E	Q:T��9�Vǔ��pL`�"OrԚ�.Utd�g��|�y)"O�i3B�Ї[܃�c�!D�eB�"O<|y!�C�	0����9Jo1��"On��AYP�>� �Ѱ6j��r"O�I���M�|5�fJV�[[>���"O�+\�L9��'`�`8��>3�!�$��	|��CCD��n�D4�3Mؒs!�dA��T�����	B����î��d!�d�M������u�plHҍA�M�!�U2��z��$qU��C���YQ!�D@M�*@3c�3ss��
���	Q�!�DL�)^F���B8b��z��T7{!��B��>E2�D���z�C͗�!�DX�[p�䡞7*�>1��ᕋv!�$�c�]�ˢtz�	��O�!�䌚6
P�ꇌ]����*�:o�!�E�e�B�C]��)`�p�Qt"Oi��O[�
���ɱ��cU�(8a"O�`p�[=�~��p�L�MLt9��"OX�r5̐�h�}��,T""�s�"Ol� �j�5�.\�U��)�A�A"Ole(eG��|`-��đZ�T"Ox�Q��d�r�a��F��-�T"O�J��F�D"쟈x�p���"O�`C�#e�2v���(m�!�d��BD�*#\�\��p��f�!��(gm���w`�B���K��U��!�F<ڧ ���a�����!�X6r�x����� �^���͚4�!��_�@ �n'8�88� ҹ{{!�6rP���_\�� ���S0y!��Oy|��ш	���da�C�_!�D%?U�)�P�L�V�S��ZW!��%�@D`���ej���s�Z�%q!�K!�N $�#d��[��L�<�!�$��q8.��c����ڄ"ˁp�!�0���X���6���OJ�t!��KJ    ��     �  �  S  #*  �2  �:  �@  6G  �M  �S  Z  R`  �f  �l  s  _y  �  ޅ  "�  f�  ��  �  7�  ��  ޱ  +�  �  a�  ��  ��  ��  ��  "�  c�  3�   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p Gx*=�S����l
��P/��9�W�&�y�  BMV@���B���( (ў"~Γ8��u���E ����Ϗ<��\��I͟t��n�Pj��{�iP�)fɔ�8A�=D��k�`O0XN}�Q�G�&5g:D�T;2�	��V'Y(&�
%i!O8D��x��Z!�x-2e�[uĔ�37D�Xq��ڍp7����֏Z�d�5D�h 'j�4I��T� ��0.���=D���I�'�(	 aoX� �ܙ��;��ȟ���fFM���u#��N*:� h� "O�1�P��-M����D��,�@� �R�xG{��Ƀ�
���&N�h2��V��r#!�d]=�� !��J!fw��2�mD�!�$�<X�EP"T�Φ@�� �!�Ă�Y_NؚFK��p�aj "/!�$˗�p�勁�h�PQ#g�%�z"�DU�|}�5IR �T�kU&U��_y��|ʟ�'�ࠐU���l�����J� '�긐��N5c�t(맮;�d�l�? б`�mL6p��*D��zM��"�|b�'P$�Z?@��ҕ�F�3�2�RM��i�e��0���s?�'��)a>Yӄ,)pa��`��ߔZlܐ"�E4�O��	�+9�@I3~��C�˟�b�|�⋓6�p<�B��	k�αhp���q��9�"l�PDxr��(�P H//]���Dɑ�<^D�E�O|�=E���/!Z��/�~t(�M��P�@��'��R��N4|���ըGM3�5p�'p�(:B	�.o^���H�>`F�:�'�FU�d�b�E�-Mk���	�'���ҡ�� �)�E؈niʭ�'�H@& �
�� �+�2}�n�)
�'^jP�R
Z���e+� r�	�'�(0����	H����N��$�"����O\�~��&�9eݞ	�U&E[�^XPf��I�<a0-�%i�ĭ�"�����c�G�<���-k䔤�W�TZh��ÎL�<j��0�\C��ي:�^m� ��F~��'�N�B���MW:P�` �m�T��'窠i6��)$JPD�a���W���'6���ˏV��<�P�R0R�ȳ�'	JU�#C�~�t5��eԢ4��
�'�d��t��si,uB�G+�@M 	�'�^ V-NY�p�!ڨe
�'��x0��ynl�9�H&f�����'�9�)�.2,st(�[N�	�'��!��ŉ��z��(T�l��']XE�2���>�����ѝJ��
�'8��r)H�1�L��A	̛=˖�P�'�~|a�i�;�Tݒ�F7�.��
�'��]YR)M�{�yd$06��	�'@�RH�O��A�ヂxP �
�'���i˼I�]�`�I�XK�'I�:3L]�KiV8����$٢�'���!D ��DA�4'H�t|�q9�'��9sw�ȟC[Љ�Ao�	�2�'���&�	�8�Fa֤wmy�'|ԅ�Q
҈2��t���&)`d��'���`蘍'�&�Rp�3�t�3�'@��!�1 @��R��<���'.���i�"��&k�� ����'��A�
��;�n�:�#\�*��}�
�'Z�ҷE�+7; A��%Ժ�S
�'n`����TxثU-�g����'~PՑ���R:�sF,�W�@���'����o�+J�}k���9R�6u�'�~��q
^8Y�4`��I�2p��'1���/���ݚ�$�;>�\��
�'���Sv�м1/T1��$1H��Ey	�'rDX`�-ȸ-@$��7(�p���'��C�F�25�ǂ�V$q)	�'��<��J�=^�A��K9���J	�'��x�g_>oL	�ᓂE�h,p�'��l�@�S�
J"5J���*iIĭ��'����bEH�, �I�n�R,��'|�M�«U�Sa)���;=���' 
l*�Ӂ{P��KVዦ4�=��'� �s�W�m18#h	�4��9�'���
S��,C���nW�=���*
�'�b�1Rc�+��Y�B'�(:]���	�':�SC�;�tTj�o[?2ؼ��'5�1WC޴<�'��&;�lJ�'z*9�d"��Cߨ
��D�:*ȑ�'�$�S��<* �(Ʈ�=&������ x�Q+B�+n` �X�kj�"O�܁��@=tM򍸀��RU�Е"OlHq�Ǥw�����/7R��3"O8�(p�� s���t�D�j3Z@ô"OX�ۂeǝy;d2 #A"=(ZU��"O1���ؘ��L�U�/f!(�+"OԠyǩ�E���Y�nJ7�u��"O�P���i�	�S-��>�FL��"O*;6g$)jVI����5!�~�s�"O��Ҥ���5l��T�ѰvC�܁"O�I�#	g��åZ2-(��b"O��"NքD�P,C���6#JqSU"O�`J5L��2��񣥢c�)��١�y��6^.�U�����p��B��y2(�+V�XU��l�+R�NDR0H؊�y2��jS��@BW,y�X H�G	�y���a�(`�3'Ŗv20�` F��y��F�(Մx�%�όbz义�nS��y�D�q��i+���a�AO˼�yB�RB�"B�
*���xaM��yr X6����o�AT�;��ybjV�Sh��;w��E�|��o^��yR�ڢB�t���M^�hs�Y��K(�y� C�"HHd̜<g����?�yb+�
hP��ٶ�� Zv�$!S鍁�y�/�{q8��Z1E85�ˤcuTC�I�j���2�m'%�����J�5"C䉓&V$Ț�B�m@5���	4XD8B�ɥZ��0��ʕ%� iQ�4[�RB�;w"`8�!�&��C��j��B�ɋ9z��(s.�?Q!�8�dkPW�B�+wm��Z$�0vv,�C��]�B�I'2zY�$M[/S��P�+�2�rC�	0#�i�iI,}��Y �i�,C�I�S�^h�� G�V��m��F&M�VB�?Ia�����,F�y���lorB�	*V�e3Ta��� @����m�ZB�	:M)�m���_!:J0�
DN��W�C� �����$9�1j��ȕ$]<B�I<Af�\9��'%
 ��o�8n�B�I?{����O�5��,��mW"TR<B�ɷ|��딂K>P�>ug�{A0B��m����NFo�J�`Eڑ8B�I� [�0��KY����%�f�B�	�MF���ˡN^����.��B�ɸ02����\�@q�DO:U�4B�f��$�.ӫ{Itŀ!��?VNC�I�kj`���#"}49Sб	�^C�	+���#j�i�$�1��Q3b�tC�IU� �[&�V-/�����
8�8C�I<%v�%�E)$\���ᣁ-\��B�ɜ���7h��O��)��80ɞB�I�I���׊�!CR���!E �B�f�)�e��>h��u��ErB�I�H=���I��_�Z�R��OOjB�ɪw�+ �I�?�����{�C�'�$���Ӛ7�ʔI���2�VC�I ��4*D�)5?��kge�0�>C䉧k�d^j��B���P_f�@4"Of���MQ��Y��VSCZ�"O"�ƦA�A�x8��"ҚU�v�F"O8��3F�ft4Rro��n��"O�I��OOi�U�B+B��<��"O~p2Q�ɃNʤ�{�f߼~��B"O� �l�t�C�!β���Ŋ�^�"�9D"O\�!���1׈�1e.� ye��&"O8��[�O�,p�&���g,�9z""OT$ۦ%_.u���0O֫V$�@��"O�6
E�/��S�d�L�2��'�b�'	�'vB�'o"�'3��'���h[�J"ɢ֡;(��Գ�'�b�'J��'n��'b�'�B�'��QQR�� @1P��W ��{u�����'��'��'a�'8��'*��'�h�qt"�PV��'�ҽh�)�Q�'!��'�b�'N��'>2�'wb�' ���q�^�*��q�X�?6<�6�'eb�'�b�'-��'��'y��'P��Q�q����K�P�^M;V�'/"�'���'"��'9��'���'!�s�H
q����쟚4{(��'R�'���'�r�'���'q��'\D����eQ<Pz��#E��b��'���'j��'B�'Gr�'�"�'�pi����2/�F倅���3l�8+2�'D�'#��'��'��'f��'Jr��'kDF6ΝYs ��:��6�'���'�'���' �'���'�N��]�f<X�·�_4f��P��'v�'���'M2�'
��'��'x��˓a_��|`Â�ش:�����'"�'���'�2�'���'�r�'����g�<P�N0Z��ͼT���'���'���'���'JL6��O��DM5:b��晊wi�$k�%8H�vЕ'+�\�b>�M�V�L�/�X�
"������Wl��Uʠ��O�dlq��|ΓJd�v�&l��y`ï�Da	��J���7��O�8�snӖ�O�|�!T�Z�3�&�O2&d�B�;!���Ξ4RZ��҈y��'[�IJ�Oi�}�F1y��0j��H�XuX��Ӹ��d�-����Mϻ>:j;�����=�WD�i�P뵳i��7�f�է�Ow$�I��iC�D�5U�l�0�W�HDeb�S�Y�ӺQ<��; �ԧN�<�=ͧ�?�Saܰc���+b&Rca/	��qy��|�~��aV��'Q1<%S�o����T,�/kj���O� oڔ�M�'���4p&"�h�,ڑTd�F��d���6�� �j����|±��u�o�O�wF��@�i oC�f�w.�<	)Od��s������N����H�o�
 �Ly���ݴC ��'D7&�i>�!��ټc@�8: #�4���w�t��0�4'�f�'��P2t�iX�	4y��׉ql�m�Sl�P(�	�U&��~E^�2�
���|�.O��$����8�����/�*7��� �JΓF*���&"B
Ӳ ���c�SШ��� S�$�.m#!�J�7B�9��ٺ�*ch�;&�����G��;qT-

���C�
\X)�\�0�B�'�rL���sG��H[�����.>n��@F�&C��iu�Y�%`\�"$�R,N����M�JC���-
�L�͋�%Q�(4Bף�.o�.]m���@��ğ$����� �yV��v$���S��D�f=�&�'�hTr��O��9}r��0=f��RD�r���
ۿ�M Ll^���'z��'���+���O������]��S�@� �j��"JƦ��E�D���$�"|��	(Tx#�ڍT�FH�%C���ǿiq��'��'<�Or�d�O<�I�*���*VN.tQ����]����?�����/Oh�d�O����Õ���$�Ty&+ʩ � IU�}���ƻ9�˓'�����<�W-�@��BnH���	hJ39��6Y7 ă��2?I��?q��?��~0� )!B 1��hb��D:@��F�O����<	�����?����sÈ
�'q� Ѣ� �`|H�JѰHsV=�'	��'���'%��	ki�!""� ���(--TL�5@�>v}�6��O����O&�O����ONxSN�/<�����=8d�H'�5Q��$	G���$�O����O����O�80í�O�$�O���u�ݍi
���'��T���ŎȦ5��V�I�0����Ֆ`����~- 7K�P�l�)P��#ɺl����My�YW�����^-��-��,�좗+֌bs6�!0-v�	�h�ɠ^S�#<�OКE�C��l�:ux�8b����4�?	�4謵����?���?��'�?a��;`��?^�Ҝ�t�K�Ѽź�*��U�	ڟ�)�U'Ȭb�b?-��Bɗ f�`���b�� CxӶ4JB��Ob��<9����d�<1��K'Ŗ�P�0X
-����l�&�5�E�y��)�O�b�EN��Yu�]Y��U�RC ��	�	���;)@@@�����O��O�������LrP�ʠ�&;o��HOVt̓fD�����T�'���'���O[�(�p��k����*�I�����5�x��'�B�|Zc`T8����VHF��S���,ߴ�?�����$�O(���O���?�ajT,��q�T<AT����B��
1@+O���OL��?�	_y2�V�
.V8j�"F5�x4Õ��Ai����Z��d�O����ORʓF�|Y
�=�rT���S�8C =���gt.ժR���	�0�	]y2�'���J���iL0lхc�:,J��E�=����&�.��[1kf�[#��C�Թ��<��O�,�p�ٿUz��Ѥԟ��8��'q`��ޟ��[�h&p��'����G\#G�"Q�c��x�1NM�da�E�t��7���*�JvhD�)��b�6d`
�@$�#J8�]�ꐦ\ޙ�E!�~�����6Z�d�,P8�����u�? J`1�%^�I�����k��,�R�hȊ�p58�G�� Hż`AS�Z���lZ�{�Ͳ Y֟|��͟�Sa��HJ�[���Y{�La�L�<������Ug�a���Ďb�a�O�1�bL�&�$iy���56���gE�j��aaA��I>yY��åV>���%�O����a�B��슷�S1���8��o�����ˮy�:��I�M;���?�M~���?��C�$lz�E��6ځ�b��d;)���?1�eE��sKT	P=X@�~>��<1������;�4�?��D�9v�up�䇵��}���]��?����T�˔����?y���?������O��D��G0�M�QL /�N׎�g�fp����Oofh�P�-d�2�S�ȈZ��	6!� �T�V�ұJ4B�X����F^���Ȗk�0#D���?=���$˒f�0D���'�����Dh�����	
 ��O��ԟ�I̟t�'ל\�hՕ�F��CO�,���X�'DyC5��NϮe`sC6"�^�ⷫ/��|����d�6� nZT ̘FfZ�T���𮑚d���	ğ�����ءBa^Οt��ן���]q� B����I�Ñ�z�8G ���i3n	D@���8I��V���e~ʅ�E�KLصS��.2��	[��^�{x�F/�'J��q�f�޴Q�6&�t�f��O
�D�u[�,Ѡ)��*P�D2�O�|*�H$�,�Iڟ��?�OH��!�ώd��Ѐ�(F1q �"�yRǙ����8ڧB|X���H�?[10\�B���U?|M�E����'�I1PZ9��4�?����I#h����C�*��@8��U�d�Q&�O*���O��XF��O��O��'x^�*a�B�R4J�ᣌH�ZDyR��B;�]#�L2eR
}�ЊK����In�se�I�F܌$��i4�(OpIc��'k)�i�O��0�F� l(��[U�i�b�O&�"~�,`UI�ũzQ<�bw�	�����D*��\�S��|`'ϴZ`ԩ5芳E��``\���3���M����?����"F����?���?�w�:EB�`�D�CN^�k��utTZ��i��'��3W���c��PQ�x)�����C4y5(V�F'L�!�	ژ_��S��?A%+Q.BAX�)GZ�X�/�8T�EH��?iCT��	+��d��&݄~𬨗�i��������<�����>)P: �ŋVc�4|�`�V�<�K>I�i��#}"��!��M֡��f,{�卧h����?���B�=� L��?��?9�U?��	+ aܼ Vȗ�U2T�]� ݦ%s@�~�^d�Qŝ�t��[���?M���E�1OZ��&F�t(l[��+8����<}l�Tx�G�1r���!�
��IO ?f^-����u�u�<�f�cTxCQ�Jq���;��Vßh"!F�矴�I���<9�����<
�5:c`��_�H-[�+�1FQ!�d�O�}(�/B/`�l��c�G��h�DCx�'���'D�	y�jT��4y��EP��ޠ>�H1y�+
�`�*)����?����?)3J�!�?�����χ?�p�+D��Qk�����`����!a0u�BՓm���Ó�Е���߽.�T�H���I�BL�SG��(����pI�CdI�v�ɉ?bx�an�;�YXK>�qn͟�C�4y'��أ���M@� �Av�	�@�izRR�4�	J�S�T�+Oy2�;�͋�^�%A��>�0<�����E�d!K7+&�<IۂN�L��dʍj���$�<yP�J�"6�N�O\���|r�h������R+D�z�F(9��5@���?A��h�,A��OT3b����^�R��|�.�ҵ	W�U�öyr�� �6�d���P�yTO؜�t�{��θ7Uj�@�c�B�4|�&�F>P�5�C  Q)� �m�_<�(&�<���O�-F��o�4j���A"��t�n)P��%�y⯏J��=j��D�"��=���!��|��x��	��y�d�	�����ή�yR�Z?7B6m�O@��|2w� �?���?��Ƈ������
IH�9��,�@.��XFP(Ԭ�'B.[��Q@7 �?��|��K�2�cȩp�^Y�q�,QD���F�]$p���D��,.r�Ŭ�l�v��8`�!�LTQ��;l`9�!E).�a� �/8~"D#���?q��i�6M�Oz"~��5!N����/�Y{�l�a
�F������X���!7J�D��eQ(���` J!g��b������HO����O��!a�Rr�ĘWg׬T�A���Of���6$MN�&J�O����O��d��s��?yG��{%�� �H��|�s��B8E�h���`��iގ��s�èU��\�'3Q����1$�p���)��"�@@8(�ĸ"�)�ސ��!-V9}��ӂ�(Ov����yf����JO�X2D�OK��?���䓍?Y���Ės�"A�_r��i(4IC	�'���Cb�C�H��eC�U��؍x�� ��|:����EfŚl�<���/��r��\`�-�i�<y'��9?��	"!.�=]x2,X���a�<���ػ:{�q�O7l*)�SB�<I���$��}0!"[e����g�<	�� , �ۘ�ԅSc�O|�<��i�k��<�����p� ���	�M�<� ��kgMߞ_��`F�[�>���E"O�D�r(��]W򍳦��%z ���"O�<k�� KD ��eń�Z���ض"Oa��蒢Q�Ƭ�ЦE�e�<(�1"O���� |�`���U��!#t*O��95T�ul�3Db���'Q"����)dX[�J]-�ȑ�'� ##�1VǖR�ļX+&��'�xe�bGQ8m���3�
�H��T`�'��P�ot�<�yDA�9?��'�d-����oo���0$�;2�^;�',��+�ML*-T\�p�R= ��qr�'�2�6hH2}��Z f&pj����'��ă�F��"��(��'��a�ȩ�	�'��$��QvU%R�B�mzjh�
�'�*x�G�T5R�@2Eѳc��R
�'�\�V#_&#�� � +Կ\'|4�
�'s
P�$�)w�Eېh��q+
�'� ��ƗZ���#�#+U��Y�'4��;CKݫl?X�8FF�(�8�{�'���#�O�����b�)�=j �J�'L2�J�f�t�x� �lܼ�ܭ��'���k�(�)I����F�Ӡ|׬���'wn�	R����mӯS�q%vUQ�'آMk��A�L���A�Ɵ ����'#��3�DF�@����]1#�>=�'X&qP�G_Yx�t�&
f�c�G�|E򑍗�>h�d=,O~ Y�ʳ' ��0�w�t���'F"�P䦁zB���.@��{4h�W;��!D�; Z���
O�S�$E
��4ƍ�G�h0�����ZLj�Z�FɳT�|���((��=��I��	��w$�Ru[7Nz�B�	�r���	�'W���*�)M�@ *��a��zvm�	 *�4�g}��P�-�ԴS��(m�D� �C��y�
�>`[T�Q�"m�m�C���MCG��',
4�S���-�H��ǓS�N�3 ��)luy7�Է([J��퉍noƝ�m[�?'�
S��k3B��:#��!뇌�wu<=�_x�����W�a&	܅N�>��>s��n~�S�,�^�����kȖcdJ�p�i�3*�D��l�	�y���=L�<���ƌ"q����k�z����S:1n�*���(���Y�0�%Z���Q`��a�̙DM(�O�1�-�`�P�V���	"�:0�T�$�h��)�\�x�(��CL�H˓����쌃Ga=`u��f�$|E~� %�='����1"�ۭ�M��F�36zr��r��&Y�^���oY9�dB�If��m��j�f�:�[G��3
e��[�5�!�:<�P*�z6]�Sܧ\��X�I���A��SV�)��Z�(�&�)b��E�pAȡy����͘�+`� B�O��w�/��I�K���'�6�Hª	/,Z�y�ԋ:'jʽʋ�$�f<�i;�Brh��+�"_���}Zf��trIK�`E�o���Ḋ%�O���|i$吒�Ѫl_�8	�Q�;���(\Zͩ��fP�e�#a�>��`^-7�1��&�?Is�P�`N�'���h޼k���,��+�l����dΕ�r@wʔ{2�۱���>I�'��% �����%Wʾ9�V$Ќ��Zj	OQ�Xp��x򁕯~��]3gh��
��jv���J�X�����U��(��w��0�s-��

�Š�ꏯ4��������p�'�0D�H߷VE���7GM�N�lԫ��ن%FZ"?)��ݝy�tha�N=O6-3��K˦y��۹}O�Hk������m�<��'D�1p۴^Bl�rf�3zR%���f��d�S�2 XR��S�����.͘Q8�'�� ��G�6��͊�ɐ�� -�����-4�tM�G	B� �^���t��6퉎i(@���;[ pA�b���Q��Y��;kM2�[��Y�:��)x1LҸE�轱�,���0=$m�O�2�ԍR��8zv��)O� F �a��+	� ���3N��;�2D�f�P�m��<�P�ҸCW���ؕ%�5K�
l���*��&�ǽ=�z(b�&Oe�n��0/V�J��D#w��)rk5&�x���E(����ڴ;����� qk����L�8���E�@��ZA�G�FJDYswe�=HH�uRe��uT�Ei�H��@��Jb�څ�%!��vof�cA�>��&�I��y7�8K���Ag-Q�'(���ft6�EPah8y' \��&�1��0Cc+L$uFv��qڕ:���G}
� ^l���T/�Ȝ����L ��ն
ZH�����Y���Y�nS���ĨG�0N��X��x��9B��U�(L�����^�օ˵k2!�%�BȜ��s�2��O.]��A7�`C�h�; �X����\�*]�P�JO7��B��9&W�F~Rᒧj��y�u%*m�0�6d ��M3p��0+f̩�%΍#����ey��(7N(CR�˞+5Ě93�p�q�ȘD�:�:�'�B�ӫ
6����Ux*j�ӨOP�[��?V.��QU�&%!H����ɾ��ѓj�Q	X��b�b���@�HD��0N��k�+��O 	���Fa�ɳ�G>&m��ʓ��\<b�q�'{|�%��Y�#J�}���j4C����(𭂸E���ڃ�'_*�]�� s!�#dM��Ù,R�8�A��$Qv���9
��m���]�B��<� /��O(���֟7
�����H��@)c�R6')&�Q�nF�<�*钔"�%��dq��do�L� ͬV��T�!!U���ɪ(�uR�C�<b'OA<~4"?A5��_"��B�9����i�黎��b^H��1끍@�"#���o��8����A�2d�R�%8G�dʡ� ^�ɴ:t(�;�,C.-N �V�Ѐ.���)���D ���$�DT
!	�?m��B�I5��tSS�^?v���ˇ��U��]uU��a�'��aʳ��4ŀ:1�X�1D.?^��kEFIAְą�I���0	�K�^X ���� �F*�zu�A�09�p��.}�Ak��Ҏ'ay-�4��u�n��f�¬���ҍ�y��n��*��D�_�"�
0�>�y��P]��A�a?Rif3'gП�y�I�"Gx�e�EmD�I��ģAE0�yK��8Ȟ$z6JX�w�2���J�y�@���|�ڲ�b�&����	��y"l@������1K[0T�$L�yh� 	2��3&��A���"���y���$�&FW#]���&�y��<P��)��0��0Au�C�y�O��%��Z�u<�0�n\��y2i��Y��9bAL@����D7�y��P�C|F".]�5m���J���yҫ�.$=Ҡjŀ&9�Hj��ּ�y� �>I��%p�N�+5���4*Ѹ�y�� *yȀ��D�'�<�b�d�+�yRc�a^BI�p̓p�p�rB��yB#��P���׋{�2mR���y⪛� Op�AV�m��H��
V.�yR̝?r��k�D�l��3�b�y��S�ol�AB��g���	���y2e $M�v�C�ʎ�c]�hR���?�y��͟*9�d��dOU/D�*���yR�F�%+���W�� _�Hs�I9�y�W�?W(= �� `<��إDڝ�y�EV�U����뜡&�@��ĎT��y��z����A���ł��y��Q��U�d߾@X�J��L'�y�K�~�ȭ�g�	�e�Thc�Ӑ�y���vGpUQ�HE�IԺDRp&3�yb��pԼ��
^�+%�5�F腬�yb%�$�֩`���� h���Q��yrm��� �xf%�1A���;�⋲�y�֏<�X�6� P�QJC�yB�N�|/txz	�B� �r ��y"Ű���2t�T	Mj����NQ�y���8��J�M�, zAA�	;�y._�I��!Yv��=�t�X���y�@�eOfӏ��Pm���	]�yB����4kl�D��d��Y��y2nM5f � ���D� š�E��y�f)- .��� G�S���B5,�+�yRK\�b�	��ػ{�R�KĊ ��y�f�9Pv�,�G��"�AI���#�y��Č;���K�� ���ĵ�y
� mi��z�9C7��E\FL*A"O$-��$z����ޢP��"O0��Q�W�xR)B�S:@��t"O,��ck�^�����'��1�g"O�q9���{V���3�D��ɢG"OVh��G�_K��0�N�Y-f�"O�z�lGl�Z��#燢%��Z�"O���]�( ~�(�Q ��hQ"Oj��d$Ǜ��(�'�J(���"O�@�%��)��0��9�"Oe)�₣0�4����`��Ѣ�"Oĝ��#N,��!c�ʢZ�:��w"O29����ʐ���&'����"O.�b�ĕh�n���"Y._'�<�"O�ucTdD�Ad����6��ʣ"O8҅mޮG��dR�%r/�!�"O�XX���S�2)R �\2Z'(�q"O���B�C(&��Y����%Ā �"O�aЛoQh�#v�=�y��"O��&.�9G�*�{��A�;���8"O0L���N�,��!�w�L68�v�a�"O�uH�ȯ_����l�S�x�2�"O8�+��R�jH���<��5�"O�B�m�2�f�jB���!����"O��%�f3R�JP��؁"OV��S+CM�X"�*�lou�c"O:���-M�>u���ޖL�6 #""O��Z�`)��I�ޭ����b"On<!�G�m+�9Bg%�5
�����"O �x'�C�^�t��	��Z�ڔb�"O<�[���;|<$� d��+mw"�q�"OʕX��'ZHy�4%Ђ q~bS"O�,9���8�2L�B���jfT}S�"O�P��k�͐�b��٦X_�D��"O��h5����N���� Jy��"O��h&�Ԅk-���+�D��{$"ON����N..�$��ĩ�-�x�"O�� e چ�r��E�@�4�Q"O�<3Ů�W촶R�Y�k���R�"O��H�b�OT����>7W "O�L�ׁ���*aā=�ݸ�"O����� iz� V��u,����"O�dH��9(Ҵ�&O=w"=��"O�D����&�a�X�tY��`"O�ܺ3���D���1��bS|�@"O���aՋ[�T  ��U5�P5"O�<T%�Ws����f^�Hx���"O�,�u"ۉQ���A���|��@�"O��Q��.*� Ț���2� �s�"OD�(N��
Y;D��Zͬ�8�"O"�C���K3
�	�Ɨ"?!"U�w"O�� ��9�L����)+�Ef"O�M��ړ@�ZJ��=��`"O!���FcF�<[w)R=o���b�"O^���4�fѡD��*̅!"Oʙ�`�_-��p��Е/�i�0"Ot��é�:<��gDZ�	=����"O�Q�ќ4F����#��R����"OdH��Xۢ��W;���v"O^]s$����a1���^8iÆ"O��S6 	�.DDX���-R�z��'"Ox=Ѧ�P��Eق$As��)K�"Ov�cGO��rހ@r��O�)��l@�"O�d�G� �o�fL9�f��iwТ�"O� ���燐7e���q��6V^�d�P"O,e3V)MX]��aqD4+C@I�C"O�p�G)�>�ȡ#����j4"O\��R�j?��{Fb�.z�F=P"O
tAe�=NU �A8�8B"O�#��X&H Y,d)����#�!�DԐ^�>=��\�`Z�8³JQS�!�Ě0Q����"�R;�hC`�^�!�q�����"R���O� �!�$Z���][��P.0^A�.6)�!򤌆IX��A�(b�Mi�MP�n�!�$�3\A�v���0�`�z@J!�R�O�X���-C��.�2����P�!�$!�Ƚ�� �'\Κ�c	۟!�!�R�jx���,x�`�ZC�N*	6!�$E��ؼ �)�$8�8��M�=�!�,4�ݺ0��7�,�T��Sb!�dL�o� �t!�) ���[f�Qy�!�d��G�r ���ш"��uQr�u�!򤅕e��}n.Z��Y򓍙KTC�I-m|� �QLA�P���K��Y_"C�������=/�4@��V&N�C��8X�fkM�a�>�e�S��C�ɿs�
T�WI��a��������.B�	"ЀI�j�5���a@��E�BB�I�>��|�u%�s���	Fi3B�ɪb�:� �jT�n���X���:b�B��9j
5�cI�>h��4I�(F�E�@B� p D32�-j�~���!>�B�p8�@iAN�# `ȹ�I]� ��B�	��bs-nI�S�H�1&�B��4h�0��V=N���(n��DO|~�[�(�����ޙ��1�s�؃�y�Y�d��D(y�����A&�(O�=�ON�(2P�R5l�ѹ��-s��h��'ﺹk�h+h����Q�n�4��'���ⱅƮ��=����{)Ti+�'����P��$JR��`��*{�~���'�L���'@�N�!#�L�@����'$f��	�~貘���Ht%��'~�	E/&�jm��̔	�L�'�"����u��{D�t�>�	�'�:(�5S�=K�<��$�*o�T��'�6՘S*�%8�y���b72���'�X1U P�^��U{Q4n�,��	�'�*�P�gU�EV���#�b�y	�'s��"�F����+��8�`�yR��+]�L�eZ�Tؓ�o��y�E_�c�.͉���G�J<�.C�əL�2�,F�d����@���6b:C�	�r�,QـF�]���	��T<CD
C�	�#�h�t�T�&y��Q�\��B�I�s�.5������#cώ6p��B�	:�P�k��;輝�#��x��C�I�+�U+f���Å�� !pB�	�M0�2 �ǅ?A��a�
C�� ���+����xRL��+X�]�B䉺C���qGٖ'�(A�uD��	�C�	,>K��B�|Q�"�+\�C�ɬgP����>p�ГҬ�'w��C䉁:Zz���f�+��@#��lfB�ɡ<�:��/٨,=Խx���#z##=���T?Ͳ�-C�d��c_]
��%�1D�,��kņRrԽ���� 9�6E�eq��E{��� ����c��HI��mN⬴��"ObѠEI�>K0h:��6g���T��l�g8�4�sA@0*�zҢ�"D)`,˓	)�Ob=�'3���BJE # N\ 1.�#s�pj��d<O��*q��*ŚR�Y�dW��0"O��I�hT��)BP#�NV�Ѓ"O&��ŤԎi�	Rg��'���"O����΍���us$��RJ�9�"O���D���t��-�8z��"O�H��з~/ĴI����2��'"O�0�NLl֕�G1:�t��"OޘY�/��h���w�����
3"O�����8`5�����t9E"O�mص�K�J��{�f�1�m��"OjH��)�2G�(J&[��)p"O�S�ҶiC�xH$�U��J!"O�mP��<}p���C^���X�7"O�� n�߄��#bP̺ۨC"O�y+��]`x���Q��Α�$"O
�Q5���F�|)�u�A�5��h��"OZ<�̟�Q}*��u�U���4�"O��� �8m��X7�N,kC "Or↏�;���Ӗ��aA�"O�X@R�~V��Y�D,��"OЅxՁ���hrF-ן�ƍ�3"O$m���
l�RyC"_�7�B �""O\�t��3���(��J5&���8�"O�S`D���8S"D&��I[�"OlUceLZ�x��(��k��@S� :w"O>�ƨ�+Ḙ���N*;Fyh'"OLp��C���.�2qCЋ.5�e�"O �S��+;��!,X;#�f���"O�	��ː�G��T
X�_�I�T"O���f��$E���q���N.NI;�"O\p����f��\
���MD�u�"O~��FdM�2�åh�dJ\�"O�qz�(D*H,��d��+/�a3$"O�mJpoQ�wk�}�R�"v2��"O>�ro��)�`Ȓc˰r�]�"O(�D��,�����!�P��uZ�"O���S\�;�4D���DCp"ar�"O*����=I0=�/�
W�8�"O�I�T��)P�T�7�P�1~��"O��YgcA�qD�� 1#�`�Mѥ"O(ZP��:j����@� )�|x�"O��$����$�c���9B�ăG"O�-c,�vyJyR��E_���f"Opd��.�j�d���#dH�U��"OL�M^!"2ୈw�>U��r"O(��v ^?����נ:�BY�'"O���TfO���Y�jB����"ON� oא���jk.2��	�s"O�9A% ˨M���Ң�����T!�"OH����+�]sC
]=r)�(��"O�,*�^�?�]����0>*���D"O!Pa��
X����èP�A�"OleS )�=���@')�-E����"O)*@�)l��'�y	�"O��������	�b�Vz���B"O.�W����̉b��"�R�c�"OL�
`�YV��0���a���Z�"O�1��١\y�I��b�R���"Oȸ�Ї9up�02&c]�]��9A"O�I�6�U}y>@�# 40�.��"O� Tt[怂!d��HB/0p߸���"Oh���a�d3*���I�0Ĩ4�u"O|�s�n[]���&���M��| �"O�ٓa��8g���W�ПpE持"O�IH��@(hUrgE�'����"Op鳗��$1�mk�,�Q�RG"O�A;#�Y+��I;�k��cV1[�"O�4�eϋ�(�  !��gY�`ۧ"Or��á� ����QO�7B����"Oܴa�	���΂;y&�+�"O��[?g~��B��|�X��"OTQA�ŸcӔz`垌ߔyb�"OV�k� K%����
s��Ia"O��h��FK�|��� �e��a�"O$=1`ꓦK�F�A�eL�a%^���"Opa�diƥY�xQR"�G�_@F��&"O���"e���A�D19�h�"O�|c���/h�>A���
5]P�rA"O�,��A�6�8䱒`%kB��"Ol���M�)V?L!{�o�/����"O��9�J�����W ����B�"O�i���P��ժ#n0U����"O@h*Q�ks�H3rn��wȐ�"O<��"	{�DP&�חs��=[�"O���fM�7_,$ȣ,3$�fxG"OVh�	̣Fk�rA�8�.83�"O�d��aJ5e,D¢� Y'V�A"O�}7
N%Ϫ�3F�#v���7"O�Ɉ�Ʉ�.�\d�ElպV���"O�%��l� h���F��kGN���"O��
��V'OLq�#V�Y,���%"Oԕ���]��B�['����ɔ"O4��4!�xOd���fD-m�,��"O\����� j�B-�7��w�\U҄"On�
QfY:O��Fo��f��ɥ"O<����!=(j �2a��nyt��"O�p�h_<>/�� �(s�R�{�"OP|�T�Ƴ�*�Jf��x��"O*��,�r�����iÄ�J#"O�,��I�ym���d(
��=Z�"O���Λc�6݀��F�t��"ObE��X�lഔp�nƱ2��`4"O@M;�Lٚ+���#�M��[x2`��"O�#��ݗMTɑ�,A)lt�B�"O�1Q��n��)9�$"dS����"O��+�̼F�>�x�5[a<-�e"O,U욼q���b�_&bJ�૳"O��KT�FUiΨ���[�c>��"O�pbg���j`2��#��6'��I3"O�+TJ�%Z�i �Hc�E	4"O�h�B�O����.S���XT"O�(�d/�-(	 }{pM��D���x�"O��KSD���(1�ܗ��<R�"O�d���K�3� L���*?�p��"O�%��Z�
Y8�cS*����"O�E�Ō[t�T�A3�_3���D"O������f	��OV.l,�%"Or��Ԍ�:r�
Hsa�[g"H�҂"Ohd;���<J�~��mC�{���"O��"5���]DpE5� =U@D�g"O
�Y �[�
�Yw���R�B�˶"OhzP%�UY$9��ɓ�u4���"O�L�e�Q�3�	������Z�"O�Q�w��l'�`��G �%��P"O� `����� X��I���_�S��xV"O��x$��+1\5��T�e^��c�"OJHCC�5j���Ch�]`u)!"O"A:F.��Wvt�R3�^�B(V�B�"O�(V�s2|�(�0�xw"O�IZ�܌WT��C�X�C"ON��Ce�7k0�@��0d�*�"O��f���ҥ�b��iU�`��"O�0�$DJ�y�J�Q�;�"O�@�Ι&&�x5p2h&F�5"O��E]9DY��f��D�rm�"ONw�S�U6�{�duj���"O`�� �.��a�������Ȃ"O����˙?K��P"C�Q�vT�G"On��Un��!W�3R�@}�"O@���kQ-*4�1����ZX��B"O�� 3)ϒo�R�@ ��/G���E"O���M�bXp��Ah²T-@$0�"OaY�%�
[z$i�懏(����"OJ�A�!p �8�a�ѓ���3g"Oj}�&���^���Aq/��D"ON����͜� H����4 �&�IS"O�����G� ���{CF4�
<y�"OlL��C0=d�a��L+z��8)"Oꁣ��	�n�fL��21���bv"O`��F�[�g}��1����%h�"O�m0C&�6.uh� 犿ujz4T"O^���fF�~��pwƂ�#1V�3�"O-9��ķ'�H�a��Ѝ0>�e"O�L�\
���I$#]�Y���"Op��g��P�8��B߹X�"O��
�:;�I3D��"$]yT"O�ti���.h�̬�#k�����S"OBQZ��>Fr��2�j �'"O@,�c�[�&�L+�@�tm��"O��i׾Qf�TX�֑_�.y��"OtuB$��$=� �р�O4�
% 3"Ox�K1�'nI�!���ׯ#�6��'"O�����^�{Ę�u��m��1R�"O a
�-��st�X�F��~�4u�""O�� sI�	��%��ə�l��u"O�xⴧ�3 ׄ�x�̑�H�:l��"O���Ã��n��Eȕd�r"O�Ա5eˎa�`+b�_,,q�"O$��մ\�+$�&h��* "O��P�[=Y��`���rdR�s"O��x�ᐂj��\Rq^%K_N�K"O�Uc�.��I0�d�F�.B�=�&"O���ϝ�Y$��M͒7�,�&"OvYP�mB�N�:}����$~*|�"O�LH�C�1%�ޡ &�P
Ѐ�q"OJ��ᯊ]��!!ÂܛP��% "O��E�X��,]����7��\""O<m�������T���2��Lr�"O@�F�!
�� �Z�{ �c�"OJH�&��?U����i�dyV]�"O��q�JF�k�4eYf��E Q�"O�!����*Ȉ�V�A����"O�����D����C�?���"OJ��U@�J���7v�Y[3"O,��Dq�m�d��vl�ȚT"OT�SEV��M��O$
]�a��"O�}A1*@�89�,R6|GH��"O�Q#��*D�J� s`�.p��"O� Vi�K��.��Tp��Hd9�q"O!�wm�e�ei0o�#Ұ8U"O�x�a�w𴳄��! t.`��"O6�Z��:V{���2=h�m�t"Olu���� ���;��">L&�z$"O�ɠ/��@+�����҆mE��#�"OLt�D��t),*ê	[�1"O���wk�B���x�
_�NF����"Obm#w�W�w�v�z$� c=��q"O�d���V��QC�ES�X8��
T"O�	��ʵ)_��#�9%MXd(�"O�uc��I��*2��jzX;�"O�=f�Ҋ,�Д ���V����"O�p�rkɁq�]�EՀ"�x�"O�Đ�
�Ot%�qn��n)����"O��3�r�"�Ɩ(H�3�"On �u��-���_CuZ �"O�i�͎=}}�t6/�%8lh"O8d�2�L(
�MZq.�
�����"O��"U�Ҩ,�r�x�!<�z�Ó"O�]���[��p�SNn�|3"O�|I����F�Ȩi�	RE�R"Oru�BK�Bfe��<�Pa�"O���%$�)bER���'\ j�"O9r�D�db�9#��ȣb�f]��"O�뤢��qa��9S��f�����"O*�*A#����[`�!L^�5q"O�1���:5{H$e�*{R>L*�"O�'풕{x�H�b��,��w"O�Z�dZ ��Y4oH-m,Z	r�"O�U���Qxp��/��Q)2��"O��+e�'�� ��� ��p=K�"O�b��	#�4ѐC�X�A�t$*�"O���a'��x�>�c�[�Җ"O�L����
O����Ѝ�p%�q"O ��%^�49P�`Y�<+�|Q�"O~��}���gkS� �ح"b����yMė/�6y�@A�`pu�G:�y��H�fAP�	
�L԰��տ�yI�(Wo�h�FF�4!D�y��B$j2��D*�"���f�1�y�kT~'�3E#Çi�<I�-@��y��E�D;��O_�Q`��k[��yR���o\��#Q��'Q������y���]a<	��y��Eh���y���8`VQ{bGB/phV���Н�y�KS�)3�/�z���@���yb)9�� � �	\i	�7�_��y%�)~a@q��L�W��٫w㟰�yr���x-�U`S��4@N䈷�/�y�芽G�Ƭ�PA�=��p���2�yB	SU�!�H�'�y@"[�yRk�i�p��0��T��<�C�Y��y�B�Q(��ɰ�G�W�ҧ©�y�$C�(���ȵ"I�Z=dI�"(��y2��2`�&�
�g�=Ur���ɖ,�y�jP�S��x��dȪ�6G�%�yBjLP�Ĵ��[�[��X⩍�yR�N�W�Y#@BXc�H�!��y�b�e�]�dDT*?Ki��A��yb�_�d6�JG�>�(�4*[/�y2�ˍ-�8 �UFи-�TQ	h���y�A@�O���BS6f��D�y�,^,&=���ȁ9��Uq��y
� f!�"�&8Jf�/x=.��"O.I�� _"y�"��:2���p"O(T�㬕�mg\	Ԉܐu��P�"O�5��C_(`p�${�&����(W"Oʉ���^?{�E�U�6X���"O-W���jiT�(`c]�8�"O���BQ"3�<�y6��n�E�R"Ox�С��\� ��!Mj��y��"Oza[�c��X{�ɀ��� 5	t��"O�%(�CD-S��Ź�KŠih�}��"Ob,h�;��؂Jۦ@wj5PS"ORi��1V0�8bj�qe��"O�%QC�[~K8t��)�~�pMQQ"O)��i.P���#����i��x�u"O�����@,C��0JӅl��@��"OD٦#F%E6�d�*=�x�ɂ"O�yW���A�rP�I�B~n� �"O����!^�>�T8;.K(}&��6"O���$���L&�zR̄�4`8�"O�����ʰ߶�w��=_M�i��"ON0� -��(�^��+N�8@fl�"O�x�Ɇ���bJ�G��,�C"O��q�گ@iR�(����Se"OZ`��?!f�ɳ��L�2�
!"O2�C�l�?L�n�����|�z��T"O�}:���*1��k��i���XB"O�#g��,A���8f$��-��C�"O�ñ��3P��lj�@�aE9�"O�$���v�`��7��/G����"O�� �Ϡ|���d��m�-�"O��[��J�o;Rq ��"t�Qh�"O���r�ĜL4�I��˨.���"OJ�k�ρ�1x%M<P�� 
A"O���f��ZԒYx�,��ɋ"O��C�g�>s=bh�q���+o�%"O~ڔ�� K��r�ZN��"O�4�;=B��AI2H�	*�"O�T�$��Zψ)��b�:�����"OzM��"Ǉ}sr9)&b��(�~p�"O���7��<�>�Ҁ�H:s���"O*�� �!���1`���N�F}2�"O=�E��;�8�9��R�k	Y�"OZ`�Q�B�N�@S���Y[8#�"O\ �'�"f
�4(V8V����"O�@��iZ�fX-�e��A� qyP"O��`�W�0��Г��%1����T"O^���(Քs�*��b*H����"O�8c=S=�K؄%���A"OH-�!��-6#ص�$o�3c���"O"��cf�*m��%��οE�F�"OЕAV3S���A�LM���p"O
�Ӡ��n�hE[$�ݱIv�EF"O>�8��«{` �B��8cY�%"O����Gص%��#� Y9f� "�"O| rsh��6&���s *����"O6�Y#��z�X ��/��W|hY�"OL8+g��	 ��G�F�hƕ�"O��Z�`�f�KP��=}�"O"��bÂ�u�$�h�+U� �"H�A"Of�����l���ҥVp��j7"O0�I-2�b�8@��L��s"O:�����rl��$�:��P�"O̱3�)ߞc:��&�9$֎̱d"O�h�bD"G��� ��_�9�V��"O� 0i���;��i�I�e�b]�"Obl�5c��^8x��=Y�0�`�"OD�� �4y��ɴ+B�9�>�	"O�ң�T12�D��ՄU�e��d"Or|"Q�-).� �)t^����"O��
�Ȗ_�pEJ�-�35�A�P"O���0����|x��[4" !�-
@��R��5{Y�R��=O�!�'�$�V"�	�R�� ޞr,!��ќ&���"�D����@NݲD=!�
<�-�-��F�i��T� Z!�ċ<���������e��hE!� �C\�=b�iC1Yy�I�¢A�F1!���tt�@v�Q*LZEۗË�8�!�$̇I�Uic�Ɔ12�Qb�H�E!�P(�jQ���� ��O,r!�]�D�6�'�;5�4Q����z�!�DQ�&3��K k�5�^ �ؽj�!�d�)�� N�U��`�r��')�!�7iq%���O�>�hf	�(m�!����L���K�/�������w�!�ą)e�x��g��L�At�I�!�L�U������
wF4-��F�s�!��N-pS4�/3�� U$�:Q!��V�|4�4�K�w�`�`T9<A!��A���iC��4d��qD��>!�DԴYD�yJ�E�D��� I!�������ӯ_�| 
%k�G;W!���~��a"�ׯP�ƍX��� L!������4�I����j©7�!�$�%`��,�Bo���,|s��G>�!�d�%�l�с�j�>����O�!��K"�Р޼%n�8E-֧&!�Q'�"=�VJ�7:`T�����/!�	?���Qw���	)~Pq��)#�!��>XM�Q�fLGk8XL1c�0�!�d�Q]��a�k�?��g�Û.�!�D�6�z��b'��FBt%2��˥*g!�7;xr&�	O?@@:��y�!�IV@��zj������g�!��p+�l�d'<(�Y�&�Q}!�dD�>�2��4=��@+�%��|i!�ӱi�h,�pΜ�4$�Y���V�!�ĕ��V�0u���X�� S!�	�R�!���Bː	��l
�<�rAͻ�!�ߗ)7Ȕ��ĕ�����=J�!�D8(κD�L�@.���oT
q!��Ėw
�Kff�5V_�	�$1!� @�4�ʆ�'p��dA�!�F��B�!$�<5%vYC� �%�!�$�	R܄8���?�x&��@�!���YrfA���X=VL[�MK=
7!���}�U���:b4�R˘�O!�,&xp�G!�%''0�@��!�X�<ڬ���V�@�R��a�
$g!�D�&��X��<lq�$-�Mc!�D��l���S��T;585��R�d�!��C�1�&d��"ι �٥,�<o�!���AA��pB�0L	��u��e��'L ��5t^6�[6�ܴ<*Tt�'�\xɁх^��83�Ă�H.z,��'����� �5�I�K��x�
�'�L� 4�ܼG{��h����L�H�K
�'F�(Q��,m��Is����	��� ��k��?i�� �LE94�l)�`"O]�C�#�`��ˍ�	ɨ]�U"O6���N��Z5�'J@8.��M�"O�!���E�1���%�(kE"O�8���ؙU!������l �|�!"O�0�i�>nS���$���-�"O�4y�E�=��"dĩ`���
�"OT�h�ÑS7h����O�7
�Z�"OrT	v�Y7�0c'�L>g�L�R�"O�}IUɀ�L��s��RMd0�"O���@��"	y��2t��>2�(���"O���!��H�"�7G�0��"O����T-�� ʣ\���""O�|�W�� ��L���F���ہ"O��Z7br�͈�3����"O�,����[�t��ə=|@0��"Oƨ�wn��ș+��3&�吗"O�%�Ԉ[�~-��8dḩ&�uZ�"Oz@J���=0��ȃQG	�	j���b"OH�8%�DŴ,��޽J����"O���,7����+�)��"Oa
����	��E�!l��æ"O��JaÁ�$�\b���Z��p"O ��T/�_plԑ4�
A�"OV��,�0yX����4ȴ�"O�5���^�K�������3��"O�ђ嘜q���+; ��81"O���	N�����	ƭN����w"O����D		
J1A��D?�� ��"Ob���<FB1�c��-�0��"O�)��a�>�m4�ғ�<*U"O؋�Oڌ%��ja�ɦS�Vx1"O�%�s�Y8)�A	�ǲ�D��"O��f�<���Bq���Ơ���"Obˠ�Q�:�hSFN[#����"O�q�A��u�����Ԁ!Pm1"OT��4�"��VA��G2��K�"Oz񩔃9��@�*� g"OV��Ƃ��4���W$���"O\�
t�ߑ>v������xq"O����*��
�j��F!9�t�92"O$Hb����H��!�o
!ld4{"Oj�HF�ڐ7Ҧp���Ώ*fP��"O^���Y�J��1���pK�""O��G�4�N<�q'=-r��"O$Հ��,�$�u(ô%��2"O����ܢ��$��扨�8��u"Oh�ȅ�@ˈ����C#�H��"O�m�!�S��Ȼ��ύ�(��"Oq��	�$���"$D"�<��"O�}�2n�01�}CD��[��X�"O4ᒔ�]�S,,WA��q �	Q"O6Mq�'Ɂ٪�ѧ�/F�5*$"O^l��E[C&aR�.C�4��"Ob5)dDQ
���/G ^X��"O��!/�.:
��2fo�dFh��"OF�Ç��&&�8b/tS��+Em"D� � DS�+�}�ӭ6Ɇ���!D�0�"FH:*��D�)�-[����dI?D��fL��ZVd�;�f�m82y�Q�>D�, T�"gCX	�@ә�4�cra D�X�� H�:<�%A4\� o�3í>D�H5+�HnH{&�.P{�l���<D�y$Łh��DR�S29DhPAB<D�� �ȋ�I°("~���=)�d�"O.Tb�k��3
��"R�z�@��"O���EM�Q���&���H�
	��"O��!�@��TpȺV�U�K�D��"O.�١�[T�L!�r�J)�Q�#"OV�	�!�1H���!M¡a�¼�"OdPC�*#�R��wK��=x2�A�"O ���Ί�;v�<���]f�E["O�F`L� AD H��W?Q�q�"OY�+MB��,S��a�
���"O�PĂ�q���HdZ��l���"O����Z6'^=��,A��5[�"O>�`֙W�T��dI��t*��1�"O��	�`�&^�P�C�ľ7��b"O������*� ��ꖅ_�~��f"O��[Dgƹ&�V	���F���p�"OZ�HǦ��kD2���/�2���"O�a"ō  Z.��j�d����"OpdJ��4���.-j�dx"O�գ3l�R�lÅ,߼?���8"OH���,�Єk�v�L�n"O��!�Uc�{�	��A��"Of���B]>�d颳���4��"OB�+��Â?$Ȅj���U���"OԱ%aG��!Y���&Ts�)1"O�4�%��b�0��6'ZUD,M��"O�����[�kw`�B�&��+��Z "O L:q�h�0�+�,��[�b�"Oj�`���=����V=J��Lu�<i�B^-
ش�p�FN�(.������i�<��I�Ftaf�_�jD����n�<�e�R��H/T�'��SQ�<a�����~	��F:?��i�F� O�<���-�phQ�mѵ[;�,r��U�<i���~��$��j�.E��)�w��g�<�q�U�07�P1��F�t�����D\�<��#��E�f�Y�[I�AP��q�<a��K#qR�}�",Ҩl�JI�@� c�<v/n(�NX��1,�w�<�WBS&.5p�2bC��0�nv�<񇪇1���s�o�� ���
&Ón�<�6�w�@�Qv͒�8�F$�Bh�<�˓�z4�4I�� 
�<F��e�<���6q���K6杊r'��0�@a�<�� �;U�^l�.[�wG� �/�_�<�C��C
�]1���<E��*U�Hc�<�2��q^Q�`\�+$X�BcI@H�<�A?�f��ѭ�<Pn���k�N�<����4
�}����r>	���A�<9�#S36QX�U!�,���#A�<�b
�'��+S��7�Ԕ���u�<��E�,Q�1Hpf�9D���sA,K�<��	�*66�T��e�e�g�VE�<1��|'�܈T)�W���W�J~�<Q��W�cD<-�F�&���Zf�~�<yAk �r("��\�-<��)eUu�<���%]����S ׄL��%)Ms�<�5���d,;��j>��+�Jr�<a�h�I��l�N�(X�3刐q�<�RO� 4�x��f�_�J�^^B�,Hz\���F�S�T��ț���C�I�{����,ٍ70`��a��=��C�I4=Q�mYgL��(��ש;\C䉋)^�A��d8D����,C�)� q�H�AD�*��D�A[l���"O�5A��U(��]�#aO0Kb"O6<i��<�@(y􀓰g1P(��"O�����\�d9��ϞH�Ͳ�"Of�� %�������G_"P:r"O|��LX�pQia�6W&�A�V"OB���6 ��2D���t��"O8tf�9��s���o9(�Zw"O��)�!��9k*s�>0���"OX����h�t���)4��ܐW"O��	�>��	�"%Ɣhv���g"O�����(��㈵J�ra"O���
g��ȃC�X��|"OT��EX�q~d5ku�
�j�bц"Ob��фO� ��.OT��o�!�D�@)�ͩG'H1oF&�i&̒�U�!��M��g�E&��E�J�t!���>��LHq�X|y
�	 =
o!���a�n�UJ`_B(�5n�8b�!���:���Su�y��(#��<�!��K//z�)���k�r,�#+�D�!�d����xl�Hj��㑊�S4!�Γ<K�A��X�b�I�T��	�'�еPt �:@��Kw�\[6���'^HIӒ(	4Cr��3[�8��ʓ6נT�B�v�
� V#͟Li��ȓcJE��JB�o� ��P��5WN܅� 7����E >v��#˕�D^P���$�b�Ef���q
�*@�V̅�og�
���o��Y'���n�����~ x3�ӧQb����!�|�����j�T{�j%X��,���|)��"O�Ux����7J�L��Cǐ,?8!�$C���D�4�M�����ň�%@!��ǮU��I낛��k
4@>!�$ָh��x�GI�B�d\J�(��%B!��2k{�ȣ��Վ	D�ً���)(!��@�j��al�34�Ѣ�(�v!��Ԓ)���'*	�,��#
�&){!�$ފ;����R!A�<tr����!��2M�м�Ҡ�l�����(�5�!�D۷a4�auc�,|��TqƈD7s�!�Ě!Ҹ��eI�'{�j8@��[�!�dC�N}��L�5i���G
&SG!��W�=�Ԭ2&j\SXVA�&E:9;!��P�Kjd��&B��v씌3��n/!�N�v��$�gW>nݲ�Yʐ(�!�d��p�ڬ���ι��ȇnu!�$�n�fm���-DQԔ�c��0(�!�$�1B�zX@�nғ���c��4cq!�DN7I8��+@�W�#��
��ihC�/��: ���Y o�2�fC䉂S����iQ(x�l��(�g B䉮\i���B-�>4S L�`��/+ŚB�ɫRe����1L$Q��
Z�dB�I����dȁ�%��;��ڽEI>B䉪I�Ukю��L,�[��>�TB䉑a����R�!Oհ 2���0&�B�I�g�5Æ'ʾ��0SP�U�E�nB��%m��h��l�tH���=#|�C�I�����0J��0^�I�l��C�	
sS2a��$��HuL�SteܱrhB�	�F�i����T�F���,)u0B䉍E[��R�@�4�F��	�B�)� v�r-�4j/JQ)�%�4G �r�"O�8@��Һ^��tb��B?�2�g"Ov��	�.HH��AΎ5s�eʓ"O�X�O",P��1�
e �](�"O�0�"��*S�DI&��j �|z�"O��2��%�P,#�E���B�"O(L���4)v�5ۥf�dh\�"Oޑ��E�8xR��h۲rf����"O�� ��ȷm�4s�E�o��D�T"O�!��������� ��"O\�sA웸"Z�����M��ـ"O�uZ��-`(b��
i����"Oh�jŎ�!f�P��+�+Ag���"O����
Ǳ6r���SK�*�l�"O�1c��:TW�y�@DR?:�lkb"O���Þ o$%Ñ�V29���"O��ÂI
�+���-y t-Y�"O�$��K1vl]�pK� ]�đ�&"O�(�ǁt���k�`��n�H)y�"O�\��ʆ)b��a��w�����"O`%J��s�.q/L���f��JW!�D���Ѐ;���>.v~�B&�;^W!��Ӗ+��呎(_�ա�G�==E!�D�.B�\S�$ԓ.}��� �J�9�!�DLv��e��E:C��k3дH�!�$B�1���GoX�)L@IũV<H�!�$�6_V���\	���H�a�"t�!��ػ;]F��j@�%h�]
Q�Θ3!�<����hV[~q���/"!�DD+_�m��,�Hb*�k���!�D�s�)e�%A󌈐��L%O!�$�!%��=��mS2|n�EY9
 !�$��"i�"�R,}!@��<ȞQ�ȓ27�C2,ٓAD�(t�c�q�4D���&&�"�^�U �:Rt�"��6D���I�!� ���*3O:�	�
1D��1q�,6�b�K`���%�@��C
%D��z���hN�E�aMQ�'*vM��L.D�@衎�&xQ�8H��@�pͰ�-D��P�S��B]���dH���)*D��	�IT�"���Z�R�+��@>!�$�'k(�:� ��d�L�/!�$ʻ[}�сE�.`HD�o�@�B!�I+`���x��޲Kό�:�31�!�{`��eް/�x\Ӈ*'2(!��B�g����ѺET*���ˎ�!��T����fYOp��+��5J!��P�q��yP��6&�}�3e��iH!��\�شƤx�m�p&�?'!�d��;���X�f^�c�x��CD�d�!�D��g �Ey%O��W���pޭ{9!��_ҼRR�˭ez��7Bÿw0!�$���j�:iN���>`�!�$�/��97��YL�A)'o�>�!�d>_pt�CS>$�!V'�&v)!��Y�, cQ�HZ���"�>9!򄘘Z��)��	]̕`�e��N%!�d��*�ҐF���Dq�D�T�!�$�:�T�%��*��l�գ�!�����ԡ���B�$P�Λ!�$��L������(�Е�g�6_a!�$X<��P��$���_;@T���
�'���;A�	6��W��78لY�'b��V@W�N�8������(M<���� �xg�
�X ��9EIQ!3J��C�"O�8�� żl��y"��ݶ|HlH�r"O<9�u
����B߿<�)g"O�ݒ4�v��Lc���&|:���"O8�Yώ3��{�O�U�<�ڡ"O�B`ܗX ��fN�0p0�h�"O!���]$�!�d�_,Dn�5aR"O����m[1BMj9R�#���DI�"OB2U�A5Tu:)(RG x��R�"O��h$�(y�h�į�+���"O
�KŌV�w�p�(c/%�^!D"O�0Ir��9_K��-�>	�t{4"O���#��4r�ݱSM������A"O�hDH�2#��<�&̊Yܔ9�"O2$���� ��a LU)V��1�"Odqy�j^4X�Ҽ뗩ɾOȬ�17"O 8q��.c��g)�~K
8�"ObQ�tC�R��`����	iF�[7"O:U�u�԰<��!��-ƀg.���"OdH�笔�9�b��a����(�e"Ob(������K��q�]��"O���F��G�-#P�C�^B��`"O�諥$��d��(���;$T-�0"O4���&ӂ6@<l8�o�|`���"O�ede���ȓ��OQ��2�"O4�A�*�00�՘��H�C��J�"O�d�"�M��:!��EN�ˎlJc"O�@k� �6��� A�h%r�"O���s�'t�B(81KC0\��@q�"O4�i�#-H� Uqr�"O�ّCe�>���gkƑWn.�7"O��ap�M'B�Xx��*��xa6Q� "O�(��P-*ᶬ P	��O?�a��"O�}1ׂK�uC�E� H�U�mj�"Oެ��;P�X�(4�����"Od���Y� ��mr�*�ʜc�"O�B����Hy��]���"O��%m/�*u)�hU�N��"O��1�!Z;Q<�X�G�x�Ta&"OZqYs�\06�
5)����e�"O(�D�k4\��%(3Iʔ��"O`��b/�T��y��ǣD���"O!貀�A���#��h&�A"O:�Kӷ"����S@��Y
U�"O=2b@G1��PK2���dm��"O���g�H� ���?Ю��"O6e����H�Se웊U�.���"O�%�c�НX�P��d̆�@�"O���_1j���*�ꓩǾ��1"O`J�H�P��:a�3/Ȱ� �"O8��UU���
Յ�G��2"O��3��qKr5N6�Y�"O�ه!܄{9��IςzHୢ�"Ou`�
�tj�I���ݤq0� �g"O�QDȋQ%́�7�9c+����"O��C��Q.�걃acV�o��]Ps"OPɻR�k:Y��(��n��1r�"O
�Rk�{��|Z2'ɘ1�:�K�"O������)LCD�aыuCb��"O�P�p�ί}a0� *B�83���W"O��{�,��T0���b�<@X�""O����C�e���"Hu�D�"O�r&�ڑD����/� E��t�P"OԵ(�3@E ���g5�"��"O� T`c^c\&�5��?� ���"O8U�%%¸E�tPKE�5����"OT9k�k��A��K5�u�^%��"O�dB��ϻ�j�ؒ���F<�"O��Rv@��0�! ��Σ�<�IB"O�ݺk�y��(g��b�iQ�"O8�Z�nJg&�h��"� ��%�#"O6�0��O�Q�:�7��.��y��"O�CC)�(�|��χ�>����"OR��O�� x%Q ����b"O����C�9��(����	�"O|Z [X_�l�G�Y�xt�ݪ2"O��C/��T�����B�t"a�p"O���4	Q;��|�!G��2]I"O�-*юR�b0Flx�E�(]��1A"OJ��0"�`���
 }��y�"O�h�����7�"8���)u� ��G"O�]�(a�(�'��z���"Od��w��:s�X�gnU�W� ��#"O�y�^l�J�,͂M�N��"O�Ժ*�& I���B�Z�.��#"O|)��)A+=���"�Q�zgzmQ�"O�=kq�C�+i2%c�. �����"O:�[�H�]��M��a�0�ʙr"O�0듉
 za `��)���r"Of�je�J�x�/[�OĄ��"OaZ�
�"��/� O´�3"O�����;y�".��RD"O�(H���J�^%(�풠3�${D"Oj����5h���۷U�I'(%At"O�1��ʀ*�f��B˞+E����"O�tS��Q$dR�5����H=��s2"O��§��&b�'_�W�l��"O��C[�!r��"h˶i��,`�"O�A�N�>xF��t`E!�"dl,D���ÇܞQ�^�w���C׺Mh!�5D��C1C�'�$�(�/��D�aQ0D�4�݈&�Ex - �9�i��3D�(y"M�[�@*�`�N�Fh��!=D�8!���OdJ�H%bۼC����-D�8"�
]l��v+1	�&	��`,D� ӵM�\dM{$�D21Y�,D��ӧeE!,�:��2���B�ꈘD!)D��Je��� ����5�_�l��%D��`�1�YJ����n|:E?D�P��n8j6����$�T�dd>D�$91�:�,m:&�(0@s!!D� �d✆��l�s���)�� D�0Ң��9��,p�D��/�権G�:D�4 �㏟2�|9C�Ҧ0���8D��H�A�?h��-�TA�3;�0����+D�i`�T�D���2O�=N����E)D�`�1��>̰�i�C�����!&D��e�NI���G��l�$E �%D�dB&�ԇS&�qqI[-��h���"D� �c�
b�bs��'�¼yA�3D� �,J"Xp��d��?=X��#&D�l�"����iyEN % l9�F�%D�H�&��oW���#14,92�.!D�h��M�0�"��cLٌ+���U� D��"�%��(���kY�A����$:D���sn֡z�p�*� �n�$�w�<D�4���4s���T�M���sp�6D����#���f�sd`^Y��ʷ�3D�� H����xW|8��̑{1�=�&"O��g��[�b�YD+r�"O�h�&�:6qp�+�v���"O�ؐ��*Akx�**�=*�`Q�e"O�UX�'���&�[S*+a,�"O�U[�Ɓ�2-ؼjV�M�k���Q"O(��Ǭ�: `f�c��A�|��4"O&�0�˓�)�8��VE��6`�U�"O\ݢ��JdNP���I#	A判"ODbg�4��fRT=X��"O���r������ǻN0VT��"O�� �ɟ_#Tܓ�'D�w �xʄ"Ođ����"Κ��5G�!;�d#�"O���CAU�nhE+G�b�څ�A"O���dJǳzɊt�'%�5>S:	��"Olہ���=h��Cۂ
4i "O�[C�?;h����j3(�CQ"O`��`A�6i��Aӡ&d4�%"O���#��d�"ݓ���hN��@"O�ƕ�+0&�S�G&f��-#B"O�����H!b��@)��f�j��"O�Hf&�W�6�÷
��L���
"O�%�E�ӄ�|��$��*
U�E"O8��q�8@TM�'쌁f.�h�D"O��Z��L+jR(��j6=	�p&"O�9lH�zA�S��8 �JPz"OBDє�J�P$��2#�-h\YB"OT�aC�8
}��ȋ1-���b"O�yA
�}޾�h�"ߟq�4*`"O�e���&T�
%(���z�{�"O�K��	/u;�|�ā�x�.�"Oh$S �ʗ*�$�C
��9n��d"O P#�`O([��`�g��-���p�"Ov�D@�2��
���� �Di�R"O&a#ң�*0'��w�V�`r"O�xHT�ՙq�^�p��4��a7"O����,]�'
f�@���*M�F���"OtA�r)�p�p8��C�3�nB"OR���X�,���Y�E�x{ "O�!�5�H�\�zdP���<ol*��"O$hrt��>e`��P���12���y��=Br��#�֔y�`t2F.܆�y�
g��Q#�%i($yyV(C��yb�J�N$ŀ@㌊K(�aY��y�ɞ��&�x&�&8�61��� �yR
3B��a1�؊*EH����_��y���>�M�*,)Z���v$]�y��
�@A��EVjԳV۲�y�LW=}.��呣D�T�a�H�y��R�B�,�!�R�xβ�4N>�y�#��%\����[鰵��&�y�L�(��D4DQ �P�[��ڸ�y� Q_$�����rA�BM*�y�#�1 b��&Ù��J���
�yr�]��I���7}�|���I[��y��Z+�q�B�n��8���I��y��ٻ|��YK2j@�b�𘊃B��y��D%/�=kA(#Z+,�2H��y��2]���B�Rl����*�+�y����=*`���Qc.��e U�y�  �D-��#�"%Q�����˰�yBb� J0�p�#�u�h����L�y��R�C"\�ak��n��$K����y���mM"��D��0]��U�d�M3�y
� �Eʷ	,rD�D�\#~$I�"O����g��QОHBRj@�+[Tq�"O4u!��
/�t��\A$qy�"Op�1��9*ڑ0$�ό@P��"O����IW���cƍ4b�VX"O�#@�A�ln<T� �}O�Q��"O�dK0��s �P�g��E 2"Oȅ�� �23�.�2A�3�"O�Q���E�T2��0nH�O4��Bq"OIQ���!���2'��{Ҡ�	"O�( ꎫ~.���_1Dܖ!@"OV��q�V��6q[S�ҩ�D0ae"O���)�O¤�s�V����H�"O�	��$N(kc����꜆%}��&"Oy0�dBG��޲r�b!"O\HZ�%��v����K�UZ�9#�"O2h��MR�NRtK�
؋iJȀ�"O �s�NCN��s�d>$D��"O�B��R�zE�2�W�#Eb�YR"O�D�u#A�b��i2BEߓk�  �"O����A��bn���a�.VVYIB"Ov`���G�s��/� @�"Of`ۇ�Q�p�&����<D�"e"O�T:���61��e� n��R�"O�M��ȁh����`��C�^Y"a"O�D�F�M�*���r����}�fy�4"O�MHB���I�1�F=	� 0�!"O���&��9b0�̞�!i�"O0ʶ�
���Zfv�p�a0"O���������q#8*j�(�"OZ�8���["�Y�6u$.M�"O���H�#�����?o	�"O�D�G슺B�6�P����	���87"O��ֵK�P �bOV	#�-pE"O6|�A*�s���gG��8���"O�9R�&P<`����s����"O�8:E��Bf���󉙑�D�X�"O�=x��H�$���z�����y�"O�PaG�jw�B�HҼ[lEXu"O��)D�S�3�z03V��T� )(�"OmPEcE�7i��q'D_.)��kV"Oxh`3eAB<�C*�{�eI�"O��2����Y�D"�I�q�����"O�(���xi8� �����"O&XAQ$�L%HХӺ:�ڤI�"O���JV�8<�ER�D
�s��8��"OR%���d�bc�&��!ۡ"O���n˩M]@��#c�;E�<�ɷ"O�I����g����0��
i�z�"O� �E�� ��8�"Oܝ�&���"O�����ȣ@���"�M^�y՘���"Op}XG�T�L�*��S-,�>5��"O���QI��~�(��RT�"�"O���)îg�Py������6"O��GH�"%��p�眇Bl��*E"Od����-%�V������])�"O�r�I(T�<�sP���@����"OZ5���1Xg^��6ڼH�*�{�"OF�/��	h��T�p��H�c'ݻ�!���(0Ƭc�_�6���!g��0�!�d�T���2/O*�Ҽ+�جMr!�Z�>6D=ɲ��"r��uޯ�!�H�]. ��mD�)^���'gk�!�3q��Ї�"CV������+@!�� *HADW�_N(��S=���G"OM*���R��%swÓc��aZ�"O�U��c�*U�D�ɥ!�~��:S"O[�
�A��aKP�1��Cf"OQI6H�{R�L�ɋ�MT���"O�p�&��6a���H�jRp�@"O^\����� <@�E�+؅A"Oꄊ�#E����19 i��"O�����ǫa�wd�E"�鸷"O�耈����X��aԻ9�h9�"O�HZ�`��V��`��/A�"O.�:"O�ó�D/II&P['L1:3"@�"O�ũ�!�;sK<�5��!��"OR�іa�-j̒�K�ܪUf�pC"O���O��'�&�{f&��&���"O���h�>g��j�n���	y�"OT
�%];C8Y�O�;k��m��"O�ui�K�f���Q'$X2x�Y��"O��@�e� =�l��"�	
�6�+�"O ����9VD���	A�H�	�"OPd`�N�&GY
Tb�yd�
p"O*��@D2(bak�BJ�}��İA"O�(��d��X�H� G���;'"O4��䦖�1FL�[F]�&�͠�"Ol�	� �1�l�'��7x��� "O>&��lI�IܖO�P ��"O�D{�� B�<5YÍ��P�+�"O@�i�"S+轋+�0�� "O�iۄiJ�X�:|�B	?\V({�"O�-Q`�̛�Jh��.| ĭ�"O�d�a��> 1]g	G
��"O�Ī��!?��y�D�=MjMK#"Oj�����S�ZU*��"-um<D�0BE�۷vWZ4�"�>)��8$ 5D�D��ͨ�e��B�LK����%D�$�� +3H��ZR���E�H0/D�C�I�H�T=��X|m��g���$HC�I2$�lz�,ےkG�e��&�/2ZnC��.�$<�sF�1*7~e���A�~B�1|���ìsS�"�U�E�^B��`p��`ʛ�'�T�"F��K��C�I�
��� �V?A����s�/#[�C�I�"rx����4JV���ׯ��}�C����Ƞ�ImbR�H䨏	l�C�+�(B\�
:��M�R|C��@�B�vkP��0(�7��	�fC�	v:fы�aU�	��A	�B� &� C䉴
H�H2*\�ҹR�l٥Y��B�I0HxE���97�2�K�B�	�:"I�7�XI��S��!P�B�ɐ	�聈��z/H��C��;��B��5Y=����B35�6����-�$B�	�l�z�b1�X���i2�,E&�C�ɤxK�!�6ZI� ��w��#=i�O�"}bGP�PO�Ցe��/#N�BZ}�<�CI�T�
�I�%��y�>�A��w�<!f�+�]�B��)34u9��v�<��ɶ_��M1�·}���gH[�<��ޖl�� �/D��U �	Z�<y���P� t��k�W[��F�a�<�)9eB<Ȕ�0"��9å�G�<Q�i�z����OժFZ����~�<�UO#�L՘���&KX��k�$�~�<��䐇I�S'�2�Jl����C�<� 
H����d�$�̻t��0i�"O6�#f��_��8"%�6'���"�"O�'`�x'|,��J;*k^\��"O�u c �ZtӤo�uK�Z�"O�{��\�T(��/2.���3�"Oԝ����̄�b6���M`h���"O|��1lF��	��
8G>Q�
O�7��:a$�8�-@a����F�^��^���	#�	<FBQX��:M�j H`�<�{��S�[x�R�	�Zt ��� >��C�B%0� e�*W�#��N�NѢC䉳t� }!1& {�- w�M�R�hC�	�:�`Xi2�	�`DD ����? tB�	yM���Ųs�"�˧�Jl6B��<$�ND��Ƀ5�PB�����C�	5%�Z �ֱP��@m�7"~(C��Qrg��Hnh<h����\�q��'�r��p�X/+��q�䀂B^��'n2�S!�_���T�t�D�D��Y�'S�a:�g��4w�t:�f��"O�c�/�O�u�㛫m�d+0"O�e��J�jB�SC[U��0Ðx��'�X�D�C>~X�
Q�L�QD��'a�F'�L9P��E��y�J�3�'{�����L�:9��7p����'��Ջ6��Ă���,j�v	��'ഈ�7�_�p< �V�D�`s~-�O<����閠,5�5u�У������ǵF�!�Y�a����"�1b��uIV!�F=���QB�Ry��\�+�!��f�:�s.·PnĲ��üo�!�$��/yT��D
I:G������
.]!򄆡&�x�� �?)��Ű�q���8O؁C���<f�Q�s���8������>�]Lx�Q���0xґ oұ2DI��M�p�ڽ ����2.
�3���@O�<A��D��9Qb>��hp��� "p��\�D�YeN[j"\���^�$��D�x��&(����0�G��_��I��QL��@�XNE��#�Ɇ�y�ȓB�a���u�����Ff�z��C�f9�@Q��H;q�20�ȓ�d��a�'n�hd�iA:BU�ȓI�hM�Px�HU��4��$�ȓX�@�I��2���pe��*���ȓ0o\1SM�#F&8�� *|�De��E|6D��EW�}�ք�f�ʤ"�z���e*lbe �E�- .�N\}�ȓ_�~��f�o,x� �j��ȓ ��y��)�5S3��3�*�6`c��ȓl�l����C�tz���1U��e�ȓ{9b/�2�9 �G�P�0q�ȓylE� �G�e�u�C�D�oQU�ȓ*��*eo٣`8x�i�-��deV=��!�ޕ3�kF7��ᄥ D����f�����e_�t���[�FsH���?�~d"֥� v��)�9xH���a�@�d�1�.�RsI�=�ܼ��O�H��o�]��qa�I�O��]��S9V��% ��wD9JdB�m����ȓj�$�N���Vܩ�Ԑ���cܢ�C¥)S,�ɗ�Ő�\$��jt�d���ρ{f%� M��>�ņ�?I� ڢ(�*��iW���X���S�? ���2�ƝKB�<-Fn�1C"Of���J;1��-"���-H�}��"OMj2�??~�� @�U��*�"O��d`E�&K�Af�x`3� ��ybC�_�uJd*	�@	CE�?�yRᔵ#�Ҩq�M�kMԍK#F��y���&_&�)�75� ᇊD��y��O�F�r��*'"v�b��"�y��^�_��m#�++ɼ4y�
N/�y�%B-��Yڱ��(d�:�#�y�d��4�`�hG ��S�|*�@[�y�ȬXxiv����:�ؑ�ü�y�S�2#�ѱE��#A� ��yB���~;N�J�ˋ�c5j�Bف�y2�_�4�&�)mMI� �zr�T��yb��� ���V߆�kQ�;�y���z�"x���M(;!^9B!���y�h�6O�1�R�T	3�^ai�œ&�y�B4M�
I��NY;L
���F��y���*Q�ʨ��^ے<�uFQ��yr�/o5
�ѷH R�J�I��Y��yb�	�O1�iXt-]�?^qUd��y�O�8E:}a4��</`J�̏��y�1-����G�O�9�(�s.�>�y�*�&8��r6�ɺ�-�����y��4 �;�/�>M�v�(�y��::�sáM�
�Q�!&J�y��5���GM��$y��S�y���h[#̴r�z����A��y2�ҿ�����"8��2�$�&�y�N	9�p
���=~�i�P�'�y�F�>\_@頉�1�f����3�y�hH)ת�QǍ*uJp���X��y"��%4���1�%Տk���t�B��y���apF�YS��gM����Q�y�@>.�(��gF2�HR��߫�y�$�Sz-�El�"a��#����yS�"�4P�%*O�i��;4C�"�y+O�a��H+����HA����yB�7:��J�l��5>���V��y�	�IV`��F�P�/��E�a�B�yGE��LOżs��K$ȥ�y�"�<����EK9(�ٻ�"î�y�<K`��c�ᙳ#^����7�y2"�3G����0��������y��+��8y�A°��������y"�7�`�Z(�pB�j
��yBk=�B�F��Բ0��L���yG��B��K�'��L�RE��$�yr�O�F�,��"�E�I3���$��y�JC@�����ՠF @l�$f��ybf@$W�T�*�C�h�zՉ�/�*�yR@�)�(0����Y�v�@��?�yrH�.wD4z�� Bn���A ��y�7h�J��P��H��;�y���6_8�@q��:H��5y�J��y��ҫH%��_����q(��y��\0Ph� R�[�$@)p���y�N�TW���&�ʔ��2�gг�yↈ i
`C�y��8�ׅ� �y�NCE�%bk�v�AϤ�y��ؐ,�8$�M�*gz@r lY��y���J�t@�ׯ7�l3q�
4�yҎ�0xn�s��q&8��2�y
� �����|)�<�u��- Πd"O��8�
U�>p8�k�W��PB�"On�C �P8!�J����;o�5!�"OF��:�*�m�*x�,�q"O�];$B��(��1�&-�@�x<ے"O�8i���I�´�I�-��)�"Oq�sO�}��p�クObV��g"O�$��A��O���F?l^`�D"Ov���$��1������G;�Ƞ"O��6%Ӈ+���C-���`�1F"O d�(��9HH�2U*K�����"O���pkѕ{����˚�S�~50�"O�9�4`A� g���6ꐄM�|�I�"O�q��@�2V	�b��7@N�(F"O��2��NP��0H@���V"O"Y����t��3�拂6��d"O�3P�د{W"�cc݃kz>�)T"O����IC�̺"��t��e�c"O~�իJ��()�A 1K���"O�}#6FðO�|��ѪK�piYQ"O 5"�3i�>�D�*p��L+d"O"�s� �Gu��#������'�|� �)_�x���EG9os<0h掎B��Q��'..�S0�Ή~�����6U�1��'�̹ȷKƂ��D��H����	�'�옻L Q���2UR7�<�	�'��Y�e
��[]��쀧�BL[	�'~T|B�O� %b�!����b	�'���Y��L�v���总4���Q	�'�
i &��&�,Ջ��=��`��'P9Åi�-_���B	Z&@p�5��'8H��KA Y�u��J��B-��B�'�l�f҇e"���$��.9���'!@����Ky����
��t�H�'��9�M�8y2�m	�@)L�l��'�8%2vK\8?�A�#ޞᄥ�'����3@R��TƨW�n}��'L�P!���4@t�O̷E�6�z	�'y�չG�9@�
��q�M#�' 52R�U�A �i
���4�`}��')F9��%��W�!�g��q��}��'O,m�7�G a�z��%a	t��'��W*�4[�P2tFʸo���+
�'�i��[�E�����]�lB
�',d��J�{mx���g� Q�.(�	�'���Z4�Ɉ2���W�q�~8��'}�5�$�_����J�q�j���'j��1̐�a��t`��#r�#�'�ջ�J�/�a1�k��|���'(*��i��Z}��bbJ�FȬ�'�����K^LS��#H�.ܠ�'���'����@o� �b�'=t
C썠-a,l⠭����'����T���aj���;����'��M��I�c=���� ^�����'7<��D9I���fŔ'���{�'F*|�#��8�iv�'96���'���DĤ}V������1w� �'�pq01J&rH����e�@�S�'}ִb4Mā3/V�Yq�R<Y}��x	�'��1�W��GF�I���9��'�����)®��5��G�� ���'P����ڊ#���D��6�	c�'d> �&�`X��B/�GYޱY��� �:��G'�Vi��.<�5��"O�]j0�&�r������b��"O�{��B�1&��X���:{� ���ϰ&�(@�=���ON�#��8z�)��$��%0��)F��S� �7l����-�;:`z�HY�5*~<����Ms'�G-@�!#�@�^%��-��i�R��--k��U�	2\ۘ<�hE|?y�/!I������B+���g�u�(�-.^F�1$�ȌF�a"ŧV"pD�C䉄Z}���!K��ЃV�;��_a�fe�!M��!��>��i��ep�E�#�Ӧ�a���
 �$5�Vʜd�]�J��H�a}¥9;���a ߯b�T�%$:L���Bˇ�NŲ�J��N�XA6���� /���	����b�Hf�'����N�Tf0h��M�)�ny���S�C^H�hn+�?�v	�W�$�:E�@���Vb2�"�a�9[��}
T��Dr�pV�*���U�'PR;^
nʶ�I�fžsp��zݴcB��+1�X�9���D0V���J��X��u�-��0'��#�U+*��	�b�Ӕp4T
˥z&�[���.$<�K�*Dp�l3,O|�
_*��Q���n,� N�
���\�If�@.�\4���A[��i�����M����e�&��˔8n�r,���� X)�	*N6���jG�̰=Q��$3N�x�I �_M�-9���QQ����
Y)y<åD��r�L6m��v�P!#�B e���SB��
��lYGOu� ��*���#����V�V�:LA��#=1 ��H��	�@a�OP�"��� �J\�$nC�&�� as,�7�^�isoDPS��d�'m�m��b�(?e�xP*�O��i�FXn)X��f_
��D�X���3�S+6�ͳ�n_� 8�Iȿ�2U�r�O��q�B-LB��Ӎp�h�����|~A�Ӂ��v(�e���8�#I
9�0�� SXz�(a��'8��������$}��ጰC�LiA ��<�6M�T4�V),* �	�*U�BaM2A�IE !��<:pcC8L�D�0�
_�2H�+�:lCbIE�Q����	�(9v�;d��;[�6�IB�I/h�I!1���B��J���F�+1d�c���_�:��~z��1p�z�e�%:$d�u�AI�<i��^%{�L��A��\�88��b�ަѳ4o�+x�&�A���Z,�K?y,r��mH �EB?YC���j}d�Iq�!� c�*^X����wf��S�ЍI�i�g���,]�MW21z���������2t��#@IK%C'��+���9HS��
҉�?
j����0{��6M�VC>ّ���3<��IV��j	O�=j7��b�LIi��KE�����h�=� 9���+ Hl	
�;����$I!�"%��0=wPɺօ#LI^H��E3op��SG,jZ��4�d� òiq���'�nS��D�E�H`�Ii��b�� �HB�y
����Ra c�.0�t�d�Z�ӥ#�>���)2
�-swH��r�����m�nI©�6��Q8sW�`C�K�H�֜��,�M��`��o�fA0���0��M�'xڠ��kܠmR��BS$�r�ܚ�4u�p�K˽Rl����X[��׹�u�/T�!�:��weV�M��E���#��]�Y�2xP��5�T�#8Э��-�a��q3%�z칐�M
����K�J ���A���@�a�*7f�8��`�~���`͊�M[�L�d�4!�>���oQwX
GbY[��=��H� �����,V������� +b�B��P5��Z�		.�>�Kp��-`�Z�@�#�.D��6��uR����[��|���(�R?�;J,��R��"B�DBы�+!��Gz��$zhqi�џ������w�MJA��<��T����K�#L}�r��(�	N��Z���ٰ_�tRF
~v���1���(Pń�i�� �Ā���L�CtӮ� c�Ȑ���hRl�"���"=�֝�% �%[����K�Q��ܓ����ceO((��'��CEhX��3�-�>�ҡ@�:6{�`*�Ҁ=����pi*ʱC��J�Wq4)�s�m�A�ԊGæ��3%���"-��� ѭ �Z�J��dn8��}r.�	��9�������$}��E�t�ŨkT�h����ҿ\W �d���Tu�' �񘆢P�83�)�J�n%t����$@=�Tb*O�x;�k���*v)�!xu�#O3G��(�����aqt$@.,q�͇�	���MaĊêN|���"§]8����
{,&tҭOp(�Õ<g<U��盘n'N�""O��J��-'�]� &�*��IE"O6qH�❐3h��R�O�~`C�"OΠIQ �%�R$�t�����'"O܀�o;t�]�!��]����"O��ڰ�_	��8#�*nۨ1�"O�)��g,*�h�Oߥd��PC��'��mڃ���g�* �]�T�X�f8C�	\�Z@�@P��1Y��Y�a�C䉰2.l[�$VA�YR��B�ɻ9t��7'�(0�&���Fƕin�B�ɼCȈU���;Z)mց*sټB�� ��!S+�0vD�೑�խ9hO���w?\O��j1 G��V�+�c�C�Hp{Q"O�-���X��i�(@�`��l��"OT�!�	��AitE�^��2�"O� �y"�oM�y��M�;�Mr�"O$����ݎN�v�!�R�vd��R"Op�;'��7)n�( ��ەK�����"O����?w�q�F��M!��x�"Ojp"kE��h��%p� %�"O�r��-Ka��b�ş3�ڈ�"OrH�c��B�:��w�?�Xp��"O����Z�Z��j�B����"O�(yW�W���a��+;"���C"Oāy���
i�N�*�ҏM��I�t"ON��m�&caN|#a�I�q� �	G"O~���� Jڬ���DG��P݀�"O.P:bbK
v'(kD��>~6V�!"O�A���A�R �@AZY�ܢ�"O"����O7�a�V�Ӟ&Ld��"OD���L&��ȈC'n��#"Od�@�*� Y�l�%ٕ[$fuj�"O��`��3>�v�y�G�%L ��6"O������Hl2@Q��-!tSV"O�P���2)'b+�ˏz�(:�"O��Rj��0�&�����1^�T�+v"O���b %@YH��RP��s"OZi3�K�/�h+� �fٰ �v"O��e�*!;n����R$p�V���"O(t�$���1'��B�!0����b"O<�!�O�b���ġ�|t�a"O���U,G3�ᵅ�{jEIp"O�)�ׅ�Pؠ�ԃ�ek$�%"Oʴ��98%��S5�Q�Mz��p"Om��OS'u�Q`�A76m��I�"O�1��υ9C9b��ޮ!]X�k�"O`y�@�Lq$<j �=X���1"Oh�#3"��`\#�ȅO�}�&"O A�Tl��4�v�@�X�R��"O�3b$��%Z=cs�Ϊ���C�"O��!%K@R��y���Bx�A9R"O8k7꙽Rі��,�?z�p�8�"O�� ŝi��|��
]��~�Ac"O �3�X�g"᪱iMT� e��"O�p�#��Q�z3�	 N��""OB���Ig]�E)��FX�ډ9"O�us���EH���0KO�H�+3"OR�����N�l4�t�ݘ$F4X�"O���D��[N0���5���"OL��$��	���6+F�<� ��r"O2x���%@�QШ�g�X���"O`�+ �G:?洀2�,�Z� ��"OrE{�,��`����䄱Or�Iڄ"O6�BW�G%�r��p#�_h�S"O�]�LV"�<a �@�/Z����"O�!kc&�^�>���Ɔ
��S�"OĴ�S�z���Dwd�xw"O�T��B0j��B�J�g�
��2"O�$ u�ͬ��ģ��a��!q"O�c�T����"�QY�"O|��7��PJ>������"O��0f�6K��⅚.nkԐ�"O���OuΜ��֥52�����"O��` A�o���	cƕ�#����`"O$e�S��=LTv�0�"�LtrQ"OpptHγK�񳤡�5h����"O�}�ԓxl���OC�w�2f"O⽻��Օ���ag��Lh{�"OҤ�!�&��T��:;��8�F"O� `uJ��݈U�p������"r"O�(�#)W	=J��p1
ätZl�x�"O�Z �@�'�ؕh��iJ�(a�"O�=Af#3����r+�-:�P�J�"Od�"3��de>Ճ��/Rw��C"O^�"C�I��H#㌷T>�@�"O:9{�,L�s6CM�
8�c"O"�1lZ,k2u��cɨt��Ţ6"O^m�ԇ،2��u"q�=���"O�5s��Y���R�Z�F�� "O���B"R�Q���]��vQ� "O\)���� =���pJ(a8�"OX��Fϊ0���P�˕�}���Kq"Oh��RJ��X�ֈ��,��RR�1B"Of0����x��M�
C��A�"O���'?U���:��ք^�� "O<��bo��l���6r�2 �F"O�``��xHg�Q�"i�`"OR�a&BD�`$�*�
��	�"O̰����¤��A�d])WKB�i�!�$R*l$��� �̞3�Uq�
�&/B!���'�\2� Y�	��p!���K�!�4Xa`�ۗ+I�7�)��2~!�D�1j��D���)PU�P�W�Ћ-!��2"~ପ솆
Jh��+Z�t�!�d�;��elB�4�" j���!���s~�0mn%.,8�@K��!�čO�ܵ0c����X�� h !�D�*�.݊��M�B��z���%w!��]�֝�SlǞ~��B�OR�!�!�"/\xC�P� -�c.��M�!�D�*+�[�[��<K���i�!򤗴PT�Ȣ��Rb�Q��A^�!��I�*�R�'�y��[�%�!�DF�Mh�㌆8�Z\���X�!�0Pf����?�Jգ�h�?C�!�LQ���re�O0��-���ގ#�!�$�5~��d؛	͆��D�Лd�!������"�`�Fm�7aA��!�D\�N��BC g�,h��S\�!���34���iv��.l"�R��@T!�*@߲�a��{��1�T�1!��˴I�T4��!� I�w�J�S+:C�ɉ@M�ؠ��;S��p/���
C�	'n���Q#AӅAv邕@�!~@
C�	>`�P�=c���3��7"�B�1b欑h�,i� Pk�B�	�s�����Z���y��uC�Ƀm��J��R��=�B�P;�B�8]\P���_
5��:��T��lB�ɕ_�yJ��ӄI=�y��E�="CZB�I( #�C!	�|I��P>< B�ɘ&��m�"єƒ�8�@N�	DB��	i�<QȔ�r|`��R�<T�C䉤Ǻ(�Ѕ�-+�"���+1��C��nTT���k.$Ȑ�}[�C�-p6���./O���DP(M�C� r���nSl��+�h8��B�	
�(��֠���+���4�B�I�1�����S�'a���P!K;�B䉋H4艑�HE��h�U
z�B�	�o�bP�A_�P8��M�&B䉨~���r�� _�2�	[R��B��
T�T*q얰z�:e	 f��B�)� ��`���
А�!d֟���K�"O���a�;Z*y��#Aڸ@�"O���3(�������ܫ~z��"O�I�4Ό�S�6I�fE �!�*�u"O�KǃH�P��%C32��y�V"Ozd���
�fW��!%�7�f"O�܋�&�;�0X�n�"]瀱�0KL�9nF��=����O�s��ű
Ӓ���T�d�P�@#�I���E1��Y39�����4���!��*U����fBkµm�39@pi� �Jp8�`�0��me�đ��D�x�ڹ�¯�O
��	k�L��y:H����?M�'b�=O��I��7�T�1 Ưo����R�L�@7FX8"O�T�##|ҙ9��$o-��Y�
�,?\�'��@�]���L�0��Lɲ���ap�*m{���y�k@�z	4��_h�U:�����>�4�C5-`�sB��"���J����4��ײJ�iJ���,%.X ��I��MK���?��d �{T��
P�\(�ͪQ�R~[,Dz��A</�\5�2��� 2i�+ċ�M��R�عq�a�6b�]ak��z��:�nA�@�nQ��Ґ�˓a��9BkH�vi��C�2)���oZ2>@|=�n��9A%�4w+��$Vк[� N���a���2��h�7�Ͻ.�"����?]F���}R���#[xia�.�2�v!c�W�G�D	�!�#��0�j�(�!^tuI�zӸ�BfP�?��2=~!X�K#w'�Ek�EN�0�^��䋝yit�
&g�. ��1�����@,����+#R�#��܂=
�`ܴc��8csE�*~���/�L�ivȋ2��?mr��������i����4đ��1VA_5�Bi�B�'t� z���a��h�EC46��a���Vl0p�Y��M��C�28Ixk�� Bt$Cp�'i�p(@�������_�5�صP��F)ؗ蚞�~��+6k20gڟf��w'+w(Z�3!��k���Pz�c#��np�F�!��z�A) ��J�,#���i|�8�2%���_K���EĢ>i���+&��b�$}�;�=�&��_�� ��SUBV���>����� ��XpF��$��d�����˂0��ӧh���@�J�hq`�g��k�l�hA"Ov髠�J�>���9'F�'w(8Dj�>�S��L�^h��$8O���
ΫzZ��8����q���'^�i��ߨc��С%�߼&�&1I%���[�,�yFΏ]<iP��($"�yq�
i��cbԦ��"��$4/
\Q �@t}r!-(:�!!@
B��w�~8���J] �8�OK.�"�&�
�jn�ƉRf�"MPX4ّcΥ��up�-(!g 1���đ1�H�����$(��*)���!ן���Bdt*� �'Vy|}�G���� � #Π1=�x �'�:���2�"��,>��KFK5���ط�ї�M��@z�`�H�F��B ���'FlP@�%&C�UR+)0H|�ߴ$��d$I�INf�D�L��� @��u��ғ[�F�b��M�B�L�9xQM['lʨ)sE�s�,4��'.
�*&�1�F�;փr�R0��x=j�C_��-���M* ��01��36b���4e1<�y���y_75�|b��sqnEm�t���d�%
��eFF�w�H�eǅa���d�ˢI��H:w���0\r|8�F_�O��6-қJ���f���õi�W��������c	����u͛�z�����u�V�zPF���'�b��&MX�Y'v��'�X3V��u(7�ؙd���i�˛-b�![,��ty��YhK�w����dØ	���1f�i֔y�����a�#0҄�AM��# ]�4.9⁳�z\�L�>b.��w$����]t�V������	�'}��tI�E��S�`Uz7�iAƇ��B�ZpaPğ�v^1���au��\w[ ᷾i�س����h�$��F�J�@*h�s��Ex��3,ڄC��
��%'h)�6�-%Gl\C�A��DB�F�i&��Bb�'0���4��"<91.J!d�f�F!K��z�fG|b"ܔCʾɖ'ц����O4	 %%H�Q�!�n�,�{�4&c
t���#�p>�fD+�p��1��s;��V���
���BA�	�]�\��s��=q�&�1ᧂ�`_�B�.T6Na寔�z0"��d΍�E��B�	�7��8��� �$�,�r��	,�C�I>~�x`I�Z�A���!�<�HC䉽=>rh�Vʜ�X@�d���evhC�I�5���=~<��!�=\�C䉢R�����j	�S"���C�q?�B�I���Zt��._��E��ߥ!B�	�C��0*7�W�u��ؔň�?�
B�	�716��e�I5c|�J�N��C䉉���acߙ>��\x���@�C䉇C|��)M�$����ǪBP�B�)� ��p!H���<��(�D=��"Oj�Q���!K��eG��]x���"O�M��ă�w�T4K����h Zv"O��ӆCR���9���ї_��=2A"Od�A%L�)ޞ}�` \}���a�"O�xsՋlȤ���ح=����"Oh�����"g�lr#NG��0�"O��
#GB�8���'�V��"O��h�@��u�T&�Wkr�y�u"OR@�vЩ<Р쉱vG,A�"O�t8`�	�a
'%@m�t"O�(``�C�,O�7��X
�d:"O��"�a�@���O�m
,b�"O�����L&��@N�'����C"Oz��-��a��;�T�*%"O{��XRҼC�-+w����"O�l�r��5{z�yT
̰^��]q�"OhY�e�Q-�H����{�=H�"Oܰ�#��)��{\ _V�9"O�|2���6䝺rg��aم"Oz3c& L�Ƶòfݥ1~U�u"O�A"��n�z�ɁČ�w8\�w"O�1{`�A�R��Ģ��s�V��"Ob�J|�� uU4"O +%��pM�d�N�{ԍ�F"O��Ɠ�-��36J�.Nb���W"O�e١)��5i��ڦ�W�։c1"Olh���8BH 9�F�4m���V"O�,i'�ׇ;nX8G��=^n�y�"O�r�Hܕh�����Ü?~H	5"O�d`���b�dP C1
��yQ"O��p���
/u���C
�#�����"O@�S鋫L�V1 �D��Ӿ鸢"O�\�B��/�0��J�b��Li�"Od���D�mǨق���(.�x�P�"O�чĜ�L֢�G�F�w�ѱ�"Oh���I@7��A�"�)!"O�sdI��0	̗8��Yh`"O�Pb�@��>��DL΀�ZI�3"O�D1�ED5��r�eM:?Μ� "O1�ů^;�4�N�X�\��"O*�:׫�4i��ꓭ�..��a��"OB�{a��+TvX��]�U��h�V"O^��&�^,.�B��k��:A&�h�"O���@Mݽ>wf�j����=Nlh�p"O�P��
_���)��L�}�f�ۗ"O�8XG��V�nP�6���?�*�0�"OJd+G曠i�&��WKU�U����q"O����̜(!-Ƶy ���x1��"Od(;�KdE�!�T扫¶lj�"Oa�%�4"9�q!���?V�T��"O���#n�CE&M��;O��4K�"O⨘W@R�ܻ��1 d���"O�8c��כ	��0 EE&>���Q"O0J���fG�b*��0��b�"O�����&n�x�11���Al.�ID"ODD�c��J;�I�C��<h_�Ҥ"O�̀	�P\�i��H�p]D�br"O���H��A�B���ᕼ,����"ObMUO�3f�B�ď�	p�"O0=���{F���߯�Ĩ""O�p��5FX8� ��)B�-�t"ONI+a���	L�y��H���m�&"Or��ʍ�i�^I�G�"=���[�"O� b�2,�����VE�_�^8��"O�Y�KD�3��,���L�O�8�#E"O��C]CY�8+�n�6H�� 5"OX@�a�����bƈݔe�x�8�"O"ܻA*��z�dY��?��"O��!�e1��ax�ˈ<DĊ��#"O�X���{�P�p��1;dl��"O�kc���!@��C��	�g6]�7"O��b+S�7�ȋ�*H8T� �"O�Q��d��vC�Уs�N���Ah�"Ov�kԌ�7���9��K8P `"OH�a抜�\�x��L1(2́"O�${aL�������i�5�V"O�Z�@�F�8�#���T�����"OlX�1�-3�ՋV�^*-����B"O|1J�̚7|G��&� 3��a�"O��UÁ��<�a�
/?�9��"O��6���LLK���o���"OP%>B(�DЌ˸0�j��"O><I2�˰+�(�m�9���Х"O`\鴡:�R�)6�Ňv$䙶"Oҁ� ��2���r1�U�}��7"OJI�E��>Hs��·in���B"O���^�����i��,C�b"Or�M����0���'O�<��"O��صA��. F�B��*��U"Oָs��@��\�T��1��
 !�D�k��G�]#^Ѳ@s+E�(&!�
K~�җ�E�vx�5�ť�=8!��.H���� 'Jg@@Ie���a~B"
`�n�;�Z�v�(�LE54��,�A��y"OW
B�VPK�).���:A���F^~�� ��~%���S�y��aL<��S�fʸ��Ύ�q@��	�
�Pa��˺��Ĉ�OQ�T�T�OC�@�r斛n�t�TH$%�h�z&Ĩ>)���&ZA -1TK��E�b�����M��"[�)x.�HR���t�@���j�v~��T�褅��y��	�6
�TM�}�(�k!�F�{d󄞉A�VIه���(sX���a��=�T�H�e�7C1؉:�����<b���ɂ�Oh�eI&��!��(����;�.��󄑻�a����<>^�����RLp�^��'�PHx�#��0|��=Z�TI3R�\	"=�xQ@M~r�T9Ex ��yʟFXQc�<���au�	 \��̊Ն�$�rׁ��V�����,Xl:�ԧ0|:���!�n��S�Q��DE���<A�?)Z�HZ�lQ
�&-�Wϗ~�<V��;��p�������R�<Q�[/dTm�b�� m�T@�#�GC�<��-M�lz�s� �E�|�Ys��Y�<��aۃp�,u)p郕yd�y�(QU��hO�Oq,4җ�r�U����-��[�':TUia��x��[��ҳ&�8�Z�'����G�;?����G�$�x��'���S�D����]8!J�.!�"�C�'`)��Q�'r��K@#��m7\���'|�Vi k`��3� 	�c�*%��'�2� ���p��x�A��oI>xX�'���C��֑z����ưl=���'��|�ŀ>?����FG�f�����'���If���Yl�|�#Y+�h��';�-""�̯c���U,a��a��'��5�qk�?b��m�s�]E�!�
�'"L�3�Զ2(��R�
�7�dH��'�� U�,�jiS"n��dd�3�'�>����M�@7����ϣTzU��'��SӃ�!
h��.8V����'�tp�v�V.c�� ��4q � ��� ֭z§�&!�<���Tʈh"ON4[ ��&���i�Ol%��"O�����6�$Ru��6e^�T��"O�%駇�x�L�b��
4"O�82��5z�#���[��d�0"O�	[���#}��	9�� ��f"O�Tˇf�v�(����/���y�"O���FRb@~7C�Z�b=�3"O�D.�9�r�Bu�͒]>�a;3"O����үs�z�@�HÛq Ω�"OL)!�c� #�B��B6�M2"O���`�'	����I�!��(Jp"O�%�� �)n��:T�'�X���"O�2`@mN���G���XZ"O���D�q��[��^���"O~(���GʘU !�N���@�"O�1�6���@R��f��&�*""O޼��
/8L�CfA����B�"O�*�"�/XK�thǥT(�\�	u"Ov$����^���A+8¶��a"O�X�/S9=��al�=U �U�`"OH!"�KV�y�~t8�@Ϗs����"O"4�D�D>�F�B��s9�U�s"O���Tc�i�
!� ��w�tr�"OnQ�dh 	ߨd�dD8���"O���1*�p�J�@�#��!3C"O�|*@fY�C쀩��B��B��T;�"O��
�6r XE]m�f<�"O��A�[�g���a*\�Z�Ƶr�"ORy�p�� f��d�`�<}��m��"O�mxGgG)=Qh���j*x�`"O�=�h�T�b��F�H*f9<qV"O�Y�a���X��7�/<tI�"O��� Т�bh��ҍ,'Qz�"O��1`�	9S7��ѡ#֕&�tc�"O� ����|��0���-E��2"O�a��h��|��l�����"O�p֎&t��=��gU'>�r��#"O�1��0!(�U�W�� �b�qF"O�A�Ѕ6W�@��.W1.<a�"Oj��t�HUn(hwR??��M#"O�؈�l��/��pK�9��QR�"OR5����W_�̊��8{�p y�"O�EA`��p/:쓑��&3���A"Op�s�>�n}��GM� t�0�"O6�HcDڜi�Ŋ��]%?�]1�"OJ]00N˛4r��@@G0+4�Q2"O�L�MM�O��!�r��rh H�"O�� 2�5
!|��U��>s����"O��cWb� -v"���MF�r����"OBE�CG2�	xr�N�+` �b�"OP�񈙴l`�0�WBJb���"O��C���KQʠ�`�%	�pEI�"O(Tk �]=!ʴ��8��|J�"O�u�P�׹4�́����{m��"Oh���$\�1��X�̇.#f��t"O�(	�/ǍgJ��QMH���Р"O�٧���̢�����tmXa"O,�����.�xX뀯ȁg��]��"O�1����0�6�i�`�e�l��"O�-y�`�~����!	�ڨ��"O�T�����ЀE@�|��"O*�{+Ⱦ'�������B雂"Oj,�,U�%f��e	0<��呑"O� 
�c�/�:��PT�F5�����"O��r�ҟ�
��ŁGNؑ"O��:��A�b��i�rN��$Y&��"O�郀�E7qI!qí	�]Xr]#�"O4]��Ý5=��kf�:Z�T)e"O<����M '����v��6vS����"O԰�u�]+|��]��C��;��e�G"O���k��*z���℗��|�"OfM���9E�`�ʣ�)K$�c�"O�P�aA�E�x�	��Zg����"O�s,O�V\#�L�1; 4��c"OT��c��)�x[� Q&��B"O\��
ܝ!.̩�G�%��H8�"O�l�v�L�:!�Q�Gfݨ���7"OAp�S�=Kl�2�B1w6z,�t"OT�1AI3��݋gA%
��"O���Qc��	G�I�o��v���2t"Ol��tJP'���P�ݧ]E.PX�"O�:���>)&m��͏�A?!� "O��9�H�GZ�Ѫ�lW?d��T�@"OmASm�qi����7����"OT��B� j5I�)ެ�R7"O���q�&u�T��H�(~e����y�� V&h��Æ�<x}Cs�&�yR*KU�*��(��9�lt����=�y����z�.}��'կ.�T"ѨE��yr�^"����!�7%�*�8��ǧ�y"_�U�)���E����拔��yrM�X����:I��聦'Q��y",� ��e#1B]F�XUB�͍��y"���N.��C��6@�(�j��I��y��B1u!y�姅�)~�� �y2e�~�"�P=x��=���G �y���%v��gS0a��F��y��1-O����CZm*�+���yr��3/[�]��+B;zx�c�Î�y"-P�l�d1�E��7�� ��y�b��{��4���M�1^.��6���y�E@:&da�9���g��/�yR`�*,�� ��:!�<9��ˍ��y@Ŏ�����d�5$@�%9f����yb�dX��J\�f4���1M�����Z0@��
#jT��{p⑑7�Ԇ���'	Z��ur��X��8�ȓW�,I(!gQ1ҼfN!:*V��� ��d��ַH-8�T�Q̭��C�Q"'��ؠ���#Y�S���ȓj	�w 6S�"�,0q�؄ȓ.�$��C1��5+�aF�=9:Єȓ��y#��
2&�(ۆ��PIh�ȓ ��p�/�MR,�3��"k������Ź^y_���� ��E"A"O�l�"��
hX�� Ĵc�Y�"Oր�tK�1Z���N�hH$���"O��B��T�$u(��� ��;����/!�� ��ٛ�t�Vaߩh�t��ȓ�a�.��[�3eb� g�<u�ȓt�bx96 ��xxly3d앚<�ƕ��gS*a�"+Op�~Q��`�|29��pR��k�g�k��P�ě
��)�� ��9CL� ��!Y���L����xY�1p�]>r��dk��Ƚ	��,�ȓ~�P�eF�7�|��2 ��a�`��@�`<���]�W��iԌ���:��S�? �	 ��_��N�z����k�vy["Oe��̦8�>h��JÛy'�=�"O�[���1'4M�˜/�)�E"O敁%G)r�iU,� e�R"O���l��*�a� ���)�"OP�cv�?����S�ׂ��$"O�- �?;x�4�w�B�̚�"Ob�{q��E���+���i8"O:��Ą�v���5�"*�ظ�"O�ڥIǫ.hV��Tș�1���3�"OhuZg��1K:j���ӼF�n�c'"O���C��7��I���ط8��"OĬ��.���(�%H�?��"O���E��?�����	�R�k$"O$����WY� �(B�{Q"On�0�.�'j�}�/Re�"OP]��W�p���X(� "O�,zˇ�.�$�r��:{%Ц"O&�A�Q4J���q���s5"Oʸ���.���c,�:&Ҕ�"O e�<[d�Ia,D"�胥"O�(��)�?p�L;�X�9r9;�"O�h�F�:+��������XP"O�ͪ4���6�)Q�aM
*_4��"O&������+��JҬ{�"OnQCōC�O���`tI�o=�$xQ"O&��F�F�+W�d�1f�$�`42D"O��Éq��Ѐ�Ŝ"w���E"O�A�c ڃT�m��gV+'��9e"OnD[���2A8lµ��-c��P�"O�9s�'�
fa��Z��U�4��� "O�tB�H]��J�C��.��Y+�"O�%�����A�D�t���"O@���!F�|YSTC�<��qc5"O�˂e�}'���AcڂUf�=�s"O��d��2Yt,,Y�!^�Y}�,p�"ON��ĎE��� 򮜜0i���"O�x�1��0I�dp��Έ�Sdxu`�"O���Sk�.m�����:X���"ON���D���K9zQ�"O��J׃@�~ �p���(>R��"OB��ÏͶS7z�Ə;^��۷"O���MƲqpr��b탻5H 0"O��
�lHiDl�ا̃�-4�J4"Ol}��L�&bet,��Q9�m�#"O�-P�`�T��
]�_+L}�$"Oxi[���� c��9����"O�B۞7�DX�)�)��ٖ"O�� ��ԡi��9B��[��<�e"O�I#�H�$Ap4�]	Q��8 @"O�iA�CI'K���tj�,U��:3"OJ���
^r�1GL2^��,b0"O4q��'���8�*�3�0l	C"O�Lc�]�5H���������:U"O<���X?UT^�	И �FEa1"O2�cVg�*K���ڀ�^X��s�"Oa+�K�&Ў��wC4�j�q"Ox�z�MI�x��yX�I ]q(HP"O�X�.A1�.M�UaG43l�HJq"O��Y�   �